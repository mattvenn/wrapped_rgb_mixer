magic
tech sky130A
magscale 1 2
timestamp 1671027758
<< viali >>
rect 23949 39593 23983 39627
rect 27261 39593 27295 39627
rect 28089 39593 28123 39627
rect 29837 39593 29871 39627
rect 9965 39525 9999 39559
rect 1593 39457 1627 39491
rect 1777 39457 1811 39491
rect 7113 39457 7147 39491
rect 14841 39457 14875 39491
rect 21373 39457 21407 39491
rect 32689 39457 32723 39491
rect 3985 39389 4019 39423
rect 5365 39389 5399 39423
rect 6009 39389 6043 39423
rect 6561 39389 6595 39423
rect 9321 39389 9355 39423
rect 13277 39389 13311 39423
rect 13737 39389 13771 39423
rect 14289 39389 14323 39423
rect 16865 39389 16899 39423
rect 17601 39389 17635 39423
rect 18889 39389 18923 39423
rect 19625 39389 19659 39423
rect 20269 39389 20303 39423
rect 21289 39389 21323 39423
rect 22201 39389 22235 39423
rect 23397 39389 23431 39423
rect 23857 39389 23891 39423
rect 24593 39389 24627 39423
rect 25421 39389 25455 39423
rect 26065 39389 26099 39423
rect 27261 39389 27295 39423
rect 27445 39389 27479 39423
rect 28549 39389 28583 39423
rect 29745 39389 29779 39423
rect 29929 39389 29963 39423
rect 30573 39389 30607 39423
rect 31217 39389 31251 39423
rect 32505 39389 32539 39423
rect 3433 39321 3467 39355
rect 6745 39321 6779 39355
rect 14473 39321 14507 39355
rect 34345 39321 34379 39355
rect 4077 39253 4111 39287
rect 13553 39253 13587 39287
rect 16957 39253 16991 39287
rect 17693 39253 17727 39287
rect 18705 39253 18739 39287
rect 22293 39253 22327 39287
rect 24685 39253 24719 39287
rect 28641 39253 28675 39287
rect 30389 39253 30423 39287
rect 31033 39253 31067 39287
rect 1961 38981 1995 39015
rect 17049 38981 17083 39015
rect 22201 38981 22235 39015
rect 24593 38981 24627 39015
rect 29653 38981 29687 39015
rect 32597 38981 32631 39015
rect 4169 38913 4203 38947
rect 7113 38913 7147 38947
rect 10885 38913 10919 38947
rect 14013 38913 14047 38947
rect 19165 38913 19199 38947
rect 24409 38913 24443 38947
rect 29469 38913 29503 38947
rect 32413 38913 32447 38947
rect 1777 38845 1811 38879
rect 2789 38845 2823 38879
rect 4353 38845 4387 38879
rect 5825 38845 5859 38879
rect 7941 38845 7975 38879
rect 8401 38845 8435 38879
rect 8585 38845 8619 38879
rect 9045 38845 9079 38879
rect 14473 38845 14507 38879
rect 14657 38845 14691 38879
rect 16129 38845 16163 38879
rect 16865 38845 16899 38879
rect 18245 38845 18279 38879
rect 19349 38845 19383 38879
rect 19993 38845 20027 38879
rect 22017 38845 22051 38879
rect 22569 38845 22603 38879
rect 25145 38845 25179 38879
rect 27169 38845 27203 38879
rect 27353 38845 27387 38879
rect 27629 38845 27663 38879
rect 29929 38845 29963 38879
rect 32873 38845 32907 38879
rect 7205 38709 7239 38743
rect 10701 38709 10735 38743
rect 5549 38505 5583 38539
rect 9229 38505 9263 38539
rect 14381 38505 14415 38539
rect 15209 38505 15243 38539
rect 18797 38505 18831 38539
rect 22477 38505 22511 38539
rect 24041 38505 24075 38539
rect 9965 38437 9999 38471
rect 1593 38369 1627 38403
rect 1777 38369 1811 38403
rect 7757 38369 7791 38403
rect 16589 38369 16623 38403
rect 17417 38369 17451 38403
rect 19993 38369 20027 38403
rect 20729 38369 20763 38403
rect 24961 38369 24995 38403
rect 26341 38369 26375 38403
rect 29837 38369 29871 38403
rect 32689 38369 32723 38403
rect 34161 38369 34195 38403
rect 3985 38301 4019 38335
rect 4813 38301 4847 38335
rect 5457 38301 5491 38335
rect 6285 38301 6319 38335
rect 6745 38301 6779 38335
rect 9137 38301 9171 38335
rect 14289 38301 14323 38335
rect 15117 38301 15151 38335
rect 15945 38301 15979 38335
rect 16405 38301 16439 38335
rect 18705 38301 18739 38335
rect 23397 38301 23431 38335
rect 27445 38301 27479 38335
rect 27997 38301 28031 38335
rect 28825 38301 28859 38335
rect 31677 38301 31711 38335
rect 32505 38301 32539 38335
rect 3433 38233 3467 38267
rect 6929 38233 6963 38267
rect 20177 38233 20211 38267
rect 25145 38233 25179 38267
rect 30021 38233 30055 38267
rect 4077 38165 4111 38199
rect 28089 38165 28123 38199
rect 28641 38165 28675 38199
rect 5549 37961 5583 37995
rect 7205 37961 7239 37995
rect 20177 37961 20211 37995
rect 24501 37961 24535 37995
rect 3249 37893 3283 37927
rect 8125 37893 8159 37927
rect 25145 37893 25179 37927
rect 32689 37893 32723 37927
rect 34345 37893 34379 37927
rect 1685 37825 1719 37859
rect 2513 37825 2547 37859
rect 5457 37825 5491 37859
rect 7113 37825 7147 37859
rect 15669 37825 15703 37859
rect 16313 37825 16347 37859
rect 17141 37825 17175 37859
rect 17785 37825 17819 37859
rect 18981 37825 19015 37859
rect 20085 37825 20119 37859
rect 22469 37825 22503 37859
rect 23121 37825 23155 37859
rect 23765 37825 23799 37859
rect 24409 37825 24443 37859
rect 25053 37825 25087 37859
rect 26157 37825 26191 37859
rect 27169 37825 27203 37859
rect 28549 37825 28583 37859
rect 31585 37825 31619 37859
rect 3065 37757 3099 37791
rect 3525 37757 3559 37791
rect 7941 37757 7975 37791
rect 9413 37757 9447 37791
rect 28733 37757 28767 37791
rect 29009 37757 29043 37791
rect 31401 37757 31435 37791
rect 32505 37757 32539 37791
rect 19625 37689 19659 37723
rect 22569 37689 22603 37723
rect 27261 37689 27295 37723
rect 27997 37689 28031 37723
rect 16129 37621 16163 37655
rect 16957 37621 16991 37655
rect 21465 37621 21499 37655
rect 23213 37621 23247 37655
rect 23857 37621 23891 37655
rect 25973 37621 26007 37655
rect 31769 37621 31803 37655
rect 6285 37417 6319 37451
rect 20177 37417 20211 37451
rect 21373 37417 21407 37451
rect 30297 37417 30331 37451
rect 8217 37349 8251 37383
rect 2053 37281 2087 37315
rect 18245 37281 18279 37315
rect 30389 37281 30423 37315
rect 31677 37281 31711 37315
rect 33057 37281 33091 37315
rect 1593 37213 1627 37247
rect 3985 37213 4019 37247
rect 5641 37213 5675 37247
rect 6929 37213 6963 37247
rect 7389 37213 7423 37247
rect 7481 37213 7515 37247
rect 17417 37213 17451 37247
rect 18889 37213 18923 37247
rect 20637 37213 20671 37247
rect 21281 37213 21315 37247
rect 22109 37213 22143 37247
rect 22569 37213 22603 37247
rect 23397 37213 23431 37247
rect 24041 37213 24075 37247
rect 24685 37213 24719 37247
rect 25329 37213 25363 37247
rect 26525 37213 26559 37247
rect 27077 37213 27111 37247
rect 28181 37213 28215 37247
rect 29193 37213 29227 37247
rect 30113 37213 30147 37247
rect 30205 37213 30239 37247
rect 30941 37213 30975 37247
rect 31033 37213 31067 37247
rect 31861 37213 31895 37247
rect 32505 37213 32539 37247
rect 1777 37145 1811 37179
rect 4813 37145 4847 37179
rect 22661 37145 22695 37179
rect 32689 37145 32723 37179
rect 6745 37077 6779 37111
rect 17509 37077 17543 37111
rect 18705 37077 18739 37111
rect 20729 37077 20763 37111
rect 24777 37077 24811 37111
rect 25421 37077 25455 37111
rect 26341 37077 26375 37111
rect 27169 37077 27203 37111
rect 27997 37077 28031 37111
rect 29009 37077 29043 37111
rect 31217 37077 31251 37111
rect 32045 37077 32079 37111
rect 7297 36873 7331 36907
rect 1961 36805 1995 36839
rect 5641 36805 5675 36839
rect 31217 36805 31251 36839
rect 1777 36737 1811 36771
rect 4077 36737 4111 36771
rect 5549 36737 5583 36771
rect 6561 36737 6595 36771
rect 7205 36737 7239 36771
rect 17601 36737 17635 36771
rect 18245 36737 18279 36771
rect 18705 36737 18739 36771
rect 19349 36737 19383 36771
rect 20177 36737 20211 36771
rect 21465 36737 21499 36771
rect 22385 36737 22419 36771
rect 23857 36737 23891 36771
rect 24501 36737 24535 36771
rect 25145 36737 25179 36771
rect 25881 36737 25915 36771
rect 26433 36737 26467 36771
rect 27353 36737 27387 36771
rect 27997 36737 28031 36771
rect 28641 36737 28675 36771
rect 29101 36737 29135 36771
rect 29285 36737 29319 36771
rect 30113 36737 30147 36771
rect 31033 36737 31067 36771
rect 32505 36737 32539 36771
rect 2789 36669 2823 36703
rect 4445 36669 4479 36703
rect 6653 36669 6687 36703
rect 20637 36669 20671 36703
rect 21005 36669 21039 36703
rect 30849 36669 30883 36703
rect 32689 36669 32723 36703
rect 33517 36669 33551 36703
rect 18797 36601 18831 36635
rect 21281 36601 21315 36635
rect 26617 36601 26651 36635
rect 29193 36601 29227 36635
rect 17417 36533 17451 36567
rect 18061 36533 18095 36567
rect 19441 36533 19475 36567
rect 22201 36533 22235 36567
rect 23213 36533 23247 36567
rect 23673 36533 23707 36567
rect 24317 36533 24351 36567
rect 24961 36533 24995 36567
rect 25697 36533 25731 36567
rect 27169 36533 27203 36567
rect 27813 36533 27847 36567
rect 28457 36533 28491 36567
rect 30113 36533 30147 36567
rect 22937 36329 22971 36363
rect 26065 36329 26099 36363
rect 26709 36329 26743 36363
rect 27721 36329 27755 36363
rect 30205 36329 30239 36363
rect 31033 36329 31067 36363
rect 31861 36329 31895 36363
rect 29009 36261 29043 36295
rect 3249 36193 3283 36227
rect 29193 36193 29227 36227
rect 32689 36193 32723 36227
rect 34345 36193 34379 36227
rect 1961 36125 1995 36159
rect 2421 36125 2455 36159
rect 3985 36125 4019 36159
rect 5457 36125 5491 36159
rect 18429 36125 18463 36159
rect 19809 36125 19843 36159
rect 19993 36125 20027 36159
rect 20637 36125 20671 36159
rect 21281 36125 21315 36159
rect 21925 36125 21959 36159
rect 22661 36125 22695 36159
rect 22753 36125 22787 36159
rect 23397 36125 23431 36159
rect 23581 36125 23615 36159
rect 23765 36125 23799 36159
rect 24777 36125 24811 36159
rect 25789 36125 25823 36159
rect 25881 36125 25915 36159
rect 27353 36125 27387 36159
rect 27537 36125 27571 36159
rect 28181 36125 28215 36159
rect 28365 36125 28399 36159
rect 28917 36125 28951 36159
rect 29929 36125 29963 36159
rect 30021 36125 30055 36159
rect 30665 36125 30699 36159
rect 30849 36125 30883 36159
rect 31493 36125 31527 36159
rect 31677 36125 31711 36159
rect 32505 36125 32539 36159
rect 4813 36057 4847 36091
rect 6285 36057 6319 36091
rect 26525 36057 26559 36091
rect 26741 36057 26775 36091
rect 18245 35989 18279 36023
rect 19901 35989 19935 36023
rect 20453 35989 20487 36023
rect 21097 35989 21131 36023
rect 21741 35989 21775 36023
rect 24593 35989 24627 36023
rect 26893 35989 26927 36023
rect 28273 35989 28307 36023
rect 29193 35989 29227 36023
rect 21189 35785 21223 35819
rect 22477 35785 22511 35819
rect 26433 35785 26467 35819
rect 28365 35785 28399 35819
rect 29285 35785 29319 35819
rect 30113 35785 30147 35819
rect 34253 35785 34287 35819
rect 18398 35717 18432 35751
rect 23664 35717 23698 35751
rect 30573 35717 30607 35751
rect 34069 35717 34103 35751
rect 1777 35649 1811 35683
rect 3065 35649 3099 35683
rect 4537 35649 4571 35683
rect 17509 35649 17543 35683
rect 20177 35649 20211 35683
rect 21005 35649 21039 35683
rect 22293 35649 22327 35683
rect 25237 35649 25271 35683
rect 26249 35649 26283 35683
rect 27169 35649 27203 35683
rect 28181 35649 28215 35683
rect 29101 35649 29135 35683
rect 29929 35649 29963 35683
rect 30757 35649 30791 35683
rect 31571 35649 31605 35683
rect 32597 35649 32631 35683
rect 33241 35649 33275 35683
rect 33425 35649 33459 35683
rect 34345 35649 34379 35683
rect 2053 35581 2087 35615
rect 3893 35581 3927 35615
rect 5365 35581 5399 35615
rect 18153 35581 18187 35615
rect 20821 35581 20855 35615
rect 22109 35581 22143 35615
rect 23397 35581 23431 35615
rect 25329 35581 25363 35615
rect 26065 35581 26099 35615
rect 27261 35581 27295 35615
rect 27997 35581 28031 35615
rect 28917 35581 28951 35615
rect 29745 35581 29779 35615
rect 30941 35581 30975 35615
rect 31401 35581 31435 35615
rect 32413 35581 32447 35615
rect 17601 35445 17635 35479
rect 19533 35445 19567 35479
rect 19993 35445 20027 35479
rect 24777 35445 24811 35479
rect 25421 35445 25455 35479
rect 25605 35445 25639 35479
rect 27169 35445 27203 35479
rect 27537 35445 27571 35479
rect 31769 35445 31803 35479
rect 32781 35445 32815 35479
rect 33609 35445 33643 35479
rect 34069 35445 34103 35479
rect 18521 35241 18555 35275
rect 21281 35241 21315 35275
rect 22477 35241 22511 35275
rect 22937 35241 22971 35275
rect 26801 35241 26835 35275
rect 30113 35173 30147 35207
rect 2789 35105 2823 35139
rect 18153 35105 18187 35139
rect 24593 35105 24627 35139
rect 32689 35105 32723 35139
rect 1593 35037 1627 35071
rect 3985 35037 4019 35071
rect 17417 35037 17451 35071
rect 17509 35037 17543 35071
rect 18337 35037 18371 35071
rect 19533 35037 19567 35071
rect 19625 35037 19659 35071
rect 21281 35037 21315 35071
rect 21373 35037 21407 35071
rect 22201 35037 22235 35071
rect 22293 35037 22327 35071
rect 23121 35037 23155 35071
rect 23253 35037 23287 35071
rect 24041 35037 24075 35071
rect 24860 35037 24894 35071
rect 26525 35037 26559 35071
rect 26617 35037 26651 35071
rect 27629 35037 27663 35071
rect 29837 35037 29871 35071
rect 29929 35037 29963 35071
rect 30665 35037 30699 35071
rect 30921 35037 30955 35071
rect 32505 35037 32539 35071
rect 1777 34969 1811 35003
rect 4813 34969 4847 35003
rect 20269 34969 20303 35003
rect 20545 34969 20579 35003
rect 22937 34969 22971 35003
rect 27896 34969 27930 35003
rect 34345 34969 34379 35003
rect 17693 34901 17727 34935
rect 19809 34901 19843 34935
rect 20453 34901 20487 34935
rect 20637 34901 20671 34935
rect 20821 34901 20855 34935
rect 21649 34901 21683 34935
rect 23397 34901 23431 34935
rect 23857 34901 23891 34935
rect 25973 34901 26007 34935
rect 29009 34901 29043 34935
rect 32045 34901 32079 34935
rect 18797 34697 18831 34731
rect 20637 34697 20671 34731
rect 21465 34697 21499 34731
rect 23397 34697 23431 34731
rect 28549 34697 28583 34731
rect 29469 34697 29503 34731
rect 31585 34697 31619 34731
rect 19524 34629 19558 34663
rect 24102 34629 24136 34663
rect 26065 34629 26099 34663
rect 27414 34629 27448 34663
rect 30472 34629 30506 34663
rect 32689 34629 32723 34663
rect 34345 34629 34379 34663
rect 1777 34561 1811 34595
rect 17417 34561 17451 34595
rect 17684 34561 17718 34595
rect 19257 34561 19291 34595
rect 21097 34561 21131 34595
rect 21281 34561 21315 34595
rect 22017 34561 22051 34595
rect 22284 34561 22318 34595
rect 23857 34561 23891 34595
rect 25697 34561 25731 34595
rect 25881 34561 25915 34595
rect 29285 34561 29319 34595
rect 30205 34561 30239 34595
rect 32505 34561 32539 34595
rect 1961 34493 1995 34527
rect 2789 34493 2823 34527
rect 27169 34493 27203 34527
rect 29101 34493 29135 34527
rect 25237 34425 25271 34459
rect 1869 34153 1903 34187
rect 18705 34153 18739 34187
rect 22293 34153 22327 34187
rect 25973 34153 26007 34187
rect 28825 34153 28859 34187
rect 31125 34153 31159 34187
rect 31677 34153 31711 34187
rect 22845 34085 22879 34119
rect 20085 34017 20119 34051
rect 20177 34017 20211 34051
rect 26433 34017 26467 34051
rect 31677 34017 31711 34051
rect 32505 34017 32539 34051
rect 1777 33949 1811 33983
rect 2513 33949 2547 33983
rect 18153 33949 18187 33983
rect 18889 33949 18923 33983
rect 20269 33949 20303 33983
rect 20361 33949 20395 33983
rect 20913 33949 20947 33983
rect 21180 33949 21214 33983
rect 24041 33949 24075 33983
rect 24593 33949 24627 33983
rect 24849 33949 24883 33983
rect 28457 33949 28491 33983
rect 29745 33949 29779 33983
rect 30001 33949 30035 33983
rect 31585 33949 31619 33983
rect 31861 33949 31895 33983
rect 3065 33881 3099 33915
rect 23121 33881 23155 33915
rect 23397 33881 23431 33915
rect 26678 33881 26712 33915
rect 28273 33881 28307 33915
rect 32689 33881 32723 33915
rect 34345 33881 34379 33915
rect 17969 33813 18003 33847
rect 19901 33813 19935 33847
rect 23029 33813 23063 33847
rect 23213 33813 23247 33847
rect 23857 33813 23891 33847
rect 27813 33813 27847 33847
rect 28549 33813 28583 33847
rect 28641 33813 28675 33847
rect 32045 33813 32079 33847
rect 2145 33609 2179 33643
rect 20177 33609 20211 33643
rect 21373 33609 21407 33643
rect 31309 33609 31343 33643
rect 22284 33541 22318 33575
rect 24768 33541 24802 33575
rect 26617 33541 26651 33575
rect 30174 33541 30208 33575
rect 32689 33541 32723 33575
rect 34345 33541 34379 33575
rect 2053 33473 2087 33507
rect 2881 33473 2915 33507
rect 18153 33473 18187 33507
rect 18420 33473 18454 33507
rect 20361 33473 20395 33507
rect 20453 33473 20487 33507
rect 20637 33473 20671 33507
rect 21281 33473 21315 33507
rect 22017 33473 22051 33507
rect 24041 33473 24075 33507
rect 26433 33473 26467 33507
rect 27353 33473 27387 33507
rect 27813 33473 27847 33507
rect 28080 33473 28114 33507
rect 32505 33473 32539 33507
rect 20545 33405 20579 33439
rect 24501 33405 24535 33439
rect 29929 33405 29963 33439
rect 19533 33269 19567 33303
rect 23397 33269 23431 33303
rect 23857 33269 23891 33303
rect 25881 33269 25915 33303
rect 27169 33269 27203 33303
rect 29193 33269 29227 33303
rect 1593 33065 1627 33099
rect 18705 33065 18739 33099
rect 21741 33065 21775 33099
rect 23121 33065 23155 33099
rect 29193 33065 29227 33099
rect 25053 32997 25087 33031
rect 19533 32929 19567 32963
rect 31493 32929 31527 32963
rect 31861 32929 31895 32963
rect 1777 32861 1811 32895
rect 18889 32861 18923 32895
rect 19800 32861 19834 32895
rect 21465 32861 21499 32895
rect 21557 32861 21591 32895
rect 22845 32861 22879 32895
rect 22937 32861 22971 32895
rect 24777 32861 24811 32895
rect 24869 32861 24903 32895
rect 25513 32861 25547 32895
rect 27813 32861 27847 32895
rect 29745 32861 29779 32895
rect 29929 32861 29963 32895
rect 30665 32861 30699 32895
rect 30941 32861 30975 32895
rect 23673 32793 23707 32827
rect 24041 32793 24075 32827
rect 25758 32793 25792 32827
rect 28080 32793 28114 32827
rect 30849 32793 30883 32827
rect 32106 32793 32140 32827
rect 33701 32793 33735 32827
rect 33885 32793 33919 32827
rect 20913 32725 20947 32759
rect 26893 32725 26927 32759
rect 30113 32725 30147 32759
rect 31033 32725 31067 32759
rect 31217 32725 31251 32759
rect 33241 32725 33275 32759
rect 34069 32725 34103 32759
rect 20545 32521 20579 32555
rect 25605 32521 25639 32555
rect 30297 32521 30331 32555
rect 31769 32521 31803 32555
rect 18398 32453 18432 32487
rect 22928 32453 22962 32487
rect 28181 32453 28215 32487
rect 29101 32453 29135 32487
rect 29301 32453 29335 32487
rect 31309 32453 31343 32487
rect 32689 32453 32723 32487
rect 18153 32385 18187 32419
rect 20361 32385 20395 32419
rect 21097 32385 21131 32419
rect 21189 32385 21223 32419
rect 22201 32385 22235 32419
rect 24593 32385 24627 32419
rect 24685 32385 24719 32419
rect 25789 32385 25823 32419
rect 25881 32385 25915 32419
rect 25973 32385 26007 32419
rect 26111 32385 26145 32419
rect 27169 32385 27203 32419
rect 27353 32385 27387 32419
rect 27445 32385 27479 32419
rect 27629 32385 27663 32419
rect 28457 32385 28491 32419
rect 30113 32385 30147 32419
rect 31493 32385 31527 32419
rect 31585 32385 31619 32419
rect 32505 32385 32539 32419
rect 20177 32317 20211 32351
rect 22661 32317 22695 32351
rect 26249 32317 26283 32351
rect 28365 32317 28399 32351
rect 29929 32317 29963 32351
rect 34345 32317 34379 32351
rect 27537 32249 27571 32283
rect 28641 32249 28675 32283
rect 19533 32181 19567 32215
rect 21373 32181 21407 32215
rect 22017 32181 22051 32215
rect 24041 32181 24075 32215
rect 24869 32181 24903 32215
rect 28181 32181 28215 32215
rect 29285 32181 29319 32215
rect 29469 32181 29503 32215
rect 31309 32181 31343 32215
rect 17417 31977 17451 32011
rect 20177 31977 20211 32011
rect 23121 31977 23155 32011
rect 24041 31977 24075 32011
rect 24593 31977 24627 32011
rect 30113 31977 30147 32011
rect 33793 31977 33827 32011
rect 25881 31909 25915 31943
rect 31677 31909 31711 31943
rect 18429 31841 18463 31875
rect 19809 31841 19843 31875
rect 24685 31841 24719 31875
rect 25513 31841 25547 31875
rect 29745 31841 29779 31875
rect 31217 31841 31251 31875
rect 32413 31841 32447 31875
rect 2053 31773 2087 31807
rect 17601 31773 17635 31807
rect 18153 31773 18187 31807
rect 18265 31773 18299 31807
rect 19993 31773 20027 31807
rect 20913 31773 20947 31807
rect 22845 31773 22879 31807
rect 23673 31773 23707 31807
rect 23857 31773 23891 31807
rect 24869 31773 24903 31807
rect 25697 31773 25731 31807
rect 26617 31773 26651 31807
rect 29009 31773 29043 31807
rect 29929 31773 29963 31807
rect 30573 31773 30607 31807
rect 30758 31773 30792 31807
rect 30849 31773 30883 31807
rect 31677 31773 31711 31807
rect 31953 31773 31987 31807
rect 32680 31773 32714 31807
rect 21158 31705 21192 31739
rect 24593 31705 24627 31739
rect 26884 31705 26918 31739
rect 28641 31705 28675 31739
rect 30941 31705 30975 31739
rect 31059 31705 31093 31739
rect 22293 31637 22327 31671
rect 25053 31637 25087 31671
rect 27997 31637 28031 31671
rect 31861 31637 31895 31671
rect 17049 31433 17083 31467
rect 21005 31433 21039 31467
rect 31585 31433 31619 31467
rect 31769 31433 31803 31467
rect 21097 31365 21131 31399
rect 22376 31365 22410 31399
rect 24860 31365 24894 31399
rect 27414 31365 27448 31399
rect 31493 31365 31527 31399
rect 32689 31365 32723 31399
rect 1777 31297 1811 31331
rect 17233 31297 17267 31331
rect 17877 31297 17911 31331
rect 18604 31297 18638 31331
rect 20913 31297 20947 31331
rect 22109 31297 22143 31331
rect 24133 31297 24167 31331
rect 26433 31297 26467 31331
rect 26617 31297 26651 31331
rect 27169 31297 27203 31331
rect 29377 31297 29411 31331
rect 29644 31297 29678 31331
rect 31401 31297 31435 31331
rect 32505 31297 32539 31331
rect 34345 31297 34379 31331
rect 1961 31229 1995 31263
rect 2789 31229 2823 31263
rect 18337 31229 18371 31263
rect 24593 31229 24627 31263
rect 31217 31229 31251 31263
rect 20729 31161 20763 31195
rect 23489 31161 23523 31195
rect 17693 31093 17727 31127
rect 19717 31093 19751 31127
rect 21281 31093 21315 31127
rect 23949 31093 23983 31127
rect 25973 31093 26007 31127
rect 26433 31093 26467 31127
rect 28549 31093 28583 31127
rect 30757 31093 30791 31127
rect 2145 30889 2179 30923
rect 18705 30889 18739 30923
rect 19533 30889 19567 30923
rect 21741 30889 21775 30923
rect 22201 30889 22235 30923
rect 24961 30889 24995 30923
rect 30205 30889 30239 30923
rect 33425 30889 33459 30923
rect 18889 30821 18923 30855
rect 23489 30821 23523 30855
rect 24041 30821 24075 30855
rect 31309 30821 31343 30855
rect 18061 30753 18095 30787
rect 19533 30753 19567 30787
rect 20361 30753 20395 30787
rect 22385 30753 22419 30787
rect 30021 30753 30055 30787
rect 30849 30753 30883 30787
rect 32045 30753 32079 30787
rect 2053 30685 2087 30719
rect 17233 30685 17267 30719
rect 17785 30685 17819 30719
rect 17877 30685 17911 30719
rect 19441 30685 19475 30719
rect 20628 30685 20662 30719
rect 22201 30685 22235 30719
rect 22477 30685 22511 30719
rect 23673 30685 23707 30719
rect 23765 30685 23799 30719
rect 24685 30685 24719 30719
rect 24777 30685 24811 30719
rect 28457 30685 28491 30719
rect 28733 30685 28767 30719
rect 29929 30685 29963 30719
rect 30941 30685 30975 30719
rect 33885 30685 33919 30719
rect 34069 30685 34103 30719
rect 18521 30617 18555 30651
rect 18737 30617 18771 30651
rect 23857 30617 23891 30651
rect 26065 30617 26099 30651
rect 28273 30617 28307 30651
rect 32290 30617 32324 30651
rect 17049 30549 17083 30583
rect 19809 30549 19843 30583
rect 22661 30549 22695 30583
rect 27353 30549 27387 30583
rect 28641 30549 28675 30583
rect 34253 30549 34287 30583
rect 17509 30345 17543 30379
rect 21373 30345 21407 30379
rect 23397 30345 23431 30379
rect 18409 30277 18443 30311
rect 22262 30277 22296 30311
rect 25044 30277 25078 30311
rect 27804 30277 27838 30311
rect 32413 30277 32447 30311
rect 33232 30277 33266 30311
rect 17693 30209 17727 30243
rect 18153 30209 18187 30243
rect 20249 30209 20283 30243
rect 24041 30209 24075 30243
rect 24777 30209 24811 30243
rect 29837 30209 29871 30243
rect 30849 30209 30883 30243
rect 32321 30209 32355 30243
rect 32505 30209 32539 30243
rect 32965 30209 32999 30243
rect 19993 30141 20027 30175
rect 22017 30141 22051 30175
rect 23857 30141 23891 30175
rect 27537 30141 27571 30175
rect 29745 30141 29779 30175
rect 30205 30141 30239 30175
rect 30941 30141 30975 30175
rect 26157 30073 26191 30107
rect 28917 30073 28951 30107
rect 19533 30005 19567 30039
rect 24225 30005 24259 30039
rect 31217 30005 31251 30039
rect 34345 30005 34379 30039
rect 16221 29801 16255 29835
rect 23029 29801 23063 29835
rect 29745 29801 29779 29835
rect 17509 29733 17543 29767
rect 20085 29733 20119 29767
rect 20177 29733 20211 29767
rect 23857 29733 23891 29767
rect 25973 29733 26007 29767
rect 27721 29733 27755 29767
rect 33241 29733 33275 29767
rect 24593 29665 24627 29699
rect 26065 29665 26099 29699
rect 27077 29665 27111 29699
rect 30205 29665 30239 29699
rect 33701 29665 33735 29699
rect 16405 29597 16439 29631
rect 16865 29597 16899 29631
rect 17233 29597 17267 29631
rect 17509 29597 17543 29631
rect 17785 29597 17819 29631
rect 18429 29597 18463 29631
rect 18521 29597 18555 29631
rect 18613 29597 18647 29631
rect 18889 29597 18923 29631
rect 19993 29597 20027 29631
rect 20269 29597 20303 29631
rect 20821 29597 20855 29631
rect 22661 29597 22695 29631
rect 22845 29597 22879 29631
rect 23581 29597 23615 29631
rect 23673 29597 23707 29631
rect 24777 29597 24811 29631
rect 24961 29597 24995 29631
rect 25237 29597 25271 29631
rect 25881 29597 25915 29631
rect 26157 29597 26191 29631
rect 27353 29597 27387 29631
rect 27562 29597 27596 29631
rect 28825 29575 28859 29609
rect 28917 29597 28951 29631
rect 29101 29597 29135 29631
rect 29193 29597 29227 29631
rect 29929 29597 29963 29631
rect 30021 29597 30055 29631
rect 30297 29597 30331 29631
rect 30941 29597 30975 29631
rect 31401 29597 31435 29631
rect 33425 29597 33459 29631
rect 33609 29597 33643 29631
rect 34161 29597 34195 29631
rect 34345 29597 34379 29631
rect 18245 29529 18279 29563
rect 18731 29529 18765 29563
rect 19809 29529 19843 29563
rect 21088 29529 21122 29563
rect 24869 29529 24903 29563
rect 25099 29529 25133 29563
rect 25697 29529 25731 29563
rect 31646 29529 31680 29563
rect 16681 29461 16715 29495
rect 17693 29461 17727 29495
rect 22201 29461 22235 29495
rect 27445 29461 27479 29495
rect 28641 29461 28675 29495
rect 30757 29461 30791 29495
rect 32781 29461 32815 29495
rect 34253 29461 34287 29495
rect 20545 29257 20579 29291
rect 21373 29257 21407 29291
rect 24593 29257 24627 29291
rect 31125 29257 31159 29291
rect 33701 29257 33735 29291
rect 19410 29189 19444 29223
rect 21097 29189 21131 29223
rect 22385 29189 22419 29223
rect 25237 29189 25271 29223
rect 28641 29189 28675 29223
rect 32689 29189 32723 29223
rect 17325 29121 17359 29155
rect 17592 29121 17626 29155
rect 19165 29121 19199 29155
rect 22109 29121 22143 29155
rect 22201 29121 22235 29155
rect 23480 29121 23514 29155
rect 26157 29121 26191 29155
rect 27445 29121 27479 29155
rect 27629 29121 27663 29155
rect 27813 29121 27847 29155
rect 27997 29121 28031 29155
rect 31355 29121 31389 29155
rect 31490 29124 31524 29158
rect 31585 29121 31619 29155
rect 31769 29121 31803 29155
rect 32321 29121 32355 29155
rect 32505 29121 32539 29155
rect 32781 29121 32815 29155
rect 33517 29121 33551 29155
rect 33793 29121 33827 29155
rect 23213 29053 23247 29087
rect 27721 29053 27755 29087
rect 25605 28985 25639 29019
rect 25697 28985 25731 29019
rect 26433 28985 26467 29019
rect 26617 28985 26651 29019
rect 28181 28985 28215 29019
rect 33333 28985 33367 29019
rect 18705 28917 18739 28951
rect 29929 28917 29963 28951
rect 16129 28713 16163 28747
rect 22293 28713 22327 28747
rect 25973 28713 26007 28747
rect 27813 28713 27847 28747
rect 33885 28713 33919 28747
rect 17417 28645 17451 28679
rect 23857 28645 23891 28679
rect 19809 28577 19843 28611
rect 28825 28577 28859 28611
rect 29009 28577 29043 28611
rect 32781 28577 32815 28611
rect 32965 28577 32999 28611
rect 33517 28577 33551 28611
rect 16313 28509 16347 28543
rect 16957 28509 16991 28543
rect 17601 28509 17635 28543
rect 18153 28509 18187 28543
rect 18245 28509 18279 28543
rect 19533 28509 19567 28543
rect 19625 28509 19659 28543
rect 24041 28509 24075 28543
rect 24593 28509 24627 28543
rect 24860 28509 24894 28543
rect 26433 28509 26467 28543
rect 26700 28509 26734 28543
rect 28917 28509 28951 28543
rect 29101 28509 29135 28543
rect 29745 28509 29779 28543
rect 31585 28509 31619 28543
rect 32689 28509 32723 28543
rect 33609 28509 33643 28543
rect 18429 28441 18463 28475
rect 20821 28441 20855 28475
rect 23029 28441 23063 28475
rect 23213 28441 23247 28475
rect 30012 28441 30046 28475
rect 32321 28441 32355 28475
rect 16773 28373 16807 28407
rect 23397 28373 23431 28407
rect 28641 28373 28675 28407
rect 31125 28373 31159 28407
rect 31769 28373 31803 28407
rect 23489 28169 23523 28203
rect 27537 28169 27571 28203
rect 31217 28169 31251 28203
rect 17601 28101 17635 28135
rect 20453 28101 20487 28135
rect 30021 28101 30055 28135
rect 32689 28101 32723 28135
rect 16129 28033 16163 28067
rect 16313 28033 16347 28067
rect 17141 28033 17175 28067
rect 18521 28033 18555 28067
rect 18777 28033 18811 28067
rect 21189 28033 21223 28067
rect 21281 28033 21315 28067
rect 22109 28033 22143 28067
rect 22365 28033 22399 28067
rect 24133 28033 24167 28067
rect 24593 28033 24627 28067
rect 24849 28033 24883 28067
rect 26617 28033 26651 28067
rect 27353 28033 27387 28067
rect 28457 28033 28491 28067
rect 29285 28033 29319 28067
rect 29469 28031 29503 28065
rect 29555 28033 29589 28067
rect 29848 28033 29882 28067
rect 30481 28033 30515 28067
rect 30665 28033 30699 28067
rect 30757 28033 30791 28067
rect 31493 28033 31527 28067
rect 32505 28033 32539 28067
rect 20637 27965 20671 27999
rect 27169 27965 27203 27999
rect 28365 27965 28399 27999
rect 28825 27965 28859 27999
rect 29653 27965 29687 27999
rect 31401 27965 31435 27999
rect 31585 27965 31619 27999
rect 31677 27965 31711 27999
rect 34345 27965 34379 27999
rect 16957 27897 16991 27931
rect 17969 27897 18003 27931
rect 26433 27897 26467 27931
rect 16129 27829 16163 27863
rect 18061 27829 18095 27863
rect 19901 27829 19935 27863
rect 21465 27829 21499 27863
rect 23949 27829 23983 27863
rect 25973 27829 26007 27863
rect 30481 27829 30515 27863
rect 24777 27625 24811 27659
rect 34345 27625 34379 27659
rect 16865 27557 16899 27591
rect 23121 27557 23155 27591
rect 25973 27557 26007 27591
rect 26709 27557 26743 27591
rect 27813 27557 27847 27591
rect 6469 27489 6503 27523
rect 7849 27489 7883 27523
rect 17693 27489 17727 27523
rect 17902 27489 17936 27523
rect 29929 27489 29963 27523
rect 30205 27489 30239 27523
rect 31309 27489 31343 27523
rect 31769 27489 31803 27523
rect 32321 27489 32355 27523
rect 32965 27489 32999 27523
rect 16037 27421 16071 27455
rect 16497 27421 16531 27455
rect 17417 27421 17451 27455
rect 17785 27421 17819 27455
rect 18613 27421 18647 27455
rect 18705 27421 18739 27455
rect 19441 27421 19475 27455
rect 21281 27421 21315 27455
rect 23489 27421 23523 27455
rect 24685 27421 24719 27455
rect 25329 27421 25363 27455
rect 26433 27421 26467 27455
rect 27997 27421 28031 27455
rect 28273 27421 28307 27455
rect 28917 27421 28951 27455
rect 29193 27421 29227 27455
rect 30021 27421 30055 27455
rect 30113 27421 30147 27455
rect 31401 27421 31435 27455
rect 32045 27421 32079 27455
rect 32137 27421 32171 27455
rect 6653 27353 6687 27387
rect 19686 27353 19720 27387
rect 21548 27353 21582 27387
rect 23673 27353 23707 27387
rect 25814 27353 25848 27387
rect 33210 27353 33244 27387
rect 15853 27285 15887 27319
rect 16957 27285 16991 27319
rect 18061 27285 18095 27319
rect 18889 27285 18923 27319
rect 20821 27285 20855 27319
rect 22661 27285 22695 27319
rect 23305 27285 23339 27319
rect 23397 27285 23431 27319
rect 25605 27285 25639 27319
rect 25697 27285 25731 27319
rect 26893 27285 26927 27319
rect 28181 27285 28215 27319
rect 28733 27285 28767 27319
rect 29101 27285 29135 27319
rect 29745 27285 29779 27319
rect 32321 27285 32355 27319
rect 32597 27285 32631 27319
rect 6653 27081 6687 27115
rect 8769 27081 8803 27115
rect 20821 27081 20855 27115
rect 28457 27081 28491 27115
rect 19708 27013 19742 27047
rect 23949 27013 23983 27047
rect 6561 26945 6595 26979
rect 8953 26945 8987 26979
rect 16129 26945 16163 26979
rect 16313 26945 16347 26979
rect 16865 26945 16899 26979
rect 17049 26945 17083 26979
rect 17693 26945 17727 26979
rect 17785 26945 17819 26979
rect 17969 26945 18003 26979
rect 18061 26945 18095 26979
rect 18521 26945 18555 26979
rect 18705 26945 18739 26979
rect 19441 26945 19475 26979
rect 21465 26945 21499 26979
rect 22017 26945 22051 26979
rect 22284 26945 22318 26979
rect 24225 26945 24259 26979
rect 25237 26945 25271 26979
rect 25493 26945 25527 26979
rect 27169 26945 27203 26979
rect 29653 26945 29687 26979
rect 29745 26945 29779 26979
rect 29837 26945 29871 26979
rect 30021 26945 30055 26979
rect 31401 26945 31435 26979
rect 31490 26948 31524 26982
rect 31585 26945 31619 26979
rect 31769 26945 31803 26979
rect 32505 26945 32539 26979
rect 33517 26945 33551 26979
rect 33701 26945 33735 26979
rect 33793 26945 33827 26979
rect 24041 26877 24075 26911
rect 32413 26877 32447 26911
rect 32873 26877 32907 26911
rect 17509 26809 17543 26843
rect 24409 26809 24443 26843
rect 16129 26741 16163 26775
rect 16865 26741 16899 26775
rect 18889 26741 18923 26775
rect 21281 26741 21315 26775
rect 23397 26741 23431 26775
rect 24133 26741 24167 26775
rect 26617 26741 26651 26775
rect 29377 26741 29411 26775
rect 31125 26741 31159 26775
rect 33333 26741 33367 26775
rect 26157 26537 26191 26571
rect 29009 26537 29043 26571
rect 30113 26537 30147 26571
rect 31585 26537 31619 26571
rect 19441 26469 19475 26503
rect 24961 26469 24995 26503
rect 28549 26469 28583 26503
rect 30481 26469 30515 26503
rect 32045 26469 32079 26503
rect 17877 26401 17911 26435
rect 22477 26401 22511 26435
rect 23673 26401 23707 26435
rect 24685 26401 24719 26435
rect 25145 26401 25179 26435
rect 26249 26401 26283 26435
rect 30573 26401 30607 26435
rect 16773 26333 16807 26367
rect 17049 26333 17083 26367
rect 17509 26333 17543 26367
rect 17693 26333 17727 26367
rect 17785 26333 17819 26367
rect 18061 26333 18095 26367
rect 18245 26333 18279 26367
rect 18705 26333 18739 26367
rect 18889 26333 18923 26367
rect 19625 26333 19659 26367
rect 20177 26333 20211 26367
rect 20821 26333 20855 26367
rect 23213 26333 23247 26367
rect 23515 26333 23549 26367
rect 25881 26333 25915 26367
rect 25973 26333 26007 26367
rect 27169 26333 27203 26367
rect 29009 26333 29043 26367
rect 29193 26333 29227 26367
rect 30297 26333 30331 26367
rect 31769 26333 31803 26367
rect 31861 26333 31895 26367
rect 32137 26333 32171 26367
rect 32781 26333 32815 26367
rect 33037 26333 33071 26367
rect 16589 26265 16623 26299
rect 16957 26265 16991 26299
rect 20269 26265 20303 26299
rect 23305 26265 23339 26299
rect 23397 26265 23431 26299
rect 27436 26265 27470 26299
rect 18797 26197 18831 26231
rect 23029 26197 23063 26231
rect 25697 26197 25731 26231
rect 34161 26197 34195 26231
rect 26525 25993 26559 26027
rect 17417 25925 17451 25959
rect 22928 25925 22962 25959
rect 24746 25925 24780 25959
rect 27537 25925 27571 25959
rect 31309 25925 31343 25959
rect 15669 25857 15703 25891
rect 17601 25857 17635 25891
rect 17693 25857 17727 25891
rect 17969 25857 18003 25891
rect 18613 25857 18647 25891
rect 18797 25857 18831 25891
rect 18889 25857 18923 25891
rect 19349 25857 19383 25891
rect 19605 25857 19639 25891
rect 21189 25857 21223 25891
rect 21373 25857 21407 25891
rect 21465 25857 21499 25891
rect 22201 25857 22235 25891
rect 22661 25857 22695 25891
rect 26341 25857 26375 25891
rect 27813 25857 27847 25891
rect 27905 25860 27939 25894
rect 27997 25857 28031 25891
rect 28181 25857 28215 25891
rect 28641 25857 28675 25891
rect 28908 25857 28942 25891
rect 31033 25857 31067 25891
rect 31181 25857 31215 25891
rect 31401 25857 31435 25891
rect 31498 25857 31532 25891
rect 32505 25857 32539 25891
rect 34345 25857 34379 25891
rect 17877 25789 17911 25823
rect 24501 25789 24535 25823
rect 32689 25789 32723 25823
rect 16313 25721 16347 25755
rect 22017 25721 22051 25755
rect 24041 25721 24075 25755
rect 25881 25721 25915 25755
rect 2053 25653 2087 25687
rect 18429 25653 18463 25687
rect 20729 25653 20763 25687
rect 21189 25653 21223 25687
rect 30021 25653 30055 25687
rect 31677 25653 31711 25687
rect 16589 25449 16623 25483
rect 19441 25449 19475 25483
rect 23397 25449 23431 25483
rect 24961 25449 24995 25483
rect 27905 25449 27939 25483
rect 32045 25449 32079 25483
rect 29193 25381 29227 25415
rect 1593 25313 1627 25347
rect 2789 25313 2823 25347
rect 16037 25313 16071 25347
rect 18429 25313 18463 25347
rect 22845 25313 22879 25347
rect 25973 25313 26007 25347
rect 26433 25313 26467 25347
rect 31585 25313 31619 25347
rect 31677 25313 31711 25347
rect 32505 25313 32539 25347
rect 32689 25313 32723 25347
rect 15301 25245 15335 25279
rect 15945 25245 15979 25279
rect 16589 25245 16623 25279
rect 16773 25245 16807 25279
rect 17417 25245 17451 25279
rect 18337 25245 18371 25279
rect 19717 25245 19751 25279
rect 19809 25245 19843 25279
rect 19906 25245 19940 25279
rect 20085 25245 20119 25279
rect 20821 25245 20855 25279
rect 23121 25245 23155 25279
rect 23857 25245 23891 25279
rect 25697 25245 25731 25279
rect 25881 25245 25915 25279
rect 26065 25245 26099 25279
rect 26249 25245 26283 25279
rect 27077 25245 27111 25279
rect 27169 25245 27203 25279
rect 27353 25245 27387 25279
rect 27445 25245 27479 25279
rect 28089 25245 28123 25279
rect 28365 25245 28399 25279
rect 28825 25245 28859 25279
rect 29009 25245 29043 25279
rect 30297 25245 30331 25279
rect 30665 25245 30699 25279
rect 31309 25245 31343 25279
rect 31493 25245 31527 25279
rect 31861 25245 31895 25279
rect 1777 25177 1811 25211
rect 17233 25177 17267 25211
rect 21088 25177 21122 25211
rect 23213 25177 23247 25211
rect 24685 25177 24719 25211
rect 30481 25177 30515 25211
rect 30573 25177 30607 25211
rect 34345 25177 34379 25211
rect 15393 25109 15427 25143
rect 17601 25109 17635 25143
rect 18705 25109 18739 25143
rect 22201 25109 22235 25143
rect 23029 25109 23063 25143
rect 23949 25109 23983 25143
rect 26893 25109 26927 25143
rect 28273 25109 28307 25143
rect 30849 25109 30883 25143
rect 2145 24905 2179 24939
rect 16221 24905 16255 24939
rect 25697 24905 25731 24939
rect 26525 24905 26559 24939
rect 27905 24905 27939 24939
rect 17417 24837 17451 24871
rect 17617 24837 17651 24871
rect 18981 24837 19015 24871
rect 33609 24837 33643 24871
rect 2053 24769 2087 24803
rect 16037 24769 16071 24803
rect 18245 24769 18279 24803
rect 18429 24769 18463 24803
rect 18889 24769 18923 24803
rect 19073 24769 19107 24803
rect 19717 24769 19751 24803
rect 20361 24769 20395 24803
rect 20453 24769 20487 24803
rect 21281 24769 21315 24803
rect 21465 24769 21499 24803
rect 22477 24769 22511 24803
rect 22744 24769 22778 24803
rect 24317 24769 24351 24803
rect 24573 24769 24607 24803
rect 26341 24769 26375 24803
rect 26617 24769 26651 24803
rect 27721 24769 27755 24803
rect 27997 24769 28031 24803
rect 28724 24769 28758 24803
rect 30297 24769 30331 24803
rect 30481 24769 30515 24803
rect 31309 24769 31343 24803
rect 31401 24769 31435 24803
rect 31677 24769 31711 24803
rect 32321 24769 32355 24803
rect 32505 24769 32539 24803
rect 32597 24769 32631 24803
rect 32689 24769 32723 24803
rect 33333 24769 33367 24803
rect 33517 24769 33551 24803
rect 33701 24769 33735 24803
rect 20637 24701 20671 24735
rect 21097 24701 21131 24735
rect 27537 24701 27571 24735
rect 28457 24701 28491 24735
rect 19533 24633 19567 24667
rect 31585 24633 31619 24667
rect 33885 24633 33919 24667
rect 17601 24565 17635 24599
rect 17785 24565 17819 24599
rect 18337 24565 18371 24599
rect 20545 24565 20579 24599
rect 23857 24565 23891 24599
rect 26157 24565 26191 24599
rect 29837 24565 29871 24599
rect 30665 24565 30699 24599
rect 31125 24565 31159 24599
rect 32873 24565 32907 24599
rect 16773 24361 16807 24395
rect 17233 24361 17267 24395
rect 22017 24361 22051 24395
rect 22937 24361 22971 24395
rect 23121 24361 23155 24395
rect 23949 24361 23983 24395
rect 30113 24361 30147 24395
rect 30941 24361 30975 24395
rect 31585 24361 31619 24395
rect 16313 24225 16347 24259
rect 23581 24225 23615 24259
rect 24961 24225 24995 24259
rect 27077 24225 27111 24259
rect 27353 24225 27387 24259
rect 28457 24225 28491 24259
rect 28549 24225 28583 24259
rect 30205 24225 30239 24259
rect 15577 24157 15611 24191
rect 15761 24157 15795 24191
rect 16405 24157 16439 24191
rect 17417 24157 17451 24191
rect 17693 24157 17727 24191
rect 18475 24157 18509 24191
rect 18613 24157 18647 24191
rect 18726 24157 18760 24191
rect 18889 24157 18923 24191
rect 19441 24157 19475 24191
rect 22845 24157 22879 24191
rect 22937 24157 22971 24191
rect 23765 24157 23799 24191
rect 24869 24157 24903 24191
rect 25881 24157 25915 24191
rect 26065 24157 26099 24191
rect 26157 24157 26191 24191
rect 26985 24157 27019 24191
rect 28365 24157 28399 24191
rect 28641 24157 28675 24191
rect 29745 24157 29779 24191
rect 29929 24157 29963 24191
rect 30665 24157 30699 24191
rect 31769 24157 31803 24191
rect 32045 24157 32079 24191
rect 32505 24157 32539 24191
rect 15669 24089 15703 24123
rect 18245 24089 18279 24123
rect 19686 24089 19720 24123
rect 21833 24089 21867 24123
rect 22049 24089 22083 24123
rect 22661 24089 22695 24123
rect 31953 24089 31987 24123
rect 32689 24089 32723 24123
rect 34345 24089 34379 24123
rect 17601 24021 17635 24055
rect 20821 24021 20855 24055
rect 22201 24021 22235 24055
rect 25237 24021 25271 24055
rect 25697 24021 25731 24055
rect 28181 24021 28215 24055
rect 31125 24021 31159 24055
rect 22477 23817 22511 23851
rect 18613 23749 18647 23783
rect 19318 23749 19352 23783
rect 28641 23749 28675 23783
rect 34345 23749 34379 23783
rect 15945 23681 15979 23715
rect 17049 23681 17083 23715
rect 17233 23681 17267 23715
rect 17877 23681 17911 23715
rect 18061 23681 18095 23715
rect 18153 23681 18187 23715
rect 18429 23681 18463 23715
rect 19073 23681 19107 23715
rect 21281 23681 21315 23715
rect 22017 23681 22051 23715
rect 22937 23681 22971 23715
rect 23121 23681 23155 23715
rect 23581 23681 23615 23715
rect 23848 23681 23882 23715
rect 25697 23681 25731 23715
rect 25789 23681 25823 23715
rect 25881 23681 25915 23715
rect 26065 23681 26099 23715
rect 27353 23681 27387 23715
rect 31033 23681 31067 23715
rect 16037 23613 16071 23647
rect 16313 23613 16347 23647
rect 17141 23613 17175 23647
rect 17325 23613 17359 23647
rect 18245 23613 18279 23647
rect 21097 23613 21131 23647
rect 27261 23613 27295 23647
rect 30389 23613 30423 23647
rect 31309 23613 31343 23647
rect 32505 23613 32539 23647
rect 32689 23613 32723 23647
rect 21465 23545 21499 23579
rect 16865 23477 16899 23511
rect 20453 23477 20487 23511
rect 22293 23477 22327 23511
rect 23029 23477 23063 23511
rect 24961 23477 24995 23511
rect 25421 23477 25455 23511
rect 27721 23477 27755 23511
rect 30849 23477 30883 23511
rect 31217 23477 31251 23511
rect 16681 23273 16715 23307
rect 17877 23273 17911 23307
rect 19809 23273 19843 23307
rect 22109 23273 22143 23307
rect 32045 23273 32079 23307
rect 18613 23205 18647 23239
rect 26893 23205 26927 23239
rect 31309 23205 31343 23239
rect 17601 23137 17635 23171
rect 19901 23137 19935 23171
rect 28733 23137 28767 23171
rect 28825 23137 28859 23171
rect 34345 23137 34379 23171
rect 16589 23069 16623 23103
rect 16773 23069 16807 23103
rect 17693 23069 17727 23103
rect 18889 23069 18923 23103
rect 19625 23069 19659 23103
rect 20821 23069 20855 23103
rect 23213 23069 23247 23103
rect 23489 23069 23523 23103
rect 24777 23069 24811 23103
rect 24961 23069 24995 23103
rect 25053 23069 25087 23103
rect 25513 23069 25547 23103
rect 28457 23069 28491 23103
rect 28641 23069 28675 23103
rect 29020 23069 29054 23103
rect 29653 23069 29687 23103
rect 31677 23069 31711 23103
rect 31861 23069 31895 23103
rect 32505 23069 32539 23103
rect 17233 23001 17267 23035
rect 18613 23001 18647 23035
rect 23397 23001 23431 23035
rect 25758 23001 25792 23035
rect 27445 23001 27479 23035
rect 29920 23001 29954 23035
rect 32689 23001 32723 23035
rect 18797 22933 18831 22967
rect 19441 22933 19475 22967
rect 23029 22933 23063 22967
rect 24593 22933 24627 22967
rect 27721 22933 27755 22967
rect 29193 22933 29227 22967
rect 31033 22933 31067 22967
rect 17049 22729 17083 22763
rect 19809 22729 19843 22763
rect 21189 22729 21223 22763
rect 25881 22729 25915 22763
rect 26617 22729 26651 22763
rect 29101 22729 29135 22763
rect 31401 22729 31435 22763
rect 34253 22729 34287 22763
rect 20821 22661 20855 22695
rect 22284 22661 22318 22695
rect 30288 22661 30322 22695
rect 17233 22593 17267 22627
rect 18429 22593 18463 22627
rect 18696 22593 18730 22627
rect 20637 22593 20671 22627
rect 20913 22593 20947 22627
rect 21005 22593 21039 22627
rect 24124 22593 24158 22627
rect 25697 22593 25731 22627
rect 25973 22593 26007 22627
rect 26433 22593 26467 22627
rect 26617 22593 26651 22627
rect 28917 22593 28951 22627
rect 29193 22593 29227 22627
rect 30021 22593 30055 22627
rect 32321 22593 32355 22627
rect 32588 22593 32622 22627
rect 34161 22593 34195 22627
rect 34345 22593 34379 22627
rect 17509 22525 17543 22559
rect 22017 22525 22051 22559
rect 23857 22525 23891 22559
rect 27629 22525 27663 22559
rect 27997 22525 28031 22559
rect 28089 22525 28123 22559
rect 17417 22457 17451 22491
rect 25697 22457 25731 22491
rect 23397 22389 23431 22423
rect 25237 22389 25271 22423
rect 28273 22389 28307 22423
rect 28733 22389 28767 22423
rect 33701 22389 33735 22423
rect 19717 22185 19751 22219
rect 24593 22185 24627 22219
rect 28825 22185 28859 22219
rect 31125 22185 31159 22219
rect 17601 22117 17635 22151
rect 18705 22117 18739 22151
rect 23857 22117 23891 22151
rect 16221 22049 16255 22083
rect 16497 22049 16531 22083
rect 17325 22049 17359 22083
rect 20361 22049 20395 22083
rect 20821 22049 20855 22083
rect 24041 22049 24075 22083
rect 24961 22049 24995 22083
rect 29745 22049 29779 22083
rect 16129 21981 16163 22015
rect 17233 21981 17267 22015
rect 18429 21981 18463 22015
rect 18613 21981 18647 22015
rect 18797 21981 18831 22015
rect 20545 21981 20579 22015
rect 20637 21981 20671 22015
rect 20913 21981 20947 22015
rect 21649 21981 21683 22015
rect 21742 21981 21776 22015
rect 22155 21981 22189 22015
rect 22753 21981 22787 22015
rect 23121 21981 23155 22015
rect 23765 21981 23799 22015
rect 24777 21981 24811 22015
rect 25053 21981 25087 22015
rect 26065 21981 26099 22015
rect 26433 21981 26467 22015
rect 27629 21981 27663 22015
rect 27721 21981 27755 22015
rect 27813 21981 27847 22015
rect 27997 21981 28031 22015
rect 30001 21981 30035 22015
rect 31769 21981 31803 22015
rect 31953 21981 31987 22015
rect 32045 21981 32079 22015
rect 32781 21981 32815 22015
rect 18889 21913 18923 21947
rect 19533 21913 19567 21947
rect 21925 21913 21959 21947
rect 22017 21913 22051 21947
rect 22937 21913 22971 21947
rect 23029 21913 23063 21947
rect 26249 21913 26283 21947
rect 26341 21913 26375 21947
rect 28641 21913 28675 21947
rect 31585 21913 31619 21947
rect 33026 21913 33060 21947
rect 19733 21845 19767 21879
rect 19901 21845 19935 21879
rect 22293 21845 22327 21879
rect 23305 21845 23339 21879
rect 24041 21845 24075 21879
rect 26617 21845 26651 21879
rect 27353 21845 27387 21879
rect 28841 21845 28875 21879
rect 29009 21845 29043 21879
rect 34161 21845 34195 21879
rect 15301 21641 15335 21675
rect 17141 21641 17175 21675
rect 17785 21641 17819 21675
rect 21465 21641 21499 21675
rect 22569 21641 22603 21675
rect 22293 21573 22327 21607
rect 25513 21573 25547 21607
rect 27690 21573 27724 21607
rect 29285 21573 29319 21607
rect 29485 21573 29519 21607
rect 30297 21573 30331 21607
rect 30513 21573 30547 21607
rect 15117 21505 15151 21539
rect 15301 21505 15335 21539
rect 16037 21505 16071 21539
rect 17601 21505 17635 21539
rect 18972 21505 19006 21539
rect 20729 21505 20763 21539
rect 20913 21505 20947 21539
rect 21005 21505 21039 21539
rect 21281 21505 21315 21539
rect 22017 21505 22051 21539
rect 22201 21505 22235 21539
rect 22385 21505 22419 21539
rect 23745 21505 23779 21539
rect 25329 21505 25363 21539
rect 25605 21505 25639 21539
rect 26249 21505 26283 21539
rect 26341 21505 26375 21539
rect 26617 21505 26651 21539
rect 27445 21505 27479 21539
rect 31309 21505 31343 21539
rect 32873 21505 32907 21539
rect 33140 21505 33174 21539
rect 15945 21437 15979 21471
rect 16129 21437 16163 21471
rect 16221 21437 16255 21471
rect 17509 21437 17543 21471
rect 18705 21437 18739 21471
rect 21097 21437 21131 21471
rect 23489 21437 23523 21471
rect 31125 21437 31159 21471
rect 25329 21369 25363 21403
rect 29653 21369 29687 21403
rect 30665 21369 30699 21403
rect 15761 21301 15795 21335
rect 20085 21301 20119 21335
rect 24869 21301 24903 21335
rect 26065 21301 26099 21335
rect 26525 21301 26559 21335
rect 28825 21301 28859 21335
rect 29469 21301 29503 21335
rect 30481 21301 30515 21335
rect 31493 21301 31527 21335
rect 34253 21301 34287 21335
rect 16681 21097 16715 21131
rect 23581 21097 23615 21131
rect 30113 21097 30147 21131
rect 31861 21097 31895 21131
rect 17785 21029 17819 21063
rect 20085 21029 20119 21063
rect 16405 20961 16439 20995
rect 17509 20961 17543 20995
rect 28733 20961 28767 20995
rect 29009 20961 29043 20995
rect 30573 20961 30607 20995
rect 16313 20893 16347 20927
rect 17601 20893 17635 20927
rect 18475 20893 18509 20927
rect 18626 20887 18660 20921
rect 18726 20893 18760 20927
rect 18889 20893 18923 20927
rect 19441 20893 19475 20927
rect 20269 20893 20303 20927
rect 20361 20893 20395 20927
rect 20821 20893 20855 20927
rect 23765 20893 23799 20927
rect 23949 20893 23983 20927
rect 24041 20893 24075 20927
rect 26065 20893 26099 20927
rect 28641 20893 28675 20927
rect 29745 20893 29779 20927
rect 29929 20893 29963 20927
rect 30757 20893 30791 20927
rect 32505 20893 32539 20927
rect 20085 20825 20119 20859
rect 22569 20825 22603 20859
rect 24685 20825 24719 20859
rect 31677 20825 31711 20859
rect 32689 20825 32723 20859
rect 34345 20825 34379 20859
rect 17141 20757 17175 20791
rect 18245 20757 18279 20791
rect 19533 20757 19567 20791
rect 24961 20757 24995 20791
rect 27537 20757 27571 20791
rect 30941 20757 30975 20791
rect 31877 20757 31911 20791
rect 32045 20757 32079 20791
rect 17141 20553 17175 20587
rect 18429 20553 18463 20587
rect 21373 20553 21407 20587
rect 24317 20553 24351 20587
rect 25513 20553 25547 20587
rect 34253 20553 34287 20587
rect 18061 20485 18095 20519
rect 19686 20485 19720 20519
rect 26249 20485 26283 20519
rect 16037 20417 16071 20451
rect 16221 20417 16255 20451
rect 17325 20417 17359 20451
rect 18245 20417 18279 20451
rect 19441 20417 19475 20451
rect 21281 20417 21315 20451
rect 22017 20417 22051 20451
rect 22284 20417 22318 20451
rect 23857 20417 23891 20451
rect 25329 20417 25363 20451
rect 25605 20417 25639 20451
rect 26065 20417 26099 20451
rect 26341 20417 26375 20451
rect 26433 20417 26467 20451
rect 27169 20417 27203 20451
rect 27425 20417 27459 20451
rect 29193 20417 29227 20451
rect 30205 20417 30239 20451
rect 31217 20417 31251 20451
rect 31401 20417 31435 20451
rect 32321 20417 32355 20451
rect 32588 20417 32622 20451
rect 34161 20417 34195 20451
rect 34345 20417 34379 20451
rect 17601 20349 17635 20383
rect 29285 20349 29319 20383
rect 29377 20349 29411 20383
rect 29469 20349 29503 20383
rect 30113 20349 30147 20383
rect 31493 20349 31527 20383
rect 17509 20281 17543 20315
rect 20821 20281 20855 20315
rect 26617 20281 26651 20315
rect 28549 20281 28583 20315
rect 30573 20281 30607 20315
rect 16037 20213 16071 20247
rect 23397 20213 23431 20247
rect 23949 20213 23983 20247
rect 25145 20213 25179 20247
rect 29009 20213 29043 20247
rect 31033 20213 31067 20247
rect 33701 20213 33735 20247
rect 21281 20009 21315 20043
rect 26525 20009 26559 20043
rect 31769 20009 31803 20043
rect 17785 19941 17819 19975
rect 20821 19941 20855 19975
rect 21741 19941 21775 19975
rect 19441 19873 19475 19907
rect 28089 19873 28123 19907
rect 29193 19873 29227 19907
rect 32505 19873 32539 19907
rect 2053 19805 2087 19839
rect 16037 19805 16071 19839
rect 16221 19805 16255 19839
rect 16865 19805 16899 19839
rect 17049 19805 17083 19839
rect 17141 19805 17175 19839
rect 17693 19805 17727 19839
rect 18613 19805 18647 19839
rect 18705 19805 18739 19839
rect 21465 19805 21499 19839
rect 21557 19805 21591 19839
rect 21833 19805 21867 19839
rect 22385 19805 22419 19839
rect 24593 19805 24627 19839
rect 26801 19805 26835 19839
rect 26893 19805 26927 19839
rect 26985 19805 27019 19839
rect 27169 19805 27203 19839
rect 28181 19805 28215 19839
rect 29745 19805 29779 19839
rect 34345 19805 34379 19839
rect 16129 19737 16163 19771
rect 18337 19737 18371 19771
rect 18797 19737 18831 19771
rect 19686 19737 19720 19771
rect 22652 19737 22686 19771
rect 24860 19737 24894 19771
rect 28365 19737 28399 19771
rect 28825 19737 28859 19771
rect 29009 19737 29043 19771
rect 30012 19737 30046 19771
rect 31585 19737 31619 19771
rect 32689 19737 32723 19771
rect 2145 19669 2179 19703
rect 16681 19669 16715 19703
rect 18429 19669 18463 19703
rect 23765 19669 23799 19703
rect 25973 19669 26007 19703
rect 27721 19669 27755 19703
rect 31125 19669 31159 19703
rect 31785 19669 31819 19703
rect 31953 19669 31987 19703
rect 16313 19465 16347 19499
rect 18613 19465 18647 19499
rect 19901 19465 19935 19499
rect 22477 19465 22511 19499
rect 22937 19465 22971 19499
rect 27721 19465 27755 19499
rect 29101 19465 29135 19499
rect 1961 19397 1995 19431
rect 15393 19397 15427 19431
rect 24961 19397 24995 19431
rect 25161 19397 25195 19431
rect 32689 19397 32723 19431
rect 15301 19329 15335 19363
rect 15485 19329 15519 19363
rect 16129 19329 16163 19363
rect 17049 19329 17083 19363
rect 18429 19329 18463 19363
rect 19165 19329 19199 19363
rect 19349 19329 19383 19363
rect 19809 19329 19843 19363
rect 20637 19329 20671 19363
rect 20821 19329 20855 19363
rect 20913 19329 20947 19363
rect 23121 19329 23155 19363
rect 24041 19329 24075 19363
rect 24225 19329 24259 19363
rect 26065 19329 26099 19363
rect 26157 19329 26191 19363
rect 26433 19329 26467 19363
rect 27169 19329 27203 19363
rect 27353 19329 27387 19363
rect 27445 19329 27479 19363
rect 27561 19329 27595 19363
rect 28457 19329 28491 19363
rect 29561 19329 29595 19363
rect 30656 19329 30690 19363
rect 32505 19329 32539 19363
rect 1777 19261 1811 19295
rect 2237 19261 2271 19295
rect 15945 19261 15979 19295
rect 16957 19261 16991 19295
rect 22017 19261 22051 19295
rect 23397 19261 23431 19295
rect 23857 19261 23891 19295
rect 26341 19261 26375 19295
rect 28825 19261 28859 19295
rect 28917 19261 28951 19295
rect 30389 19261 30423 19295
rect 34345 19261 34379 19295
rect 17417 19193 17451 19227
rect 19165 19193 19199 19227
rect 22385 19193 22419 19227
rect 31769 19193 31803 19227
rect 20637 19125 20671 19159
rect 23305 19125 23339 19159
rect 25145 19125 25179 19159
rect 25329 19125 25363 19159
rect 25881 19125 25915 19159
rect 29745 19125 29779 19159
rect 2053 18921 2087 18955
rect 16957 18921 16991 18955
rect 17693 18921 17727 18955
rect 21097 18921 21131 18955
rect 21741 18921 21775 18955
rect 22569 18921 22603 18955
rect 22753 18921 22787 18955
rect 29101 18921 29135 18955
rect 29745 18921 29779 18955
rect 32965 18921 32999 18955
rect 33701 18921 33735 18955
rect 23765 18853 23799 18887
rect 24869 18853 24903 18887
rect 30113 18853 30147 18887
rect 32505 18853 32539 18887
rect 16681 18785 16715 18819
rect 19717 18785 19751 18819
rect 25789 18785 25823 18819
rect 26985 18785 27019 18819
rect 28181 18785 28215 18819
rect 28457 18785 28491 18819
rect 29193 18785 29227 18819
rect 30205 18785 30239 18819
rect 33793 18785 33827 18819
rect 2697 18717 2731 18751
rect 16589 18717 16623 18751
rect 17601 18717 17635 18751
rect 17785 18717 17819 18751
rect 18475 18717 18509 18751
rect 18613 18717 18647 18751
rect 18705 18717 18739 18751
rect 18889 18717 18923 18751
rect 23765 18717 23799 18751
rect 24041 18717 24075 18751
rect 25973 18717 26007 18751
rect 26157 18717 26191 18751
rect 26249 18717 26283 18751
rect 26709 18717 26743 18751
rect 26893 18717 26927 18751
rect 27077 18717 27111 18751
rect 27261 18717 27295 18751
rect 28089 18717 28123 18751
rect 28917 18717 28951 18751
rect 29009 18717 29043 18751
rect 29929 18717 29963 18751
rect 31125 18717 31159 18751
rect 33149 18717 33183 18751
rect 33241 18717 33275 18751
rect 33701 18717 33735 18751
rect 19984 18649 20018 18683
rect 21557 18649 21591 18683
rect 22385 18649 22419 18683
rect 23949 18649 23983 18683
rect 24685 18649 24719 18683
rect 31370 18649 31404 18683
rect 32965 18649 32999 18683
rect 33977 18649 34011 18683
rect 18245 18581 18279 18615
rect 21757 18581 21791 18615
rect 21925 18581 21959 18615
rect 22585 18581 22619 18615
rect 27445 18581 27479 18615
rect 17417 18377 17451 18411
rect 19809 18377 19843 18411
rect 20269 18377 20303 18411
rect 21373 18377 21407 18411
rect 27997 18377 28031 18411
rect 33057 18377 33091 18411
rect 21189 18309 21223 18343
rect 27629 18309 27663 18343
rect 32321 18309 32355 18343
rect 32505 18309 32539 18343
rect 33333 18309 33367 18343
rect 1777 18241 1811 18275
rect 17049 18241 17083 18275
rect 18429 18241 18463 18275
rect 18685 18241 18719 18275
rect 20453 18241 20487 18275
rect 20729 18241 20763 18275
rect 21465 18241 21499 18275
rect 22284 18241 22318 18275
rect 23857 18241 23891 18275
rect 24113 18241 24147 18275
rect 25881 18241 25915 18275
rect 27353 18241 27387 18275
rect 27501 18241 27535 18275
rect 27721 18241 27755 18275
rect 27859 18241 27893 18275
rect 28713 18241 28747 18275
rect 30297 18241 30331 18275
rect 30389 18241 30423 18275
rect 31493 18241 31527 18275
rect 31677 18241 31711 18275
rect 31769 18241 31803 18275
rect 32597 18241 32631 18275
rect 33057 18241 33091 18275
rect 33793 18241 33827 18275
rect 1961 18173 1995 18207
rect 2789 18173 2823 18207
rect 17141 18173 17175 18207
rect 20637 18173 20671 18207
rect 22017 18173 22051 18207
rect 25697 18173 25731 18207
rect 28457 18173 28491 18207
rect 30573 18173 30607 18207
rect 33885 18173 33919 18207
rect 34069 18173 34103 18207
rect 21189 18105 21223 18139
rect 25237 18105 25271 18139
rect 30481 18105 30515 18139
rect 32321 18105 32355 18139
rect 33149 18105 33183 18139
rect 23397 18037 23431 18071
rect 26065 18037 26099 18071
rect 29837 18037 29871 18071
rect 31493 18037 31527 18071
rect 33977 18037 34011 18071
rect 2145 17833 2179 17867
rect 20821 17833 20855 17867
rect 23857 17833 23891 17867
rect 28365 17833 28399 17867
rect 31677 17833 31711 17867
rect 19441 17697 19475 17731
rect 29837 17697 29871 17731
rect 32689 17697 32723 17731
rect 34345 17697 34379 17731
rect 2053 17629 2087 17663
rect 21557 17629 21591 17663
rect 23673 17629 23707 17663
rect 23949 17629 23983 17663
rect 24593 17629 24627 17663
rect 26433 17629 26467 17663
rect 28641 17629 28675 17663
rect 28733 17629 28767 17663
rect 28825 17629 28859 17663
rect 29009 17629 29043 17663
rect 31677 17629 31711 17663
rect 31953 17629 31987 17663
rect 32505 17629 32539 17663
rect 19686 17561 19720 17595
rect 21802 17561 21836 17595
rect 24860 17561 24894 17595
rect 26700 17561 26734 17595
rect 30082 17561 30116 17595
rect 22937 17493 22971 17527
rect 23489 17493 23523 17527
rect 25973 17493 26007 17527
rect 27813 17493 27847 17527
rect 31217 17493 31251 17527
rect 31861 17493 31895 17527
rect 19349 17289 19383 17323
rect 21465 17289 21499 17323
rect 30297 17289 30331 17323
rect 23112 17221 23146 17255
rect 24869 17221 24903 17255
rect 25085 17221 25119 17255
rect 26157 17221 26191 17255
rect 27414 17221 27448 17255
rect 31677 17221 31711 17255
rect 32689 17221 32723 17255
rect 19257 17153 19291 17187
rect 19441 17153 19475 17187
rect 20085 17153 20119 17187
rect 20352 17153 20386 17187
rect 22201 17153 22235 17187
rect 22845 17153 22879 17187
rect 26341 17153 26375 17187
rect 27169 17153 27203 17187
rect 29193 17153 29227 17187
rect 30021 17153 30055 17187
rect 30767 17175 30801 17209
rect 31493 17153 31527 17187
rect 31769 17153 31803 17187
rect 1777 17085 1811 17119
rect 1961 17085 1995 17119
rect 2789 17085 2823 17119
rect 22017 17085 22051 17119
rect 26617 17085 26651 17119
rect 29101 17085 29135 17119
rect 30113 17085 30147 17119
rect 30297 17085 30331 17119
rect 31033 17085 31067 17119
rect 32505 17085 32539 17119
rect 34345 17085 34379 17119
rect 29561 17017 29595 17051
rect 30941 17017 30975 17051
rect 31493 17017 31527 17051
rect 22385 16949 22419 16983
rect 24225 16949 24259 16983
rect 25053 16949 25087 16983
rect 25237 16949 25271 16983
rect 26525 16949 26559 16983
rect 28549 16949 28583 16983
rect 30849 16949 30883 16983
rect 2053 16745 2087 16779
rect 2605 16745 2639 16779
rect 20637 16745 20671 16779
rect 21649 16745 21683 16779
rect 22385 16745 22419 16779
rect 24777 16745 24811 16779
rect 27537 16745 27571 16779
rect 28825 16745 28859 16779
rect 29745 16745 29779 16779
rect 20729 16677 20763 16711
rect 24685 16677 24719 16711
rect 31677 16677 31711 16711
rect 20913 16609 20947 16643
rect 22569 16609 22603 16643
rect 24041 16609 24075 16643
rect 28365 16609 28399 16643
rect 32505 16609 32539 16643
rect 2513 16541 2547 16575
rect 20637 16541 20671 16575
rect 21649 16541 21683 16575
rect 21833 16541 21867 16575
rect 22293 16541 22327 16575
rect 23029 16541 23063 16575
rect 23765 16541 23799 16575
rect 23857 16541 23891 16575
rect 24593 16541 24627 16575
rect 25513 16541 25547 16575
rect 25605 16541 25639 16575
rect 26157 16541 26191 16575
rect 26341 16541 26375 16575
rect 27353 16541 27387 16575
rect 28457 16541 28491 16575
rect 30021 16541 30055 16575
rect 30757 16541 30791 16575
rect 30941 16541 30975 16575
rect 31585 16541 31619 16575
rect 31769 16541 31803 16575
rect 23121 16473 23155 16507
rect 24869 16473 24903 16507
rect 25329 16473 25363 16507
rect 29745 16473 29779 16507
rect 32689 16473 32723 16507
rect 34345 16473 34379 16507
rect 22569 16405 22603 16439
rect 24041 16405 24075 16439
rect 25427 16405 25461 16439
rect 26525 16405 26559 16439
rect 27813 16405 27847 16439
rect 29929 16405 29963 16439
rect 30849 16405 30883 16439
rect 22385 16201 22419 16235
rect 23029 16201 23063 16235
rect 24501 16201 24535 16235
rect 25329 16201 25363 16235
rect 29929 16201 29963 16235
rect 30665 16201 30699 16235
rect 31493 16201 31527 16235
rect 32413 16201 32447 16235
rect 33057 16201 33091 16235
rect 33793 16201 33827 16235
rect 23673 16133 23707 16167
rect 23857 16133 23891 16167
rect 29285 16133 29319 16167
rect 22109 16065 22143 16099
rect 22937 16065 22971 16099
rect 23121 16065 23155 16099
rect 23949 16065 23983 16099
rect 24409 16065 24443 16099
rect 25329 16065 25363 16099
rect 25421 16065 25455 16099
rect 26065 16065 26099 16099
rect 27445 16065 27479 16099
rect 27537 16065 27571 16099
rect 28365 16065 28399 16099
rect 29193 16065 29227 16099
rect 29377 16065 29411 16099
rect 29837 16065 29871 16099
rect 30021 16065 30055 16099
rect 30481 16065 30515 16099
rect 30665 16065 30699 16099
rect 31401 16065 31435 16099
rect 32321 16065 32355 16099
rect 32965 16065 32999 16099
rect 33701 16065 33735 16099
rect 33885 16065 33919 16099
rect 22201 15997 22235 16031
rect 22385 15997 22419 16031
rect 25605 15997 25639 16031
rect 26341 15997 26375 16031
rect 28457 15997 28491 16031
rect 23673 15929 23707 15963
rect 26157 15929 26191 15963
rect 28733 15929 28767 15963
rect 2053 15861 2087 15895
rect 26249 15861 26283 15895
rect 27721 15861 27755 15895
rect 23029 15657 23063 15691
rect 23857 15657 23891 15691
rect 25145 15657 25179 15691
rect 26617 15657 26651 15691
rect 27445 15657 27479 15691
rect 28273 15657 28307 15691
rect 30665 15657 30699 15691
rect 31401 15657 31435 15691
rect 32045 15657 32079 15691
rect 32597 15657 32631 15691
rect 33885 15657 33919 15691
rect 25789 15589 25823 15623
rect 1593 15521 1627 15555
rect 2789 15521 2823 15555
rect 23029 15453 23063 15487
rect 23213 15453 23247 15487
rect 23857 15453 23891 15487
rect 24041 15453 24075 15487
rect 25145 15453 25179 15487
rect 25329 15453 25363 15487
rect 25789 15453 25823 15487
rect 25973 15453 26007 15487
rect 26893 15453 26927 15487
rect 27353 15453 27387 15487
rect 28457 15453 28491 15487
rect 28733 15453 28767 15487
rect 29745 15453 29779 15487
rect 29929 15453 29963 15487
rect 30665 15453 30699 15487
rect 30849 15453 30883 15487
rect 31309 15453 31343 15487
rect 31953 15453 31987 15487
rect 32597 15453 32631 15487
rect 32781 15453 32815 15487
rect 33793 15453 33827 15487
rect 1777 15385 1811 15419
rect 26617 15385 26651 15419
rect 26801 15385 26835 15419
rect 28641 15317 28675 15351
rect 29837 15317 29871 15351
rect 2237 15113 2271 15147
rect 24869 15113 24903 15147
rect 25605 15113 25639 15147
rect 26157 15113 26191 15147
rect 27261 15113 27295 15147
rect 28089 15113 28123 15147
rect 29377 15113 29411 15147
rect 30021 15113 30055 15147
rect 32413 15113 32447 15147
rect 33057 15113 33091 15147
rect 28733 15045 28767 15079
rect 31309 15045 31343 15079
rect 2145 14977 2179 15011
rect 2789 14977 2823 15011
rect 24777 14977 24811 15011
rect 25421 14977 25455 15011
rect 25605 14977 25639 15011
rect 26065 14977 26099 15011
rect 27169 14977 27203 15011
rect 27997 14977 28031 15011
rect 28641 14977 28675 15011
rect 28825 14977 28859 15011
rect 29285 14977 29319 15011
rect 29929 14977 29963 15011
rect 31217 14977 31251 15011
rect 32321 14977 32355 15011
rect 32965 14977 32999 15011
rect 33793 14977 33827 15011
rect 30757 14909 30791 14943
rect 2881 14773 2915 14807
rect 26617 14569 26651 14603
rect 31033 14569 31067 14603
rect 31769 14569 31803 14603
rect 26065 14501 26099 14535
rect 1777 14433 1811 14467
rect 2789 14433 2823 14467
rect 30481 14433 30515 14467
rect 32505 14433 32539 14467
rect 1593 14365 1627 14399
rect 25145 14365 25179 14399
rect 25973 14365 26007 14399
rect 26617 14365 26651 14399
rect 26801 14365 26835 14399
rect 30941 14365 30975 14399
rect 34345 14365 34379 14399
rect 25237 14297 25271 14331
rect 32689 14297 32723 14331
rect 30389 14025 30423 14059
rect 31677 14025 31711 14059
rect 31033 13957 31067 13991
rect 32689 13957 32723 13991
rect 30297 13889 30331 13923
rect 30941 13889 30975 13923
rect 31585 13889 31619 13923
rect 1777 13821 1811 13855
rect 1961 13821 1995 13855
rect 2789 13821 2823 13855
rect 32505 13821 32539 13855
rect 34345 13821 34379 13855
rect 2697 13481 2731 13515
rect 31217 13481 31251 13515
rect 31861 13481 31895 13515
rect 32597 13481 32631 13515
rect 33609 13481 33643 13515
rect 2053 13413 2087 13447
rect 31125 13277 31159 13311
rect 31769 13277 31803 13311
rect 33793 13277 33827 13311
rect 2145 12937 2179 12971
rect 34345 12869 34379 12903
rect 2053 12801 2087 12835
rect 31401 12733 31435 12767
rect 32505 12733 32539 12767
rect 32689 12733 32723 12767
rect 32045 12393 32079 12427
rect 32505 12257 32539 12291
rect 34345 12257 34379 12291
rect 2053 12189 2087 12223
rect 31217 12189 31251 12223
rect 31309 12121 31343 12155
rect 32689 12121 32723 12155
rect 2145 12053 2179 12087
rect 1961 11781 1995 11815
rect 32689 11713 32723 11747
rect 33333 11713 33367 11747
rect 33977 11713 34011 11747
rect 1777 11645 1811 11679
rect 2789 11645 2823 11679
rect 2053 11305 2087 11339
rect 33241 11305 33275 11339
rect 33977 11305 34011 11339
rect 2697 11101 2731 11135
rect 33149 11101 33183 11135
rect 33885 10761 33919 10795
rect 1777 10625 1811 10659
rect 33333 10625 33367 10659
rect 33793 10625 33827 10659
rect 1961 10557 1995 10591
rect 2789 10557 2823 10591
rect 2053 10217 2087 10251
rect 34253 10217 34287 10251
rect 1961 10013 1995 10047
rect 34069 10013 34103 10047
rect 2513 9537 2547 9571
rect 2053 9333 2087 9367
rect 2605 9333 2639 9367
rect 1593 8993 1627 9027
rect 1777 8993 1811 9027
rect 2789 8993 2823 9027
rect 33977 8925 34011 8959
rect 34345 8517 34379 8551
rect 32505 8449 32539 8483
rect 1777 8381 1811 8415
rect 1961 8381 1995 8415
rect 2789 8381 2823 8415
rect 32689 8381 32723 8415
rect 2053 8041 2087 8075
rect 2605 8041 2639 8075
rect 33885 8041 33919 8075
rect 2513 7837 2547 7871
rect 3341 7837 3375 7871
rect 33333 7837 33367 7871
rect 33793 7837 33827 7871
rect 1777 7361 1811 7395
rect 33149 7361 33183 7395
rect 1961 7293 1995 7327
rect 2789 7293 2823 7327
rect 4261 7157 4295 7191
rect 33241 7157 33275 7191
rect 33977 7157 34011 7191
rect 2145 6953 2179 6987
rect 32689 6817 32723 6851
rect 34345 6817 34379 6851
rect 2053 6749 2087 6783
rect 2697 6749 2731 6783
rect 4169 6749 4203 6783
rect 4629 6749 4663 6783
rect 5457 6749 5491 6783
rect 9321 6749 9355 6783
rect 31861 6749 31895 6783
rect 32505 6749 32539 6783
rect 9965 6681 9999 6715
rect 2789 6613 2823 6647
rect 4721 6613 4755 6647
rect 31953 6613 31987 6647
rect 1961 6341 1995 6375
rect 31677 6341 31711 6375
rect 32689 6341 32723 6375
rect 1777 6273 1811 6307
rect 4721 6273 4755 6307
rect 31585 6273 31619 6307
rect 2881 6205 2915 6239
rect 32505 6205 32539 6239
rect 34345 6205 34379 6239
rect 5549 6137 5583 6171
rect 4261 6069 4295 6103
rect 4813 6069 4847 6103
rect 1593 5729 1627 5763
rect 1777 5729 1811 5763
rect 4077 5729 4111 5763
rect 32505 5729 32539 5763
rect 3985 5661 4019 5695
rect 4629 5661 4663 5695
rect 5273 5661 5307 5695
rect 6101 5661 6135 5695
rect 6561 5661 6595 5695
rect 7389 5661 7423 5695
rect 30757 5661 30791 5695
rect 31401 5661 31435 5695
rect 32045 5661 32079 5695
rect 3433 5593 3467 5627
rect 5365 5593 5399 5627
rect 32689 5593 32723 5627
rect 34345 5593 34379 5627
rect 4721 5525 4755 5559
rect 6653 5525 6687 5559
rect 1961 5253 1995 5287
rect 4261 5253 4295 5287
rect 7297 5253 7331 5287
rect 32689 5253 32723 5287
rect 6561 5185 6595 5219
rect 7205 5185 7239 5219
rect 29929 5185 29963 5219
rect 32505 5185 32539 5219
rect 1777 5117 1811 5151
rect 2789 5117 2823 5151
rect 4077 5117 4111 5151
rect 4997 5117 5031 5151
rect 33057 5117 33091 5151
rect 6653 4981 6687 5015
rect 30021 4981 30055 5015
rect 31217 4981 31251 5015
rect 1593 4641 1627 4675
rect 1777 4641 1811 4675
rect 2789 4641 2823 4675
rect 4169 4641 4203 4675
rect 4905 4641 4939 4675
rect 32505 4641 32539 4675
rect 32689 4641 32723 4675
rect 3985 4573 4019 4607
rect 6469 4573 6503 4607
rect 6929 4573 6963 4607
rect 7573 4573 7607 4607
rect 8401 4573 8435 4607
rect 19993 4573 20027 4607
rect 29193 4573 29227 4607
rect 30205 4573 30239 4607
rect 7665 4505 7699 4539
rect 30389 4505 30423 4539
rect 32045 4505 32079 4539
rect 34345 4505 34379 4539
rect 7021 4437 7055 4471
rect 20085 4437 20119 4471
rect 19809 4165 19843 4199
rect 2053 4097 2087 4131
rect 4997 4097 5031 4131
rect 5641 4097 5675 4131
rect 6561 4097 6595 4131
rect 8033 4097 8067 4131
rect 9137 4097 9171 4131
rect 28825 4097 28859 4131
rect 32505 4097 32539 4131
rect 2605 4029 2639 4063
rect 2789 4029 2823 4063
rect 4261 4029 4295 4063
rect 7389 4029 7423 4063
rect 13093 4029 13127 4063
rect 13277 4029 13311 4063
rect 13553 4029 13587 4063
rect 19625 4029 19659 4063
rect 20637 4029 20671 4063
rect 29929 4029 29963 4063
rect 30113 4029 30147 4063
rect 31769 4029 31803 4063
rect 32689 4029 32723 4063
rect 34345 4029 34379 4063
rect 5089 3893 5123 3927
rect 5733 3893 5767 3927
rect 6653 3893 6687 3927
rect 8125 3893 8159 3927
rect 9229 3893 9263 3927
rect 15761 3893 15795 3927
rect 17049 3893 17083 3927
rect 29469 3893 29503 3927
rect 13093 3689 13127 3723
rect 20269 3689 20303 3723
rect 27905 3689 27939 3723
rect 28457 3689 28491 3723
rect 34069 3689 34103 3723
rect 1593 3553 1627 3587
rect 2789 3553 2823 3587
rect 6101 3553 6135 3587
rect 6469 3553 6503 3587
rect 15577 3553 15611 3587
rect 16129 3553 16163 3587
rect 21281 3553 21315 3587
rect 31033 3553 31067 3587
rect 4169 3485 4203 3519
rect 4813 3485 4847 3519
rect 5457 3485 5491 3519
rect 5917 3485 5951 3519
rect 8401 3485 8435 3519
rect 9321 3485 9355 3519
rect 10057 3485 10091 3519
rect 10517 3485 10551 3519
rect 13737 3485 13771 3519
rect 14381 3485 14415 3519
rect 19625 3485 19659 3519
rect 20729 3485 20763 3519
rect 23857 3485 23891 3519
rect 24777 3485 24811 3519
rect 28365 3485 28399 3519
rect 29009 3485 29043 3519
rect 29929 3485 29963 3519
rect 30573 3485 30607 3519
rect 33517 3485 33551 3519
rect 33977 3485 34011 3519
rect 1777 3417 1811 3451
rect 15761 3417 15795 3451
rect 20913 3417 20947 3451
rect 31217 3417 31251 3451
rect 32873 3417 32907 3451
rect 10609 3349 10643 3383
rect 14473 3349 14507 3383
rect 23949 3349 23983 3383
rect 29101 3349 29135 3383
rect 13277 3145 13311 3179
rect 22109 3145 22143 3179
rect 27813 3145 27847 3179
rect 2053 3077 2087 3111
rect 4353 3077 4387 3111
rect 7205 3077 7239 3111
rect 9505 3077 9539 3111
rect 14473 3077 14507 3111
rect 24041 3077 24075 3111
rect 29101 3077 29135 3111
rect 29837 3077 29871 3111
rect 32505 3077 32539 3111
rect 7021 3009 7055 3043
rect 13185 3009 13219 3043
rect 14289 3009 14323 3043
rect 16865 3009 16899 3043
rect 19441 3009 19475 3043
rect 22017 3009 22051 3043
rect 23857 3009 23891 3043
rect 27721 3009 27755 3043
rect 28365 3009 28399 3043
rect 29009 3009 29043 3043
rect 29653 3009 29687 3043
rect 1869 2941 1903 2975
rect 3249 2941 3283 2975
rect 4169 2941 4203 2975
rect 5089 2941 5123 2975
rect 8401 2941 8435 2975
rect 9321 2941 9355 2975
rect 10333 2941 10367 2975
rect 14841 2941 14875 2975
rect 17049 2941 17083 2975
rect 17417 2941 17451 2975
rect 19625 2941 19659 2975
rect 19993 2941 20027 2975
rect 24501 2941 24535 2975
rect 30297 2941 30331 2975
rect 32321 2941 32355 2975
rect 33701 2941 33735 2975
rect 28457 2805 28491 2839
rect 15761 2601 15795 2635
rect 17049 2601 17083 2635
rect 18153 2601 18187 2635
rect 19533 2601 19567 2635
rect 21005 2601 21039 2635
rect 27813 2601 27847 2635
rect 28457 2533 28491 2567
rect 1593 2465 1627 2499
rect 2605 2465 2639 2499
rect 4169 2465 4203 2499
rect 4629 2465 4663 2499
rect 6561 2465 6595 2499
rect 6745 2465 6779 2499
rect 7021 2465 7055 2499
rect 9137 2465 9171 2499
rect 9781 2465 9815 2499
rect 29929 2465 29963 2499
rect 30941 2465 30975 2499
rect 32321 2465 32355 2499
rect 32873 2465 32907 2499
rect 15669 2397 15703 2431
rect 16957 2397 16991 2431
rect 18337 2397 18371 2431
rect 19441 2397 19475 2431
rect 27721 2397 27755 2431
rect 28365 2397 28399 2431
rect 29009 2397 29043 2431
rect 1777 2329 1811 2363
rect 4353 2329 4387 2363
rect 9321 2329 9355 2363
rect 29101 2329 29135 2363
rect 30113 2329 30147 2363
rect 32505 2329 32539 2363
<< metal1 >>
rect 20346 39992 20352 40044
rect 20404 40032 20410 40044
rect 32490 40032 32496 40044
rect 20404 40004 32496 40032
rect 20404 39992 20410 40004
rect 32490 39992 32496 40004
rect 32548 39992 32554 40044
rect 23934 39788 23940 39840
rect 23992 39828 23998 39840
rect 32582 39828 32588 39840
rect 23992 39800 32588 39828
rect 23992 39788 23998 39800
rect 32582 39788 32588 39800
rect 32640 39788 32646 39840
rect 1104 39738 34868 39760
rect 1104 39686 5170 39738
rect 5222 39686 5234 39738
rect 5286 39686 5298 39738
rect 5350 39686 5362 39738
rect 5414 39686 5426 39738
rect 5478 39686 13611 39738
rect 13663 39686 13675 39738
rect 13727 39686 13739 39738
rect 13791 39686 13803 39738
rect 13855 39686 13867 39738
rect 13919 39686 22052 39738
rect 22104 39686 22116 39738
rect 22168 39686 22180 39738
rect 22232 39686 22244 39738
rect 22296 39686 22308 39738
rect 22360 39686 30493 39738
rect 30545 39686 30557 39738
rect 30609 39686 30621 39738
rect 30673 39686 30685 39738
rect 30737 39686 30749 39738
rect 30801 39686 34868 39738
rect 1104 39664 34868 39686
rect 18966 39584 18972 39636
rect 19024 39624 19030 39636
rect 23934 39624 23940 39636
rect 19024 39596 22094 39624
rect 23895 39596 23940 39624
rect 19024 39584 19030 39596
rect 9953 39559 10011 39565
rect 9953 39556 9965 39559
rect 1596 39528 9965 39556
rect 1596 39497 1624 39528
rect 9953 39525 9965 39528
rect 9999 39525 10011 39559
rect 22066 39556 22094 39596
rect 23934 39584 23940 39596
rect 23992 39584 23998 39636
rect 25222 39584 25228 39636
rect 25280 39624 25286 39636
rect 27249 39627 27307 39633
rect 27249 39624 27261 39627
rect 25280 39596 27261 39624
rect 25280 39584 25286 39596
rect 27249 39593 27261 39596
rect 27295 39593 27307 39627
rect 27249 39587 27307 39593
rect 28077 39627 28135 39633
rect 28077 39593 28089 39627
rect 28123 39624 28135 39627
rect 29825 39627 29883 39633
rect 28123 39596 29776 39624
rect 28123 39593 28135 39596
rect 28077 39587 28135 39593
rect 29454 39556 29460 39568
rect 22066 39528 29460 39556
rect 9953 39519 10011 39525
rect 29454 39516 29460 39528
rect 29512 39516 29518 39568
rect 29748 39556 29776 39596
rect 29825 39593 29837 39627
rect 29871 39624 29883 39627
rect 32398 39624 32404 39636
rect 29871 39596 32404 39624
rect 29871 39593 29883 39596
rect 29825 39587 29883 39593
rect 32398 39584 32404 39596
rect 32456 39584 32462 39636
rect 31294 39556 31300 39568
rect 29748 39528 31300 39556
rect 31294 39516 31300 39528
rect 31352 39516 31358 39568
rect 1581 39491 1639 39497
rect 1581 39457 1593 39491
rect 1627 39457 1639 39491
rect 1581 39451 1639 39457
rect 1765 39491 1823 39497
rect 1765 39457 1777 39491
rect 1811 39488 1823 39491
rect 7098 39488 7104 39500
rect 1811 39460 5488 39488
rect 7059 39460 7104 39488
rect 1811 39457 1823 39460
rect 1765 39451 1823 39457
rect 3878 39380 3884 39432
rect 3936 39420 3942 39432
rect 3973 39423 4031 39429
rect 3973 39420 3985 39423
rect 3936 39392 3985 39420
rect 3936 39380 3942 39392
rect 3973 39389 3985 39392
rect 4019 39389 4031 39423
rect 3973 39383 4031 39389
rect 4154 39380 4160 39432
rect 4212 39420 4218 39432
rect 5353 39423 5411 39429
rect 5353 39420 5365 39423
rect 4212 39392 5365 39420
rect 4212 39380 4218 39392
rect 5353 39389 5365 39392
rect 5399 39389 5411 39423
rect 5353 39383 5411 39389
rect 1302 39312 1308 39364
rect 1360 39352 1366 39364
rect 3421 39355 3479 39361
rect 3421 39352 3433 39355
rect 1360 39324 3433 39352
rect 1360 39312 1366 39324
rect 3421 39321 3433 39324
rect 3467 39321 3479 39355
rect 3421 39315 3479 39321
rect 3234 39244 3240 39296
rect 3292 39284 3298 39296
rect 4065 39287 4123 39293
rect 4065 39284 4077 39287
rect 3292 39256 4077 39284
rect 3292 39244 3298 39256
rect 4065 39253 4077 39256
rect 4111 39253 4123 39287
rect 5460 39284 5488 39460
rect 7098 39448 7104 39460
rect 7156 39448 7162 39500
rect 14826 39488 14832 39500
rect 14787 39460 14832 39488
rect 14826 39448 14832 39460
rect 14884 39448 14890 39500
rect 21361 39491 21419 39497
rect 17604 39460 21220 39488
rect 5997 39423 6055 39429
rect 5997 39389 6009 39423
rect 6043 39420 6055 39423
rect 6549 39423 6607 39429
rect 6549 39420 6561 39423
rect 6043 39392 6561 39420
rect 6043 39389 6055 39392
rect 5997 39383 6055 39389
rect 6549 39389 6561 39392
rect 6595 39389 6607 39423
rect 9306 39420 9312 39432
rect 9267 39392 9312 39420
rect 6549 39383 6607 39389
rect 9306 39380 9312 39392
rect 9364 39380 9370 39432
rect 13265 39423 13323 39429
rect 13265 39389 13277 39423
rect 13311 39420 13323 39423
rect 13722 39420 13728 39432
rect 13311 39392 13728 39420
rect 13311 39389 13323 39392
rect 13265 39383 13323 39389
rect 13722 39380 13728 39392
rect 13780 39380 13786 39432
rect 13998 39380 14004 39432
rect 14056 39420 14062 39432
rect 14277 39423 14335 39429
rect 14277 39420 14289 39423
rect 14056 39392 14289 39420
rect 14056 39380 14062 39392
rect 14277 39389 14289 39392
rect 14323 39389 14335 39423
rect 16850 39420 16856 39432
rect 16763 39392 16856 39420
rect 14277 39383 14335 39389
rect 16850 39380 16856 39392
rect 16908 39420 16914 39432
rect 16908 39392 17264 39420
rect 16908 39380 16914 39392
rect 6730 39352 6736 39364
rect 6691 39324 6736 39352
rect 6730 39312 6736 39324
rect 6788 39312 6794 39364
rect 14458 39352 14464 39364
rect 14419 39324 14464 39352
rect 14458 39312 14464 39324
rect 14516 39312 14522 39364
rect 17236 39352 17264 39392
rect 17310 39380 17316 39432
rect 17368 39420 17374 39432
rect 17604 39429 17632 39460
rect 17589 39423 17647 39429
rect 17589 39420 17601 39423
rect 17368 39392 17601 39420
rect 17368 39380 17374 39392
rect 17589 39389 17601 39392
rect 17635 39389 17647 39423
rect 17589 39383 17647 39389
rect 18690 39380 18696 39432
rect 18748 39420 18754 39432
rect 18877 39423 18935 39429
rect 18877 39420 18889 39423
rect 18748 39392 18889 39420
rect 18748 39380 18754 39392
rect 18877 39389 18889 39392
rect 18923 39389 18935 39423
rect 18877 39383 18935 39389
rect 19150 39380 19156 39432
rect 19208 39420 19214 39432
rect 19613 39423 19671 39429
rect 19613 39420 19625 39423
rect 19208 39392 19625 39420
rect 19208 39380 19214 39392
rect 19613 39389 19625 39392
rect 19659 39389 19671 39423
rect 20254 39420 20260 39432
rect 20215 39392 20260 39420
rect 19613 39383 19671 39389
rect 20254 39380 20260 39392
rect 20312 39380 20318 39432
rect 21192 39420 21220 39460
rect 21361 39457 21373 39491
rect 21407 39488 21419 39491
rect 32677 39491 32735 39497
rect 32677 39488 32689 39491
rect 21407 39460 32689 39488
rect 21407 39457 21419 39460
rect 21361 39451 21419 39457
rect 32677 39457 32689 39460
rect 32723 39457 32735 39491
rect 32677 39451 32735 39457
rect 21277 39423 21335 39429
rect 21277 39420 21289 39423
rect 21192 39392 21289 39420
rect 21277 39389 21289 39392
rect 21323 39420 21335 39423
rect 21450 39420 21456 39432
rect 21323 39392 21456 39420
rect 21323 39389 21335 39392
rect 21277 39383 21335 39389
rect 21450 39380 21456 39392
rect 21508 39380 21514 39432
rect 22094 39380 22100 39432
rect 22152 39420 22158 39432
rect 22189 39423 22247 39429
rect 22189 39420 22201 39423
rect 22152 39392 22201 39420
rect 22152 39380 22158 39392
rect 22189 39389 22201 39392
rect 22235 39389 22247 39423
rect 23382 39420 23388 39432
rect 23343 39392 23388 39420
rect 22189 39383 22247 39389
rect 23382 39380 23388 39392
rect 23440 39380 23446 39432
rect 23842 39420 23848 39432
rect 23803 39392 23848 39420
rect 23842 39380 23848 39392
rect 23900 39380 23906 39432
rect 24581 39423 24639 39429
rect 24581 39420 24593 39423
rect 23952 39392 24593 39420
rect 23952 39352 23980 39392
rect 24581 39389 24593 39392
rect 24627 39389 24639 39423
rect 24581 39383 24639 39389
rect 25409 39423 25467 39429
rect 25409 39389 25421 39423
rect 25455 39389 25467 39423
rect 26050 39420 26056 39432
rect 26011 39392 26056 39420
rect 25409 39383 25467 39389
rect 17236 39324 23980 39352
rect 24394 39312 24400 39364
rect 24452 39352 24458 39364
rect 25424 39352 25452 39383
rect 26050 39380 26056 39392
rect 26108 39380 26114 39432
rect 27249 39423 27307 39429
rect 27249 39389 27261 39423
rect 27295 39389 27307 39423
rect 27249 39383 27307 39389
rect 27433 39423 27491 39429
rect 27433 39389 27445 39423
rect 27479 39420 27491 39423
rect 28442 39420 28448 39432
rect 27479 39392 28448 39420
rect 27479 39389 27491 39392
rect 27433 39383 27491 39389
rect 24452 39324 25452 39352
rect 24452 39312 24458 39324
rect 7282 39284 7288 39296
rect 5460 39256 7288 39284
rect 4065 39247 4123 39253
rect 7282 39244 7288 39256
rect 7340 39244 7346 39296
rect 13446 39244 13452 39296
rect 13504 39284 13510 39296
rect 13541 39287 13599 39293
rect 13541 39284 13553 39287
rect 13504 39256 13553 39284
rect 13504 39244 13510 39256
rect 13541 39253 13553 39256
rect 13587 39253 13599 39287
rect 13541 39247 13599 39253
rect 16574 39244 16580 39296
rect 16632 39284 16638 39296
rect 16945 39287 17003 39293
rect 16945 39284 16957 39287
rect 16632 39256 16957 39284
rect 16632 39244 16638 39256
rect 16945 39253 16957 39256
rect 16991 39253 17003 39287
rect 16945 39247 17003 39253
rect 17034 39244 17040 39296
rect 17092 39284 17098 39296
rect 17681 39287 17739 39293
rect 17681 39284 17693 39287
rect 17092 39256 17693 39284
rect 17092 39244 17098 39256
rect 17681 39253 17693 39256
rect 17727 39253 17739 39287
rect 17681 39247 17739 39253
rect 18322 39244 18328 39296
rect 18380 39284 18386 39296
rect 18693 39287 18751 39293
rect 18693 39284 18705 39287
rect 18380 39256 18705 39284
rect 18380 39244 18386 39256
rect 18693 39253 18705 39256
rect 18739 39253 18751 39287
rect 18693 39247 18751 39253
rect 22186 39244 22192 39296
rect 22244 39284 22250 39296
rect 22281 39287 22339 39293
rect 22281 39284 22293 39287
rect 22244 39256 22293 39284
rect 22244 39244 22250 39256
rect 22281 39253 22293 39256
rect 22327 39253 22339 39287
rect 22281 39247 22339 39253
rect 24578 39244 24584 39296
rect 24636 39284 24642 39296
rect 24673 39287 24731 39293
rect 24673 39284 24685 39287
rect 24636 39256 24685 39284
rect 24636 39244 24642 39256
rect 24673 39253 24685 39256
rect 24719 39253 24731 39287
rect 27264 39284 27292 39383
rect 28442 39380 28448 39392
rect 28500 39380 28506 39432
rect 28537 39423 28595 39429
rect 28537 39389 28549 39423
rect 28583 39389 28595 39423
rect 28537 39383 28595 39389
rect 28258 39312 28264 39364
rect 28316 39352 28322 39364
rect 28552 39352 28580 39383
rect 28626 39380 28632 39432
rect 28684 39420 28690 39432
rect 29733 39423 29791 39429
rect 29733 39420 29745 39423
rect 28684 39392 29745 39420
rect 28684 39380 28690 39392
rect 29733 39389 29745 39392
rect 29779 39389 29791 39423
rect 29733 39383 29791 39389
rect 29822 39380 29828 39432
rect 29880 39420 29886 39432
rect 29917 39423 29975 39429
rect 29917 39420 29929 39423
rect 29880 39392 29929 39420
rect 29880 39380 29886 39392
rect 29917 39389 29929 39392
rect 29963 39389 29975 39423
rect 30558 39420 30564 39432
rect 30519 39392 30564 39420
rect 29917 39383 29975 39389
rect 30558 39380 30564 39392
rect 30616 39380 30622 39432
rect 31205 39423 31263 39429
rect 31205 39420 31217 39423
rect 30760 39392 31217 39420
rect 28316 39324 28580 39352
rect 28316 39312 28322 39324
rect 30190 39312 30196 39364
rect 30248 39352 30254 39364
rect 30248 39324 30512 39352
rect 30248 39312 30254 39324
rect 28534 39284 28540 39296
rect 27264 39256 28540 39284
rect 24673 39247 24731 39253
rect 28534 39244 28540 39256
rect 28592 39244 28598 39296
rect 28629 39287 28687 39293
rect 28629 39253 28641 39287
rect 28675 39284 28687 39287
rect 29638 39284 29644 39296
rect 28675 39256 29644 39284
rect 28675 39253 28687 39256
rect 28629 39247 28687 39253
rect 29638 39244 29644 39256
rect 29696 39244 29702 39296
rect 30374 39284 30380 39296
rect 30335 39256 30380 39284
rect 30374 39244 30380 39256
rect 30432 39244 30438 39296
rect 30484 39284 30512 39324
rect 30760 39284 30788 39392
rect 31205 39389 31217 39392
rect 31251 39389 31263 39423
rect 32490 39420 32496 39432
rect 32451 39392 32496 39420
rect 31205 39383 31263 39389
rect 32490 39380 32496 39392
rect 32548 39380 32554 39432
rect 34330 39352 34336 39364
rect 34291 39324 34336 39352
rect 34330 39312 34336 39324
rect 34388 39312 34394 39364
rect 30484 39256 30788 39284
rect 30926 39244 30932 39296
rect 30984 39284 30990 39296
rect 31021 39287 31079 39293
rect 31021 39284 31033 39287
rect 30984 39256 31033 39284
rect 30984 39244 30990 39256
rect 31021 39253 31033 39256
rect 31067 39253 31079 39287
rect 31021 39247 31079 39253
rect 1104 39194 35027 39216
rect 1104 39142 9390 39194
rect 9442 39142 9454 39194
rect 9506 39142 9518 39194
rect 9570 39142 9582 39194
rect 9634 39142 9646 39194
rect 9698 39142 17831 39194
rect 17883 39142 17895 39194
rect 17947 39142 17959 39194
rect 18011 39142 18023 39194
rect 18075 39142 18087 39194
rect 18139 39142 26272 39194
rect 26324 39142 26336 39194
rect 26388 39142 26400 39194
rect 26452 39142 26464 39194
rect 26516 39142 26528 39194
rect 26580 39142 34713 39194
rect 34765 39142 34777 39194
rect 34829 39142 34841 39194
rect 34893 39142 34905 39194
rect 34957 39142 34969 39194
rect 35021 39142 35027 39194
rect 1104 39120 35027 39142
rect 3510 39040 3516 39092
rect 3568 39080 3574 39092
rect 3568 39052 10916 39080
rect 3568 39040 3574 39052
rect 1949 39015 2007 39021
rect 1949 38981 1961 39015
rect 1995 39012 2007 39015
rect 5074 39012 5080 39024
rect 1995 38984 5080 39012
rect 1995 38981 2007 38984
rect 1949 38975 2007 38981
rect 5074 38972 5080 38984
rect 5132 38972 5138 39024
rect 4154 38944 4160 38956
rect 4115 38916 4160 38944
rect 4154 38904 4160 38916
rect 4212 38904 4218 38956
rect 10888 38953 10916 39052
rect 23382 39040 23388 39092
rect 23440 39080 23446 39092
rect 23440 39052 31754 39080
rect 23440 39040 23446 39052
rect 17034 39012 17040 39024
rect 16995 38984 17040 39012
rect 17034 38972 17040 38984
rect 17092 38972 17098 39024
rect 22186 39012 22192 39024
rect 22147 38984 22192 39012
rect 22186 38972 22192 38984
rect 22244 38972 22250 39024
rect 24578 39012 24584 39024
rect 24539 38984 24584 39012
rect 24578 38972 24584 38984
rect 24636 38972 24642 39024
rect 26970 38972 26976 39024
rect 27028 39012 27034 39024
rect 28258 39012 28264 39024
rect 27028 38984 28264 39012
rect 27028 38972 27034 38984
rect 28258 38972 28264 38984
rect 28316 38972 28322 39024
rect 29638 39012 29644 39024
rect 29599 38984 29644 39012
rect 29638 38972 29644 38984
rect 29696 38972 29702 39024
rect 7101 38947 7159 38953
rect 7101 38913 7113 38947
rect 7147 38913 7159 38947
rect 7101 38907 7159 38913
rect 10873 38947 10931 38953
rect 10873 38913 10885 38947
rect 10919 38913 10931 38947
rect 13998 38944 14004 38956
rect 13959 38916 14004 38944
rect 10873 38907 10931 38913
rect 1765 38879 1823 38885
rect 1765 38845 1777 38879
rect 1811 38845 1823 38879
rect 2774 38876 2780 38888
rect 2735 38848 2780 38876
rect 1765 38839 1823 38845
rect 1780 38808 1808 38839
rect 2774 38836 2780 38848
rect 2832 38836 2838 38888
rect 4341 38879 4399 38885
rect 4341 38845 4353 38879
rect 4387 38876 4399 38879
rect 5534 38876 5540 38888
rect 4387 38848 5540 38876
rect 4387 38845 4399 38848
rect 4341 38839 4399 38845
rect 5534 38836 5540 38848
rect 5592 38836 5598 38888
rect 5810 38876 5816 38888
rect 5771 38848 5816 38876
rect 5810 38836 5816 38848
rect 5868 38836 5874 38888
rect 3970 38808 3976 38820
rect 1780 38780 3976 38808
rect 3970 38768 3976 38780
rect 4028 38768 4034 38820
rect 7116 38808 7144 38907
rect 13998 38904 14004 38916
rect 14056 38904 14062 38956
rect 19150 38944 19156 38956
rect 19111 38916 19156 38944
rect 19150 38904 19156 38916
rect 19208 38904 19214 38956
rect 24394 38944 24400 38956
rect 24355 38916 24400 38944
rect 24394 38904 24400 38916
rect 24452 38904 24458 38956
rect 29454 38944 29460 38956
rect 29415 38916 29460 38944
rect 29454 38904 29460 38916
rect 29512 38904 29518 38956
rect 31726 38944 31754 39052
rect 32582 39012 32588 39024
rect 32543 38984 32588 39012
rect 32582 38972 32588 38984
rect 32640 38972 32646 39024
rect 32401 38947 32459 38953
rect 32401 38944 32413 38947
rect 31726 38916 32413 38944
rect 32401 38913 32413 38916
rect 32447 38913 32459 38947
rect 32401 38907 32459 38913
rect 7929 38879 7987 38885
rect 7929 38845 7941 38879
rect 7975 38876 7987 38879
rect 8389 38879 8447 38885
rect 8389 38876 8401 38879
rect 7975 38848 8401 38876
rect 7975 38845 7987 38848
rect 7929 38839 7987 38845
rect 8389 38845 8401 38848
rect 8435 38845 8447 38879
rect 8570 38876 8576 38888
rect 8531 38848 8576 38876
rect 8389 38839 8447 38845
rect 8570 38836 8576 38848
rect 8628 38836 8634 38888
rect 9030 38876 9036 38888
rect 8991 38848 9036 38876
rect 9030 38836 9036 38848
rect 9088 38836 9094 38888
rect 14461 38879 14519 38885
rect 14461 38845 14473 38879
rect 14507 38845 14519 38879
rect 14461 38839 14519 38845
rect 14645 38879 14703 38885
rect 14645 38845 14657 38879
rect 14691 38876 14703 38879
rect 15194 38876 15200 38888
rect 14691 38848 15200 38876
rect 14691 38845 14703 38848
rect 14645 38839 14703 38845
rect 14366 38808 14372 38820
rect 6886 38780 14372 38808
rect 3878 38700 3884 38752
rect 3936 38740 3942 38752
rect 6886 38740 6914 38780
rect 14366 38768 14372 38780
rect 14424 38768 14430 38820
rect 14476 38808 14504 38839
rect 15194 38836 15200 38848
rect 15252 38836 15258 38888
rect 16114 38876 16120 38888
rect 16075 38848 16120 38876
rect 16114 38836 16120 38848
rect 16172 38836 16178 38888
rect 16853 38879 16911 38885
rect 16853 38845 16865 38879
rect 16899 38876 16911 38879
rect 17678 38876 17684 38888
rect 16899 38848 17684 38876
rect 16899 38845 16911 38848
rect 16853 38839 16911 38845
rect 17678 38836 17684 38848
rect 17736 38836 17742 38888
rect 18230 38876 18236 38888
rect 18191 38848 18236 38876
rect 18230 38836 18236 38848
rect 18288 38836 18294 38888
rect 19334 38876 19340 38888
rect 19295 38848 19340 38876
rect 19334 38836 19340 38848
rect 19392 38836 19398 38888
rect 19978 38876 19984 38888
rect 19939 38848 19984 38876
rect 19978 38836 19984 38848
rect 20036 38836 20042 38888
rect 22005 38879 22063 38885
rect 22005 38845 22017 38879
rect 22051 38876 22063 38879
rect 22370 38876 22376 38888
rect 22051 38848 22376 38876
rect 22051 38845 22063 38848
rect 22005 38839 22063 38845
rect 22370 38836 22376 38848
rect 22428 38836 22434 38888
rect 22554 38876 22560 38888
rect 22515 38848 22560 38876
rect 22554 38836 22560 38848
rect 22612 38836 22618 38888
rect 25130 38876 25136 38888
rect 25091 38848 25136 38876
rect 25130 38836 25136 38848
rect 25188 38836 25194 38888
rect 27157 38879 27215 38885
rect 27157 38845 27169 38879
rect 27203 38845 27215 38879
rect 27338 38876 27344 38888
rect 27299 38848 27344 38876
rect 27157 38839 27215 38845
rect 15654 38808 15660 38820
rect 14476 38780 15660 38808
rect 15654 38768 15660 38780
rect 15712 38768 15718 38820
rect 20530 38768 20536 38820
rect 20588 38808 20594 38820
rect 27172 38808 27200 38839
rect 27338 38836 27344 38848
rect 27396 38836 27402 38888
rect 27617 38879 27675 38885
rect 27617 38876 27629 38879
rect 27540 38848 27629 38876
rect 20588 38780 27200 38808
rect 20588 38768 20594 38780
rect 3936 38712 6914 38740
rect 7193 38743 7251 38749
rect 3936 38700 3942 38712
rect 7193 38709 7205 38743
rect 7239 38740 7251 38743
rect 8110 38740 8116 38752
rect 7239 38712 8116 38740
rect 7239 38709 7251 38712
rect 7193 38703 7251 38709
rect 8110 38700 8116 38712
rect 8168 38700 8174 38752
rect 10689 38743 10747 38749
rect 10689 38709 10701 38743
rect 10735 38740 10747 38743
rect 16666 38740 16672 38752
rect 10735 38712 16672 38740
rect 10735 38709 10747 38712
rect 10689 38703 10747 38709
rect 16666 38700 16672 38712
rect 16724 38700 16730 38752
rect 23842 38700 23848 38752
rect 23900 38740 23906 38752
rect 26970 38740 26976 38752
rect 23900 38712 26976 38740
rect 23900 38700 23906 38712
rect 26970 38700 26976 38712
rect 27028 38700 27034 38752
rect 27062 38700 27068 38752
rect 27120 38740 27126 38752
rect 27540 38740 27568 38848
rect 27617 38845 27629 38848
rect 27663 38845 27675 38879
rect 27617 38839 27675 38845
rect 29917 38879 29975 38885
rect 29917 38845 29929 38879
rect 29963 38845 29975 38879
rect 29917 38839 29975 38845
rect 28350 38768 28356 38820
rect 28408 38808 28414 38820
rect 29932 38808 29960 38839
rect 30558 38836 30564 38888
rect 30616 38876 30622 38888
rect 31846 38876 31852 38888
rect 30616 38848 31852 38876
rect 30616 38836 30622 38848
rect 31846 38836 31852 38848
rect 31904 38836 31910 38888
rect 32858 38876 32864 38888
rect 32819 38848 32864 38876
rect 32858 38836 32864 38848
rect 32916 38836 32922 38888
rect 28408 38780 29960 38808
rect 28408 38768 28414 38780
rect 27120 38712 27568 38740
rect 27120 38700 27126 38712
rect 28442 38700 28448 38752
rect 28500 38740 28506 38752
rect 32766 38740 32772 38752
rect 28500 38712 32772 38740
rect 28500 38700 28506 38712
rect 32766 38700 32772 38712
rect 32824 38700 32830 38752
rect 1104 38650 34868 38672
rect 1104 38598 5170 38650
rect 5222 38598 5234 38650
rect 5286 38598 5298 38650
rect 5350 38598 5362 38650
rect 5414 38598 5426 38650
rect 5478 38598 13611 38650
rect 13663 38598 13675 38650
rect 13727 38598 13739 38650
rect 13791 38598 13803 38650
rect 13855 38598 13867 38650
rect 13919 38598 22052 38650
rect 22104 38598 22116 38650
rect 22168 38598 22180 38650
rect 22232 38598 22244 38650
rect 22296 38598 22308 38650
rect 22360 38598 30493 38650
rect 30545 38598 30557 38650
rect 30609 38598 30621 38650
rect 30673 38598 30685 38650
rect 30737 38598 30749 38650
rect 30801 38598 34868 38650
rect 1104 38576 34868 38598
rect 5537 38539 5595 38545
rect 5537 38505 5549 38539
rect 5583 38536 5595 38539
rect 6730 38536 6736 38548
rect 5583 38508 6736 38536
rect 5583 38505 5595 38508
rect 5537 38499 5595 38505
rect 6730 38496 6736 38508
rect 6788 38496 6794 38548
rect 8570 38496 8576 38548
rect 8628 38536 8634 38548
rect 9217 38539 9275 38545
rect 9217 38536 9229 38539
rect 8628 38508 9229 38536
rect 8628 38496 8634 38508
rect 9217 38505 9229 38508
rect 9263 38505 9275 38539
rect 9217 38499 9275 38505
rect 14369 38539 14427 38545
rect 14369 38505 14381 38539
rect 14415 38536 14427 38539
rect 14458 38536 14464 38548
rect 14415 38508 14464 38536
rect 14415 38505 14427 38508
rect 14369 38499 14427 38505
rect 14458 38496 14464 38508
rect 14516 38496 14522 38548
rect 15194 38536 15200 38548
rect 15155 38508 15200 38536
rect 15194 38496 15200 38508
rect 15252 38496 15258 38548
rect 18785 38539 18843 38545
rect 18785 38505 18797 38539
rect 18831 38536 18843 38539
rect 19334 38536 19340 38548
rect 18831 38508 19340 38536
rect 18831 38505 18843 38508
rect 18785 38499 18843 38505
rect 19334 38496 19340 38508
rect 19392 38496 19398 38548
rect 22370 38496 22376 38548
rect 22428 38536 22434 38548
rect 22465 38539 22523 38545
rect 22465 38536 22477 38539
rect 22428 38508 22477 38536
rect 22428 38496 22434 38508
rect 22465 38505 22477 38508
rect 22511 38505 22523 38539
rect 22465 38499 22523 38505
rect 24029 38539 24087 38545
rect 24029 38505 24041 38539
rect 24075 38536 24087 38539
rect 29362 38536 29368 38548
rect 24075 38508 29368 38536
rect 24075 38505 24087 38508
rect 24029 38499 24087 38505
rect 29362 38496 29368 38508
rect 29420 38496 29426 38548
rect 9953 38471 10011 38477
rect 9953 38468 9965 38471
rect 1596 38440 9965 38468
rect 1596 38409 1624 38440
rect 9953 38437 9965 38440
rect 9999 38437 10011 38471
rect 9953 38431 10011 38437
rect 16022 38428 16028 38480
rect 16080 38468 16086 38480
rect 25038 38468 25044 38480
rect 16080 38440 25044 38468
rect 16080 38428 16086 38440
rect 25038 38428 25044 38440
rect 25096 38428 25102 38480
rect 25774 38428 25780 38480
rect 25832 38468 25838 38480
rect 25832 38440 26372 38468
rect 25832 38428 25838 38440
rect 1581 38403 1639 38409
rect 1581 38369 1593 38403
rect 1627 38369 1639 38403
rect 1581 38363 1639 38369
rect 1765 38403 1823 38409
rect 1765 38369 1777 38403
rect 1811 38400 1823 38403
rect 7742 38400 7748 38412
rect 1811 38372 5580 38400
rect 7703 38372 7748 38400
rect 1811 38369 1823 38372
rect 1765 38363 1823 38369
rect 3973 38335 4031 38341
rect 3973 38301 3985 38335
rect 4019 38301 4031 38335
rect 3973 38295 4031 38301
rect 658 38224 664 38276
rect 716 38264 722 38276
rect 3421 38267 3479 38273
rect 3421 38264 3433 38267
rect 716 38236 3433 38264
rect 716 38224 722 38236
rect 3421 38233 3433 38236
rect 3467 38233 3479 38267
rect 3988 38264 4016 38295
rect 4154 38292 4160 38344
rect 4212 38332 4218 38344
rect 4801 38335 4859 38341
rect 4801 38332 4813 38335
rect 4212 38304 4813 38332
rect 4212 38292 4218 38304
rect 4801 38301 4813 38304
rect 4847 38301 4859 38335
rect 4801 38295 4859 38301
rect 4890 38292 4896 38344
rect 4948 38332 4954 38344
rect 5445 38335 5503 38341
rect 5445 38332 5457 38335
rect 4948 38304 5457 38332
rect 4948 38292 4954 38304
rect 5445 38301 5457 38304
rect 5491 38301 5503 38335
rect 5445 38295 5503 38301
rect 4430 38264 4436 38276
rect 3988 38236 4436 38264
rect 3421 38227 3479 38233
rect 4430 38224 4436 38236
rect 4488 38224 4494 38276
rect 5552 38264 5580 38372
rect 7742 38360 7748 38372
rect 7800 38360 7806 38412
rect 16574 38400 16580 38412
rect 16535 38372 16580 38400
rect 16574 38360 16580 38372
rect 16632 38360 16638 38412
rect 17402 38400 17408 38412
rect 17363 38372 17408 38400
rect 17402 38360 17408 38372
rect 17460 38360 17466 38412
rect 19981 38403 20039 38409
rect 19981 38369 19993 38403
rect 20027 38400 20039 38403
rect 20254 38400 20260 38412
rect 20027 38372 20260 38400
rect 20027 38369 20039 38372
rect 19981 38363 20039 38369
rect 20254 38360 20260 38372
rect 20312 38360 20318 38412
rect 20622 38360 20628 38412
rect 20680 38400 20686 38412
rect 20717 38403 20775 38409
rect 20717 38400 20729 38403
rect 20680 38372 20729 38400
rect 20680 38360 20686 38372
rect 20717 38369 20729 38372
rect 20763 38369 20775 38403
rect 20717 38363 20775 38369
rect 24949 38403 25007 38409
rect 24949 38369 24961 38403
rect 24995 38400 25007 38403
rect 26050 38400 26056 38412
rect 24995 38372 26056 38400
rect 24995 38369 25007 38372
rect 24949 38363 25007 38369
rect 26050 38360 26056 38372
rect 26108 38360 26114 38412
rect 26344 38409 26372 38440
rect 26418 38428 26424 38480
rect 26476 38468 26482 38480
rect 26476 38440 32720 38468
rect 26476 38428 26482 38440
rect 26329 38403 26387 38409
rect 26329 38369 26341 38403
rect 26375 38369 26387 38403
rect 26329 38363 26387 38369
rect 26436 38372 28948 38400
rect 6273 38335 6331 38341
rect 6273 38301 6285 38335
rect 6319 38332 6331 38335
rect 6733 38335 6791 38341
rect 6733 38332 6745 38335
rect 6319 38304 6745 38332
rect 6319 38301 6331 38304
rect 6273 38295 6331 38301
rect 6733 38301 6745 38304
rect 6779 38301 6791 38335
rect 9122 38332 9128 38344
rect 9083 38304 9128 38332
rect 6733 38295 6791 38301
rect 9122 38292 9128 38304
rect 9180 38292 9186 38344
rect 14274 38332 14280 38344
rect 14235 38304 14280 38332
rect 14274 38292 14280 38304
rect 14332 38292 14338 38344
rect 14366 38292 14372 38344
rect 14424 38332 14430 38344
rect 15105 38335 15163 38341
rect 15105 38332 15117 38335
rect 14424 38304 15117 38332
rect 14424 38292 14430 38304
rect 15105 38301 15117 38304
rect 15151 38301 15163 38335
rect 15105 38295 15163 38301
rect 15933 38335 15991 38341
rect 15933 38301 15945 38335
rect 15979 38332 15991 38335
rect 16393 38335 16451 38341
rect 16393 38332 16405 38335
rect 15979 38304 16405 38332
rect 15979 38301 15991 38304
rect 15933 38295 15991 38301
rect 16393 38301 16405 38304
rect 16439 38301 16451 38335
rect 16393 38295 16451 38301
rect 6917 38267 6975 38273
rect 5552 38236 5672 38264
rect 4062 38196 4068 38208
rect 4023 38168 4068 38196
rect 4062 38156 4068 38168
rect 4120 38156 4126 38208
rect 5644 38196 5672 38236
rect 6917 38233 6929 38267
rect 6963 38264 6975 38267
rect 7190 38264 7196 38276
rect 6963 38236 7196 38264
rect 6963 38233 6975 38236
rect 6917 38227 6975 38233
rect 7190 38224 7196 38236
rect 7248 38224 7254 38276
rect 15120 38264 15148 38295
rect 18598 38292 18604 38344
rect 18656 38332 18662 38344
rect 18693 38335 18751 38341
rect 18693 38332 18705 38335
rect 18656 38304 18705 38332
rect 18656 38292 18662 38304
rect 18693 38301 18705 38304
rect 18739 38301 18751 38335
rect 18693 38295 18751 38301
rect 23385 38335 23443 38341
rect 23385 38301 23397 38335
rect 23431 38332 23443 38335
rect 24854 38332 24860 38344
rect 23431 38304 24860 38332
rect 23431 38301 23443 38304
rect 23385 38295 23443 38301
rect 24854 38292 24860 38304
rect 24912 38292 24918 38344
rect 16850 38264 16856 38276
rect 15120 38236 16856 38264
rect 16850 38224 16856 38236
rect 16908 38224 16914 38276
rect 20162 38264 20168 38276
rect 20123 38236 20168 38264
rect 20162 38224 20168 38236
rect 20220 38224 20226 38276
rect 25130 38224 25136 38276
rect 25188 38264 25194 38276
rect 25188 38236 25233 38264
rect 25188 38224 25194 38236
rect 7466 38196 7472 38208
rect 5644 38168 7472 38196
rect 7466 38156 7472 38168
rect 7524 38156 7530 38208
rect 18230 38156 18236 38208
rect 18288 38196 18294 38208
rect 24302 38196 24308 38208
rect 18288 38168 24308 38196
rect 18288 38156 18294 38168
rect 24302 38156 24308 38168
rect 24360 38156 24366 38208
rect 24486 38156 24492 38208
rect 24544 38196 24550 38208
rect 26436 38196 26464 38372
rect 27430 38332 27436 38344
rect 27391 38304 27436 38332
rect 27430 38292 27436 38304
rect 27488 38292 27494 38344
rect 27614 38292 27620 38344
rect 27672 38332 27678 38344
rect 27985 38335 28043 38341
rect 27985 38332 27997 38335
rect 27672 38304 27997 38332
rect 27672 38292 27678 38304
rect 27985 38301 27997 38304
rect 28031 38301 28043 38335
rect 27985 38295 28043 38301
rect 28813 38335 28871 38341
rect 28813 38301 28825 38335
rect 28859 38301 28871 38335
rect 28813 38295 28871 38301
rect 28074 38196 28080 38208
rect 24544 38168 26464 38196
rect 28035 38168 28080 38196
rect 24544 38156 24550 38168
rect 28074 38156 28080 38168
rect 28132 38156 28138 38208
rect 28350 38156 28356 38208
rect 28408 38196 28414 38208
rect 28629 38199 28687 38205
rect 28629 38196 28641 38199
rect 28408 38168 28641 38196
rect 28408 38156 28414 38168
rect 28629 38165 28641 38168
rect 28675 38165 28687 38199
rect 28828 38196 28856 38295
rect 28920 38264 28948 38372
rect 29362 38360 29368 38412
rect 29420 38400 29426 38412
rect 32692 38409 32720 38440
rect 29825 38403 29883 38409
rect 29825 38400 29837 38403
rect 29420 38372 29837 38400
rect 29420 38360 29426 38372
rect 29825 38369 29837 38372
rect 29871 38369 29883 38403
rect 29825 38363 29883 38369
rect 32677 38403 32735 38409
rect 32677 38369 32689 38403
rect 32723 38369 32735 38403
rect 34146 38400 34152 38412
rect 34107 38372 34152 38400
rect 32677 38363 32735 38369
rect 34146 38360 34152 38372
rect 34204 38360 34210 38412
rect 31665 38335 31723 38341
rect 31665 38301 31677 38335
rect 31711 38332 31723 38335
rect 32214 38332 32220 38344
rect 31711 38304 32220 38332
rect 31711 38301 31723 38304
rect 31665 38295 31723 38301
rect 32214 38292 32220 38304
rect 32272 38292 32278 38344
rect 32493 38335 32551 38341
rect 32493 38301 32505 38335
rect 32539 38301 32551 38335
rect 32493 38295 32551 38301
rect 30009 38267 30067 38273
rect 30009 38264 30021 38267
rect 28920 38236 30021 38264
rect 30009 38233 30021 38236
rect 30055 38233 30067 38267
rect 30009 38227 30067 38233
rect 30282 38224 30288 38276
rect 30340 38264 30346 38276
rect 32508 38264 32536 38295
rect 30340 38236 32536 38264
rect 30340 38224 30346 38236
rect 31202 38196 31208 38208
rect 28828 38168 31208 38196
rect 28629 38159 28687 38165
rect 31202 38156 31208 38168
rect 31260 38156 31266 38208
rect 1104 38106 35027 38128
rect 1104 38054 9390 38106
rect 9442 38054 9454 38106
rect 9506 38054 9518 38106
rect 9570 38054 9582 38106
rect 9634 38054 9646 38106
rect 9698 38054 17831 38106
rect 17883 38054 17895 38106
rect 17947 38054 17959 38106
rect 18011 38054 18023 38106
rect 18075 38054 18087 38106
rect 18139 38054 26272 38106
rect 26324 38054 26336 38106
rect 26388 38054 26400 38106
rect 26452 38054 26464 38106
rect 26516 38054 26528 38106
rect 26580 38054 34713 38106
rect 34765 38054 34777 38106
rect 34829 38054 34841 38106
rect 34893 38054 34905 38106
rect 34957 38054 34969 38106
rect 35021 38054 35027 38106
rect 1104 38032 35027 38054
rect 5534 37992 5540 38004
rect 5495 37964 5540 37992
rect 5534 37952 5540 37964
rect 5592 37952 5598 38004
rect 7190 37992 7196 38004
rect 7151 37964 7196 37992
rect 7190 37952 7196 37964
rect 7248 37952 7254 38004
rect 9122 37952 9128 38004
rect 9180 37992 9186 38004
rect 18690 37992 18696 38004
rect 9180 37964 18696 37992
rect 9180 37952 9186 37964
rect 18690 37952 18696 37964
rect 18748 37952 18754 38004
rect 20162 37992 20168 38004
rect 20123 37964 20168 37992
rect 20162 37952 20168 37964
rect 20220 37952 20226 38004
rect 23474 37992 23480 38004
rect 22066 37964 23480 37992
rect 3234 37924 3240 37936
rect 3195 37896 3240 37924
rect 3234 37884 3240 37896
rect 3292 37884 3298 37936
rect 4890 37884 4896 37936
rect 4948 37924 4954 37936
rect 8110 37924 8116 37936
rect 4948 37896 6914 37924
rect 8071 37896 8116 37924
rect 4948 37884 4954 37896
rect 1670 37856 1676 37868
rect 1631 37828 1676 37856
rect 1670 37816 1676 37828
rect 1728 37816 1734 37868
rect 2501 37859 2559 37865
rect 2501 37825 2513 37859
rect 2547 37856 2559 37859
rect 2958 37856 2964 37868
rect 2547 37828 2964 37856
rect 2547 37825 2559 37828
rect 2501 37819 2559 37825
rect 2958 37816 2964 37828
rect 3016 37816 3022 37868
rect 4798 37816 4804 37868
rect 4856 37856 4862 37868
rect 5445 37859 5503 37865
rect 5445 37856 5457 37859
rect 4856 37828 5457 37856
rect 4856 37816 4862 37828
rect 5445 37825 5457 37828
rect 5491 37856 5503 37859
rect 6362 37856 6368 37868
rect 5491 37828 6368 37856
rect 5491 37825 5503 37828
rect 5445 37819 5503 37825
rect 6362 37816 6368 37828
rect 6420 37816 6426 37868
rect 6886 37856 6914 37896
rect 8110 37884 8116 37896
rect 8168 37884 8174 37936
rect 8386 37884 8392 37936
rect 8444 37924 8450 37936
rect 8444 37896 9444 37924
rect 8444 37884 8450 37896
rect 7101 37859 7159 37865
rect 7101 37856 7113 37859
rect 6886 37828 7113 37856
rect 7101 37825 7113 37828
rect 7147 37856 7159 37859
rect 7147 37828 7880 37856
rect 7147 37825 7159 37828
rect 7101 37819 7159 37825
rect 3050 37788 3056 37800
rect 3011 37760 3056 37788
rect 3050 37748 3056 37760
rect 3108 37748 3114 37800
rect 3418 37748 3424 37800
rect 3476 37788 3482 37800
rect 3513 37791 3571 37797
rect 3513 37788 3525 37791
rect 3476 37760 3525 37788
rect 3476 37748 3482 37760
rect 3513 37757 3525 37760
rect 3559 37757 3571 37791
rect 3513 37751 3571 37757
rect 7852 37720 7880 37828
rect 7929 37791 7987 37797
rect 7929 37757 7941 37791
rect 7975 37788 7987 37791
rect 9306 37788 9312 37800
rect 7975 37760 9312 37788
rect 7975 37757 7987 37760
rect 7929 37751 7987 37757
rect 9306 37748 9312 37760
rect 9364 37748 9370 37800
rect 9416 37797 9444 37896
rect 18598 37884 18604 37936
rect 18656 37924 18662 37936
rect 22066 37924 22094 37964
rect 23474 37952 23480 37964
rect 23532 37952 23538 38004
rect 24486 37992 24492 38004
rect 24447 37964 24492 37992
rect 24486 37952 24492 37964
rect 24544 37952 24550 38004
rect 30282 37992 30288 38004
rect 24596 37964 30288 37992
rect 18656 37896 22094 37924
rect 18656 37884 18662 37896
rect 22186 37884 22192 37936
rect 22244 37924 22250 37936
rect 24596 37924 24624 37964
rect 30282 37952 30288 37964
rect 30340 37952 30346 38004
rect 25130 37924 25136 37936
rect 22244 37896 24624 37924
rect 25091 37896 25136 37924
rect 22244 37884 22250 37896
rect 25130 37884 25136 37896
rect 25188 37884 25194 37936
rect 25314 37884 25320 37936
rect 25372 37924 25378 37936
rect 30006 37924 30012 37936
rect 25372 37896 30012 37924
rect 25372 37884 25378 37896
rect 30006 37884 30012 37896
rect 30064 37884 30070 37936
rect 30098 37884 30104 37936
rect 30156 37924 30162 37936
rect 32677 37927 32735 37933
rect 32677 37924 32689 37927
rect 30156 37896 32689 37924
rect 30156 37884 30162 37896
rect 32677 37893 32689 37896
rect 32723 37893 32735 37927
rect 34330 37924 34336 37936
rect 34291 37896 34336 37924
rect 32677 37887 32735 37893
rect 34330 37884 34336 37896
rect 34388 37884 34394 37936
rect 15654 37856 15660 37868
rect 15615 37828 15660 37856
rect 15654 37816 15660 37828
rect 15712 37816 15718 37868
rect 16301 37859 16359 37865
rect 16301 37825 16313 37859
rect 16347 37856 16359 37859
rect 16390 37856 16396 37868
rect 16347 37828 16396 37856
rect 16347 37825 16359 37828
rect 16301 37819 16359 37825
rect 16390 37816 16396 37828
rect 16448 37816 16454 37868
rect 17126 37856 17132 37868
rect 17087 37828 17132 37856
rect 17126 37816 17132 37828
rect 17184 37816 17190 37868
rect 17678 37816 17684 37868
rect 17736 37856 17742 37868
rect 17773 37859 17831 37865
rect 17773 37856 17785 37859
rect 17736 37828 17785 37856
rect 17736 37816 17742 37828
rect 17773 37825 17785 37828
rect 17819 37825 17831 37859
rect 18966 37856 18972 37868
rect 18927 37828 18972 37856
rect 17773 37819 17831 37825
rect 18966 37816 18972 37828
rect 19024 37816 19030 37868
rect 20073 37859 20131 37865
rect 20073 37825 20085 37859
rect 20119 37856 20131 37859
rect 20438 37856 20444 37868
rect 20119 37828 20444 37856
rect 20119 37825 20131 37828
rect 20073 37819 20131 37825
rect 20438 37816 20444 37828
rect 20496 37816 20502 37868
rect 22457 37859 22515 37865
rect 22457 37856 22469 37859
rect 22296 37828 22469 37856
rect 9401 37791 9459 37797
rect 9401 37757 9413 37791
rect 9447 37757 9459 37791
rect 9401 37751 9459 37757
rect 18690 37748 18696 37800
rect 18748 37788 18754 37800
rect 22296 37788 22324 37828
rect 22457 37825 22469 37828
rect 22503 37856 22515 37859
rect 23109 37859 23167 37865
rect 22503 37828 23060 37856
rect 22503 37825 22515 37828
rect 22457 37819 22515 37825
rect 18748 37760 22324 37788
rect 23032 37788 23060 37828
rect 23109 37825 23121 37859
rect 23155 37856 23167 37859
rect 23474 37856 23480 37868
rect 23155 37828 23480 37856
rect 23155 37825 23167 37828
rect 23109 37819 23167 37825
rect 23474 37816 23480 37828
rect 23532 37816 23538 37868
rect 23753 37859 23811 37865
rect 23753 37825 23765 37859
rect 23799 37825 23811 37859
rect 24394 37856 24400 37868
rect 24355 37828 24400 37856
rect 23753 37819 23811 37825
rect 23768 37788 23796 37819
rect 24394 37816 24400 37828
rect 24452 37816 24458 37868
rect 25038 37856 25044 37868
rect 24999 37828 25044 37856
rect 25038 37816 25044 37828
rect 25096 37816 25102 37868
rect 26145 37859 26203 37865
rect 26145 37825 26157 37859
rect 26191 37825 26203 37859
rect 26145 37819 26203 37825
rect 25314 37788 25320 37800
rect 23032 37760 25320 37788
rect 18748 37748 18754 37760
rect 25314 37748 25320 37760
rect 25372 37748 25378 37800
rect 26160 37788 26188 37819
rect 27154 37816 27160 37868
rect 27212 37856 27218 37868
rect 27212 37828 27257 37856
rect 27212 37816 27218 37828
rect 27430 37816 27436 37868
rect 27488 37856 27494 37868
rect 28537 37859 28595 37865
rect 28537 37856 28549 37859
rect 27488 37828 28549 37856
rect 27488 37816 27494 37828
rect 28537 37825 28549 37828
rect 28583 37825 28595 37859
rect 31570 37856 31576 37868
rect 31531 37828 31576 37856
rect 28537 37819 28595 37825
rect 31570 37816 31576 37828
rect 31628 37816 31634 37868
rect 27522 37788 27528 37800
rect 26160 37760 27528 37788
rect 27522 37748 27528 37760
rect 27580 37748 27586 37800
rect 27614 37748 27620 37800
rect 27672 37788 27678 37800
rect 28721 37791 28779 37797
rect 28721 37788 28733 37791
rect 27672 37760 28733 37788
rect 27672 37748 27678 37760
rect 28721 37757 28733 37760
rect 28767 37757 28779 37791
rect 28994 37788 29000 37800
rect 28955 37760 29000 37788
rect 28721 37751 28779 37757
rect 28994 37748 29000 37760
rect 29052 37748 29058 37800
rect 29638 37748 29644 37800
rect 29696 37788 29702 37800
rect 30926 37788 30932 37800
rect 29696 37760 30932 37788
rect 29696 37748 29702 37760
rect 30926 37748 30932 37760
rect 30984 37748 30990 37800
rect 31386 37788 31392 37800
rect 31347 37760 31392 37788
rect 31386 37748 31392 37760
rect 31444 37748 31450 37800
rect 32490 37788 32496 37800
rect 31496 37760 32168 37788
rect 32451 37760 32496 37788
rect 16574 37720 16580 37732
rect 7852 37692 16580 37720
rect 16574 37680 16580 37692
rect 16632 37680 16638 37732
rect 19613 37723 19671 37729
rect 19613 37689 19625 37723
rect 19659 37720 19671 37723
rect 22186 37720 22192 37732
rect 19659 37692 22192 37720
rect 19659 37689 19671 37692
rect 19613 37683 19671 37689
rect 22186 37680 22192 37692
rect 22244 37680 22250 37732
rect 22557 37723 22615 37729
rect 22557 37689 22569 37723
rect 22603 37720 22615 37723
rect 22603 37692 24256 37720
rect 22603 37689 22615 37692
rect 22557 37683 22615 37689
rect 5718 37612 5724 37664
rect 5776 37652 5782 37664
rect 16022 37652 16028 37664
rect 5776 37624 16028 37652
rect 5776 37612 5782 37624
rect 16022 37612 16028 37624
rect 16080 37612 16086 37664
rect 16114 37612 16120 37664
rect 16172 37652 16178 37664
rect 16945 37655 17003 37661
rect 16172 37624 16217 37652
rect 16172 37612 16178 37624
rect 16945 37621 16957 37655
rect 16991 37652 17003 37655
rect 21174 37652 21180 37664
rect 16991 37624 21180 37652
rect 16991 37621 17003 37624
rect 16945 37615 17003 37621
rect 21174 37612 21180 37624
rect 21232 37612 21238 37664
rect 21450 37652 21456 37664
rect 21411 37624 21456 37652
rect 21450 37612 21456 37624
rect 21508 37612 21514 37664
rect 23201 37655 23259 37661
rect 23201 37621 23213 37655
rect 23247 37652 23259 37655
rect 23750 37652 23756 37664
rect 23247 37624 23756 37652
rect 23247 37621 23259 37624
rect 23201 37615 23259 37621
rect 23750 37612 23756 37624
rect 23808 37612 23814 37664
rect 23845 37655 23903 37661
rect 23845 37621 23857 37655
rect 23891 37652 23903 37655
rect 24118 37652 24124 37664
rect 23891 37624 24124 37652
rect 23891 37621 23903 37624
rect 23845 37615 23903 37621
rect 24118 37612 24124 37624
rect 24176 37612 24182 37664
rect 24228 37652 24256 37692
rect 24302 37680 24308 37732
rect 24360 37720 24366 37732
rect 27249 37723 27307 37729
rect 24360 37692 26096 37720
rect 24360 37680 24366 37692
rect 25774 37652 25780 37664
rect 24228 37624 25780 37652
rect 25774 37612 25780 37624
rect 25832 37612 25838 37664
rect 25958 37652 25964 37664
rect 25919 37624 25964 37652
rect 25958 37612 25964 37624
rect 26016 37612 26022 37664
rect 26068 37652 26096 37692
rect 27249 37689 27261 37723
rect 27295 37720 27307 37723
rect 27338 37720 27344 37732
rect 27295 37692 27344 37720
rect 27295 37689 27307 37692
rect 27249 37683 27307 37689
rect 27338 37680 27344 37692
rect 27396 37680 27402 37732
rect 27985 37723 28043 37729
rect 27985 37689 27997 37723
rect 28031 37720 28043 37723
rect 31496 37720 31524 37760
rect 28031 37692 31524 37720
rect 32140 37720 32168 37760
rect 32490 37748 32496 37760
rect 32548 37748 32554 37800
rect 32582 37720 32588 37732
rect 32140 37692 32588 37720
rect 28031 37689 28043 37692
rect 27985 37683 28043 37689
rect 32582 37680 32588 37692
rect 32640 37680 32646 37732
rect 31757 37655 31815 37661
rect 31757 37652 31769 37655
rect 26068 37624 31769 37652
rect 31757 37621 31769 37624
rect 31803 37621 31815 37655
rect 31757 37615 31815 37621
rect 1104 37562 34868 37584
rect 1104 37510 5170 37562
rect 5222 37510 5234 37562
rect 5286 37510 5298 37562
rect 5350 37510 5362 37562
rect 5414 37510 5426 37562
rect 5478 37510 13611 37562
rect 13663 37510 13675 37562
rect 13727 37510 13739 37562
rect 13791 37510 13803 37562
rect 13855 37510 13867 37562
rect 13919 37510 22052 37562
rect 22104 37510 22116 37562
rect 22168 37510 22180 37562
rect 22232 37510 22244 37562
rect 22296 37510 22308 37562
rect 22360 37510 30493 37562
rect 30545 37510 30557 37562
rect 30609 37510 30621 37562
rect 30673 37510 30685 37562
rect 30737 37510 30749 37562
rect 30801 37510 34868 37562
rect 1104 37488 34868 37510
rect 3050 37408 3056 37460
rect 3108 37448 3114 37460
rect 6273 37451 6331 37457
rect 6273 37448 6285 37451
rect 3108 37420 6285 37448
rect 3108 37408 3114 37420
rect 6273 37417 6285 37420
rect 6319 37417 6331 37451
rect 6273 37411 6331 37417
rect 6362 37408 6368 37460
rect 6420 37448 6426 37460
rect 6420 37420 12434 37448
rect 6420 37408 6426 37420
rect 3970 37340 3976 37392
rect 4028 37380 4034 37392
rect 8205 37383 8263 37389
rect 8205 37380 8217 37383
rect 4028 37352 8217 37380
rect 4028 37340 4034 37352
rect 8205 37349 8217 37352
rect 8251 37349 8263 37383
rect 12406 37380 12434 37420
rect 14274 37408 14280 37460
rect 14332 37448 14338 37460
rect 15286 37448 15292 37460
rect 14332 37420 15292 37448
rect 14332 37408 14338 37420
rect 15286 37408 15292 37420
rect 15344 37448 15350 37460
rect 20165 37451 20223 37457
rect 15344 37420 19380 37448
rect 15344 37408 15350 37420
rect 19242 37380 19248 37392
rect 12406 37352 19248 37380
rect 8205 37343 8263 37349
rect 19242 37340 19248 37352
rect 19300 37340 19306 37392
rect 2038 37312 2044 37324
rect 1999 37284 2044 37312
rect 2038 37272 2044 37284
rect 2096 37272 2102 37324
rect 3326 37272 3332 37324
rect 3384 37312 3390 37324
rect 18233 37315 18291 37321
rect 3384 37284 6868 37312
rect 3384 37272 3390 37284
rect 1581 37247 1639 37253
rect 1581 37213 1593 37247
rect 1627 37213 1639 37247
rect 1581 37207 1639 37213
rect 1596 37108 1624 37207
rect 2958 37204 2964 37256
rect 3016 37244 3022 37256
rect 3970 37244 3976 37256
rect 3016 37216 3976 37244
rect 3016 37204 3022 37216
rect 3970 37204 3976 37216
rect 4028 37204 4034 37256
rect 5534 37204 5540 37256
rect 5592 37244 5598 37256
rect 5629 37247 5687 37253
rect 5629 37244 5641 37247
rect 5592 37216 5641 37244
rect 5592 37204 5598 37216
rect 5629 37213 5641 37216
rect 5675 37213 5687 37247
rect 6730 37244 6736 37256
rect 5629 37207 5687 37213
rect 6656 37216 6736 37244
rect 1765 37179 1823 37185
rect 1765 37145 1777 37179
rect 1811 37176 1823 37179
rect 4062 37176 4068 37188
rect 1811 37148 4068 37176
rect 1811 37145 1823 37148
rect 1765 37139 1823 37145
rect 4062 37136 4068 37148
rect 4120 37136 4126 37188
rect 4614 37136 4620 37188
rect 4672 37176 4678 37188
rect 4801 37179 4859 37185
rect 4801 37176 4813 37179
rect 4672 37148 4813 37176
rect 4672 37136 4678 37148
rect 4801 37145 4813 37148
rect 4847 37176 4859 37179
rect 6656 37176 6684 37216
rect 6730 37204 6736 37216
rect 6788 37204 6794 37256
rect 6840 37244 6868 37284
rect 18233 37281 18245 37315
rect 18279 37312 18291 37315
rect 19150 37312 19156 37324
rect 18279 37284 19156 37312
rect 18279 37281 18291 37284
rect 18233 37275 18291 37281
rect 19150 37272 19156 37284
rect 19208 37272 19214 37324
rect 19352 37312 19380 37420
rect 20165 37417 20177 37451
rect 20211 37448 20223 37451
rect 20346 37448 20352 37460
rect 20211 37420 20352 37448
rect 20211 37417 20223 37420
rect 20165 37411 20223 37417
rect 20346 37408 20352 37420
rect 20404 37408 20410 37460
rect 21358 37448 21364 37460
rect 21319 37420 21364 37448
rect 21358 37408 21364 37420
rect 21416 37408 21422 37460
rect 24394 37448 24400 37460
rect 22066 37420 24400 37448
rect 19426 37340 19432 37392
rect 19484 37380 19490 37392
rect 22066 37380 22094 37420
rect 24394 37408 24400 37420
rect 24452 37408 24458 37460
rect 24854 37408 24860 37460
rect 24912 37448 24918 37460
rect 25682 37448 25688 37460
rect 24912 37420 25688 37448
rect 24912 37408 24918 37420
rect 25682 37408 25688 37420
rect 25740 37408 25746 37460
rect 25774 37408 25780 37460
rect 25832 37448 25838 37460
rect 30098 37448 30104 37460
rect 25832 37420 30104 37448
rect 25832 37408 25838 37420
rect 30098 37408 30104 37420
rect 30156 37408 30162 37460
rect 30285 37451 30343 37457
rect 30285 37417 30297 37451
rect 30331 37448 30343 37451
rect 34054 37448 34060 37460
rect 30331 37420 34060 37448
rect 30331 37417 30343 37420
rect 30285 37411 30343 37417
rect 34054 37408 34060 37420
rect 34112 37408 34118 37460
rect 32490 37380 32496 37392
rect 19484 37352 22094 37380
rect 23492 37352 32496 37380
rect 19484 37340 19490 37352
rect 19352 37284 20760 37312
rect 6917 37247 6975 37253
rect 6917 37244 6929 37247
rect 6840 37216 6929 37244
rect 6917 37213 6929 37216
rect 6963 37213 6975 37247
rect 7374 37244 7380 37256
rect 7335 37216 7380 37244
rect 6917 37207 6975 37213
rect 7374 37204 7380 37216
rect 7432 37204 7438 37256
rect 7466 37204 7472 37256
rect 7524 37244 7530 37256
rect 17402 37244 17408 37256
rect 7524 37216 7569 37244
rect 17363 37216 17408 37244
rect 7524 37204 7530 37216
rect 17402 37204 17408 37216
rect 17460 37244 17466 37256
rect 18598 37244 18604 37256
rect 17460 37216 18604 37244
rect 17460 37204 17466 37216
rect 18598 37204 18604 37216
rect 18656 37204 18662 37256
rect 18874 37244 18880 37256
rect 18835 37216 18880 37244
rect 18874 37204 18880 37216
rect 18932 37204 18938 37256
rect 20438 37204 20444 37256
rect 20496 37244 20502 37256
rect 20625 37247 20683 37253
rect 20625 37244 20637 37247
rect 20496 37216 20637 37244
rect 20496 37204 20502 37216
rect 20625 37213 20637 37216
rect 20671 37213 20683 37247
rect 20732 37244 20760 37284
rect 21450 37272 21456 37324
rect 21508 37312 21514 37324
rect 23492 37312 23520 37352
rect 32490 37340 32496 37352
rect 32548 37340 32554 37392
rect 29914 37312 29920 37324
rect 21508 37284 23520 37312
rect 23584 37284 29920 37312
rect 21508 37272 21514 37284
rect 21269 37247 21327 37253
rect 21269 37244 21281 37247
rect 20732 37216 21281 37244
rect 20625 37207 20683 37213
rect 21269 37213 21281 37216
rect 21315 37244 21327 37247
rect 21910 37244 21916 37256
rect 21315 37216 21916 37244
rect 21315 37213 21327 37216
rect 21269 37207 21327 37213
rect 21910 37204 21916 37216
rect 21968 37204 21974 37256
rect 22097 37247 22155 37253
rect 22097 37213 22109 37247
rect 22143 37244 22155 37247
rect 22462 37244 22468 37256
rect 22143 37216 22468 37244
rect 22143 37213 22155 37216
rect 22097 37207 22155 37213
rect 22462 37204 22468 37216
rect 22520 37204 22526 37256
rect 22557 37247 22615 37253
rect 22557 37213 22569 37247
rect 22603 37244 22615 37247
rect 22738 37244 22744 37256
rect 22603 37216 22744 37244
rect 22603 37213 22615 37216
rect 22557 37207 22615 37213
rect 22738 37204 22744 37216
rect 22796 37204 22802 37256
rect 23385 37247 23443 37253
rect 23385 37213 23397 37247
rect 23431 37244 23443 37247
rect 23584 37244 23612 37284
rect 29914 37272 29920 37284
rect 29972 37272 29978 37324
rect 30377 37315 30435 37321
rect 30377 37281 30389 37315
rect 30423 37312 30435 37315
rect 30742 37312 30748 37324
rect 30423 37284 30748 37312
rect 30423 37281 30435 37284
rect 30377 37275 30435 37281
rect 30742 37272 30748 37284
rect 30800 37272 30806 37324
rect 31478 37272 31484 37324
rect 31536 37312 31542 37324
rect 31665 37315 31723 37321
rect 31665 37312 31677 37315
rect 31536 37284 31677 37312
rect 31536 37272 31542 37284
rect 31665 37281 31677 37284
rect 31711 37281 31723 37315
rect 33042 37312 33048 37324
rect 33003 37284 33048 37312
rect 31665 37275 31723 37281
rect 33042 37272 33048 37284
rect 33100 37272 33106 37324
rect 24026 37244 24032 37256
rect 23431 37216 23612 37244
rect 23987 37216 24032 37244
rect 23431 37213 23443 37216
rect 23385 37207 23443 37213
rect 24026 37204 24032 37216
rect 24084 37204 24090 37256
rect 24670 37244 24676 37256
rect 24631 37216 24676 37244
rect 24670 37204 24676 37216
rect 24728 37204 24734 37256
rect 25314 37244 25320 37256
rect 25275 37216 25320 37244
rect 25314 37204 25320 37216
rect 25372 37204 25378 37256
rect 26050 37204 26056 37256
rect 26108 37244 26114 37256
rect 26513 37247 26571 37253
rect 26513 37244 26525 37247
rect 26108 37216 26525 37244
rect 26108 37204 26114 37216
rect 26513 37213 26525 37216
rect 26559 37213 26571 37247
rect 26513 37207 26571 37213
rect 26970 37204 26976 37256
rect 27028 37244 27034 37256
rect 27065 37247 27123 37253
rect 27065 37244 27077 37247
rect 27028 37216 27077 37244
rect 27028 37204 27034 37216
rect 27065 37213 27077 37216
rect 27111 37213 27123 37247
rect 28166 37244 28172 37256
rect 28127 37216 28172 37244
rect 27065 37207 27123 37213
rect 28166 37204 28172 37216
rect 28224 37204 28230 37256
rect 29178 37244 29184 37256
rect 29139 37216 29184 37244
rect 29178 37204 29184 37216
rect 29236 37204 29242 37256
rect 30098 37244 30104 37256
rect 30059 37216 30104 37244
rect 30098 37204 30104 37216
rect 30156 37204 30162 37256
rect 30193 37247 30251 37253
rect 30193 37213 30205 37247
rect 30239 37244 30251 37247
rect 30282 37244 30288 37256
rect 30239 37216 30288 37244
rect 30239 37213 30251 37216
rect 30193 37207 30251 37213
rect 30282 37204 30288 37216
rect 30340 37204 30346 37256
rect 30929 37247 30987 37253
rect 30929 37213 30941 37247
rect 30975 37213 30987 37247
rect 30929 37207 30987 37213
rect 31021 37247 31079 37253
rect 31021 37213 31033 37247
rect 31067 37244 31079 37247
rect 31570 37244 31576 37256
rect 31067 37216 31576 37244
rect 31067 37213 31079 37216
rect 31021 37207 31079 37213
rect 22649 37179 22707 37185
rect 4847 37148 6684 37176
rect 6748 37148 22094 37176
rect 4847 37145 4859 37148
rect 4801 37139 4859 37145
rect 4154 37108 4160 37120
rect 1596 37080 4160 37108
rect 4154 37068 4160 37080
rect 4212 37068 4218 37120
rect 6748 37117 6776 37148
rect 6733 37111 6791 37117
rect 6733 37077 6745 37111
rect 6779 37077 6791 37111
rect 6733 37071 6791 37077
rect 6822 37068 6828 37120
rect 6880 37108 6886 37120
rect 14274 37108 14280 37120
rect 6880 37080 14280 37108
rect 6880 37068 6886 37080
rect 14274 37068 14280 37080
rect 14332 37068 14338 37120
rect 17494 37108 17500 37120
rect 17455 37080 17500 37108
rect 17494 37068 17500 37080
rect 17552 37068 17558 37120
rect 18693 37111 18751 37117
rect 18693 37077 18705 37111
rect 18739 37108 18751 37111
rect 19058 37108 19064 37120
rect 18739 37080 19064 37108
rect 18739 37077 18751 37080
rect 18693 37071 18751 37077
rect 19058 37068 19064 37080
rect 19116 37068 19122 37120
rect 20714 37108 20720 37120
rect 20675 37080 20720 37108
rect 20714 37068 20720 37080
rect 20772 37068 20778 37120
rect 22066 37108 22094 37148
rect 22649 37145 22661 37179
rect 22695 37176 22707 37179
rect 30006 37176 30012 37188
rect 22695 37148 30012 37176
rect 22695 37145 22707 37148
rect 22649 37139 22707 37145
rect 30006 37136 30012 37148
rect 30064 37136 30070 37188
rect 30944 37176 30972 37207
rect 31570 37204 31576 37216
rect 31628 37244 31634 37256
rect 31849 37247 31907 37253
rect 31849 37244 31861 37247
rect 31628 37216 31861 37244
rect 31628 37204 31634 37216
rect 31849 37213 31861 37216
rect 31895 37213 31907 37247
rect 32490 37244 32496 37256
rect 32451 37216 32496 37244
rect 31849 37207 31907 37213
rect 32490 37204 32496 37216
rect 32548 37204 32554 37256
rect 31110 37176 31116 37188
rect 30944 37148 31116 37176
rect 31110 37136 31116 37148
rect 31168 37136 31174 37188
rect 32674 37176 32680 37188
rect 32635 37148 32680 37176
rect 32674 37136 32680 37148
rect 32732 37136 32738 37188
rect 23566 37108 23572 37120
rect 22066 37080 23572 37108
rect 23566 37068 23572 37080
rect 23624 37068 23630 37120
rect 24762 37108 24768 37120
rect 24723 37080 24768 37108
rect 24762 37068 24768 37080
rect 24820 37068 24826 37120
rect 25406 37108 25412 37120
rect 25367 37080 25412 37108
rect 25406 37068 25412 37080
rect 25464 37068 25470 37120
rect 26329 37111 26387 37117
rect 26329 37077 26341 37111
rect 26375 37108 26387 37111
rect 26970 37108 26976 37120
rect 26375 37080 26976 37108
rect 26375 37077 26387 37080
rect 26329 37071 26387 37077
rect 26970 37068 26976 37080
rect 27028 37068 27034 37120
rect 27154 37108 27160 37120
rect 27115 37080 27160 37108
rect 27154 37068 27160 37080
rect 27212 37068 27218 37120
rect 27982 37108 27988 37120
rect 27943 37080 27988 37108
rect 27982 37068 27988 37080
rect 28040 37068 28046 37120
rect 28997 37111 29055 37117
rect 28997 37077 29009 37111
rect 29043 37108 29055 37111
rect 29362 37108 29368 37120
rect 29043 37080 29368 37108
rect 29043 37077 29055 37080
rect 28997 37071 29055 37077
rect 29362 37068 29368 37080
rect 29420 37068 29426 37120
rect 29730 37068 29736 37120
rect 29788 37108 29794 37120
rect 30558 37108 30564 37120
rect 29788 37080 30564 37108
rect 29788 37068 29794 37080
rect 30558 37068 30564 37080
rect 30616 37068 30622 37120
rect 30926 37068 30932 37120
rect 30984 37108 30990 37120
rect 31205 37111 31263 37117
rect 31205 37108 31217 37111
rect 30984 37080 31217 37108
rect 30984 37068 30990 37080
rect 31205 37077 31217 37080
rect 31251 37077 31263 37111
rect 32030 37108 32036 37120
rect 31991 37080 32036 37108
rect 31205 37071 31263 37077
rect 32030 37068 32036 37080
rect 32088 37068 32094 37120
rect 1104 37018 35027 37040
rect 1104 36966 9390 37018
rect 9442 36966 9454 37018
rect 9506 36966 9518 37018
rect 9570 36966 9582 37018
rect 9634 36966 9646 37018
rect 9698 36966 17831 37018
rect 17883 36966 17895 37018
rect 17947 36966 17959 37018
rect 18011 36966 18023 37018
rect 18075 36966 18087 37018
rect 18139 36966 26272 37018
rect 26324 36966 26336 37018
rect 26388 36966 26400 37018
rect 26452 36966 26464 37018
rect 26516 36966 26528 37018
rect 26580 36966 34713 37018
rect 34765 36966 34777 37018
rect 34829 36966 34841 37018
rect 34893 36966 34905 37018
rect 34957 36966 34969 37018
rect 35021 36966 35027 37018
rect 1104 36944 35027 36966
rect 5534 36904 5540 36916
rect 1780 36876 5540 36904
rect 1780 36777 1808 36876
rect 5534 36864 5540 36876
rect 5592 36864 5598 36916
rect 7282 36904 7288 36916
rect 7243 36876 7288 36904
rect 7282 36864 7288 36876
rect 7340 36864 7346 36916
rect 20714 36864 20720 36916
rect 20772 36904 20778 36916
rect 32674 36904 32680 36916
rect 20772 36876 32680 36904
rect 20772 36864 20778 36876
rect 32674 36864 32680 36876
rect 32732 36864 32738 36916
rect 1949 36839 2007 36845
rect 1949 36805 1961 36839
rect 1995 36836 2007 36839
rect 5629 36839 5687 36845
rect 5629 36836 5641 36839
rect 1995 36808 5641 36836
rect 1995 36805 2007 36808
rect 1949 36799 2007 36805
rect 5629 36805 5641 36808
rect 5675 36805 5687 36839
rect 27614 36836 27620 36848
rect 5629 36799 5687 36805
rect 20916 36808 27620 36836
rect 1765 36771 1823 36777
rect 1765 36737 1777 36771
rect 1811 36737 1823 36771
rect 1765 36731 1823 36737
rect 3970 36728 3976 36780
rect 4028 36768 4034 36780
rect 4065 36771 4123 36777
rect 4065 36768 4077 36771
rect 4028 36740 4077 36768
rect 4028 36728 4034 36740
rect 4065 36737 4077 36740
rect 4111 36737 4123 36771
rect 5534 36768 5540 36780
rect 5447 36740 5540 36768
rect 4065 36731 4123 36737
rect 5534 36728 5540 36740
rect 5592 36768 5598 36780
rect 5718 36768 5724 36780
rect 5592 36740 5724 36768
rect 5592 36728 5598 36740
rect 5718 36728 5724 36740
rect 5776 36728 5782 36780
rect 6546 36768 6552 36780
rect 6507 36740 6552 36768
rect 6546 36728 6552 36740
rect 6604 36728 6610 36780
rect 7193 36771 7251 36777
rect 7193 36737 7205 36771
rect 7239 36768 7251 36771
rect 7374 36768 7380 36780
rect 7239 36740 7380 36768
rect 7239 36737 7251 36740
rect 7193 36731 7251 36737
rect 7374 36728 7380 36740
rect 7432 36768 7438 36780
rect 17310 36768 17316 36780
rect 7432 36740 17316 36768
rect 7432 36728 7438 36740
rect 17310 36728 17316 36740
rect 17368 36728 17374 36780
rect 17586 36768 17592 36780
rect 17547 36740 17592 36768
rect 17586 36728 17592 36740
rect 17644 36728 17650 36780
rect 18230 36768 18236 36780
rect 18191 36740 18236 36768
rect 18230 36728 18236 36740
rect 18288 36728 18294 36780
rect 18690 36768 18696 36780
rect 18651 36740 18696 36768
rect 18690 36728 18696 36740
rect 18748 36728 18754 36780
rect 19334 36768 19340 36780
rect 19295 36740 19340 36768
rect 19334 36728 19340 36740
rect 19392 36728 19398 36780
rect 20165 36771 20223 36777
rect 20165 36737 20177 36771
rect 20211 36768 20223 36771
rect 20530 36768 20536 36780
rect 20211 36740 20536 36768
rect 20211 36737 20223 36740
rect 20165 36731 20223 36737
rect 20530 36728 20536 36740
rect 20588 36728 20594 36780
rect 2774 36700 2780 36712
rect 2735 36672 2780 36700
rect 2774 36660 2780 36672
rect 2832 36660 2838 36712
rect 4430 36700 4436 36712
rect 4391 36672 4436 36700
rect 4430 36660 4436 36672
rect 4488 36700 4494 36712
rect 4982 36700 4988 36712
rect 4488 36672 4988 36700
rect 4488 36660 4494 36672
rect 4982 36660 4988 36672
rect 5040 36660 5046 36712
rect 5074 36660 5080 36712
rect 5132 36700 5138 36712
rect 6641 36703 6699 36709
rect 6641 36700 6653 36703
rect 5132 36672 6653 36700
rect 5132 36660 5138 36672
rect 6641 36669 6653 36672
rect 6687 36669 6699 36703
rect 20438 36700 20444 36712
rect 6641 36663 6699 36669
rect 6886 36672 20444 36700
rect 5000 36632 5028 36660
rect 6886 36632 6914 36672
rect 20438 36660 20444 36672
rect 20496 36660 20502 36712
rect 20622 36700 20628 36712
rect 20583 36672 20628 36700
rect 20622 36660 20628 36672
rect 20680 36660 20686 36712
rect 5000 36604 6914 36632
rect 18785 36635 18843 36641
rect 18785 36601 18797 36635
rect 18831 36632 18843 36635
rect 20916 36632 20944 36808
rect 27614 36796 27620 36808
rect 27672 36796 27678 36848
rect 30006 36836 30012 36848
rect 28644 36808 30012 36836
rect 21453 36771 21511 36777
rect 21453 36737 21465 36771
rect 21499 36737 21511 36771
rect 22370 36768 22376 36780
rect 22331 36740 22376 36768
rect 21453 36731 21511 36737
rect 20993 36703 21051 36709
rect 20993 36669 21005 36703
rect 21039 36700 21051 36703
rect 21468 36700 21496 36731
rect 22370 36728 22376 36740
rect 22428 36728 22434 36780
rect 22922 36728 22928 36780
rect 22980 36768 22986 36780
rect 23845 36771 23903 36777
rect 23845 36768 23857 36771
rect 22980 36740 23857 36768
rect 22980 36728 22986 36740
rect 23845 36737 23857 36740
rect 23891 36737 23903 36771
rect 24486 36768 24492 36780
rect 24447 36740 24492 36768
rect 23845 36731 23903 36737
rect 24486 36728 24492 36740
rect 24544 36728 24550 36780
rect 25130 36768 25136 36780
rect 25091 36740 25136 36768
rect 25130 36728 25136 36740
rect 25188 36728 25194 36780
rect 25866 36768 25872 36780
rect 25827 36740 25872 36768
rect 25866 36728 25872 36740
rect 25924 36728 25930 36780
rect 26418 36768 26424 36780
rect 26379 36740 26424 36768
rect 26418 36728 26424 36740
rect 26476 36728 26482 36780
rect 26510 36728 26516 36780
rect 26568 36768 26574 36780
rect 27341 36771 27399 36777
rect 27341 36768 27353 36771
rect 26568 36740 27353 36768
rect 26568 36728 26574 36740
rect 27341 36737 27353 36740
rect 27387 36737 27399 36771
rect 27341 36731 27399 36737
rect 27985 36771 28043 36777
rect 27985 36737 27997 36771
rect 28031 36768 28043 36771
rect 28534 36768 28540 36780
rect 28031 36740 28540 36768
rect 28031 36737 28043 36740
rect 27985 36731 28043 36737
rect 28534 36728 28540 36740
rect 28592 36728 28598 36780
rect 28644 36777 28672 36808
rect 30006 36796 30012 36808
rect 30064 36796 30070 36848
rect 30558 36796 30564 36848
rect 30616 36836 30622 36848
rect 30616 36808 31156 36836
rect 30616 36796 30622 36808
rect 28629 36771 28687 36777
rect 28629 36737 28641 36771
rect 28675 36737 28687 36771
rect 29086 36768 29092 36780
rect 29047 36740 29092 36768
rect 28629 36731 28687 36737
rect 29086 36728 29092 36740
rect 29144 36728 29150 36780
rect 29273 36771 29331 36777
rect 29273 36737 29285 36771
rect 29319 36768 29331 36771
rect 29454 36768 29460 36780
rect 29319 36740 29460 36768
rect 29319 36737 29331 36740
rect 29273 36731 29331 36737
rect 29454 36728 29460 36740
rect 29512 36728 29518 36780
rect 29546 36728 29552 36780
rect 29604 36768 29610 36780
rect 30101 36771 30159 36777
rect 30101 36768 30113 36771
rect 29604 36740 30113 36768
rect 29604 36728 29610 36740
rect 30101 36737 30113 36740
rect 30147 36737 30159 36771
rect 31021 36771 31079 36777
rect 31021 36768 31033 36771
rect 30101 36731 30159 36737
rect 30208 36740 31033 36768
rect 25314 36700 25320 36712
rect 21039 36672 25320 36700
rect 21039 36669 21051 36672
rect 20993 36663 21051 36669
rect 25314 36660 25320 36672
rect 25372 36660 25378 36712
rect 30208 36700 30236 36740
rect 31021 36737 31033 36740
rect 31067 36737 31079 36771
rect 31128 36768 31156 36808
rect 31202 36796 31208 36848
rect 31260 36836 31266 36848
rect 31260 36808 31305 36836
rect 31260 36796 31266 36808
rect 32493 36771 32551 36777
rect 32493 36768 32505 36771
rect 31128 36740 32505 36768
rect 31021 36731 31079 36737
rect 32493 36737 32505 36740
rect 32539 36737 32551 36771
rect 32493 36731 32551 36737
rect 30834 36700 30840 36712
rect 26528 36672 30236 36700
rect 30795 36672 30840 36700
rect 18831 36604 20944 36632
rect 21269 36635 21327 36641
rect 18831 36601 18843 36604
rect 18785 36595 18843 36601
rect 21269 36601 21281 36635
rect 21315 36632 21327 36635
rect 26528 36632 26556 36672
rect 30834 36660 30840 36672
rect 30892 36660 30898 36712
rect 31938 36660 31944 36712
rect 31996 36700 32002 36712
rect 32677 36703 32735 36709
rect 32677 36700 32689 36703
rect 31996 36672 32689 36700
rect 31996 36660 32002 36672
rect 32677 36669 32689 36672
rect 32723 36669 32735 36703
rect 33502 36700 33508 36712
rect 33463 36672 33508 36700
rect 32677 36663 32735 36669
rect 33502 36660 33508 36672
rect 33560 36660 33566 36712
rect 21315 36604 26556 36632
rect 26605 36635 26663 36641
rect 21315 36601 21327 36604
rect 21269 36595 21327 36601
rect 26605 36601 26617 36635
rect 26651 36632 26663 36635
rect 27890 36632 27896 36644
rect 26651 36604 27896 36632
rect 26651 36601 26663 36604
rect 26605 36595 26663 36601
rect 27890 36592 27896 36604
rect 27948 36592 27954 36644
rect 29181 36635 29239 36641
rect 29181 36601 29193 36635
rect 29227 36632 29239 36635
rect 30926 36632 30932 36644
rect 29227 36604 30932 36632
rect 29227 36601 29239 36604
rect 29181 36595 29239 36601
rect 30926 36592 30932 36604
rect 30984 36592 30990 36644
rect 17405 36567 17463 36573
rect 17405 36533 17417 36567
rect 17451 36564 17463 36567
rect 17678 36564 17684 36576
rect 17451 36536 17684 36564
rect 17451 36533 17463 36536
rect 17405 36527 17463 36533
rect 17678 36524 17684 36536
rect 17736 36524 17742 36576
rect 18049 36567 18107 36573
rect 18049 36533 18061 36567
rect 18095 36564 18107 36567
rect 18966 36564 18972 36576
rect 18095 36536 18972 36564
rect 18095 36533 18107 36536
rect 18049 36527 18107 36533
rect 18966 36524 18972 36536
rect 19024 36524 19030 36576
rect 19429 36567 19487 36573
rect 19429 36533 19441 36567
rect 19475 36564 19487 36567
rect 20530 36564 20536 36576
rect 19475 36536 20536 36564
rect 19475 36533 19487 36536
rect 19429 36527 19487 36533
rect 20530 36524 20536 36536
rect 20588 36524 20594 36576
rect 22189 36567 22247 36573
rect 22189 36533 22201 36567
rect 22235 36564 22247 36567
rect 22554 36564 22560 36576
rect 22235 36536 22560 36564
rect 22235 36533 22247 36536
rect 22189 36527 22247 36533
rect 22554 36524 22560 36536
rect 22612 36524 22618 36576
rect 23201 36567 23259 36573
rect 23201 36533 23213 36567
rect 23247 36564 23259 36567
rect 23382 36564 23388 36576
rect 23247 36536 23388 36564
rect 23247 36533 23259 36536
rect 23201 36527 23259 36533
rect 23382 36524 23388 36536
rect 23440 36524 23446 36576
rect 23658 36564 23664 36576
rect 23619 36536 23664 36564
rect 23658 36524 23664 36536
rect 23716 36524 23722 36576
rect 24302 36564 24308 36576
rect 24263 36536 24308 36564
rect 24302 36524 24308 36536
rect 24360 36524 24366 36576
rect 24854 36524 24860 36576
rect 24912 36564 24918 36576
rect 24949 36567 25007 36573
rect 24949 36564 24961 36567
rect 24912 36536 24961 36564
rect 24912 36524 24918 36536
rect 24949 36533 24961 36536
rect 24995 36533 25007 36567
rect 25682 36564 25688 36576
rect 25643 36536 25688 36564
rect 24949 36527 25007 36533
rect 25682 36524 25688 36536
rect 25740 36524 25746 36576
rect 26142 36524 26148 36576
rect 26200 36564 26206 36576
rect 26510 36564 26516 36576
rect 26200 36536 26516 36564
rect 26200 36524 26206 36536
rect 26510 36524 26516 36536
rect 26568 36524 26574 36576
rect 27154 36564 27160 36576
rect 27115 36536 27160 36564
rect 27154 36524 27160 36536
rect 27212 36524 27218 36576
rect 27246 36524 27252 36576
rect 27304 36564 27310 36576
rect 27801 36567 27859 36573
rect 27801 36564 27813 36567
rect 27304 36536 27813 36564
rect 27304 36524 27310 36536
rect 27801 36533 27813 36536
rect 27847 36533 27859 36567
rect 28442 36564 28448 36576
rect 28403 36536 28448 36564
rect 27801 36527 27859 36533
rect 28442 36524 28448 36536
rect 28500 36524 28506 36576
rect 28534 36524 28540 36576
rect 28592 36564 28598 36576
rect 29270 36564 29276 36576
rect 28592 36536 29276 36564
rect 28592 36524 28598 36536
rect 29270 36524 29276 36536
rect 29328 36524 29334 36576
rect 29914 36524 29920 36576
rect 29972 36564 29978 36576
rect 30101 36567 30159 36573
rect 30101 36564 30113 36567
rect 29972 36536 30113 36564
rect 29972 36524 29978 36536
rect 30101 36533 30113 36536
rect 30147 36533 30159 36567
rect 30101 36527 30159 36533
rect 30282 36524 30288 36576
rect 30340 36564 30346 36576
rect 32950 36564 32956 36576
rect 30340 36536 32956 36564
rect 30340 36524 30346 36536
rect 32950 36524 32956 36536
rect 33008 36524 33014 36576
rect 1104 36474 34868 36496
rect 1104 36422 5170 36474
rect 5222 36422 5234 36474
rect 5286 36422 5298 36474
rect 5350 36422 5362 36474
rect 5414 36422 5426 36474
rect 5478 36422 13611 36474
rect 13663 36422 13675 36474
rect 13727 36422 13739 36474
rect 13791 36422 13803 36474
rect 13855 36422 13867 36474
rect 13919 36422 22052 36474
rect 22104 36422 22116 36474
rect 22168 36422 22180 36474
rect 22232 36422 22244 36474
rect 22296 36422 22308 36474
rect 22360 36422 30493 36474
rect 30545 36422 30557 36474
rect 30609 36422 30621 36474
rect 30673 36422 30685 36474
rect 30737 36422 30749 36474
rect 30801 36422 34868 36474
rect 1104 36400 34868 36422
rect 22738 36360 22744 36372
rect 19352 36332 22744 36360
rect 19352 36304 19380 36332
rect 22738 36320 22744 36332
rect 22796 36320 22802 36372
rect 22922 36360 22928 36372
rect 22883 36332 22928 36360
rect 22922 36320 22928 36332
rect 22980 36320 22986 36372
rect 26050 36360 26056 36372
rect 26011 36332 26056 36360
rect 26050 36320 26056 36332
rect 26108 36320 26114 36372
rect 26697 36363 26755 36369
rect 26697 36329 26709 36363
rect 26743 36360 26755 36363
rect 27062 36360 27068 36372
rect 26743 36332 27068 36360
rect 26743 36329 26755 36332
rect 26697 36323 26755 36329
rect 27062 36320 27068 36332
rect 27120 36320 27126 36372
rect 27522 36320 27528 36372
rect 27580 36360 27586 36372
rect 27709 36363 27767 36369
rect 27709 36360 27721 36363
rect 27580 36332 27721 36360
rect 27580 36320 27586 36332
rect 27709 36329 27721 36332
rect 27755 36329 27767 36363
rect 30190 36360 30196 36372
rect 30151 36332 30196 36360
rect 27709 36323 27767 36329
rect 30190 36320 30196 36332
rect 30248 36320 30254 36372
rect 31018 36360 31024 36372
rect 30979 36332 31024 36360
rect 31018 36320 31024 36332
rect 31076 36320 31082 36372
rect 31754 36320 31760 36372
rect 31812 36360 31818 36372
rect 31849 36363 31907 36369
rect 31849 36360 31861 36363
rect 31812 36332 31861 36360
rect 31812 36320 31818 36332
rect 31849 36329 31861 36332
rect 31895 36329 31907 36363
rect 31849 36323 31907 36329
rect 32214 36320 32220 36372
rect 32272 36360 32278 36372
rect 32272 36332 32720 36360
rect 32272 36320 32278 36332
rect 19334 36292 19340 36304
rect 3252 36264 19340 36292
rect 3252 36236 3280 36264
rect 19334 36252 19340 36264
rect 19392 36252 19398 36304
rect 25222 36292 25228 36304
rect 19996 36264 25228 36292
rect 3234 36224 3240 36236
rect 3147 36196 3240 36224
rect 3234 36184 3240 36196
rect 3292 36184 3298 36236
rect 4798 36224 4804 36236
rect 3804 36196 4804 36224
rect 1762 36116 1768 36168
rect 1820 36156 1826 36168
rect 1949 36159 2007 36165
rect 1949 36156 1961 36159
rect 1820 36128 1961 36156
rect 1820 36116 1826 36128
rect 1949 36125 1961 36128
rect 1995 36125 2007 36159
rect 1949 36119 2007 36125
rect 2038 36116 2044 36168
rect 2096 36156 2102 36168
rect 2409 36159 2467 36165
rect 2409 36156 2421 36159
rect 2096 36128 2421 36156
rect 2096 36116 2102 36128
rect 2409 36125 2421 36128
rect 2455 36156 2467 36159
rect 3804 36156 3832 36196
rect 4798 36184 4804 36196
rect 4856 36184 4862 36236
rect 3970 36156 3976 36168
rect 2455 36128 3832 36156
rect 3931 36128 3976 36156
rect 2455 36125 2467 36128
rect 2409 36119 2467 36125
rect 3970 36116 3976 36128
rect 4028 36156 4034 36168
rect 5445 36159 5503 36165
rect 5445 36156 5457 36159
rect 4028 36128 5457 36156
rect 4028 36116 4034 36128
rect 5445 36125 5457 36128
rect 5491 36125 5503 36159
rect 9122 36156 9128 36168
rect 5445 36119 5503 36125
rect 5552 36128 9128 36156
rect 4798 36088 4804 36100
rect 4759 36060 4804 36088
rect 4798 36048 4804 36060
rect 4856 36088 4862 36100
rect 5552 36088 5580 36128
rect 9122 36116 9128 36128
rect 9180 36116 9186 36168
rect 18414 36156 18420 36168
rect 18375 36128 18420 36156
rect 18414 36116 18420 36128
rect 18472 36116 18478 36168
rect 19794 36156 19800 36168
rect 19755 36128 19800 36156
rect 19794 36116 19800 36128
rect 19852 36116 19858 36168
rect 19996 36165 20024 36264
rect 25222 36252 25228 36264
rect 25280 36252 25286 36304
rect 25314 36252 25320 36304
rect 25372 36292 25378 36304
rect 28718 36292 28724 36304
rect 25372 36264 28724 36292
rect 25372 36252 25378 36264
rect 28718 36252 28724 36264
rect 28776 36252 28782 36304
rect 28997 36295 29055 36301
rect 28997 36261 29009 36295
rect 29043 36292 29055 36295
rect 30282 36292 30288 36304
rect 29043 36264 30288 36292
rect 29043 36261 29055 36264
rect 28997 36255 29055 36261
rect 30282 36252 30288 36264
rect 30340 36252 30346 36304
rect 30834 36292 30840 36304
rect 30576 36264 30840 36292
rect 26602 36224 26608 36236
rect 23032 36196 26608 36224
rect 19981 36159 20039 36165
rect 19981 36125 19993 36159
rect 20027 36125 20039 36159
rect 20622 36156 20628 36168
rect 20583 36128 20628 36156
rect 19981 36119 20039 36125
rect 20622 36116 20628 36128
rect 20680 36116 20686 36168
rect 21266 36156 21272 36168
rect 21227 36128 21272 36156
rect 21266 36116 21272 36128
rect 21324 36116 21330 36168
rect 21910 36156 21916 36168
rect 21871 36128 21916 36156
rect 21910 36116 21916 36128
rect 21968 36116 21974 36168
rect 22646 36156 22652 36168
rect 22607 36128 22652 36156
rect 22646 36116 22652 36128
rect 22704 36116 22710 36168
rect 22738 36116 22744 36168
rect 22796 36156 22802 36168
rect 23032 36156 23060 36196
rect 22796 36128 23060 36156
rect 22796 36116 22802 36128
rect 23290 36116 23296 36168
rect 23348 36156 23354 36168
rect 23385 36159 23443 36165
rect 23385 36156 23397 36159
rect 23348 36128 23397 36156
rect 23348 36116 23354 36128
rect 23385 36125 23397 36128
rect 23431 36125 23443 36159
rect 23566 36156 23572 36168
rect 23527 36128 23572 36156
rect 23385 36119 23443 36125
rect 23566 36116 23572 36128
rect 23624 36116 23630 36168
rect 23753 36159 23811 36165
rect 23753 36125 23765 36159
rect 23799 36156 23811 36159
rect 24765 36159 24823 36165
rect 24765 36156 24777 36159
rect 23799 36128 24777 36156
rect 23799 36125 23811 36128
rect 23753 36119 23811 36125
rect 24765 36125 24777 36128
rect 24811 36125 24823 36159
rect 25774 36156 25780 36168
rect 25735 36128 25780 36156
rect 24765 36119 24823 36125
rect 25774 36116 25780 36128
rect 25832 36116 25838 36168
rect 25884 36165 25912 36196
rect 26602 36184 26608 36196
rect 26660 36224 26666 36236
rect 29178 36224 29184 36236
rect 26660 36196 27568 36224
rect 29139 36196 29184 36224
rect 26660 36184 26666 36196
rect 25869 36159 25927 36165
rect 25869 36125 25881 36159
rect 25915 36125 25927 36159
rect 27338 36156 27344 36168
rect 25869 36119 25927 36125
rect 26528 36128 27344 36156
rect 4856 36060 5580 36088
rect 6273 36091 6331 36097
rect 4856 36048 4862 36060
rect 6273 36057 6285 36091
rect 6319 36057 6331 36091
rect 17402 36088 17408 36100
rect 6273 36051 6331 36057
rect 6886 36060 17408 36088
rect 6288 36020 6316 36051
rect 6546 36020 6552 36032
rect 6288 35992 6552 36020
rect 6546 35980 6552 35992
rect 6604 36020 6610 36032
rect 6886 36020 6914 36060
rect 17402 36048 17408 36060
rect 17460 36048 17466 36100
rect 26528 36097 26556 36128
rect 27338 36116 27344 36128
rect 27396 36116 27402 36168
rect 27540 36165 27568 36196
rect 29178 36184 29184 36196
rect 29236 36224 29242 36236
rect 30576 36224 30604 36264
rect 30834 36252 30840 36264
rect 30892 36252 30898 36304
rect 31110 36224 31116 36236
rect 29236 36196 30604 36224
rect 30668 36196 31116 36224
rect 29236 36184 29242 36196
rect 27525 36159 27583 36165
rect 27525 36125 27537 36159
rect 27571 36125 27583 36159
rect 27525 36119 27583 36125
rect 27798 36116 27804 36168
rect 27856 36156 27862 36168
rect 28169 36159 28227 36165
rect 28169 36156 28181 36159
rect 27856 36128 28181 36156
rect 27856 36116 27862 36128
rect 28169 36125 28181 36128
rect 28215 36125 28227 36159
rect 28169 36119 28227 36125
rect 28258 36116 28264 36168
rect 28316 36156 28322 36168
rect 28353 36159 28411 36165
rect 28353 36156 28365 36159
rect 28316 36128 28365 36156
rect 28316 36116 28322 36128
rect 28353 36125 28365 36128
rect 28399 36125 28411 36159
rect 28902 36156 28908 36168
rect 28863 36128 28908 36156
rect 28353 36119 28411 36125
rect 28902 36116 28908 36128
rect 28960 36116 28966 36168
rect 29914 36156 29920 36168
rect 29875 36128 29920 36156
rect 29914 36116 29920 36128
rect 29972 36116 29978 36168
rect 30668 36165 30696 36196
rect 31110 36184 31116 36196
rect 31168 36184 31174 36236
rect 32692 36233 32720 36332
rect 32677 36227 32735 36233
rect 31220 36196 31616 36224
rect 30009 36159 30067 36165
rect 30009 36125 30021 36159
rect 30055 36125 30067 36159
rect 30009 36119 30067 36125
rect 30653 36159 30711 36165
rect 30653 36125 30665 36159
rect 30699 36125 30711 36159
rect 30653 36119 30711 36125
rect 30837 36159 30895 36165
rect 30837 36125 30849 36159
rect 30883 36156 30895 36159
rect 31220 36156 31248 36196
rect 31588 36168 31616 36196
rect 32677 36193 32689 36227
rect 32723 36193 32735 36227
rect 34330 36224 34336 36236
rect 34291 36196 34336 36224
rect 32677 36187 32735 36193
rect 34330 36184 34336 36196
rect 34388 36184 34394 36236
rect 30883 36128 31248 36156
rect 31481 36159 31539 36165
rect 30883 36125 30895 36128
rect 30837 36119 30895 36125
rect 31481 36125 31493 36159
rect 31527 36125 31539 36159
rect 31481 36119 31539 36125
rect 26513 36091 26571 36097
rect 26513 36057 26525 36091
rect 26559 36057 26571 36091
rect 26513 36051 26571 36057
rect 26729 36091 26787 36097
rect 26729 36057 26741 36091
rect 26775 36088 26787 36091
rect 26775 36060 27200 36088
rect 26775 36057 26787 36060
rect 26729 36051 26787 36057
rect 18230 36020 18236 36032
rect 6604 35992 6914 36020
rect 18191 35992 18236 36020
rect 6604 35980 6610 35992
rect 18230 35980 18236 35992
rect 18288 35980 18294 36032
rect 19886 36020 19892 36032
rect 19847 35992 19892 36020
rect 19886 35980 19892 35992
rect 19944 35980 19950 36032
rect 20162 35980 20168 36032
rect 20220 36020 20226 36032
rect 20441 36023 20499 36029
rect 20441 36020 20453 36023
rect 20220 35992 20453 36020
rect 20220 35980 20226 35992
rect 20441 35989 20453 35992
rect 20487 35989 20499 36023
rect 21082 36020 21088 36032
rect 21043 35992 21088 36020
rect 20441 35983 20499 35989
rect 21082 35980 21088 35992
rect 21140 35980 21146 36032
rect 21729 36023 21787 36029
rect 21729 35989 21741 36023
rect 21775 36020 21787 36023
rect 22462 36020 22468 36032
rect 21775 35992 22468 36020
rect 21775 35989 21787 35992
rect 21729 35983 21787 35989
rect 22462 35980 22468 35992
rect 22520 35980 22526 36032
rect 24581 36023 24639 36029
rect 24581 35989 24593 36023
rect 24627 36020 24639 36023
rect 24670 36020 24676 36032
rect 24627 35992 24676 36020
rect 24627 35989 24639 35992
rect 24581 35983 24639 35989
rect 24670 35980 24676 35992
rect 24728 35980 24734 36032
rect 26878 35980 26884 36032
rect 26936 36020 26942 36032
rect 27172 36020 27200 36060
rect 29086 36048 29092 36100
rect 29144 36088 29150 36100
rect 30024 36088 30052 36119
rect 30190 36088 30196 36100
rect 29144 36060 29500 36088
rect 30024 36060 30196 36088
rect 29144 36048 29150 36060
rect 27430 36020 27436 36032
rect 26936 35992 26981 36020
rect 27172 35992 27436 36020
rect 26936 35980 26942 35992
rect 27430 35980 27436 35992
rect 27488 35980 27494 36032
rect 28261 36023 28319 36029
rect 28261 35989 28273 36023
rect 28307 36020 28319 36023
rect 28718 36020 28724 36032
rect 28307 35992 28724 36020
rect 28307 35989 28319 35992
rect 28261 35983 28319 35989
rect 28718 35980 28724 35992
rect 28776 35980 28782 36032
rect 29181 36023 29239 36029
rect 29181 35989 29193 36023
rect 29227 36020 29239 36023
rect 29362 36020 29368 36032
rect 29227 35992 29368 36020
rect 29227 35989 29239 35992
rect 29181 35983 29239 35989
rect 29362 35980 29368 35992
rect 29420 35980 29426 36032
rect 29472 36020 29500 36060
rect 30190 36048 30196 36060
rect 30248 36088 30254 36100
rect 30852 36088 30880 36119
rect 30248 36060 30880 36088
rect 31493 36088 31521 36119
rect 31570 36116 31576 36168
rect 31628 36156 31634 36168
rect 31665 36159 31723 36165
rect 31665 36156 31677 36159
rect 31628 36128 31677 36156
rect 31628 36116 31634 36128
rect 31665 36125 31677 36128
rect 31711 36125 31723 36159
rect 31665 36119 31723 36125
rect 32493 36159 32551 36165
rect 32493 36125 32505 36159
rect 32539 36125 32551 36159
rect 32493 36119 32551 36125
rect 32030 36088 32036 36100
rect 31493 36060 32036 36088
rect 30248 36048 30254 36060
rect 32030 36048 32036 36060
rect 32088 36048 32094 36100
rect 32508 36020 32536 36119
rect 29472 35992 32536 36020
rect 1104 35930 35027 35952
rect 1104 35878 9390 35930
rect 9442 35878 9454 35930
rect 9506 35878 9518 35930
rect 9570 35878 9582 35930
rect 9634 35878 9646 35930
rect 9698 35878 17831 35930
rect 17883 35878 17895 35930
rect 17947 35878 17959 35930
rect 18011 35878 18023 35930
rect 18075 35878 18087 35930
rect 18139 35878 26272 35930
rect 26324 35878 26336 35930
rect 26388 35878 26400 35930
rect 26452 35878 26464 35930
rect 26516 35878 26528 35930
rect 26580 35878 34713 35930
rect 34765 35878 34777 35930
rect 34829 35878 34841 35930
rect 34893 35878 34905 35930
rect 34957 35878 34969 35930
rect 35021 35878 35027 35930
rect 1104 35856 35027 35878
rect 21177 35819 21235 35825
rect 21177 35785 21189 35819
rect 21223 35816 21235 35819
rect 21266 35816 21272 35828
rect 21223 35788 21272 35816
rect 21223 35785 21235 35788
rect 21177 35779 21235 35785
rect 21266 35776 21272 35788
rect 21324 35776 21330 35828
rect 22370 35776 22376 35828
rect 22428 35816 22434 35828
rect 22465 35819 22523 35825
rect 22465 35816 22477 35819
rect 22428 35788 22477 35816
rect 22428 35776 22434 35788
rect 22465 35785 22477 35788
rect 22511 35785 22523 35819
rect 22465 35779 22523 35785
rect 25130 35776 25136 35828
rect 25188 35816 25194 35828
rect 26421 35819 26479 35825
rect 26421 35816 26433 35819
rect 25188 35788 26433 35816
rect 25188 35776 25194 35788
rect 26421 35785 26433 35788
rect 26467 35785 26479 35819
rect 26421 35779 26479 35785
rect 28166 35776 28172 35828
rect 28224 35816 28230 35828
rect 28353 35819 28411 35825
rect 28353 35816 28365 35819
rect 28224 35788 28365 35816
rect 28224 35776 28230 35788
rect 28353 35785 28365 35788
rect 28399 35785 28411 35819
rect 28353 35779 28411 35785
rect 29178 35776 29184 35828
rect 29236 35816 29242 35828
rect 29273 35819 29331 35825
rect 29273 35816 29285 35819
rect 29236 35788 29285 35816
rect 29236 35776 29242 35788
rect 29273 35785 29285 35788
rect 29319 35785 29331 35819
rect 29273 35779 29331 35785
rect 30006 35776 30012 35828
rect 30064 35816 30070 35828
rect 30101 35819 30159 35825
rect 30101 35816 30113 35819
rect 30064 35788 30113 35816
rect 30064 35776 30070 35788
rect 30101 35785 30113 35788
rect 30147 35785 30159 35819
rect 34241 35819 34299 35825
rect 34241 35816 34253 35819
rect 30101 35779 30159 35785
rect 31588 35788 31984 35816
rect 18230 35708 18236 35760
rect 18288 35748 18294 35760
rect 18386 35751 18444 35757
rect 18386 35748 18398 35751
rect 18288 35720 18398 35748
rect 18288 35708 18294 35720
rect 18386 35717 18398 35720
rect 18432 35717 18444 35751
rect 18386 35711 18444 35717
rect 23652 35751 23710 35757
rect 23652 35717 23664 35751
rect 23698 35748 23710 35751
rect 24302 35748 24308 35760
rect 23698 35720 24308 35748
rect 23698 35717 23710 35720
rect 23652 35711 23710 35717
rect 24302 35708 24308 35720
rect 24360 35708 24366 35760
rect 25774 35708 25780 35760
rect 25832 35748 25838 35760
rect 25832 35720 27200 35748
rect 25832 35708 25838 35720
rect 1765 35683 1823 35689
rect 1765 35649 1777 35683
rect 1811 35680 1823 35683
rect 2498 35680 2504 35692
rect 1811 35652 2504 35680
rect 1811 35649 1823 35652
rect 1765 35643 1823 35649
rect 2498 35640 2504 35652
rect 2556 35680 2562 35692
rect 3053 35683 3111 35689
rect 3053 35680 3065 35683
rect 2556 35652 3065 35680
rect 2556 35640 2562 35652
rect 3053 35649 3065 35652
rect 3099 35649 3111 35683
rect 3053 35643 3111 35649
rect 3970 35640 3976 35692
rect 4028 35680 4034 35692
rect 4525 35683 4583 35689
rect 4525 35680 4537 35683
rect 4028 35652 4537 35680
rect 4028 35640 4034 35652
rect 4525 35649 4537 35652
rect 4571 35649 4583 35683
rect 4525 35643 4583 35649
rect 16574 35640 16580 35692
rect 16632 35680 16638 35692
rect 17497 35683 17555 35689
rect 17497 35680 17509 35683
rect 16632 35652 17509 35680
rect 16632 35640 16638 35652
rect 17497 35649 17509 35652
rect 17543 35649 17555 35683
rect 17497 35643 17555 35649
rect 17678 35640 17684 35692
rect 17736 35680 17742 35692
rect 20165 35683 20223 35689
rect 17736 35652 20116 35680
rect 17736 35640 17742 35652
rect 2038 35612 2044 35624
rect 1999 35584 2044 35612
rect 2038 35572 2044 35584
rect 2096 35572 2102 35624
rect 3878 35612 3884 35624
rect 3839 35584 3884 35612
rect 3878 35572 3884 35584
rect 3936 35572 3942 35624
rect 5353 35615 5411 35621
rect 5353 35581 5365 35615
rect 5399 35612 5411 35615
rect 6546 35612 6552 35624
rect 5399 35584 6552 35612
rect 5399 35581 5411 35584
rect 5353 35575 5411 35581
rect 6546 35572 6552 35584
rect 6604 35572 6610 35624
rect 18141 35615 18199 35621
rect 18141 35581 18153 35615
rect 18187 35581 18199 35615
rect 18141 35575 18199 35581
rect 17586 35476 17592 35488
rect 17547 35448 17592 35476
rect 17586 35436 17592 35448
rect 17644 35436 17650 35488
rect 18156 35476 18184 35575
rect 19242 35476 19248 35488
rect 18156 35448 19248 35476
rect 19242 35436 19248 35448
rect 19300 35436 19306 35488
rect 19518 35476 19524 35488
rect 19479 35448 19524 35476
rect 19518 35436 19524 35448
rect 19576 35436 19582 35488
rect 19978 35476 19984 35488
rect 19939 35448 19984 35476
rect 19978 35436 19984 35448
rect 20036 35436 20042 35488
rect 20088 35476 20116 35652
rect 20165 35649 20177 35683
rect 20211 35680 20223 35683
rect 20714 35680 20720 35692
rect 20211 35652 20720 35680
rect 20211 35649 20223 35652
rect 20165 35643 20223 35649
rect 20714 35640 20720 35652
rect 20772 35640 20778 35692
rect 20990 35680 20996 35692
rect 20903 35652 20996 35680
rect 20990 35640 20996 35652
rect 21048 35680 21054 35692
rect 21266 35680 21272 35692
rect 21048 35652 21272 35680
rect 21048 35640 21054 35652
rect 21266 35640 21272 35652
rect 21324 35680 21330 35692
rect 22281 35683 22339 35689
rect 22281 35680 22293 35683
rect 21324 35652 22293 35680
rect 21324 35640 21330 35652
rect 22281 35649 22293 35652
rect 22327 35680 22339 35683
rect 22738 35680 22744 35692
rect 22327 35652 22744 35680
rect 22327 35649 22339 35652
rect 22281 35643 22339 35649
rect 22738 35640 22744 35652
rect 22796 35640 22802 35692
rect 25222 35680 25228 35692
rect 23032 35652 24440 35680
rect 25183 35652 25228 35680
rect 20622 35572 20628 35624
rect 20680 35612 20686 35624
rect 20809 35615 20867 35621
rect 20809 35612 20821 35615
rect 20680 35584 20821 35612
rect 20680 35572 20686 35584
rect 20809 35581 20821 35584
rect 20855 35581 20867 35615
rect 20809 35575 20867 35581
rect 22097 35615 22155 35621
rect 22097 35581 22109 35615
rect 22143 35612 22155 35615
rect 22922 35612 22928 35624
rect 22143 35584 22928 35612
rect 22143 35581 22155 35584
rect 22097 35575 22155 35581
rect 22922 35572 22928 35584
rect 22980 35572 22986 35624
rect 23032 35476 23060 35652
rect 23382 35612 23388 35624
rect 23343 35584 23388 35612
rect 23382 35572 23388 35584
rect 23440 35572 23446 35624
rect 24412 35544 24440 35652
rect 25222 35640 25228 35652
rect 25280 35640 25286 35692
rect 26237 35683 26295 35689
rect 26237 35649 26249 35683
rect 26283 35680 26295 35683
rect 26602 35680 26608 35692
rect 26283 35652 26608 35680
rect 26283 35649 26295 35652
rect 26237 35643 26295 35649
rect 26602 35640 26608 35652
rect 26660 35640 26666 35692
rect 27062 35680 27068 35692
rect 26712 35652 27068 35680
rect 25130 35572 25136 35624
rect 25188 35612 25194 35624
rect 25317 35615 25375 35621
rect 25317 35612 25329 35615
rect 25188 35584 25329 35612
rect 25188 35572 25194 35584
rect 25317 35581 25329 35584
rect 25363 35581 25375 35615
rect 25317 35575 25375 35581
rect 26053 35615 26111 35621
rect 26053 35581 26065 35615
rect 26099 35612 26111 35615
rect 26712 35612 26740 35652
rect 27062 35640 27068 35652
rect 27120 35640 27126 35692
rect 27172 35689 27200 35720
rect 27890 35708 27896 35760
rect 27948 35748 27954 35760
rect 30561 35751 30619 35757
rect 27948 35720 28212 35748
rect 27948 35708 27954 35720
rect 28184 35689 28212 35720
rect 30561 35717 30573 35751
rect 30607 35748 30619 35751
rect 31588 35748 31616 35788
rect 31956 35760 31984 35788
rect 33244 35788 34253 35816
rect 30607 35720 31616 35748
rect 30607 35717 30619 35720
rect 30561 35711 30619 35717
rect 31938 35708 31944 35760
rect 31996 35708 32002 35760
rect 27157 35683 27215 35689
rect 27157 35649 27169 35683
rect 27203 35649 27215 35683
rect 27157 35643 27215 35649
rect 28169 35683 28227 35689
rect 28169 35649 28181 35683
rect 28215 35680 28227 35683
rect 29089 35683 29147 35689
rect 29089 35680 29101 35683
rect 28215 35652 29101 35680
rect 28215 35649 28227 35652
rect 28169 35643 28227 35649
rect 29089 35649 29101 35652
rect 29135 35680 29147 35683
rect 29914 35680 29920 35692
rect 29135 35652 29920 35680
rect 29135 35649 29147 35652
rect 29089 35643 29147 35649
rect 29914 35640 29920 35652
rect 29972 35680 29978 35692
rect 30190 35680 30196 35692
rect 29972 35652 30196 35680
rect 29972 35640 29978 35652
rect 30190 35640 30196 35652
rect 30248 35640 30254 35692
rect 30745 35683 30803 35689
rect 30745 35649 30757 35683
rect 30791 35680 30803 35683
rect 31559 35683 31617 35689
rect 30791 35678 31156 35680
rect 31220 35678 31524 35680
rect 30791 35652 31524 35678
rect 30791 35649 30803 35652
rect 31128 35650 31248 35652
rect 30745 35643 30803 35649
rect 26099 35584 26740 35612
rect 26099 35581 26111 35584
rect 26053 35575 26111 35581
rect 26786 35572 26792 35624
rect 26844 35612 26850 35624
rect 27249 35615 27307 35621
rect 27249 35612 27261 35615
rect 26844 35584 27261 35612
rect 26844 35572 26850 35584
rect 27249 35581 27261 35584
rect 27295 35612 27307 35615
rect 27338 35612 27344 35624
rect 27295 35584 27344 35612
rect 27295 35581 27307 35584
rect 27249 35575 27307 35581
rect 27338 35572 27344 35584
rect 27396 35572 27402 35624
rect 27985 35615 28043 35621
rect 27985 35581 27997 35615
rect 28031 35612 28043 35615
rect 28074 35612 28080 35624
rect 28031 35584 28080 35612
rect 28031 35581 28043 35584
rect 27985 35575 28043 35581
rect 28074 35572 28080 35584
rect 28132 35612 28138 35624
rect 28534 35612 28540 35624
rect 28132 35584 28540 35612
rect 28132 35572 28138 35584
rect 28534 35572 28540 35584
rect 28592 35572 28598 35624
rect 28810 35572 28816 35624
rect 28868 35612 28874 35624
rect 28905 35615 28963 35621
rect 28905 35612 28917 35615
rect 28868 35584 28917 35612
rect 28868 35572 28874 35584
rect 28905 35581 28917 35584
rect 28951 35581 28963 35615
rect 28905 35575 28963 35581
rect 29178 35572 29184 35624
rect 29236 35612 29242 35624
rect 29733 35615 29791 35621
rect 29733 35612 29745 35615
rect 29236 35584 29745 35612
rect 29236 35572 29242 35584
rect 29733 35581 29745 35584
rect 29779 35581 29791 35615
rect 29733 35575 29791 35581
rect 30929 35615 30987 35621
rect 30929 35581 30941 35615
rect 30975 35612 30987 35615
rect 31018 35612 31024 35624
rect 30975 35584 31024 35612
rect 30975 35581 30987 35584
rect 30929 35575 30987 35581
rect 31018 35572 31024 35584
rect 31076 35572 31082 35624
rect 31389 35615 31447 35621
rect 31389 35581 31401 35615
rect 31435 35581 31447 35615
rect 31496 35612 31524 35652
rect 31559 35649 31571 35683
rect 31605 35680 31617 35683
rect 31662 35680 31668 35692
rect 31605 35652 31668 35680
rect 31605 35649 31617 35652
rect 31559 35643 31617 35649
rect 31662 35640 31668 35652
rect 31720 35640 31726 35692
rect 31754 35640 31760 35692
rect 31812 35680 31818 35692
rect 32585 35683 32643 35689
rect 32585 35680 32597 35683
rect 31812 35652 32597 35680
rect 31812 35640 31818 35652
rect 32585 35649 32597 35652
rect 32631 35649 32643 35683
rect 32585 35643 32643 35649
rect 32950 35640 32956 35692
rect 33008 35680 33014 35692
rect 33244 35689 33272 35788
rect 34241 35785 34253 35788
rect 34287 35785 34299 35819
rect 34241 35779 34299 35785
rect 34054 35748 34060 35760
rect 34015 35720 34060 35748
rect 34054 35708 34060 35720
rect 34112 35708 34118 35760
rect 33229 35683 33287 35689
rect 33229 35680 33241 35683
rect 33008 35652 33241 35680
rect 33008 35640 33014 35652
rect 33229 35649 33241 35652
rect 33275 35649 33287 35683
rect 33229 35643 33287 35649
rect 33413 35683 33471 35689
rect 33413 35649 33425 35683
rect 33459 35649 33471 35683
rect 33413 35643 33471 35649
rect 34333 35683 34391 35689
rect 34333 35649 34345 35683
rect 34379 35649 34391 35683
rect 34333 35643 34391 35649
rect 31846 35612 31852 35624
rect 31496 35584 31852 35612
rect 31389 35575 31447 35581
rect 28626 35544 28632 35556
rect 24412 35516 28632 35544
rect 28626 35504 28632 35516
rect 28684 35504 28690 35556
rect 30834 35504 30840 35556
rect 30892 35544 30898 35556
rect 31404 35544 31432 35575
rect 31846 35572 31852 35584
rect 31904 35572 31910 35624
rect 32401 35615 32459 35621
rect 32401 35581 32413 35615
rect 32447 35612 32459 35615
rect 32858 35612 32864 35624
rect 32447 35584 32864 35612
rect 32447 35581 32459 35584
rect 32401 35575 32459 35581
rect 32858 35572 32864 35584
rect 32916 35612 32922 35624
rect 33428 35612 33456 35643
rect 32916 35584 33456 35612
rect 32916 35572 32922 35584
rect 33502 35572 33508 35624
rect 33560 35612 33566 35624
rect 34348 35612 34376 35643
rect 33560 35584 34376 35612
rect 33560 35572 33566 35584
rect 30892 35516 31432 35544
rect 30892 35504 30898 35516
rect 20088 35448 23060 35476
rect 23106 35436 23112 35488
rect 23164 35476 23170 35488
rect 24765 35479 24823 35485
rect 24765 35476 24777 35479
rect 23164 35448 24777 35476
rect 23164 35436 23170 35448
rect 24765 35445 24777 35448
rect 24811 35445 24823 35479
rect 24765 35439 24823 35445
rect 25409 35479 25467 35485
rect 25409 35445 25421 35479
rect 25455 35476 25467 35479
rect 25498 35476 25504 35488
rect 25455 35448 25504 35476
rect 25455 35445 25467 35448
rect 25409 35439 25467 35445
rect 25498 35436 25504 35448
rect 25556 35436 25562 35488
rect 25593 35479 25651 35485
rect 25593 35445 25605 35479
rect 25639 35476 25651 35479
rect 26050 35476 26056 35488
rect 25639 35448 26056 35476
rect 25639 35445 25651 35448
rect 25593 35439 25651 35445
rect 26050 35436 26056 35448
rect 26108 35436 26114 35488
rect 26510 35436 26516 35488
rect 26568 35476 26574 35488
rect 27157 35479 27215 35485
rect 27157 35476 27169 35479
rect 26568 35448 27169 35476
rect 26568 35436 26574 35448
rect 27157 35445 27169 35448
rect 27203 35445 27215 35479
rect 27522 35476 27528 35488
rect 27483 35448 27528 35476
rect 27157 35439 27215 35445
rect 27522 35436 27528 35448
rect 27580 35436 27586 35488
rect 27614 35436 27620 35488
rect 27672 35476 27678 35488
rect 30926 35476 30932 35488
rect 27672 35448 30932 35476
rect 27672 35436 27678 35448
rect 30926 35436 30932 35448
rect 30984 35436 30990 35488
rect 31754 35476 31760 35488
rect 31715 35448 31760 35476
rect 31754 35436 31760 35448
rect 31812 35436 31818 35488
rect 32766 35476 32772 35488
rect 32727 35448 32772 35476
rect 32766 35436 32772 35448
rect 32824 35436 32830 35488
rect 33134 35436 33140 35488
rect 33192 35476 33198 35488
rect 33597 35479 33655 35485
rect 33597 35476 33609 35479
rect 33192 35448 33609 35476
rect 33192 35436 33198 35448
rect 33597 35445 33609 35448
rect 33643 35445 33655 35479
rect 33597 35439 33655 35445
rect 33686 35436 33692 35488
rect 33744 35476 33750 35488
rect 34057 35479 34115 35485
rect 34057 35476 34069 35479
rect 33744 35448 34069 35476
rect 33744 35436 33750 35448
rect 34057 35445 34069 35448
rect 34103 35445 34115 35479
rect 34057 35439 34115 35445
rect 1104 35386 34868 35408
rect 1104 35334 5170 35386
rect 5222 35334 5234 35386
rect 5286 35334 5298 35386
rect 5350 35334 5362 35386
rect 5414 35334 5426 35386
rect 5478 35334 13611 35386
rect 13663 35334 13675 35386
rect 13727 35334 13739 35386
rect 13791 35334 13803 35386
rect 13855 35334 13867 35386
rect 13919 35334 22052 35386
rect 22104 35334 22116 35386
rect 22168 35334 22180 35386
rect 22232 35334 22244 35386
rect 22296 35334 22308 35386
rect 22360 35334 30493 35386
rect 30545 35334 30557 35386
rect 30609 35334 30621 35386
rect 30673 35334 30685 35386
rect 30737 35334 30749 35386
rect 30801 35334 34868 35386
rect 1104 35312 34868 35334
rect 18414 35232 18420 35284
rect 18472 35272 18478 35284
rect 18509 35275 18567 35281
rect 18509 35272 18521 35275
rect 18472 35244 18521 35272
rect 18472 35232 18478 35244
rect 18509 35241 18521 35244
rect 18555 35241 18567 35275
rect 18509 35235 18567 35241
rect 20622 35232 20628 35284
rect 20680 35272 20686 35284
rect 21269 35275 21327 35281
rect 21269 35272 21281 35275
rect 20680 35244 21281 35272
rect 20680 35232 20686 35244
rect 21269 35241 21281 35244
rect 21315 35241 21327 35275
rect 21269 35235 21327 35241
rect 22370 35232 22376 35284
rect 22428 35272 22434 35284
rect 22465 35275 22523 35281
rect 22465 35272 22477 35275
rect 22428 35244 22477 35272
rect 22428 35232 22434 35244
rect 22465 35241 22477 35244
rect 22511 35241 22523 35275
rect 22922 35272 22928 35284
rect 22883 35244 22928 35272
rect 22465 35235 22523 35241
rect 22922 35232 22928 35244
rect 22980 35232 22986 35284
rect 23290 35272 23296 35284
rect 23032 35244 23296 35272
rect 21358 35204 21364 35216
rect 18156 35176 21364 35204
rect 2774 35136 2780 35148
rect 2735 35108 2780 35136
rect 2774 35096 2780 35108
rect 2832 35096 2838 35148
rect 16666 35096 16672 35148
rect 16724 35136 16730 35148
rect 18156 35145 18184 35176
rect 21358 35164 21364 35176
rect 21416 35204 21422 35216
rect 23032 35204 23060 35244
rect 23290 35232 23296 35244
rect 23348 35232 23354 35284
rect 25866 35232 25872 35284
rect 25924 35272 25930 35284
rect 26789 35275 26847 35281
rect 26789 35272 26801 35275
rect 25924 35244 26801 35272
rect 25924 35232 25930 35244
rect 26789 35241 26801 35244
rect 26835 35241 26847 35275
rect 26789 35235 26847 35241
rect 27154 35232 27160 35284
rect 27212 35272 27218 35284
rect 27212 35244 30144 35272
rect 27212 35232 27218 35244
rect 21416 35176 23060 35204
rect 21416 35164 21422 35176
rect 23106 35164 23112 35216
rect 23164 35164 23170 35216
rect 28994 35164 29000 35216
rect 29052 35204 29058 35216
rect 29362 35204 29368 35216
rect 29052 35176 29368 35204
rect 29052 35164 29058 35176
rect 29362 35164 29368 35176
rect 29420 35164 29426 35216
rect 29638 35164 29644 35216
rect 29696 35204 29702 35216
rect 29822 35204 29828 35216
rect 29696 35176 29828 35204
rect 29696 35164 29702 35176
rect 29822 35164 29828 35176
rect 29880 35164 29886 35216
rect 30116 35213 30144 35244
rect 30101 35207 30159 35213
rect 30101 35173 30113 35207
rect 30147 35173 30159 35207
rect 30101 35167 30159 35173
rect 18141 35139 18199 35145
rect 16724 35108 17540 35136
rect 16724 35096 16730 35108
rect 1581 35071 1639 35077
rect 1581 35037 1593 35071
rect 1627 35037 1639 35071
rect 3970 35068 3976 35080
rect 3883 35040 3976 35068
rect 1581 35031 1639 35037
rect 1596 34932 1624 35031
rect 3970 35028 3976 35040
rect 4028 35028 4034 35080
rect 17512 35077 17540 35108
rect 18141 35105 18153 35139
rect 18187 35105 18199 35139
rect 21450 35136 21456 35148
rect 18141 35099 18199 35105
rect 21284 35108 21456 35136
rect 17405 35071 17463 35077
rect 17405 35037 17417 35071
rect 17451 35037 17463 35071
rect 17405 35031 17463 35037
rect 17497 35071 17555 35077
rect 17497 35037 17509 35071
rect 17543 35037 17555 35071
rect 17497 35031 17555 35037
rect 1765 35003 1823 35009
rect 1765 34969 1777 35003
rect 1811 35000 1823 35003
rect 2130 35000 2136 35012
rect 1811 34972 2136 35000
rect 1811 34969 1823 34972
rect 1765 34963 1823 34969
rect 2130 34960 2136 34972
rect 2188 34960 2194 35012
rect 2498 34960 2504 35012
rect 2556 35000 2562 35012
rect 3988 35000 4016 35028
rect 2556 34972 4016 35000
rect 2556 34960 2562 34972
rect 4706 34960 4712 35012
rect 4764 35000 4770 35012
rect 4801 35003 4859 35009
rect 4801 35000 4813 35003
rect 4764 34972 4813 35000
rect 4764 34960 4770 34972
rect 4801 34969 4813 34972
rect 4847 35000 4859 35003
rect 5534 35000 5540 35012
rect 4847 34972 5540 35000
rect 4847 34969 4859 34972
rect 4801 34963 4859 34969
rect 5534 34960 5540 34972
rect 5592 34960 5598 35012
rect 17420 35000 17448 35031
rect 18156 35000 18184 35099
rect 18322 35068 18328 35080
rect 18283 35040 18328 35068
rect 18322 35028 18328 35040
rect 18380 35028 18386 35080
rect 19518 35068 19524 35080
rect 19431 35040 19524 35068
rect 19518 35028 19524 35040
rect 19576 35028 19582 35080
rect 19613 35071 19671 35077
rect 19613 35037 19625 35071
rect 19659 35068 19671 35071
rect 20990 35068 20996 35080
rect 19659 35040 20996 35068
rect 19659 35037 19671 35040
rect 19613 35031 19671 35037
rect 20990 35028 20996 35040
rect 21048 35028 21054 35080
rect 21284 35077 21312 35108
rect 21450 35096 21456 35108
rect 21508 35096 21514 35148
rect 22738 35136 22744 35148
rect 22296 35108 22744 35136
rect 21269 35071 21327 35077
rect 21269 35037 21281 35071
rect 21315 35037 21327 35071
rect 21269 35031 21327 35037
rect 21361 35071 21419 35077
rect 21361 35037 21373 35071
rect 21407 35037 21419 35071
rect 22186 35068 22192 35080
rect 22147 35040 22192 35068
rect 21361 35031 21419 35037
rect 17420 34972 18184 35000
rect 19536 35000 19564 35028
rect 20254 35000 20260 35012
rect 19536 34972 19932 35000
rect 20215 34972 20260 35000
rect 2866 34932 2872 34944
rect 1596 34904 2872 34932
rect 2866 34892 2872 34904
rect 2924 34892 2930 34944
rect 17681 34935 17739 34941
rect 17681 34901 17693 34935
rect 17727 34932 17739 34935
rect 18322 34932 18328 34944
rect 17727 34904 18328 34932
rect 17727 34901 17739 34904
rect 17681 34895 17739 34901
rect 18322 34892 18328 34904
rect 18380 34892 18386 34944
rect 19794 34932 19800 34944
rect 19755 34904 19800 34932
rect 19794 34892 19800 34904
rect 19852 34892 19858 34944
rect 19904 34932 19932 34972
rect 20254 34960 20260 34972
rect 20312 34960 20318 35012
rect 20533 35003 20591 35009
rect 20533 34969 20545 35003
rect 20579 35000 20591 35003
rect 21376 35000 21404 35031
rect 22186 35028 22192 35040
rect 22244 35028 22250 35080
rect 22296 35077 22324 35108
rect 22738 35096 22744 35108
rect 22796 35096 22802 35148
rect 23124 35077 23152 35164
rect 24578 35136 24584 35148
rect 24539 35108 24584 35136
rect 24578 35096 24584 35108
rect 24636 35096 24642 35148
rect 28626 35096 28632 35148
rect 28684 35136 28690 35148
rect 32677 35139 32735 35145
rect 32677 35136 32689 35139
rect 28684 35108 30788 35136
rect 28684 35096 28690 35108
rect 23290 35077 23296 35080
rect 22281 35071 22339 35077
rect 22281 35037 22293 35071
rect 22327 35037 22339 35071
rect 22281 35031 22339 35037
rect 23109 35071 23167 35077
rect 23109 35037 23121 35071
rect 23155 35037 23167 35071
rect 23109 35031 23167 35037
rect 23241 35071 23296 35077
rect 23241 35037 23253 35071
rect 23287 35037 23296 35071
rect 23241 35031 23296 35037
rect 23290 35028 23296 35031
rect 23348 35028 23354 35080
rect 24854 35077 24860 35080
rect 24029 35071 24087 35077
rect 24029 35037 24041 35071
rect 24075 35068 24087 35071
rect 24848 35068 24860 35077
rect 24075 35040 24716 35068
rect 24815 35040 24860 35068
rect 24075 35037 24087 35040
rect 24029 35031 24087 35037
rect 22370 35000 22376 35012
rect 20579 34972 22376 35000
rect 20579 34969 20591 34972
rect 20533 34963 20591 34969
rect 22370 34960 22376 34972
rect 22428 34960 22434 35012
rect 22925 35003 22983 35009
rect 22925 35000 22937 35003
rect 22480 34972 22937 35000
rect 20438 34932 20444 34944
rect 19904 34904 20444 34932
rect 20438 34892 20444 34904
rect 20496 34892 20502 34944
rect 20622 34932 20628 34944
rect 20583 34904 20628 34932
rect 20622 34892 20628 34904
rect 20680 34892 20686 34944
rect 20806 34932 20812 34944
rect 20767 34904 20812 34932
rect 20806 34892 20812 34904
rect 20864 34892 20870 34944
rect 21634 34932 21640 34944
rect 21595 34904 21640 34932
rect 21634 34892 21640 34904
rect 21692 34892 21698 34944
rect 22186 34892 22192 34944
rect 22244 34932 22250 34944
rect 22480 34932 22508 34972
rect 22925 34969 22937 34972
rect 22971 35000 22983 35003
rect 23566 35000 23572 35012
rect 22971 34972 23572 35000
rect 22971 34969 22983 34972
rect 22925 34963 22983 34969
rect 23566 34960 23572 34972
rect 23624 34960 23630 35012
rect 24688 35000 24716 35040
rect 24848 35031 24860 35040
rect 24854 35028 24860 35031
rect 24912 35028 24918 35080
rect 26510 35068 26516 35080
rect 26471 35040 26516 35068
rect 26510 35028 26516 35040
rect 26568 35028 26574 35080
rect 26605 35071 26663 35077
rect 26605 35037 26617 35071
rect 26651 35037 26663 35071
rect 26605 35031 26663 35037
rect 26620 35000 26648 35031
rect 27154 35028 27160 35080
rect 27212 35068 27218 35080
rect 27617 35071 27675 35077
rect 27617 35068 27629 35071
rect 27212 35040 27629 35068
rect 27212 35028 27218 35040
rect 27617 35037 27629 35040
rect 27663 35068 27675 35071
rect 29822 35068 29828 35080
rect 27663 35040 28304 35068
rect 29783 35040 29828 35068
rect 27663 35037 27675 35040
rect 27617 35031 27675 35037
rect 27706 35000 27712 35012
rect 24688 34972 26556 35000
rect 26620 34972 27712 35000
rect 22244 34904 22508 34932
rect 22244 34892 22250 34904
rect 22738 34892 22744 34944
rect 22796 34932 22802 34944
rect 23385 34935 23443 34941
rect 23385 34932 23397 34935
rect 22796 34904 23397 34932
rect 22796 34892 22802 34904
rect 23385 34901 23397 34904
rect 23431 34901 23443 34935
rect 23385 34895 23443 34901
rect 23845 34935 23903 34941
rect 23845 34901 23857 34935
rect 23891 34932 23903 34935
rect 24854 34932 24860 34944
rect 23891 34904 24860 34932
rect 23891 34901 23903 34904
rect 23845 34895 23903 34901
rect 24854 34892 24860 34904
rect 24912 34892 24918 34944
rect 25866 34892 25872 34944
rect 25924 34932 25930 34944
rect 25961 34935 26019 34941
rect 25961 34932 25973 34935
rect 25924 34904 25973 34932
rect 25924 34892 25930 34904
rect 25961 34901 25973 34904
rect 26007 34901 26019 34935
rect 26528 34932 26556 34972
rect 27706 34960 27712 34972
rect 27764 34960 27770 35012
rect 27884 35003 27942 35009
rect 27884 34969 27896 35003
rect 27930 35000 27942 35003
rect 27982 35000 27988 35012
rect 27930 34972 27988 35000
rect 27930 34969 27942 34972
rect 27884 34963 27942 34969
rect 27982 34960 27988 34972
rect 28040 34960 28046 35012
rect 28276 35000 28304 35040
rect 29822 35028 29828 35040
rect 29880 35028 29886 35080
rect 29914 35028 29920 35080
rect 29972 35068 29978 35080
rect 30653 35071 30711 35077
rect 30653 35068 30665 35071
rect 29972 35040 30017 35068
rect 30116 35040 30665 35068
rect 29972 35028 29978 35040
rect 30116 35012 30144 35040
rect 30653 35037 30665 35040
rect 30699 35037 30711 35071
rect 30760 35068 30788 35108
rect 31726 35108 32689 35136
rect 30909 35071 30967 35077
rect 30909 35068 30921 35071
rect 30760 35040 30921 35068
rect 30653 35031 30711 35037
rect 30909 35037 30921 35040
rect 30955 35037 30967 35071
rect 30909 35031 30967 35037
rect 30098 35000 30104 35012
rect 28276 34972 30104 35000
rect 30098 34960 30104 34972
rect 30156 34960 30162 35012
rect 31726 35000 31754 35108
rect 32677 35105 32689 35108
rect 32723 35105 32735 35139
rect 32677 35099 32735 35105
rect 32122 35028 32128 35080
rect 32180 35068 32186 35080
rect 32493 35071 32551 35077
rect 32493 35068 32505 35071
rect 32180 35040 32505 35068
rect 32180 35028 32186 35040
rect 32493 35037 32505 35040
rect 32539 35037 32551 35071
rect 32493 35031 32551 35037
rect 30392 34972 31754 35000
rect 34333 35003 34391 35009
rect 27614 34932 27620 34944
rect 26528 34904 27620 34932
rect 25961 34895 26019 34901
rect 27614 34892 27620 34904
rect 27672 34892 27678 34944
rect 28258 34892 28264 34944
rect 28316 34932 28322 34944
rect 28810 34932 28816 34944
rect 28316 34904 28816 34932
rect 28316 34892 28322 34904
rect 28810 34892 28816 34904
rect 28868 34932 28874 34944
rect 28997 34935 29055 34941
rect 28997 34932 29009 34935
rect 28868 34904 29009 34932
rect 28868 34892 28874 34904
rect 28997 34901 29009 34904
rect 29043 34901 29055 34935
rect 28997 34895 29055 34901
rect 29362 34892 29368 34944
rect 29420 34932 29426 34944
rect 30392 34932 30420 34972
rect 34333 34969 34345 35003
rect 34379 35000 34391 35003
rect 34606 35000 34612 35012
rect 34379 34972 34612 35000
rect 34379 34969 34391 34972
rect 34333 34963 34391 34969
rect 34606 34960 34612 34972
rect 34664 34960 34670 35012
rect 29420 34904 30420 34932
rect 29420 34892 29426 34904
rect 31662 34892 31668 34944
rect 31720 34932 31726 34944
rect 32030 34932 32036 34944
rect 31720 34904 32036 34932
rect 31720 34892 31726 34904
rect 32030 34892 32036 34904
rect 32088 34892 32094 34944
rect 1104 34842 35027 34864
rect 1104 34790 9390 34842
rect 9442 34790 9454 34842
rect 9506 34790 9518 34842
rect 9570 34790 9582 34842
rect 9634 34790 9646 34842
rect 9698 34790 17831 34842
rect 17883 34790 17895 34842
rect 17947 34790 17959 34842
rect 18011 34790 18023 34842
rect 18075 34790 18087 34842
rect 18139 34790 26272 34842
rect 26324 34790 26336 34842
rect 26388 34790 26400 34842
rect 26452 34790 26464 34842
rect 26516 34790 26528 34842
rect 26580 34790 34713 34842
rect 34765 34790 34777 34842
rect 34829 34790 34841 34842
rect 34893 34790 34905 34842
rect 34957 34790 34969 34842
rect 35021 34790 35027 34842
rect 1104 34768 35027 34790
rect 17126 34688 17132 34740
rect 17184 34728 17190 34740
rect 18785 34731 18843 34737
rect 17184 34700 18736 34728
rect 17184 34688 17190 34700
rect 18230 34660 18236 34672
rect 17420 34632 18236 34660
rect 1762 34592 1768 34604
rect 1723 34564 1768 34592
rect 1762 34552 1768 34564
rect 1820 34552 1826 34604
rect 17420 34601 17448 34632
rect 18230 34620 18236 34632
rect 18288 34620 18294 34672
rect 18708 34660 18736 34700
rect 18785 34697 18797 34731
rect 18831 34728 18843 34731
rect 20254 34728 20260 34740
rect 18831 34700 20260 34728
rect 18831 34697 18843 34700
rect 18785 34691 18843 34697
rect 20254 34688 20260 34700
rect 20312 34688 20318 34740
rect 20622 34728 20628 34740
rect 20583 34700 20628 34728
rect 20622 34688 20628 34700
rect 20680 34688 20686 34740
rect 20714 34688 20720 34740
rect 20772 34728 20778 34740
rect 21453 34731 21511 34737
rect 21453 34728 21465 34731
rect 20772 34700 21465 34728
rect 20772 34688 20778 34700
rect 21453 34697 21465 34700
rect 21499 34697 21511 34731
rect 21453 34691 21511 34697
rect 22646 34688 22652 34740
rect 22704 34728 22710 34740
rect 23290 34728 23296 34740
rect 22704 34700 23296 34728
rect 22704 34688 22710 34700
rect 23290 34688 23296 34700
rect 23348 34728 23354 34740
rect 23385 34731 23443 34737
rect 23385 34728 23397 34731
rect 23348 34700 23397 34728
rect 23348 34688 23354 34700
rect 23385 34697 23397 34700
rect 23431 34697 23443 34731
rect 23385 34691 23443 34697
rect 23934 34688 23940 34740
rect 23992 34728 23998 34740
rect 24578 34728 24584 34740
rect 23992 34700 24584 34728
rect 23992 34688 23998 34700
rect 24578 34688 24584 34700
rect 24636 34688 24642 34740
rect 25406 34688 25412 34740
rect 25464 34728 25470 34740
rect 28534 34728 28540 34740
rect 25464 34700 28028 34728
rect 28495 34700 28540 34728
rect 25464 34688 25470 34700
rect 19334 34660 19340 34672
rect 18708 34632 19340 34660
rect 19334 34620 19340 34632
rect 19392 34620 19398 34672
rect 19512 34663 19570 34669
rect 19512 34629 19524 34663
rect 19558 34660 19570 34663
rect 19978 34660 19984 34672
rect 19558 34632 19984 34660
rect 19558 34629 19570 34632
rect 19512 34623 19570 34629
rect 19978 34620 19984 34632
rect 20036 34620 20042 34672
rect 20272 34660 20300 34688
rect 20272 34632 20392 34660
rect 17405 34595 17463 34601
rect 17405 34561 17417 34595
rect 17451 34561 17463 34595
rect 17405 34555 17463 34561
rect 17672 34595 17730 34601
rect 17672 34561 17684 34595
rect 17718 34592 17730 34595
rect 18690 34592 18696 34604
rect 17718 34564 18696 34592
rect 17718 34561 17730 34564
rect 17672 34555 17730 34561
rect 18690 34552 18696 34564
rect 18748 34552 18754 34604
rect 19242 34592 19248 34604
rect 19203 34564 19248 34592
rect 19242 34552 19248 34564
rect 19300 34552 19306 34604
rect 20364 34592 20392 34632
rect 22020 34632 23428 34660
rect 21085 34595 21143 34601
rect 21085 34592 21097 34595
rect 20364 34564 21097 34592
rect 21085 34561 21097 34564
rect 21131 34561 21143 34595
rect 21266 34592 21272 34604
rect 21227 34564 21272 34592
rect 21085 34555 21143 34561
rect 21266 34552 21272 34564
rect 21324 34592 21330 34604
rect 21450 34592 21456 34604
rect 21324 34564 21456 34592
rect 21324 34552 21330 34564
rect 21450 34552 21456 34564
rect 21508 34552 21514 34604
rect 21726 34552 21732 34604
rect 21784 34592 21790 34604
rect 22020 34601 22048 34632
rect 23400 34604 23428 34632
rect 23658 34620 23664 34672
rect 23716 34660 23722 34672
rect 24090 34663 24148 34669
rect 24090 34660 24102 34663
rect 23716 34632 24102 34660
rect 23716 34620 23722 34632
rect 24090 34629 24102 34632
rect 24136 34629 24148 34663
rect 24090 34623 24148 34629
rect 24210 34620 24216 34672
rect 24268 34660 24274 34672
rect 26053 34663 26111 34669
rect 26053 34660 26065 34663
rect 24268 34632 26065 34660
rect 24268 34620 24274 34632
rect 26053 34629 26065 34632
rect 26099 34629 26111 34663
rect 26053 34623 26111 34629
rect 26970 34620 26976 34672
rect 27028 34660 27034 34672
rect 27402 34663 27460 34669
rect 27402 34660 27414 34663
rect 27028 34632 27414 34660
rect 27028 34620 27034 34632
rect 27402 34629 27414 34632
rect 27448 34629 27460 34663
rect 27402 34623 27460 34629
rect 22005 34595 22063 34601
rect 22005 34592 22017 34595
rect 21784 34564 22017 34592
rect 21784 34552 21790 34564
rect 22005 34561 22017 34564
rect 22051 34561 22063 34595
rect 22005 34555 22063 34561
rect 22272 34595 22330 34601
rect 22272 34561 22284 34595
rect 22318 34592 22330 34595
rect 22554 34592 22560 34604
rect 22318 34564 22560 34592
rect 22318 34561 22330 34564
rect 22272 34555 22330 34561
rect 22554 34552 22560 34564
rect 22612 34552 22618 34604
rect 23382 34552 23388 34604
rect 23440 34592 23446 34604
rect 23845 34595 23903 34601
rect 23845 34592 23857 34595
rect 23440 34564 23857 34592
rect 23440 34552 23446 34564
rect 23845 34561 23857 34564
rect 23891 34592 23903 34595
rect 23934 34592 23940 34604
rect 23891 34564 23940 34592
rect 23891 34561 23903 34564
rect 23845 34555 23903 34561
rect 23934 34552 23940 34564
rect 23992 34552 23998 34604
rect 24394 34552 24400 34604
rect 24452 34592 24458 34604
rect 25685 34595 25743 34601
rect 25685 34592 25697 34595
rect 24452 34564 25697 34592
rect 24452 34552 24458 34564
rect 25685 34561 25697 34564
rect 25731 34561 25743 34595
rect 25685 34555 25743 34561
rect 25774 34552 25780 34604
rect 25832 34592 25838 34604
rect 25869 34595 25927 34601
rect 25869 34592 25881 34595
rect 25832 34564 25881 34592
rect 25832 34552 25838 34564
rect 25869 34561 25881 34564
rect 25915 34561 25927 34595
rect 28000 34592 28028 34700
rect 28534 34688 28540 34700
rect 28592 34688 28598 34740
rect 29270 34688 29276 34740
rect 29328 34728 29334 34740
rect 29457 34731 29515 34737
rect 29457 34728 29469 34731
rect 29328 34700 29469 34728
rect 29328 34688 29334 34700
rect 29457 34697 29469 34700
rect 29503 34697 29515 34731
rect 29457 34691 29515 34697
rect 29822 34688 29828 34740
rect 29880 34728 29886 34740
rect 31202 34728 31208 34740
rect 29880 34700 31208 34728
rect 29880 34688 29886 34700
rect 31202 34688 31208 34700
rect 31260 34688 31266 34740
rect 31294 34688 31300 34740
rect 31352 34728 31358 34740
rect 31573 34731 31631 34737
rect 31573 34728 31585 34731
rect 31352 34700 31585 34728
rect 31352 34688 31358 34700
rect 31573 34697 31585 34700
rect 31619 34728 31631 34731
rect 31754 34728 31760 34740
rect 31619 34700 31760 34728
rect 31619 34697 31631 34700
rect 31573 34691 31631 34697
rect 31754 34688 31760 34700
rect 31812 34688 31818 34740
rect 29914 34620 29920 34672
rect 29972 34660 29978 34672
rect 30098 34660 30104 34672
rect 29972 34632 30104 34660
rect 29972 34620 29978 34632
rect 30098 34620 30104 34632
rect 30156 34660 30162 34672
rect 30460 34663 30518 34669
rect 30156 34632 30236 34660
rect 30156 34620 30162 34632
rect 28000 34564 28212 34592
rect 25869 34555 25927 34561
rect 1946 34524 1952 34536
rect 1907 34496 1952 34524
rect 1946 34484 1952 34496
rect 2004 34484 2010 34536
rect 2774 34524 2780 34536
rect 2735 34496 2780 34524
rect 2774 34484 2780 34496
rect 2832 34484 2838 34536
rect 20990 34484 20996 34536
rect 21048 34524 21054 34536
rect 21744 34524 21772 34552
rect 21048 34496 21772 34524
rect 21048 34484 21054 34496
rect 26418 34484 26424 34536
rect 26476 34524 26482 34536
rect 27154 34524 27160 34536
rect 26476 34496 27160 34524
rect 26476 34484 26482 34496
rect 27154 34484 27160 34496
rect 27212 34484 27218 34536
rect 28184 34524 28212 34564
rect 28810 34552 28816 34604
rect 28868 34592 28874 34604
rect 29273 34595 29331 34601
rect 29273 34592 29285 34595
rect 28868 34564 29285 34592
rect 28868 34552 28874 34564
rect 29273 34561 29285 34564
rect 29319 34592 29331 34595
rect 30006 34592 30012 34604
rect 29319 34564 30012 34592
rect 29319 34561 29331 34564
rect 29273 34555 29331 34561
rect 30006 34552 30012 34564
rect 30064 34552 30070 34604
rect 30208 34601 30236 34632
rect 30460 34629 30472 34663
rect 30506 34660 30518 34663
rect 30558 34660 30564 34672
rect 30506 34632 30564 34660
rect 30506 34629 30518 34632
rect 30460 34623 30518 34629
rect 30558 34620 30564 34632
rect 30616 34620 30622 34672
rect 32677 34663 32735 34669
rect 32677 34660 32689 34663
rect 31726 34632 32689 34660
rect 30193 34595 30251 34601
rect 30193 34561 30205 34595
rect 30239 34561 30251 34595
rect 31726 34592 31754 34632
rect 32677 34629 32689 34632
rect 32723 34629 32735 34663
rect 34330 34660 34336 34672
rect 34291 34632 34336 34660
rect 32677 34623 32735 34629
rect 34330 34620 34336 34632
rect 34388 34620 34394 34672
rect 32490 34592 32496 34604
rect 30193 34555 30251 34561
rect 30300 34564 31754 34592
rect 32451 34564 32496 34592
rect 29089 34527 29147 34533
rect 28184 34496 29040 34524
rect 20530 34416 20536 34468
rect 20588 34456 20594 34468
rect 21818 34456 21824 34468
rect 20588 34428 21824 34456
rect 20588 34416 20594 34428
rect 21818 34416 21824 34428
rect 21876 34416 21882 34468
rect 23750 34456 23756 34468
rect 22940 34428 23756 34456
rect 16114 34348 16120 34400
rect 16172 34388 16178 34400
rect 21266 34388 21272 34400
rect 16172 34360 21272 34388
rect 16172 34348 16178 34360
rect 21266 34348 21272 34360
rect 21324 34348 21330 34400
rect 21542 34348 21548 34400
rect 21600 34388 21606 34400
rect 22940 34388 22968 34428
rect 23750 34416 23756 34428
rect 23808 34416 23814 34468
rect 25038 34416 25044 34468
rect 25096 34456 25102 34468
rect 25225 34459 25283 34465
rect 25225 34456 25237 34459
rect 25096 34428 25237 34456
rect 25096 34416 25102 34428
rect 25225 34425 25237 34428
rect 25271 34425 25283 34459
rect 29012 34456 29040 34496
rect 29089 34493 29101 34527
rect 29135 34524 29147 34527
rect 29362 34524 29368 34536
rect 29135 34496 29368 34524
rect 29135 34493 29147 34496
rect 29089 34487 29147 34493
rect 29362 34484 29368 34496
rect 29420 34484 29426 34536
rect 30300 34524 30328 34564
rect 32490 34552 32496 34564
rect 32548 34552 32554 34604
rect 29472 34496 30328 34524
rect 29472 34456 29500 34496
rect 29012 34428 29500 34456
rect 25225 34419 25283 34425
rect 21600 34360 22968 34388
rect 21600 34348 21606 34360
rect 23014 34348 23020 34400
rect 23072 34388 23078 34400
rect 29822 34388 29828 34400
rect 23072 34360 29828 34388
rect 23072 34348 23078 34360
rect 29822 34348 29828 34360
rect 29880 34348 29886 34400
rect 30098 34348 30104 34400
rect 30156 34388 30162 34400
rect 31570 34388 31576 34400
rect 30156 34360 31576 34388
rect 30156 34348 30162 34360
rect 31570 34348 31576 34360
rect 31628 34348 31634 34400
rect 1104 34298 34868 34320
rect 1104 34246 5170 34298
rect 5222 34246 5234 34298
rect 5286 34246 5298 34298
rect 5350 34246 5362 34298
rect 5414 34246 5426 34298
rect 5478 34246 13611 34298
rect 13663 34246 13675 34298
rect 13727 34246 13739 34298
rect 13791 34246 13803 34298
rect 13855 34246 13867 34298
rect 13919 34246 22052 34298
rect 22104 34246 22116 34298
rect 22168 34246 22180 34298
rect 22232 34246 22244 34298
rect 22296 34246 22308 34298
rect 22360 34246 30493 34298
rect 30545 34246 30557 34298
rect 30609 34246 30621 34298
rect 30673 34246 30685 34298
rect 30737 34246 30749 34298
rect 30801 34246 34868 34298
rect 1104 34224 34868 34246
rect 1857 34187 1915 34193
rect 1857 34153 1869 34187
rect 1903 34184 1915 34187
rect 1946 34184 1952 34196
rect 1903 34156 1952 34184
rect 1903 34153 1915 34156
rect 1857 34147 1915 34153
rect 1946 34144 1952 34156
rect 2004 34144 2010 34196
rect 18690 34184 18696 34196
rect 18651 34156 18696 34184
rect 18690 34144 18696 34156
rect 18748 34144 18754 34196
rect 21542 34184 21548 34196
rect 18800 34156 21548 34184
rect 4430 34048 4436 34060
rect 1780 34020 4436 34048
rect 1780 33989 1808 34020
rect 4430 34008 4436 34020
rect 4488 34008 4494 34060
rect 6546 34008 6552 34060
rect 6604 34048 6610 34060
rect 18800 34048 18828 34156
rect 21542 34144 21548 34156
rect 21600 34144 21606 34196
rect 21818 34144 21824 34196
rect 21876 34144 21882 34196
rect 22002 34144 22008 34196
rect 22060 34184 22066 34196
rect 22281 34187 22339 34193
rect 22060 34156 22232 34184
rect 22060 34144 22066 34156
rect 20806 34116 20812 34128
rect 20088 34088 20812 34116
rect 20088 34057 20116 34088
rect 20806 34076 20812 34088
rect 20864 34076 20870 34128
rect 21836 34116 21864 34144
rect 22204 34116 22232 34156
rect 22281 34153 22293 34187
rect 22327 34184 22339 34187
rect 22370 34184 22376 34196
rect 22327 34156 22376 34184
rect 22327 34153 22339 34156
rect 22281 34147 22339 34153
rect 22370 34144 22376 34156
rect 22428 34144 22434 34196
rect 25961 34187 26019 34193
rect 22480 34156 25912 34184
rect 22480 34116 22508 34156
rect 21836 34088 22094 34116
rect 22204 34088 22508 34116
rect 6604 34020 18828 34048
rect 20073 34051 20131 34057
rect 6604 34008 6610 34020
rect 20073 34017 20085 34051
rect 20119 34017 20131 34051
rect 20073 34011 20131 34017
rect 20165 34051 20223 34057
rect 20165 34017 20177 34051
rect 20211 34048 20223 34051
rect 22066 34048 22094 34088
rect 22646 34076 22652 34128
rect 22704 34116 22710 34128
rect 22833 34119 22891 34125
rect 22833 34116 22845 34119
rect 22704 34088 22845 34116
rect 22704 34076 22710 34088
rect 22833 34085 22845 34088
rect 22879 34085 22891 34119
rect 22833 34079 22891 34085
rect 23014 34048 23020 34060
rect 20211 34020 20852 34048
rect 22066 34020 23020 34048
rect 20211 34017 20223 34020
rect 20165 34011 20223 34017
rect 1765 33983 1823 33989
rect 1765 33949 1777 33983
rect 1811 33949 1823 33983
rect 2498 33980 2504 33992
rect 2459 33952 2504 33980
rect 1765 33943 1823 33949
rect 2498 33940 2504 33952
rect 2556 33940 2562 33992
rect 18141 33983 18199 33989
rect 18141 33949 18153 33983
rect 18187 33980 18199 33983
rect 18322 33980 18328 33992
rect 18187 33952 18328 33980
rect 18187 33949 18199 33952
rect 18141 33943 18199 33949
rect 18322 33940 18328 33952
rect 18380 33940 18386 33992
rect 18877 33983 18935 33989
rect 18877 33949 18889 33983
rect 18923 33980 18935 33983
rect 19794 33980 19800 33992
rect 18923 33952 19800 33980
rect 18923 33949 18935 33952
rect 18877 33943 18935 33949
rect 19794 33940 19800 33952
rect 19852 33940 19858 33992
rect 20257 33983 20315 33989
rect 20257 33949 20269 33983
rect 20303 33949 20315 33983
rect 20257 33943 20315 33949
rect 3050 33912 3056 33924
rect 3011 33884 3056 33912
rect 3050 33872 3056 33884
rect 3108 33912 3114 33924
rect 4890 33912 4896 33924
rect 3108 33884 4896 33912
rect 3108 33872 3114 33884
rect 4890 33872 4896 33884
rect 4948 33872 4954 33924
rect 17957 33847 18015 33853
rect 17957 33813 17969 33847
rect 18003 33844 18015 33847
rect 18414 33844 18420 33856
rect 18003 33816 18420 33844
rect 18003 33813 18015 33816
rect 17957 33807 18015 33813
rect 18414 33804 18420 33816
rect 18472 33804 18478 33856
rect 19794 33804 19800 33856
rect 19852 33844 19858 33856
rect 19889 33847 19947 33853
rect 19889 33844 19901 33847
rect 19852 33816 19901 33844
rect 19852 33804 19858 33816
rect 19889 33813 19901 33816
rect 19935 33813 19947 33847
rect 19889 33807 19947 33813
rect 20070 33804 20076 33856
rect 20128 33844 20134 33856
rect 20272 33844 20300 33943
rect 20346 33940 20352 33992
rect 20404 33980 20410 33992
rect 20404 33952 20449 33980
rect 20404 33940 20410 33952
rect 20128 33816 20300 33844
rect 20824 33844 20852 34020
rect 23014 34008 23020 34020
rect 23072 34008 23078 34060
rect 20901 33983 20959 33989
rect 20901 33949 20913 33983
rect 20947 33980 20959 33983
rect 20990 33980 20996 33992
rect 20947 33952 20996 33980
rect 20947 33949 20959 33952
rect 20901 33943 20959 33949
rect 20990 33940 20996 33952
rect 21048 33940 21054 33992
rect 21168 33983 21226 33989
rect 21168 33949 21180 33983
rect 21214 33949 21226 33983
rect 24029 33983 24087 33989
rect 21168 33943 21226 33949
rect 22204 33952 23428 33980
rect 21082 33872 21088 33924
rect 21140 33912 21146 33924
rect 21192 33912 21220 33943
rect 21140 33884 21220 33912
rect 21140 33872 21146 33884
rect 21266 33872 21272 33924
rect 21324 33912 21330 33924
rect 22002 33912 22008 33924
rect 21324 33884 22008 33912
rect 21324 33872 21330 33884
rect 22002 33872 22008 33884
rect 22060 33872 22066 33924
rect 22204 33844 22232 33952
rect 23106 33912 23112 33924
rect 23067 33884 23112 33912
rect 23106 33872 23112 33884
rect 23164 33872 23170 33924
rect 23400 33921 23428 33952
rect 24029 33949 24041 33983
rect 24075 33980 24087 33983
rect 24210 33980 24216 33992
rect 24075 33952 24216 33980
rect 24075 33949 24087 33952
rect 24029 33943 24087 33949
rect 24210 33940 24216 33952
rect 24268 33940 24274 33992
rect 24578 33980 24584 33992
rect 24539 33952 24584 33980
rect 24578 33940 24584 33952
rect 24636 33940 24642 33992
rect 24670 33940 24676 33992
rect 24728 33980 24734 33992
rect 24837 33983 24895 33989
rect 24837 33980 24849 33983
rect 24728 33952 24849 33980
rect 24728 33940 24734 33952
rect 24837 33949 24849 33952
rect 24883 33949 24895 33983
rect 24837 33943 24895 33949
rect 23385 33915 23443 33921
rect 23385 33881 23397 33915
rect 23431 33881 23443 33915
rect 23566 33912 23572 33924
rect 23385 33875 23443 33881
rect 23483 33884 23572 33912
rect 20824 33816 22232 33844
rect 20128 33804 20134 33816
rect 22922 33804 22928 33856
rect 22980 33844 22986 33856
rect 23017 33847 23075 33853
rect 23017 33844 23029 33847
rect 22980 33816 23029 33844
rect 22980 33804 22986 33816
rect 23017 33813 23029 33816
rect 23063 33813 23075 33847
rect 23017 33807 23075 33813
rect 23201 33847 23259 33853
rect 23201 33813 23213 33847
rect 23247 33844 23259 33847
rect 23483 33844 23511 33884
rect 23566 33872 23572 33884
rect 23624 33912 23630 33924
rect 25038 33912 25044 33924
rect 23624 33884 25044 33912
rect 23624 33872 23630 33884
rect 25038 33872 25044 33884
rect 25096 33872 25102 33924
rect 23842 33844 23848 33856
rect 23247 33816 23511 33844
rect 23803 33816 23848 33844
rect 23247 33813 23259 33816
rect 23201 33807 23259 33813
rect 23842 33804 23848 33816
rect 23900 33804 23906 33856
rect 25884 33844 25912 34156
rect 25961 34153 25973 34187
rect 26007 34184 26019 34187
rect 26602 34184 26608 34196
rect 26007 34156 26608 34184
rect 26007 34153 26019 34156
rect 25961 34147 26019 34153
rect 26602 34144 26608 34156
rect 26660 34144 26666 34196
rect 27430 34144 27436 34196
rect 27488 34184 27494 34196
rect 28813 34187 28871 34193
rect 28813 34184 28825 34187
rect 27488 34156 28825 34184
rect 27488 34144 27494 34156
rect 28813 34153 28825 34156
rect 28859 34153 28871 34187
rect 30098 34184 30104 34196
rect 28813 34147 28871 34153
rect 28966 34156 30104 34184
rect 27614 34076 27620 34128
rect 27672 34116 27678 34128
rect 28966 34116 28994 34156
rect 30098 34144 30104 34156
rect 30156 34144 30162 34196
rect 31110 34184 31116 34196
rect 31071 34156 31116 34184
rect 31110 34144 31116 34156
rect 31168 34144 31174 34196
rect 31665 34187 31723 34193
rect 31665 34153 31677 34187
rect 31711 34153 31723 34187
rect 31665 34147 31723 34153
rect 27672 34088 28994 34116
rect 27672 34076 27678 34088
rect 29086 34076 29092 34128
rect 29144 34116 29150 34128
rect 29144 34088 29592 34116
rect 29144 34076 29150 34088
rect 26418 34048 26424 34060
rect 26379 34020 26424 34048
rect 26418 34008 26424 34020
rect 26476 34008 26482 34060
rect 29454 34048 29460 34060
rect 27448 34020 29460 34048
rect 27448 33980 27476 34020
rect 29454 34008 29460 34020
rect 29512 34008 29518 34060
rect 27264 33952 27476 33980
rect 25958 33872 25964 33924
rect 26016 33912 26022 33924
rect 26666 33915 26724 33921
rect 26666 33912 26678 33915
rect 26016 33884 26678 33912
rect 26016 33872 26022 33884
rect 26666 33881 26678 33884
rect 26712 33881 26724 33915
rect 27264 33912 27292 33952
rect 28074 33940 28080 33992
rect 28132 33980 28138 33992
rect 28445 33983 28503 33989
rect 28445 33980 28457 33983
rect 28132 33952 28457 33980
rect 28132 33940 28138 33952
rect 28445 33949 28457 33952
rect 28491 33949 28503 33983
rect 28445 33943 28503 33949
rect 28534 33940 28540 33992
rect 28592 33980 28598 33992
rect 28592 33952 29500 33980
rect 28592 33940 28598 33952
rect 26666 33875 26724 33881
rect 26804 33884 27292 33912
rect 26804 33844 26832 33884
rect 27338 33872 27344 33924
rect 27396 33912 27402 33924
rect 28258 33912 28264 33924
rect 27396 33884 28120 33912
rect 28219 33884 28264 33912
rect 27396 33872 27402 33884
rect 25884 33816 26832 33844
rect 27062 33804 27068 33856
rect 27120 33844 27126 33856
rect 27430 33844 27436 33856
rect 27120 33816 27436 33844
rect 27120 33804 27126 33816
rect 27430 33804 27436 33816
rect 27488 33844 27494 33856
rect 27801 33847 27859 33853
rect 27801 33844 27813 33847
rect 27488 33816 27813 33844
rect 27488 33804 27494 33816
rect 27801 33813 27813 33816
rect 27847 33813 27859 33847
rect 28092 33844 28120 33884
rect 28258 33872 28264 33884
rect 28316 33872 28322 33924
rect 29086 33912 29092 33924
rect 28368 33884 29092 33912
rect 28368 33844 28396 33884
rect 29086 33872 29092 33884
rect 29144 33872 29150 33924
rect 28534 33844 28540 33856
rect 28092 33816 28396 33844
rect 28495 33816 28540 33844
rect 27801 33807 27859 33813
rect 28534 33804 28540 33816
rect 28592 33804 28598 33856
rect 28626 33804 28632 33856
rect 28684 33844 28690 33856
rect 29178 33844 29184 33856
rect 28684 33816 29184 33844
rect 28684 33804 28690 33816
rect 29178 33804 29184 33816
rect 29236 33804 29242 33856
rect 29472 33844 29500 33952
rect 29564 33912 29592 34088
rect 29730 34076 29736 34128
rect 29788 34076 29794 34128
rect 31570 34076 31576 34128
rect 31628 34116 31634 34128
rect 31680 34116 31708 34147
rect 31628 34088 31708 34116
rect 31628 34076 31634 34088
rect 29748 34048 29776 34076
rect 29748 34020 29868 34048
rect 29730 33980 29736 33992
rect 29691 33952 29736 33980
rect 29730 33940 29736 33952
rect 29788 33940 29794 33992
rect 29840 33980 29868 34020
rect 31294 34008 31300 34060
rect 31352 34048 31358 34060
rect 31665 34051 31723 34057
rect 31665 34048 31677 34051
rect 31352 34020 31677 34048
rect 31352 34008 31358 34020
rect 31665 34017 31677 34020
rect 31711 34017 31723 34051
rect 31665 34011 31723 34017
rect 31754 34008 31760 34060
rect 31812 34048 31818 34060
rect 31812 34020 31892 34048
rect 31812 34008 31818 34020
rect 29989 33983 30047 33989
rect 29989 33980 30001 33983
rect 29840 33952 30001 33980
rect 29989 33949 30001 33952
rect 30035 33949 30047 33983
rect 29989 33943 30047 33949
rect 30926 33940 30932 33992
rect 30984 33980 30990 33992
rect 31110 33980 31116 33992
rect 30984 33952 31116 33980
rect 30984 33940 30990 33952
rect 31110 33940 31116 33952
rect 31168 33980 31174 33992
rect 31864 33989 31892 34020
rect 32030 34008 32036 34060
rect 32088 34048 32094 34060
rect 32493 34051 32551 34057
rect 32493 34048 32505 34051
rect 32088 34020 32505 34048
rect 32088 34008 32094 34020
rect 32493 34017 32505 34020
rect 32539 34017 32551 34051
rect 32493 34011 32551 34017
rect 31573 33983 31631 33989
rect 31573 33980 31585 33983
rect 31168 33952 31585 33980
rect 31168 33940 31174 33952
rect 31573 33949 31585 33952
rect 31619 33949 31631 33983
rect 31573 33943 31631 33949
rect 31849 33983 31907 33989
rect 31849 33949 31861 33983
rect 31895 33949 31907 33983
rect 31849 33943 31907 33949
rect 30098 33912 30104 33924
rect 29564 33884 30104 33912
rect 30098 33872 30104 33884
rect 30156 33872 30162 33924
rect 30834 33872 30840 33924
rect 30892 33912 30898 33924
rect 31864 33912 31892 33943
rect 30892 33884 31892 33912
rect 30892 33872 30898 33884
rect 32122 33872 32128 33924
rect 32180 33912 32186 33924
rect 32677 33915 32735 33921
rect 32677 33912 32689 33915
rect 32180 33884 32689 33912
rect 32180 33872 32186 33884
rect 32677 33881 32689 33884
rect 32723 33881 32735 33915
rect 34330 33912 34336 33924
rect 34291 33884 34336 33912
rect 32677 33875 32735 33881
rect 34330 33872 34336 33884
rect 34388 33872 34394 33924
rect 30558 33844 30564 33856
rect 29472 33816 30564 33844
rect 30558 33804 30564 33816
rect 30616 33804 30622 33856
rect 31938 33804 31944 33856
rect 31996 33844 32002 33856
rect 32033 33847 32091 33853
rect 32033 33844 32045 33847
rect 31996 33816 32045 33844
rect 31996 33804 32002 33816
rect 32033 33813 32045 33816
rect 32079 33813 32091 33847
rect 32033 33807 32091 33813
rect 1104 33754 35027 33776
rect 1104 33702 9390 33754
rect 9442 33702 9454 33754
rect 9506 33702 9518 33754
rect 9570 33702 9582 33754
rect 9634 33702 9646 33754
rect 9698 33702 17831 33754
rect 17883 33702 17895 33754
rect 17947 33702 17959 33754
rect 18011 33702 18023 33754
rect 18075 33702 18087 33754
rect 18139 33702 26272 33754
rect 26324 33702 26336 33754
rect 26388 33702 26400 33754
rect 26452 33702 26464 33754
rect 26516 33702 26528 33754
rect 26580 33702 34713 33754
rect 34765 33702 34777 33754
rect 34829 33702 34841 33754
rect 34893 33702 34905 33754
rect 34957 33702 34969 33754
rect 35021 33702 35027 33754
rect 1104 33680 35027 33702
rect 2130 33640 2136 33652
rect 2091 33612 2136 33640
rect 2130 33600 2136 33612
rect 2188 33600 2194 33652
rect 19058 33600 19064 33652
rect 19116 33640 19122 33652
rect 19978 33640 19984 33652
rect 19116 33612 19984 33640
rect 19116 33600 19122 33612
rect 19978 33600 19984 33612
rect 20036 33600 20042 33652
rect 20165 33643 20223 33649
rect 20165 33609 20177 33643
rect 20211 33640 20223 33643
rect 20346 33640 20352 33652
rect 20211 33612 20352 33640
rect 20211 33609 20223 33612
rect 20165 33603 20223 33609
rect 20346 33600 20352 33612
rect 20404 33600 20410 33652
rect 21361 33643 21419 33649
rect 21361 33609 21373 33643
rect 21407 33640 21419 33643
rect 21450 33640 21456 33652
rect 21407 33612 21456 33640
rect 21407 33609 21419 33612
rect 21361 33603 21419 33609
rect 21450 33600 21456 33612
rect 21508 33600 21514 33652
rect 21726 33600 21732 33652
rect 21784 33640 21790 33652
rect 31294 33640 31300 33652
rect 21784 33612 29868 33640
rect 31255 33612 31300 33640
rect 21784 33600 21790 33612
rect 3234 33572 3240 33584
rect 2332 33544 3240 33572
rect 2332 33516 2360 33544
rect 3234 33532 3240 33544
rect 3292 33532 3298 33584
rect 16206 33532 16212 33584
rect 16264 33572 16270 33584
rect 22272 33575 22330 33581
rect 16264 33544 22232 33572
rect 16264 33532 16270 33544
rect 2041 33507 2099 33513
rect 2041 33473 2053 33507
rect 2087 33504 2099 33507
rect 2314 33504 2320 33516
rect 2087 33476 2320 33504
rect 2087 33473 2099 33476
rect 2041 33467 2099 33473
rect 2314 33464 2320 33476
rect 2372 33464 2378 33516
rect 2866 33504 2872 33516
rect 2827 33476 2872 33504
rect 2866 33464 2872 33476
rect 2924 33464 2930 33516
rect 18141 33507 18199 33513
rect 18141 33473 18153 33507
rect 18187 33504 18199 33507
rect 18230 33504 18236 33516
rect 18187 33476 18236 33504
rect 18187 33473 18199 33476
rect 18141 33467 18199 33473
rect 18230 33464 18236 33476
rect 18288 33464 18294 33516
rect 18414 33513 18420 33516
rect 18408 33504 18420 33513
rect 18375 33476 18420 33504
rect 18408 33467 18420 33476
rect 18414 33464 18420 33467
rect 18472 33464 18478 33516
rect 18966 33464 18972 33516
rect 19024 33504 19030 33516
rect 19024 33476 19932 33504
rect 19024 33464 19030 33476
rect 19518 33300 19524 33312
rect 19479 33272 19524 33300
rect 19518 33260 19524 33272
rect 19576 33260 19582 33312
rect 19904 33300 19932 33476
rect 20254 33464 20260 33516
rect 20312 33504 20318 33516
rect 20349 33507 20407 33513
rect 20349 33504 20361 33507
rect 20312 33476 20361 33504
rect 20312 33464 20318 33476
rect 20349 33473 20361 33476
rect 20395 33473 20407 33507
rect 20349 33467 20407 33473
rect 20438 33464 20444 33516
rect 20496 33504 20502 33516
rect 20496 33476 20541 33504
rect 20496 33464 20502 33476
rect 20622 33464 20628 33516
rect 20680 33504 20686 33516
rect 21266 33504 21272 33516
rect 20680 33476 20725 33504
rect 21227 33476 21272 33504
rect 20680 33464 20686 33476
rect 21266 33464 21272 33476
rect 21324 33464 21330 33516
rect 21818 33464 21824 33516
rect 21876 33504 21882 33516
rect 22005 33507 22063 33513
rect 22005 33504 22017 33507
rect 21876 33476 22017 33504
rect 21876 33464 21882 33476
rect 22005 33473 22017 33476
rect 22051 33473 22063 33507
rect 22204 33504 22232 33544
rect 22272 33541 22284 33575
rect 22318 33572 22330 33575
rect 22462 33572 22468 33584
rect 22318 33544 22468 33572
rect 22318 33541 22330 33544
rect 22272 33535 22330 33541
rect 22462 33532 22468 33544
rect 22520 33532 22526 33584
rect 24756 33575 24814 33581
rect 22572 33544 24164 33572
rect 22572 33504 22600 33544
rect 24026 33504 24032 33516
rect 22204 33476 22600 33504
rect 23987 33476 24032 33504
rect 22005 33467 22063 33473
rect 24026 33464 24032 33476
rect 24084 33464 24090 33516
rect 24136 33504 24164 33544
rect 24756 33541 24768 33575
rect 24802 33572 24814 33575
rect 25682 33572 25688 33584
rect 24802 33544 25688 33572
rect 24802 33541 24814 33544
rect 24756 33535 24814 33541
rect 25682 33532 25688 33544
rect 25740 33532 25746 33584
rect 25774 33532 25780 33584
rect 25832 33572 25838 33584
rect 26605 33575 26663 33581
rect 26605 33572 26617 33575
rect 25832 33544 26617 33572
rect 25832 33532 25838 33544
rect 26605 33541 26617 33544
rect 26651 33541 26663 33575
rect 29730 33572 29736 33584
rect 26605 33535 26663 33541
rect 27816 33544 29736 33572
rect 26421 33507 26479 33513
rect 24136 33476 25544 33504
rect 20533 33439 20591 33445
rect 20533 33405 20545 33439
rect 20579 33436 20591 33439
rect 21634 33436 21640 33448
rect 20579 33408 21640 33436
rect 20579 33405 20591 33408
rect 20533 33399 20591 33405
rect 21634 33396 21640 33408
rect 21692 33396 21698 33448
rect 24486 33436 24492 33448
rect 24447 33408 24492 33436
rect 24486 33396 24492 33408
rect 24544 33396 24550 33448
rect 25516 33436 25544 33476
rect 26421 33473 26433 33507
rect 26467 33504 26479 33507
rect 26694 33504 26700 33516
rect 26467 33476 26700 33504
rect 26467 33473 26479 33476
rect 26421 33467 26479 33473
rect 26694 33464 26700 33476
rect 26752 33464 26758 33516
rect 27338 33504 27344 33516
rect 27299 33476 27344 33504
rect 27338 33464 27344 33476
rect 27396 33464 27402 33516
rect 27816 33513 27844 33544
rect 29730 33532 29736 33544
rect 29788 33532 29794 33584
rect 29840 33572 29868 33612
rect 31294 33600 31300 33612
rect 31352 33600 31358 33652
rect 30162 33575 30220 33581
rect 30162 33572 30174 33575
rect 29840 33544 30174 33572
rect 30162 33541 30174 33544
rect 30208 33541 30220 33575
rect 30162 33535 30220 33541
rect 30558 33532 30564 33584
rect 30616 33572 30622 33584
rect 32122 33572 32128 33584
rect 30616 33544 32128 33572
rect 30616 33532 30622 33544
rect 32122 33532 32128 33544
rect 32180 33532 32186 33584
rect 32306 33532 32312 33584
rect 32364 33572 32370 33584
rect 32677 33575 32735 33581
rect 32677 33572 32689 33575
rect 32364 33544 32689 33572
rect 32364 33532 32370 33544
rect 32677 33541 32689 33544
rect 32723 33541 32735 33575
rect 32677 33535 32735 33541
rect 34333 33575 34391 33581
rect 34333 33541 34345 33575
rect 34379 33572 34391 33575
rect 34422 33572 34428 33584
rect 34379 33544 34428 33572
rect 34379 33541 34391 33544
rect 34333 33535 34391 33541
rect 34422 33532 34428 33544
rect 34480 33532 34486 33584
rect 27801 33507 27859 33513
rect 27801 33473 27813 33507
rect 27847 33473 27859 33507
rect 27801 33467 27859 33473
rect 28068 33507 28126 33513
rect 28068 33473 28080 33507
rect 28114 33504 28126 33507
rect 29270 33504 29276 33516
rect 28114 33476 29276 33504
rect 28114 33473 28126 33476
rect 28068 33467 28126 33473
rect 29270 33464 29276 33476
rect 29328 33464 29334 33516
rect 29454 33464 29460 33516
rect 29512 33504 29518 33516
rect 32493 33507 32551 33513
rect 32493 33504 32505 33507
rect 29512 33476 32505 33504
rect 29512 33464 29518 33476
rect 32493 33473 32505 33476
rect 32539 33473 32551 33507
rect 32493 33467 32551 33473
rect 27614 33436 27620 33448
rect 25516 33408 27620 33436
rect 27614 33396 27620 33408
rect 27672 33396 27678 33448
rect 29914 33436 29920 33448
rect 29875 33408 29920 33436
rect 29914 33396 29920 33408
rect 29972 33396 29978 33448
rect 29270 33368 29276 33380
rect 23216 33340 23980 33368
rect 23216 33300 23244 33340
rect 19904 33272 23244 33300
rect 23290 33260 23296 33312
rect 23348 33300 23354 33312
rect 23385 33303 23443 33309
rect 23385 33300 23397 33303
rect 23348 33272 23397 33300
rect 23348 33260 23354 33272
rect 23385 33269 23397 33272
rect 23431 33269 23443 33303
rect 23385 33263 23443 33269
rect 23474 33260 23480 33312
rect 23532 33300 23538 33312
rect 23845 33303 23903 33309
rect 23845 33300 23857 33303
rect 23532 33272 23857 33300
rect 23532 33260 23538 33272
rect 23845 33269 23857 33272
rect 23891 33269 23903 33303
rect 23952 33300 23980 33340
rect 25792 33340 27292 33368
rect 25792 33300 25820 33340
rect 23952 33272 25820 33300
rect 25869 33303 25927 33309
rect 23845 33263 23903 33269
rect 25869 33269 25881 33303
rect 25915 33300 25927 33303
rect 26602 33300 26608 33312
rect 25915 33272 26608 33300
rect 25915 33269 25927 33272
rect 25869 33263 25927 33269
rect 26602 33260 26608 33272
rect 26660 33260 26666 33312
rect 26694 33260 26700 33312
rect 26752 33300 26758 33312
rect 27157 33303 27215 33309
rect 27157 33300 27169 33303
rect 26752 33272 27169 33300
rect 26752 33260 26758 33272
rect 27157 33269 27169 33272
rect 27203 33269 27215 33303
rect 27264 33300 27292 33340
rect 28736 33340 29276 33368
rect 28736 33300 28764 33340
rect 29270 33328 29276 33340
rect 29328 33328 29334 33380
rect 29178 33300 29184 33312
rect 27264 33272 28764 33300
rect 29139 33272 29184 33300
rect 27157 33263 27215 33269
rect 29178 33260 29184 33272
rect 29236 33260 29242 33312
rect 29822 33260 29828 33312
rect 29880 33300 29886 33312
rect 32674 33300 32680 33312
rect 29880 33272 32680 33300
rect 29880 33260 29886 33272
rect 32674 33260 32680 33272
rect 32732 33260 32738 33312
rect 1104 33210 34868 33232
rect 1104 33158 5170 33210
rect 5222 33158 5234 33210
rect 5286 33158 5298 33210
rect 5350 33158 5362 33210
rect 5414 33158 5426 33210
rect 5478 33158 13611 33210
rect 13663 33158 13675 33210
rect 13727 33158 13739 33210
rect 13791 33158 13803 33210
rect 13855 33158 13867 33210
rect 13919 33158 22052 33210
rect 22104 33158 22116 33210
rect 22168 33158 22180 33210
rect 22232 33158 22244 33210
rect 22296 33158 22308 33210
rect 22360 33158 30493 33210
rect 30545 33158 30557 33210
rect 30609 33158 30621 33210
rect 30673 33158 30685 33210
rect 30737 33158 30749 33210
rect 30801 33158 34868 33210
rect 1104 33136 34868 33158
rect 1581 33099 1639 33105
rect 1581 33065 1593 33099
rect 1627 33096 1639 33099
rect 1670 33096 1676 33108
rect 1627 33068 1676 33096
rect 1627 33065 1639 33068
rect 1581 33059 1639 33065
rect 1670 33056 1676 33068
rect 1728 33056 1734 33108
rect 18693 33099 18751 33105
rect 18693 33065 18705 33099
rect 18739 33096 18751 33099
rect 19702 33096 19708 33108
rect 18739 33068 19708 33096
rect 18739 33065 18751 33068
rect 18693 33059 18751 33065
rect 19702 33056 19708 33068
rect 19760 33096 19766 33108
rect 20622 33096 20628 33108
rect 19760 33068 20628 33096
rect 19760 33056 19766 33068
rect 20622 33056 20628 33068
rect 20680 33056 20686 33108
rect 21729 33099 21787 33105
rect 21729 33065 21741 33099
rect 21775 33096 21787 33099
rect 21910 33096 21916 33108
rect 21775 33068 21916 33096
rect 21775 33065 21787 33068
rect 21729 33059 21787 33065
rect 21910 33056 21916 33068
rect 21968 33056 21974 33108
rect 23109 33099 23167 33105
rect 23109 33065 23121 33099
rect 23155 33096 23167 33099
rect 24026 33096 24032 33108
rect 23155 33068 24032 33096
rect 23155 33065 23167 33068
rect 23109 33059 23167 33065
rect 24026 33056 24032 33068
rect 24084 33056 24090 33108
rect 26142 33056 26148 33108
rect 26200 33096 26206 33108
rect 26200 33068 28764 33096
rect 26200 33056 26206 33068
rect 13446 32988 13452 33040
rect 13504 33028 13510 33040
rect 19426 33028 19432 33040
rect 13504 33000 19432 33028
rect 13504 32988 13510 33000
rect 19426 32988 19432 33000
rect 19484 32988 19490 33040
rect 25041 33031 25099 33037
rect 25041 33028 25053 33031
rect 20548 33000 25053 33028
rect 18414 32920 18420 32972
rect 18472 32960 18478 32972
rect 19242 32960 19248 32972
rect 18472 32932 19248 32960
rect 18472 32920 18478 32932
rect 19242 32920 19248 32932
rect 19300 32960 19306 32972
rect 19521 32963 19579 32969
rect 19521 32960 19533 32963
rect 19300 32932 19533 32960
rect 19300 32920 19306 32932
rect 19521 32929 19533 32932
rect 19567 32929 19579 32963
rect 19521 32923 19579 32929
rect 1765 32895 1823 32901
rect 1765 32861 1777 32895
rect 1811 32892 1823 32895
rect 2958 32892 2964 32904
rect 1811 32864 2964 32892
rect 1811 32861 1823 32864
rect 1765 32855 1823 32861
rect 2958 32852 2964 32864
rect 3016 32852 3022 32904
rect 18874 32892 18880 32904
rect 18835 32864 18880 32892
rect 18874 32852 18880 32864
rect 18932 32852 18938 32904
rect 19794 32901 19800 32904
rect 19788 32892 19800 32901
rect 19755 32864 19800 32892
rect 19788 32855 19800 32864
rect 19794 32852 19800 32855
rect 19852 32852 19858 32904
rect 20548 32824 20576 33000
rect 25041 32997 25053 33000
rect 25087 32997 25099 33031
rect 28736 33028 28764 33068
rect 28810 33056 28816 33108
rect 28868 33096 28874 33108
rect 29181 33099 29239 33105
rect 29181 33096 29193 33099
rect 28868 33068 29193 33096
rect 28868 33056 28874 33068
rect 29181 33065 29193 33068
rect 29227 33065 29239 33099
rect 29181 33059 29239 33065
rect 29270 33056 29276 33108
rect 29328 33096 29334 33108
rect 32582 33096 32588 33108
rect 29328 33068 32588 33096
rect 29328 33056 29334 33068
rect 32582 33056 32588 33068
rect 32640 33056 32646 33108
rect 29822 33028 29828 33040
rect 28736 33000 29828 33028
rect 25041 32991 25099 32997
rect 29822 32988 29828 33000
rect 29880 32988 29886 33040
rect 29914 32988 29920 33040
rect 29972 33028 29978 33040
rect 29972 33000 31892 33028
rect 29972 32988 29978 33000
rect 20622 32920 20628 32972
rect 20680 32960 20686 32972
rect 29932 32960 29960 32988
rect 31864 32969 31892 33000
rect 31481 32963 31539 32969
rect 31481 32960 31493 32963
rect 20680 32932 24716 32960
rect 20680 32920 20686 32932
rect 21453 32895 21511 32901
rect 21453 32861 21465 32895
rect 21499 32861 21511 32895
rect 21453 32855 21511 32861
rect 19996 32796 20576 32824
rect 21468 32824 21496 32855
rect 21542 32852 21548 32904
rect 21600 32892 21606 32904
rect 22830 32892 22836 32904
rect 21600 32864 21645 32892
rect 22791 32864 22836 32892
rect 21600 32852 21606 32864
rect 22830 32852 22836 32864
rect 22888 32852 22894 32904
rect 22925 32895 22983 32901
rect 22925 32861 22937 32895
rect 22971 32861 22983 32895
rect 22925 32855 22983 32861
rect 22370 32824 22376 32836
rect 21468 32796 22376 32824
rect 16022 32716 16028 32768
rect 16080 32756 16086 32768
rect 19996 32756 20024 32796
rect 22370 32784 22376 32796
rect 22428 32784 22434 32836
rect 22462 32784 22468 32836
rect 22520 32824 22526 32836
rect 22940 32824 22968 32855
rect 23382 32824 23388 32836
rect 22520 32796 23388 32824
rect 22520 32784 22526 32796
rect 23382 32784 23388 32796
rect 23440 32784 23446 32836
rect 23658 32824 23664 32836
rect 23619 32796 23664 32824
rect 23658 32784 23664 32796
rect 23716 32784 23722 32836
rect 24029 32827 24087 32833
rect 24029 32793 24041 32827
rect 24075 32824 24087 32827
rect 24118 32824 24124 32836
rect 24075 32796 24124 32824
rect 24075 32793 24087 32796
rect 24029 32787 24087 32793
rect 24118 32784 24124 32796
rect 24176 32784 24182 32836
rect 16080 32728 20024 32756
rect 16080 32716 16086 32728
rect 20162 32716 20168 32768
rect 20220 32756 20226 32768
rect 20622 32756 20628 32768
rect 20220 32728 20628 32756
rect 20220 32716 20226 32728
rect 20622 32716 20628 32728
rect 20680 32716 20686 32768
rect 20898 32756 20904 32768
rect 20859 32728 20904 32756
rect 20898 32716 20904 32728
rect 20956 32716 20962 32768
rect 22830 32716 22836 32768
rect 22888 32756 22894 32768
rect 23290 32756 23296 32768
rect 22888 32728 23296 32756
rect 22888 32716 22894 32728
rect 23290 32716 23296 32728
rect 23348 32716 23354 32768
rect 24688 32756 24716 32932
rect 28828 32932 29960 32960
rect 30024 32932 31493 32960
rect 24765 32895 24823 32901
rect 24765 32861 24777 32895
rect 24811 32861 24823 32895
rect 24765 32855 24823 32861
rect 24857 32895 24915 32901
rect 24857 32861 24869 32895
rect 24903 32892 24915 32895
rect 24946 32892 24952 32904
rect 24903 32864 24952 32892
rect 24903 32861 24915 32864
rect 24857 32855 24915 32861
rect 24780 32824 24808 32855
rect 24946 32852 24952 32864
rect 25004 32852 25010 32904
rect 25501 32895 25559 32901
rect 25501 32861 25513 32895
rect 25547 32892 25559 32895
rect 26602 32892 26608 32904
rect 25547 32864 26608 32892
rect 25547 32861 25559 32864
rect 25501 32855 25559 32861
rect 26602 32852 26608 32864
rect 26660 32892 26666 32904
rect 27801 32895 27859 32901
rect 27801 32892 27813 32895
rect 26660 32864 27813 32892
rect 26660 32852 26666 32864
rect 27801 32861 27813 32864
rect 27847 32892 27859 32895
rect 28828 32892 28856 32932
rect 27847 32864 28856 32892
rect 27847 32861 27859 32864
rect 27801 32855 27859 32861
rect 29178 32852 29184 32904
rect 29236 32892 29242 32904
rect 29733 32895 29791 32901
rect 29733 32892 29745 32895
rect 29236 32864 29745 32892
rect 29236 32852 29242 32864
rect 29733 32861 29745 32864
rect 29779 32861 29791 32895
rect 29914 32892 29920 32904
rect 29875 32864 29920 32892
rect 29733 32855 29791 32861
rect 29914 32852 29920 32864
rect 29972 32852 29978 32904
rect 25406 32824 25412 32836
rect 24780 32796 25412 32824
rect 25406 32784 25412 32796
rect 25464 32784 25470 32836
rect 25590 32784 25596 32836
rect 25648 32824 25654 32836
rect 25746 32827 25804 32833
rect 25746 32824 25758 32827
rect 25648 32796 25758 32824
rect 25648 32784 25654 32796
rect 25746 32793 25758 32796
rect 25792 32793 25804 32827
rect 28068 32827 28126 32833
rect 25746 32787 25804 32793
rect 26804 32796 28028 32824
rect 26804 32756 26832 32796
rect 24688 32728 26832 32756
rect 26881 32759 26939 32765
rect 26881 32725 26893 32759
rect 26927 32756 26939 32759
rect 27430 32756 27436 32768
rect 26927 32728 27436 32756
rect 26927 32725 26939 32728
rect 26881 32719 26939 32725
rect 27430 32716 27436 32728
rect 27488 32716 27494 32768
rect 28000 32756 28028 32796
rect 28068 32793 28080 32827
rect 28114 32824 28126 32827
rect 28442 32824 28448 32836
rect 28114 32796 28448 32824
rect 28114 32793 28126 32796
rect 28068 32787 28126 32793
rect 28442 32784 28448 32796
rect 28500 32784 28506 32836
rect 30024 32824 30052 32932
rect 31481 32929 31493 32932
rect 31527 32929 31539 32963
rect 31481 32923 31539 32929
rect 31849 32963 31907 32969
rect 31849 32929 31861 32963
rect 31895 32929 31907 32963
rect 31849 32923 31907 32929
rect 30653 32895 30711 32901
rect 30653 32861 30665 32895
rect 30699 32892 30711 32895
rect 30742 32892 30748 32904
rect 30699 32864 30748 32892
rect 30699 32861 30711 32864
rect 30653 32855 30711 32861
rect 30742 32852 30748 32864
rect 30800 32852 30806 32904
rect 30929 32895 30987 32901
rect 30929 32861 30941 32895
rect 30975 32892 30987 32895
rect 31294 32892 31300 32904
rect 30975 32864 31300 32892
rect 30975 32861 30987 32864
rect 30929 32855 30987 32861
rect 31294 32852 31300 32864
rect 31352 32852 31358 32904
rect 31496 32892 31524 32923
rect 31496 32864 31754 32892
rect 28552 32796 30052 32824
rect 30837 32827 30895 32833
rect 28552 32756 28580 32796
rect 30837 32793 30849 32827
rect 30883 32824 30895 32827
rect 31570 32824 31576 32836
rect 30883 32796 31576 32824
rect 30883 32793 30895 32796
rect 30837 32787 30895 32793
rect 31570 32784 31576 32796
rect 31628 32784 31634 32836
rect 31726 32824 31754 32864
rect 32094 32827 32152 32833
rect 32094 32824 32106 32827
rect 31726 32796 32106 32824
rect 32094 32793 32106 32796
rect 32140 32793 32152 32827
rect 32094 32787 32152 32793
rect 33689 32827 33747 32833
rect 33689 32793 33701 32827
rect 33735 32824 33747 32827
rect 33778 32824 33784 32836
rect 33735 32796 33784 32824
rect 33735 32793 33747 32796
rect 33689 32787 33747 32793
rect 33778 32784 33784 32796
rect 33836 32784 33842 32836
rect 33873 32827 33931 32833
rect 33873 32793 33885 32827
rect 33919 32824 33931 32827
rect 34238 32824 34244 32836
rect 33919 32796 34244 32824
rect 33919 32793 33931 32796
rect 33873 32787 33931 32793
rect 34238 32784 34244 32796
rect 34296 32784 34302 32836
rect 28000 32728 28580 32756
rect 29822 32716 29828 32768
rect 29880 32756 29886 32768
rect 30101 32759 30159 32765
rect 30101 32756 30113 32759
rect 29880 32728 30113 32756
rect 29880 32716 29886 32728
rect 30101 32725 30113 32728
rect 30147 32725 30159 32759
rect 30101 32719 30159 32725
rect 30926 32716 30932 32768
rect 30984 32756 30990 32768
rect 31021 32759 31079 32765
rect 31021 32756 31033 32759
rect 30984 32728 31033 32756
rect 30984 32716 30990 32728
rect 31021 32725 31033 32728
rect 31067 32725 31079 32759
rect 31021 32719 31079 32725
rect 31110 32716 31116 32768
rect 31168 32756 31174 32768
rect 31205 32759 31263 32765
rect 31205 32756 31217 32759
rect 31168 32728 31217 32756
rect 31168 32716 31174 32728
rect 31205 32725 31217 32728
rect 31251 32725 31263 32759
rect 31205 32719 31263 32725
rect 31478 32716 31484 32768
rect 31536 32756 31542 32768
rect 33229 32759 33287 32765
rect 33229 32756 33241 32759
rect 31536 32728 33241 32756
rect 31536 32716 31542 32728
rect 33229 32725 33241 32728
rect 33275 32725 33287 32759
rect 34054 32756 34060 32768
rect 34015 32728 34060 32756
rect 33229 32719 33287 32725
rect 34054 32716 34060 32728
rect 34112 32716 34118 32768
rect 1104 32666 35027 32688
rect 1104 32614 9390 32666
rect 9442 32614 9454 32666
rect 9506 32614 9518 32666
rect 9570 32614 9582 32666
rect 9634 32614 9646 32666
rect 9698 32614 17831 32666
rect 17883 32614 17895 32666
rect 17947 32614 17959 32666
rect 18011 32614 18023 32666
rect 18075 32614 18087 32666
rect 18139 32614 26272 32666
rect 26324 32614 26336 32666
rect 26388 32614 26400 32666
rect 26452 32614 26464 32666
rect 26516 32614 26528 32666
rect 26580 32614 34713 32666
rect 34765 32614 34777 32666
rect 34829 32614 34841 32666
rect 34893 32614 34905 32666
rect 34957 32614 34969 32666
rect 35021 32614 35027 32666
rect 1104 32592 35027 32614
rect 16298 32512 16304 32564
rect 16356 32552 16362 32564
rect 16356 32524 18552 32552
rect 16356 32512 16362 32524
rect 17402 32444 17408 32496
rect 17460 32484 17466 32496
rect 18386 32487 18444 32493
rect 18386 32484 18398 32487
rect 17460 32456 18398 32484
rect 17460 32444 17466 32456
rect 18386 32453 18398 32456
rect 18432 32453 18444 32487
rect 18524 32484 18552 32524
rect 18874 32512 18880 32564
rect 18932 32552 18938 32564
rect 20533 32555 20591 32561
rect 20533 32552 20545 32555
rect 18932 32524 20545 32552
rect 18932 32512 18938 32524
rect 20533 32521 20545 32524
rect 20579 32521 20591 32555
rect 20533 32515 20591 32521
rect 20622 32512 20628 32564
rect 20680 32552 20686 32564
rect 23014 32552 23020 32564
rect 20680 32524 23020 32552
rect 20680 32512 20686 32524
rect 23014 32512 23020 32524
rect 23072 32512 23078 32564
rect 23106 32512 23112 32564
rect 23164 32552 23170 32564
rect 25590 32552 25596 32564
rect 23164 32524 25452 32552
rect 25551 32524 25596 32552
rect 23164 32512 23170 32524
rect 21266 32484 21272 32496
rect 18524 32456 21272 32484
rect 18386 32447 18444 32453
rect 21266 32444 21272 32456
rect 21324 32444 21330 32496
rect 22916 32487 22974 32493
rect 22916 32453 22928 32487
rect 22962 32484 22974 32487
rect 23842 32484 23848 32496
rect 22962 32456 23848 32484
rect 22962 32453 22974 32456
rect 22916 32447 22974 32453
rect 23842 32444 23848 32456
rect 23900 32444 23906 32496
rect 24946 32484 24952 32496
rect 24596 32456 24952 32484
rect 18141 32419 18199 32425
rect 18141 32385 18153 32419
rect 18187 32416 18199 32419
rect 18230 32416 18236 32428
rect 18187 32388 18236 32416
rect 18187 32385 18199 32388
rect 18141 32379 18199 32385
rect 18230 32376 18236 32388
rect 18288 32376 18294 32428
rect 20349 32419 20407 32425
rect 20349 32385 20361 32419
rect 20395 32416 20407 32419
rect 20438 32416 20444 32428
rect 20395 32388 20444 32416
rect 20395 32385 20407 32388
rect 20349 32379 20407 32385
rect 20438 32376 20444 32388
rect 20496 32376 20502 32428
rect 21082 32416 21088 32428
rect 21043 32388 21088 32416
rect 21082 32376 21088 32388
rect 21140 32376 21146 32428
rect 21177 32419 21235 32425
rect 21177 32385 21189 32419
rect 21223 32385 21235 32419
rect 21177 32379 21235 32385
rect 22189 32419 22247 32425
rect 22189 32385 22201 32419
rect 22235 32416 22247 32419
rect 23934 32416 23940 32428
rect 22235 32388 23940 32416
rect 22235 32385 22247 32388
rect 22189 32379 22247 32385
rect 19610 32308 19616 32360
rect 19668 32348 19674 32360
rect 20165 32351 20223 32357
rect 20165 32348 20177 32351
rect 19668 32320 20177 32348
rect 19668 32308 19674 32320
rect 20165 32317 20177 32320
rect 20211 32348 20223 32351
rect 20898 32348 20904 32360
rect 20211 32320 20904 32348
rect 20211 32317 20223 32320
rect 20165 32311 20223 32317
rect 20898 32308 20904 32320
rect 20956 32308 20962 32360
rect 21192 32348 21220 32379
rect 23934 32376 23940 32388
rect 23992 32376 23998 32428
rect 24596 32425 24624 32456
rect 24946 32444 24952 32456
rect 25004 32484 25010 32496
rect 25222 32484 25228 32496
rect 25004 32456 25228 32484
rect 25004 32444 25010 32456
rect 25222 32444 25228 32456
rect 25280 32444 25286 32496
rect 25424 32484 25452 32524
rect 25590 32512 25596 32524
rect 25648 32512 25654 32564
rect 26050 32552 26056 32564
rect 25700 32524 26056 32552
rect 25700 32484 25728 32524
rect 26050 32512 26056 32524
rect 26108 32512 26114 32564
rect 26142 32512 26148 32564
rect 26200 32552 26206 32564
rect 29454 32552 29460 32564
rect 26200 32524 28764 32552
rect 26200 32512 26206 32524
rect 26878 32484 26884 32496
rect 25424 32456 25728 32484
rect 25792 32456 26884 32484
rect 25792 32425 25820 32456
rect 26878 32444 26884 32456
rect 26936 32444 26942 32496
rect 28169 32487 28227 32493
rect 28169 32453 28181 32487
rect 28215 32484 28227 32487
rect 28626 32484 28632 32496
rect 28215 32456 28632 32484
rect 28215 32453 28227 32456
rect 28169 32447 28227 32453
rect 28626 32444 28632 32456
rect 28684 32444 28690 32496
rect 24581 32419 24639 32425
rect 24581 32385 24593 32419
rect 24627 32385 24639 32419
rect 24581 32379 24639 32385
rect 24673 32419 24731 32425
rect 24673 32385 24685 32419
rect 24719 32385 24731 32419
rect 24673 32379 24731 32385
rect 25777 32419 25835 32425
rect 25777 32385 25789 32419
rect 25823 32385 25835 32419
rect 25777 32379 25835 32385
rect 25869 32419 25927 32425
rect 25869 32385 25881 32419
rect 25915 32385 25927 32419
rect 25869 32379 25927 32385
rect 25961 32419 26019 32425
rect 25961 32385 25973 32419
rect 26007 32385 26019 32419
rect 25961 32379 26019 32385
rect 26099 32419 26157 32425
rect 26099 32385 26111 32419
rect 26145 32416 26157 32419
rect 27157 32419 27215 32425
rect 27157 32416 27169 32419
rect 26145 32388 27169 32416
rect 26145 32385 26157 32388
rect 26099 32379 26157 32385
rect 27157 32385 27169 32388
rect 27203 32385 27215 32419
rect 27338 32416 27344 32428
rect 27299 32388 27344 32416
rect 27157 32379 27215 32385
rect 22462 32348 22468 32360
rect 21192 32320 22468 32348
rect 21192 32280 21220 32320
rect 22462 32308 22468 32320
rect 22520 32308 22526 32360
rect 22646 32348 22652 32360
rect 22607 32320 22652 32348
rect 22646 32308 22652 32320
rect 22704 32308 22710 32360
rect 23842 32308 23848 32360
rect 23900 32348 23906 32360
rect 24688 32348 24716 32379
rect 23900 32320 24716 32348
rect 23900 32308 23906 32320
rect 19076 32252 21220 32280
rect 24688 32280 24716 32320
rect 25682 32308 25688 32360
rect 25740 32348 25746 32360
rect 25884 32348 25912 32379
rect 25740 32320 25912 32348
rect 25740 32308 25746 32320
rect 25774 32280 25780 32292
rect 24688 32252 25780 32280
rect 19076 32224 19104 32252
rect 25774 32240 25780 32252
rect 25832 32240 25838 32292
rect 25866 32240 25872 32292
rect 25924 32280 25930 32292
rect 25976 32280 26004 32379
rect 27338 32376 27344 32388
rect 27396 32376 27402 32428
rect 27433 32419 27491 32425
rect 27433 32385 27445 32419
rect 27479 32416 27491 32419
rect 27522 32416 27528 32428
rect 27479 32388 27528 32416
rect 27479 32385 27491 32388
rect 27433 32379 27491 32385
rect 27522 32376 27528 32388
rect 27580 32376 27586 32428
rect 27617 32419 27675 32425
rect 27617 32385 27629 32419
rect 27663 32385 27675 32419
rect 27617 32379 27675 32385
rect 26237 32351 26295 32357
rect 26237 32317 26249 32351
rect 26283 32317 26295 32351
rect 27632 32348 27660 32379
rect 28258 32376 28264 32428
rect 28316 32416 28322 32428
rect 28445 32419 28503 32425
rect 28445 32416 28457 32419
rect 28316 32388 28457 32416
rect 28316 32376 28322 32388
rect 28445 32385 28457 32388
rect 28491 32385 28503 32419
rect 28736 32416 28764 32524
rect 29104 32524 29460 32552
rect 29104 32493 29132 32524
rect 29454 32512 29460 32524
rect 29512 32512 29518 32564
rect 30190 32512 30196 32564
rect 30248 32552 30254 32564
rect 30285 32555 30343 32561
rect 30285 32552 30297 32555
rect 30248 32524 30297 32552
rect 30248 32512 30254 32524
rect 30285 32521 30297 32524
rect 30331 32521 30343 32555
rect 31570 32552 31576 32564
rect 30285 32515 30343 32521
rect 31312 32524 31576 32552
rect 31312 32496 31340 32524
rect 31570 32512 31576 32524
rect 31628 32512 31634 32564
rect 31662 32512 31668 32564
rect 31720 32512 31726 32564
rect 31754 32512 31760 32564
rect 31812 32552 31818 32564
rect 31812 32524 31857 32552
rect 31812 32512 31818 32524
rect 29089 32487 29147 32493
rect 29089 32453 29101 32487
rect 29135 32453 29147 32487
rect 29089 32447 29147 32453
rect 29178 32444 29184 32496
rect 29236 32484 29242 32496
rect 29289 32487 29347 32493
rect 29289 32484 29301 32487
rect 29236 32456 29301 32484
rect 29236 32444 29242 32456
rect 29289 32453 29301 32456
rect 29335 32453 29347 32487
rect 31294 32484 31300 32496
rect 31255 32456 31300 32484
rect 29289 32447 29347 32453
rect 31294 32444 31300 32456
rect 31352 32444 31358 32496
rect 31386 32444 31392 32496
rect 31444 32484 31450 32496
rect 31680 32484 31708 32512
rect 32674 32484 32680 32496
rect 31444 32456 31616 32484
rect 31680 32456 32536 32484
rect 32635 32456 32680 32484
rect 31444 32444 31450 32456
rect 28736 32388 29316 32416
rect 28445 32379 28503 32385
rect 26237 32311 26295 32317
rect 27448 32320 27660 32348
rect 28353 32351 28411 32357
rect 25924 32252 26004 32280
rect 25924 32240 25930 32252
rect 26050 32240 26056 32292
rect 26108 32280 26114 32292
rect 26252 32280 26280 32311
rect 27448 32292 27476 32320
rect 28353 32317 28365 32351
rect 28399 32348 28411 32351
rect 28534 32348 28540 32360
rect 28399 32320 28540 32348
rect 28399 32317 28411 32320
rect 28353 32311 28411 32317
rect 28534 32308 28540 32320
rect 28592 32308 28598 32360
rect 26108 32252 26280 32280
rect 26108 32240 26114 32252
rect 27430 32240 27436 32292
rect 27488 32240 27494 32292
rect 27525 32283 27583 32289
rect 27525 32249 27537 32283
rect 27571 32280 27583 32283
rect 28629 32283 28687 32289
rect 28629 32280 28641 32283
rect 27571 32252 28641 32280
rect 27571 32249 27583 32252
rect 27525 32243 27583 32249
rect 28629 32249 28641 32252
rect 28675 32249 28687 32283
rect 28629 32243 28687 32249
rect 19058 32172 19064 32224
rect 19116 32172 19122 32224
rect 19334 32172 19340 32224
rect 19392 32212 19398 32224
rect 19521 32215 19579 32221
rect 19521 32212 19533 32215
rect 19392 32184 19533 32212
rect 19392 32172 19398 32184
rect 19521 32181 19533 32184
rect 19567 32181 19579 32215
rect 19521 32175 19579 32181
rect 20714 32172 20720 32224
rect 20772 32212 20778 32224
rect 21361 32215 21419 32221
rect 21361 32212 21373 32215
rect 20772 32184 21373 32212
rect 20772 32172 20778 32184
rect 21361 32181 21373 32184
rect 21407 32181 21419 32215
rect 21361 32175 21419 32181
rect 21450 32172 21456 32224
rect 21508 32212 21514 32224
rect 22005 32215 22063 32221
rect 22005 32212 22017 32215
rect 21508 32184 22017 32212
rect 21508 32172 21514 32184
rect 22005 32181 22017 32184
rect 22051 32181 22063 32215
rect 24026 32212 24032 32224
rect 23939 32184 24032 32212
rect 22005 32175 22063 32181
rect 24026 32172 24032 32184
rect 24084 32212 24090 32224
rect 24670 32212 24676 32224
rect 24084 32184 24676 32212
rect 24084 32172 24090 32184
rect 24670 32172 24676 32184
rect 24728 32172 24734 32224
rect 24857 32215 24915 32221
rect 24857 32181 24869 32215
rect 24903 32212 24915 32215
rect 27982 32212 27988 32224
rect 24903 32184 27988 32212
rect 24903 32181 24915 32184
rect 24857 32175 24915 32181
rect 27982 32172 27988 32184
rect 28040 32172 28046 32224
rect 28074 32172 28080 32224
rect 28132 32212 28138 32224
rect 29288 32221 29316 32388
rect 29822 32376 29828 32428
rect 29880 32416 29886 32428
rect 30101 32419 30159 32425
rect 30101 32416 30113 32419
rect 29880 32388 30113 32416
rect 29880 32376 29886 32388
rect 30101 32385 30113 32388
rect 30147 32385 30159 32419
rect 31478 32416 31484 32428
rect 31439 32388 31484 32416
rect 30101 32379 30159 32385
rect 31478 32376 31484 32388
rect 31536 32376 31542 32428
rect 31588 32425 31616 32456
rect 32508 32425 32536 32456
rect 32674 32444 32680 32456
rect 32732 32444 32738 32496
rect 31573 32419 31631 32425
rect 31573 32385 31585 32419
rect 31619 32385 31631 32419
rect 31573 32379 31631 32385
rect 32493 32419 32551 32425
rect 32493 32385 32505 32419
rect 32539 32385 32551 32419
rect 32493 32379 32551 32385
rect 29454 32308 29460 32360
rect 29512 32348 29518 32360
rect 29917 32351 29975 32357
rect 29917 32348 29929 32351
rect 29512 32320 29929 32348
rect 29512 32308 29518 32320
rect 29917 32317 29929 32320
rect 29963 32317 29975 32351
rect 29917 32311 29975 32317
rect 30834 32308 30840 32360
rect 30892 32348 30898 32360
rect 31588 32348 31616 32379
rect 33410 32348 33416 32360
rect 30892 32320 33416 32348
rect 30892 32308 30898 32320
rect 33410 32308 33416 32320
rect 33468 32308 33474 32360
rect 34330 32348 34336 32360
rect 34291 32320 34336 32348
rect 34330 32308 34336 32320
rect 34388 32308 34394 32360
rect 29730 32240 29736 32292
rect 29788 32280 29794 32292
rect 32306 32280 32312 32292
rect 29788 32252 32312 32280
rect 29788 32240 29794 32252
rect 32306 32240 32312 32252
rect 32364 32240 32370 32292
rect 28169 32215 28227 32221
rect 28169 32212 28181 32215
rect 28132 32184 28181 32212
rect 28132 32172 28138 32184
rect 28169 32181 28181 32184
rect 28215 32181 28227 32215
rect 28169 32175 28227 32181
rect 29273 32215 29331 32221
rect 29273 32181 29285 32215
rect 29319 32181 29331 32215
rect 29454 32212 29460 32224
rect 29415 32184 29460 32212
rect 29273 32175 29331 32181
rect 29454 32172 29460 32184
rect 29512 32172 29518 32224
rect 31202 32172 31208 32224
rect 31260 32212 31266 32224
rect 31297 32215 31355 32221
rect 31297 32212 31309 32215
rect 31260 32184 31309 32212
rect 31260 32172 31266 32184
rect 31297 32181 31309 32184
rect 31343 32212 31355 32215
rect 31386 32212 31392 32224
rect 31343 32184 31392 32212
rect 31343 32181 31355 32184
rect 31297 32175 31355 32181
rect 31386 32172 31392 32184
rect 31444 32172 31450 32224
rect 1104 32122 34868 32144
rect 1104 32070 5170 32122
rect 5222 32070 5234 32122
rect 5286 32070 5298 32122
rect 5350 32070 5362 32122
rect 5414 32070 5426 32122
rect 5478 32070 13611 32122
rect 13663 32070 13675 32122
rect 13727 32070 13739 32122
rect 13791 32070 13803 32122
rect 13855 32070 13867 32122
rect 13919 32070 22052 32122
rect 22104 32070 22116 32122
rect 22168 32070 22180 32122
rect 22232 32070 22244 32122
rect 22296 32070 22308 32122
rect 22360 32070 30493 32122
rect 30545 32070 30557 32122
rect 30609 32070 30621 32122
rect 30673 32070 30685 32122
rect 30737 32070 30749 32122
rect 30801 32070 34868 32122
rect 1104 32048 34868 32070
rect 17402 32008 17408 32020
rect 17363 31980 17408 32008
rect 17402 31968 17408 31980
rect 17460 31968 17466 32020
rect 17586 31968 17592 32020
rect 17644 32008 17650 32020
rect 20165 32011 20223 32017
rect 20165 32008 20177 32011
rect 17644 31980 20177 32008
rect 17644 31968 17650 31980
rect 20165 31977 20177 31980
rect 20211 31977 20223 32011
rect 20165 31971 20223 31977
rect 21266 31968 21272 32020
rect 21324 32008 21330 32020
rect 21324 31980 22094 32008
rect 21324 31968 21330 31980
rect 17678 31900 17684 31952
rect 17736 31940 17742 31952
rect 17736 31912 19196 31940
rect 17736 31900 17742 31912
rect 18417 31875 18475 31881
rect 18417 31872 18429 31875
rect 17604 31844 18429 31872
rect 1762 31764 1768 31816
rect 1820 31804 1826 31816
rect 17604 31813 17632 31844
rect 18417 31841 18429 31844
rect 18463 31841 18475 31875
rect 18417 31835 18475 31841
rect 2041 31807 2099 31813
rect 2041 31804 2053 31807
rect 1820 31776 2053 31804
rect 1820 31764 1826 31776
rect 2041 31773 2053 31776
rect 2087 31773 2099 31807
rect 2041 31767 2099 31773
rect 17589 31807 17647 31813
rect 17589 31773 17601 31807
rect 17635 31773 17647 31807
rect 17589 31767 17647 31773
rect 18141 31807 18199 31813
rect 18141 31773 18153 31807
rect 18187 31804 18199 31807
rect 18253 31807 18311 31813
rect 18187 31776 18221 31804
rect 18187 31773 18199 31776
rect 18141 31767 18199 31773
rect 18253 31773 18265 31807
rect 18299 31804 18311 31807
rect 19058 31804 19064 31816
rect 18299 31776 19064 31804
rect 18299 31773 18311 31776
rect 18253 31767 18311 31773
rect 18156 31736 18184 31767
rect 19058 31764 19064 31776
rect 19116 31764 19122 31816
rect 19168 31804 19196 31912
rect 19242 31900 19248 31952
rect 19300 31940 19306 31952
rect 22066 31940 22094 31980
rect 23106 31968 23112 32020
rect 23164 32008 23170 32020
rect 23164 31980 23209 32008
rect 23164 31968 23170 31980
rect 23934 31968 23940 32020
rect 23992 32008 23998 32020
rect 24029 32011 24087 32017
rect 24029 32008 24041 32011
rect 23992 31980 24041 32008
rect 23992 31968 23998 31980
rect 24029 31977 24041 31980
rect 24075 31977 24087 32011
rect 24029 31971 24087 31977
rect 24486 31968 24492 32020
rect 24544 32008 24550 32020
rect 24581 32011 24639 32017
rect 24581 32008 24593 32011
rect 24544 31980 24593 32008
rect 24544 31968 24550 31980
rect 24581 31977 24593 31980
rect 24627 31977 24639 32011
rect 24581 31971 24639 31977
rect 25498 31968 25504 32020
rect 25556 32008 25562 32020
rect 25774 32008 25780 32020
rect 25556 31980 25780 32008
rect 25556 31968 25562 31980
rect 25774 31968 25780 31980
rect 25832 32008 25838 32020
rect 26142 32008 26148 32020
rect 25832 31980 26148 32008
rect 25832 31968 25838 31980
rect 26142 31968 26148 31980
rect 26200 31968 26206 32020
rect 27614 31968 27620 32020
rect 27672 32008 27678 32020
rect 29822 32008 29828 32020
rect 27672 31980 29828 32008
rect 27672 31968 27678 31980
rect 29822 31968 29828 31980
rect 29880 32008 29886 32020
rect 30098 32008 30104 32020
rect 29880 31980 29960 32008
rect 30059 31980 30104 32008
rect 29880 31968 29886 31980
rect 25869 31943 25927 31949
rect 25869 31940 25881 31943
rect 19300 31912 20392 31940
rect 22066 31912 25881 31940
rect 19300 31900 19306 31912
rect 20364 31884 20392 31912
rect 25869 31909 25881 31912
rect 25915 31909 25927 31943
rect 25869 31903 25927 31909
rect 27632 31912 29868 31940
rect 19518 31832 19524 31884
rect 19576 31872 19582 31884
rect 19797 31875 19855 31881
rect 19797 31872 19809 31875
rect 19576 31844 19809 31872
rect 19576 31832 19582 31844
rect 19797 31841 19809 31844
rect 19843 31841 19855 31875
rect 19797 31835 19855 31841
rect 20346 31832 20352 31884
rect 20404 31872 20410 31884
rect 22646 31872 22652 31884
rect 20404 31844 20944 31872
rect 20404 31832 20410 31844
rect 19610 31804 19616 31816
rect 19168 31776 19616 31804
rect 19610 31764 19616 31776
rect 19668 31764 19674 31816
rect 19981 31807 20039 31813
rect 19981 31773 19993 31807
rect 20027 31804 20039 31807
rect 20438 31804 20444 31816
rect 20027 31776 20444 31804
rect 20027 31773 20039 31776
rect 19981 31767 20039 31773
rect 20438 31764 20444 31776
rect 20496 31764 20502 31816
rect 20916 31813 20944 31844
rect 22480 31844 22652 31872
rect 20901 31807 20959 31813
rect 20901 31773 20913 31807
rect 20947 31804 20959 31807
rect 22370 31804 22376 31816
rect 20947 31776 22376 31804
rect 20947 31773 20959 31776
rect 20901 31767 20959 31773
rect 22370 31764 22376 31776
rect 22428 31804 22434 31816
rect 22480 31804 22508 31844
rect 22646 31832 22652 31844
rect 22704 31832 22710 31884
rect 23566 31872 23572 31884
rect 22848 31844 23572 31872
rect 22848 31813 22876 31844
rect 23566 31832 23572 31844
rect 23624 31872 23630 31884
rect 24210 31872 24216 31884
rect 23624 31844 24216 31872
rect 23624 31832 23630 31844
rect 24210 31832 24216 31844
rect 24268 31832 24274 31884
rect 24670 31832 24676 31884
rect 24728 31872 24734 31884
rect 25498 31872 25504 31884
rect 24728 31844 24773 31872
rect 25459 31844 25504 31872
rect 24728 31832 24734 31844
rect 25498 31832 25504 31844
rect 25556 31832 25562 31884
rect 25700 31844 26464 31872
rect 25700 31816 25728 31844
rect 22428 31776 22508 31804
rect 22833 31807 22891 31813
rect 22428 31764 22434 31776
rect 22833 31773 22845 31807
rect 22879 31773 22891 31807
rect 22833 31767 22891 31773
rect 22922 31764 22928 31816
rect 22980 31804 22986 31816
rect 23661 31807 23719 31813
rect 23661 31804 23673 31807
rect 22980 31776 23673 31804
rect 22980 31764 22986 31776
rect 23661 31773 23673 31776
rect 23707 31773 23719 31807
rect 23842 31804 23848 31816
rect 23803 31776 23848 31804
rect 23661 31767 23719 31773
rect 23842 31764 23848 31776
rect 23900 31764 23906 31816
rect 24857 31807 24915 31813
rect 24857 31804 24869 31807
rect 23952 31776 24869 31804
rect 18506 31736 18512 31748
rect 18156 31708 18512 31736
rect 18506 31696 18512 31708
rect 18564 31696 18570 31748
rect 20622 31736 20628 31748
rect 18616 31708 20628 31736
rect 17494 31628 17500 31680
rect 17552 31668 17558 31680
rect 18616 31668 18644 31708
rect 20622 31696 20628 31708
rect 20680 31696 20686 31748
rect 20806 31696 20812 31748
rect 20864 31736 20870 31748
rect 21146 31739 21204 31745
rect 21146 31736 21158 31739
rect 20864 31708 21158 31736
rect 20864 31696 20870 31708
rect 21146 31705 21158 31708
rect 21192 31705 21204 31739
rect 22462 31736 22468 31748
rect 21146 31699 21204 31705
rect 22112 31708 22468 31736
rect 17552 31640 18644 31668
rect 17552 31628 17558 31640
rect 19150 31628 19156 31680
rect 19208 31668 19214 31680
rect 22112 31668 22140 31708
rect 22462 31696 22468 31708
rect 22520 31696 22526 31748
rect 23290 31696 23296 31748
rect 23348 31736 23354 31748
rect 23952 31736 23980 31776
rect 24857 31773 24869 31776
rect 24903 31773 24915 31807
rect 25682 31804 25688 31816
rect 25643 31776 25688 31804
rect 24857 31767 24915 31773
rect 25682 31764 25688 31776
rect 25740 31764 25746 31816
rect 26436 31804 26464 31844
rect 26436 31776 26556 31804
rect 23348 31708 23980 31736
rect 23348 31696 23354 31708
rect 24394 31696 24400 31748
rect 24452 31736 24458 31748
rect 24581 31739 24639 31745
rect 24581 31736 24593 31739
rect 24452 31708 24593 31736
rect 24452 31696 24458 31708
rect 24581 31705 24593 31708
rect 24627 31705 24639 31739
rect 24581 31699 24639 31705
rect 19208 31640 22140 31668
rect 19208 31628 19214 31640
rect 22186 31628 22192 31680
rect 22244 31668 22250 31680
rect 22281 31671 22339 31677
rect 22281 31668 22293 31671
rect 22244 31640 22293 31668
rect 22244 31628 22250 31640
rect 22281 31637 22293 31640
rect 22327 31668 22339 31671
rect 22554 31668 22560 31680
rect 22327 31640 22560 31668
rect 22327 31637 22339 31640
rect 22281 31631 22339 31637
rect 22554 31628 22560 31640
rect 22612 31628 22618 31680
rect 23382 31628 23388 31680
rect 23440 31668 23446 31680
rect 23842 31668 23848 31680
rect 23440 31640 23848 31668
rect 23440 31628 23446 31640
rect 23842 31628 23848 31640
rect 23900 31628 23906 31680
rect 25038 31668 25044 31680
rect 24999 31640 25044 31668
rect 25038 31628 25044 31640
rect 25096 31628 25102 31680
rect 26528 31668 26556 31776
rect 26602 31764 26608 31816
rect 26660 31804 26666 31816
rect 27154 31804 27160 31816
rect 26660 31776 27160 31804
rect 26660 31764 26666 31776
rect 27154 31764 27160 31776
rect 27212 31764 27218 31816
rect 27632 31804 27660 31912
rect 29733 31875 29791 31881
rect 29733 31872 29745 31875
rect 27264 31776 27660 31804
rect 27724 31844 29745 31872
rect 26872 31739 26930 31745
rect 26872 31705 26884 31739
rect 26918 31736 26930 31739
rect 27264 31736 27292 31776
rect 26918 31708 27292 31736
rect 26918 31705 26930 31708
rect 26872 31699 26930 31705
rect 27430 31696 27436 31748
rect 27488 31736 27494 31748
rect 27724 31736 27752 31844
rect 29733 31841 29745 31844
rect 29779 31841 29791 31875
rect 29733 31835 29791 31841
rect 28166 31764 28172 31816
rect 28224 31804 28230 31816
rect 28442 31804 28448 31816
rect 28224 31776 28448 31804
rect 28224 31764 28230 31776
rect 28442 31764 28448 31776
rect 28500 31806 28506 31816
rect 28997 31807 29055 31813
rect 28500 31804 28672 31806
rect 28997 31804 29009 31807
rect 28500 31778 29009 31804
rect 28500 31776 28507 31778
rect 28644 31776 29009 31778
rect 28500 31764 28506 31776
rect 28997 31773 29009 31776
rect 29043 31773 29055 31807
rect 28997 31767 29055 31773
rect 27488 31708 27752 31736
rect 27488 31696 27494 31708
rect 28258 31696 28264 31748
rect 28316 31736 28322 31748
rect 28629 31739 28687 31745
rect 28629 31736 28641 31739
rect 28316 31708 28641 31736
rect 28316 31696 28322 31708
rect 28629 31705 28641 31708
rect 28675 31705 28687 31739
rect 28629 31699 28687 31705
rect 28810 31696 28816 31748
rect 28868 31736 28874 31748
rect 29362 31736 29368 31748
rect 28868 31708 29368 31736
rect 28868 31696 28874 31708
rect 29362 31696 29368 31708
rect 29420 31696 29426 31748
rect 29840 31736 29868 31912
rect 29932 31813 29960 31980
rect 30098 31968 30104 31980
rect 30156 31968 30162 32020
rect 30650 31968 30656 32020
rect 30708 32008 30714 32020
rect 31754 32008 31760 32020
rect 30708 31980 31760 32008
rect 30708 31968 30714 31980
rect 31754 31968 31760 31980
rect 31812 31968 31818 32020
rect 33781 32011 33839 32017
rect 33781 32008 33793 32011
rect 31864 31980 33793 32008
rect 31294 31900 31300 31952
rect 31352 31940 31358 31952
rect 31665 31943 31723 31949
rect 31665 31940 31677 31943
rect 31352 31912 31677 31940
rect 31352 31900 31358 31912
rect 31665 31909 31677 31912
rect 31711 31909 31723 31943
rect 31665 31903 31723 31909
rect 31110 31872 31116 31884
rect 30852 31844 31116 31872
rect 29917 31807 29975 31813
rect 29917 31773 29929 31807
rect 29963 31773 29975 31807
rect 30561 31807 30619 31813
rect 30561 31804 30573 31807
rect 29917 31767 29975 31773
rect 30208 31776 30573 31804
rect 30208 31736 30236 31776
rect 30561 31773 30573 31776
rect 30607 31773 30619 31807
rect 30561 31767 30619 31773
rect 30650 31764 30656 31816
rect 30708 31804 30714 31816
rect 30852 31813 30880 31844
rect 31110 31832 31116 31844
rect 31168 31832 31174 31884
rect 31205 31875 31263 31881
rect 31205 31841 31217 31875
rect 31251 31841 31263 31875
rect 31205 31835 31263 31841
rect 30746 31807 30804 31813
rect 30746 31804 30758 31807
rect 30708 31776 30758 31804
rect 30708 31764 30714 31776
rect 30746 31773 30758 31776
rect 30792 31773 30804 31807
rect 30746 31767 30804 31773
rect 30837 31807 30895 31813
rect 30837 31773 30849 31807
rect 30883 31773 30895 31807
rect 31220 31794 31248 31835
rect 31570 31832 31576 31884
rect 31628 31872 31634 31884
rect 31864 31872 31892 31980
rect 33781 31977 33793 31980
rect 33827 31977 33839 32011
rect 33781 31971 33839 31977
rect 32214 31872 32220 31884
rect 31628 31844 31892 31872
rect 31956 31844 32220 31872
rect 31628 31832 31634 31844
rect 31662 31804 31668 31816
rect 30837 31767 30895 31773
rect 30926 31736 30932 31748
rect 29840 31708 30236 31736
rect 30887 31708 30932 31736
rect 30926 31696 30932 31708
rect 30984 31696 30990 31748
rect 31018 31696 31024 31748
rect 31076 31745 31082 31748
rect 31076 31739 31105 31745
rect 31202 31742 31208 31794
rect 31260 31742 31266 31794
rect 31623 31776 31668 31804
rect 31662 31764 31668 31776
rect 31720 31764 31726 31816
rect 31956 31813 31984 31844
rect 32214 31832 32220 31844
rect 32272 31832 32278 31884
rect 32306 31832 32312 31884
rect 32364 31872 32370 31884
rect 32401 31875 32459 31881
rect 32401 31872 32413 31875
rect 32364 31844 32413 31872
rect 32364 31832 32370 31844
rect 32401 31841 32413 31844
rect 32447 31841 32459 31875
rect 32401 31835 32459 31841
rect 32674 31813 32680 31816
rect 31941 31807 31999 31813
rect 31941 31773 31953 31807
rect 31987 31773 31999 31807
rect 31941 31767 31999 31773
rect 32668 31767 32680 31813
rect 32732 31804 32738 31816
rect 32732 31776 32768 31804
rect 32674 31764 32680 31767
rect 32732 31764 32738 31776
rect 31093 31705 31105 31739
rect 31076 31699 31105 31705
rect 31076 31696 31082 31699
rect 27614 31668 27620 31680
rect 26528 31640 27620 31668
rect 27614 31628 27620 31640
rect 27672 31628 27678 31680
rect 27890 31628 27896 31680
rect 27948 31668 27954 31680
rect 27985 31671 28043 31677
rect 27985 31668 27997 31671
rect 27948 31640 27997 31668
rect 27948 31628 27954 31640
rect 27985 31637 27997 31640
rect 28031 31637 28043 31671
rect 27985 31631 28043 31637
rect 31849 31671 31907 31677
rect 31849 31637 31861 31671
rect 31895 31668 31907 31671
rect 32398 31668 32404 31680
rect 31895 31640 32404 31668
rect 31895 31637 31907 31640
rect 31849 31631 31907 31637
rect 32398 31628 32404 31640
rect 32456 31628 32462 31680
rect 1104 31578 35027 31600
rect 1104 31526 9390 31578
rect 9442 31526 9454 31578
rect 9506 31526 9518 31578
rect 9570 31526 9582 31578
rect 9634 31526 9646 31578
rect 9698 31526 17831 31578
rect 17883 31526 17895 31578
rect 17947 31526 17959 31578
rect 18011 31526 18023 31578
rect 18075 31526 18087 31578
rect 18139 31526 26272 31578
rect 26324 31526 26336 31578
rect 26388 31526 26400 31578
rect 26452 31526 26464 31578
rect 26516 31526 26528 31578
rect 26580 31526 34713 31578
rect 34765 31526 34777 31578
rect 34829 31526 34841 31578
rect 34893 31526 34905 31578
rect 34957 31526 34969 31578
rect 35021 31526 35027 31578
rect 1104 31504 35027 31526
rect 17037 31467 17095 31473
rect 17037 31433 17049 31467
rect 17083 31464 17095 31467
rect 20806 31464 20812 31476
rect 17083 31436 20812 31464
rect 17083 31433 17095 31436
rect 17037 31427 17095 31433
rect 20806 31424 20812 31436
rect 20864 31424 20870 31476
rect 20993 31467 21051 31473
rect 20993 31433 21005 31467
rect 21039 31464 21051 31467
rect 22094 31464 22100 31476
rect 21039 31436 22100 31464
rect 21039 31433 21051 31436
rect 20993 31427 21051 31433
rect 22094 31424 22100 31436
rect 22152 31424 22158 31476
rect 22462 31424 22468 31476
rect 22520 31464 22526 31476
rect 25130 31464 25136 31476
rect 22520 31436 25136 31464
rect 22520 31424 22526 31436
rect 25130 31424 25136 31436
rect 25188 31424 25194 31476
rect 31202 31464 31208 31476
rect 28184 31436 28672 31464
rect 20714 31396 20720 31408
rect 17236 31368 20720 31396
rect 1762 31328 1768 31340
rect 1723 31300 1768 31328
rect 1762 31288 1768 31300
rect 1820 31288 1826 31340
rect 17236 31337 17264 31368
rect 20714 31356 20720 31368
rect 20772 31356 20778 31408
rect 21082 31396 21088 31408
rect 21043 31368 21088 31396
rect 21082 31356 21088 31368
rect 21140 31356 21146 31408
rect 22364 31399 22422 31405
rect 22364 31365 22376 31399
rect 22410 31396 22422 31399
rect 23474 31396 23480 31408
rect 22410 31368 23480 31396
rect 22410 31365 22422 31368
rect 22364 31359 22422 31365
rect 23474 31356 23480 31368
rect 23532 31356 23538 31408
rect 24854 31405 24860 31408
rect 24848 31396 24860 31405
rect 24815 31368 24860 31396
rect 24848 31359 24860 31368
rect 24854 31356 24860 31359
rect 24912 31356 24918 31408
rect 27062 31356 27068 31408
rect 27120 31396 27126 31408
rect 27402 31399 27460 31405
rect 27402 31396 27414 31399
rect 27120 31368 27414 31396
rect 27120 31356 27126 31368
rect 27402 31365 27414 31368
rect 27448 31396 27460 31399
rect 28184 31396 28212 31436
rect 27448 31368 28212 31396
rect 28644 31396 28672 31436
rect 28828 31436 31208 31464
rect 28828 31396 28856 31436
rect 31202 31424 31208 31436
rect 31260 31424 31266 31476
rect 31570 31464 31576 31476
rect 31531 31436 31576 31464
rect 31570 31424 31576 31436
rect 31628 31424 31634 31476
rect 31754 31464 31760 31476
rect 31715 31436 31760 31464
rect 31754 31424 31760 31436
rect 31812 31424 31818 31476
rect 29822 31396 29828 31408
rect 28644 31368 28856 31396
rect 29380 31368 29828 31396
rect 27448 31365 27460 31368
rect 27402 31359 27460 31365
rect 17221 31331 17279 31337
rect 17221 31297 17233 31331
rect 17267 31297 17279 31331
rect 17221 31291 17279 31297
rect 17586 31288 17592 31340
rect 17644 31328 17650 31340
rect 18598 31337 18604 31340
rect 17865 31331 17923 31337
rect 17865 31328 17877 31331
rect 17644 31300 17877 31328
rect 17644 31288 17650 31300
rect 17865 31297 17877 31300
rect 17911 31297 17923 31331
rect 18592 31328 18604 31337
rect 18559 31300 18604 31328
rect 17865 31291 17923 31297
rect 18592 31291 18604 31300
rect 18598 31288 18604 31291
rect 18656 31288 18662 31340
rect 20530 31288 20536 31340
rect 20588 31328 20594 31340
rect 20901 31331 20959 31337
rect 20901 31328 20913 31331
rect 20588 31300 20913 31328
rect 20588 31288 20594 31300
rect 20901 31297 20913 31300
rect 20947 31297 20959 31331
rect 20901 31291 20959 31297
rect 22097 31331 22155 31337
rect 22097 31297 22109 31331
rect 22143 31328 22155 31331
rect 22646 31328 22652 31340
rect 22143 31300 22652 31328
rect 22143 31297 22155 31300
rect 22097 31291 22155 31297
rect 1949 31263 2007 31269
rect 1949 31229 1961 31263
rect 1995 31260 2007 31263
rect 2130 31260 2136 31272
rect 1995 31232 2136 31260
rect 1995 31229 2007 31232
rect 1949 31223 2007 31229
rect 2130 31220 2136 31232
rect 2188 31220 2194 31272
rect 2774 31260 2780 31272
rect 2735 31232 2780 31260
rect 2774 31220 2780 31232
rect 2832 31220 2838 31272
rect 18230 31220 18236 31272
rect 18288 31260 18294 31272
rect 18325 31263 18383 31269
rect 18325 31260 18337 31263
rect 18288 31232 18337 31260
rect 18288 31220 18294 31232
rect 18325 31229 18337 31232
rect 18371 31229 18383 31263
rect 20916 31260 20944 31291
rect 22646 31288 22652 31300
rect 22704 31288 22710 31340
rect 24121 31331 24179 31337
rect 24121 31297 24133 31331
rect 24167 31328 24179 31331
rect 24167 31300 26372 31328
rect 24167 31297 24179 31300
rect 24121 31291 24179 31297
rect 24578 31260 24584 31272
rect 20916 31232 22094 31260
rect 24539 31232 24584 31260
rect 18325 31223 18383 31229
rect 20717 31195 20775 31201
rect 20717 31161 20729 31195
rect 20763 31192 20775 31195
rect 21358 31192 21364 31204
rect 20763 31164 21364 31192
rect 20763 31161 20775 31164
rect 20717 31155 20775 31161
rect 21358 31152 21364 31164
rect 21416 31152 21422 31204
rect 17681 31127 17739 31133
rect 17681 31093 17693 31127
rect 17727 31124 17739 31127
rect 18598 31124 18604 31136
rect 17727 31096 18604 31124
rect 17727 31093 17739 31096
rect 17681 31087 17739 31093
rect 18598 31084 18604 31096
rect 18656 31084 18662 31136
rect 19242 31084 19248 31136
rect 19300 31124 19306 31136
rect 19705 31127 19763 31133
rect 19705 31124 19717 31127
rect 19300 31096 19717 31124
rect 19300 31084 19306 31096
rect 19705 31093 19717 31096
rect 19751 31093 19763 31127
rect 19705 31087 19763 31093
rect 19886 31084 19892 31136
rect 19944 31124 19950 31136
rect 21269 31127 21327 31133
rect 21269 31124 21281 31127
rect 19944 31096 21281 31124
rect 19944 31084 19950 31096
rect 21269 31093 21281 31096
rect 21315 31093 21327 31127
rect 21269 31087 21327 31093
rect 21910 31084 21916 31136
rect 21968 31124 21974 31136
rect 22066 31124 22094 31232
rect 24578 31220 24584 31232
rect 24636 31220 24642 31272
rect 26344 31260 26372 31300
rect 26418 31288 26424 31340
rect 26476 31328 26482 31340
rect 26605 31331 26663 31337
rect 26476 31300 26521 31328
rect 26476 31288 26482 31300
rect 26605 31297 26617 31331
rect 26651 31328 26663 31331
rect 26970 31328 26976 31340
rect 26651 31300 26976 31328
rect 26651 31297 26663 31300
rect 26605 31291 26663 31297
rect 26970 31288 26976 31300
rect 27028 31288 27034 31340
rect 27157 31331 27215 31337
rect 27157 31297 27169 31331
rect 27203 31328 27215 31331
rect 27246 31328 27252 31340
rect 27203 31300 27252 31328
rect 27203 31297 27215 31300
rect 27157 31291 27215 31297
rect 27246 31288 27252 31300
rect 27304 31288 27310 31340
rect 27798 31288 27804 31340
rect 27856 31328 27862 31340
rect 28718 31328 28724 31340
rect 27856 31300 28724 31328
rect 27856 31288 27862 31300
rect 28718 31288 28724 31300
rect 28776 31288 28782 31340
rect 29380 31337 29408 31368
rect 29822 31356 29828 31368
rect 29880 31356 29886 31408
rect 31478 31396 31484 31408
rect 31439 31368 31484 31396
rect 31478 31356 31484 31368
rect 31536 31356 31542 31408
rect 31846 31356 31852 31408
rect 31904 31396 31910 31408
rect 32677 31399 32735 31405
rect 32677 31396 32689 31399
rect 31904 31368 32689 31396
rect 31904 31356 31910 31368
rect 32677 31365 32689 31368
rect 32723 31365 32735 31399
rect 32677 31359 32735 31365
rect 29365 31331 29423 31337
rect 29365 31297 29377 31331
rect 29411 31297 29423 31331
rect 29365 31291 29423 31297
rect 29632 31331 29690 31337
rect 29632 31297 29644 31331
rect 29678 31328 29690 31331
rect 29678 31300 31340 31328
rect 29678 31297 29690 31300
rect 29632 31291 29690 31297
rect 27062 31260 27068 31272
rect 26344 31232 27068 31260
rect 27062 31220 27068 31232
rect 27120 31220 27126 31272
rect 30742 31220 30748 31272
rect 30800 31260 30806 31272
rect 31205 31263 31263 31269
rect 31205 31260 31217 31263
rect 30800 31232 31217 31260
rect 30800 31220 30806 31232
rect 31205 31229 31217 31232
rect 31251 31229 31263 31263
rect 31205 31223 31263 31229
rect 23477 31195 23535 31201
rect 23477 31161 23489 31195
rect 23523 31192 23535 31195
rect 23842 31192 23848 31204
rect 23523 31164 23848 31192
rect 23523 31161 23535 31164
rect 23477 31155 23535 31161
rect 23842 31152 23848 31164
rect 23900 31192 23906 31204
rect 24394 31192 24400 31204
rect 23900 31164 24400 31192
rect 23900 31152 23906 31164
rect 24394 31152 24400 31164
rect 24452 31152 24458 31204
rect 29362 31192 29368 31204
rect 25792 31164 27200 31192
rect 23566 31124 23572 31136
rect 21968 31096 23572 31124
rect 21968 31084 21974 31096
rect 23566 31084 23572 31096
rect 23624 31084 23630 31136
rect 23750 31084 23756 31136
rect 23808 31124 23814 31136
rect 23937 31127 23995 31133
rect 23937 31124 23949 31127
rect 23808 31096 23949 31124
rect 23808 31084 23814 31096
rect 23937 31093 23949 31096
rect 23983 31093 23995 31127
rect 23937 31087 23995 31093
rect 24762 31084 24768 31136
rect 24820 31124 24826 31136
rect 25792 31124 25820 31164
rect 24820 31096 25820 31124
rect 24820 31084 24826 31096
rect 25866 31084 25872 31136
rect 25924 31124 25930 31136
rect 25961 31127 26019 31133
rect 25961 31124 25973 31127
rect 25924 31096 25973 31124
rect 25924 31084 25930 31096
rect 25961 31093 25973 31096
rect 26007 31093 26019 31127
rect 25961 31087 26019 31093
rect 26421 31127 26479 31133
rect 26421 31093 26433 31127
rect 26467 31124 26479 31127
rect 26786 31124 26792 31136
rect 26467 31096 26792 31124
rect 26467 31093 26479 31096
rect 26421 31087 26479 31093
rect 26786 31084 26792 31096
rect 26844 31084 26850 31136
rect 27172 31124 27200 31164
rect 28460 31164 29368 31192
rect 28460 31124 28488 31164
rect 29362 31152 29368 31164
rect 29420 31152 29426 31204
rect 31312 31192 31340 31300
rect 31386 31288 31392 31340
rect 31444 31328 31450 31340
rect 32490 31328 32496 31340
rect 31444 31300 31489 31328
rect 32451 31300 32496 31328
rect 31444 31288 31450 31300
rect 32490 31288 32496 31300
rect 32548 31288 32554 31340
rect 34330 31328 34336 31340
rect 34291 31300 34336 31328
rect 34330 31288 34336 31300
rect 34388 31288 34394 31340
rect 31478 31220 31484 31272
rect 31536 31260 31542 31272
rect 33502 31260 33508 31272
rect 31536 31232 33508 31260
rect 31536 31220 31542 31232
rect 33502 31220 33508 31232
rect 33560 31220 33566 31272
rect 33686 31192 33692 31204
rect 30300 31164 31064 31192
rect 31312 31164 33692 31192
rect 27172 31096 28488 31124
rect 28537 31127 28595 31133
rect 28537 31093 28549 31127
rect 28583 31124 28595 31127
rect 28718 31124 28724 31136
rect 28583 31096 28724 31124
rect 28583 31093 28595 31096
rect 28537 31087 28595 31093
rect 28718 31084 28724 31096
rect 28776 31124 28782 31136
rect 30300 31124 30328 31164
rect 28776 31096 30328 31124
rect 28776 31084 28782 31096
rect 30374 31084 30380 31136
rect 30432 31124 30438 31136
rect 30745 31127 30803 31133
rect 30745 31124 30757 31127
rect 30432 31096 30757 31124
rect 30432 31084 30438 31096
rect 30745 31093 30757 31096
rect 30791 31124 30803 31127
rect 30926 31124 30932 31136
rect 30791 31096 30932 31124
rect 30791 31093 30803 31096
rect 30745 31087 30803 31093
rect 30926 31084 30932 31096
rect 30984 31084 30990 31136
rect 31036 31124 31064 31164
rect 33686 31152 33692 31164
rect 33744 31152 33750 31204
rect 34054 31124 34060 31136
rect 31036 31096 34060 31124
rect 34054 31084 34060 31096
rect 34112 31084 34118 31136
rect 1104 31034 34868 31056
rect 1104 30982 5170 31034
rect 5222 30982 5234 31034
rect 5286 30982 5298 31034
rect 5350 30982 5362 31034
rect 5414 30982 5426 31034
rect 5478 30982 13611 31034
rect 13663 30982 13675 31034
rect 13727 30982 13739 31034
rect 13791 30982 13803 31034
rect 13855 30982 13867 31034
rect 13919 30982 22052 31034
rect 22104 30982 22116 31034
rect 22168 30982 22180 31034
rect 22232 30982 22244 31034
rect 22296 30982 22308 31034
rect 22360 30982 30493 31034
rect 30545 30982 30557 31034
rect 30609 30982 30621 31034
rect 30673 30982 30685 31034
rect 30737 30982 30749 31034
rect 30801 30982 34868 31034
rect 1104 30960 34868 30982
rect 2130 30920 2136 30932
rect 2091 30892 2136 30920
rect 2130 30880 2136 30892
rect 2188 30880 2194 30932
rect 17770 30880 17776 30932
rect 17828 30920 17834 30932
rect 18693 30923 18751 30929
rect 18693 30920 18705 30923
rect 17828 30892 18705 30920
rect 17828 30880 17834 30892
rect 18693 30889 18705 30892
rect 18739 30920 18751 30923
rect 19518 30920 19524 30932
rect 18739 30892 19012 30920
rect 19479 30892 19524 30920
rect 18739 30889 18751 30892
rect 18693 30883 18751 30889
rect 18414 30812 18420 30864
rect 18472 30852 18478 30864
rect 18877 30855 18935 30861
rect 18877 30852 18889 30855
rect 18472 30824 18889 30852
rect 18472 30812 18478 30824
rect 18877 30821 18889 30824
rect 18923 30821 18935 30855
rect 18984 30852 19012 30892
rect 19518 30880 19524 30892
rect 19576 30880 19582 30932
rect 21082 30880 21088 30932
rect 21140 30920 21146 30932
rect 21729 30923 21787 30929
rect 21729 30920 21741 30923
rect 21140 30892 21741 30920
rect 21140 30880 21146 30892
rect 21729 30889 21741 30892
rect 21775 30889 21787 30923
rect 21729 30883 21787 30889
rect 19334 30852 19340 30864
rect 18984 30824 19340 30852
rect 18877 30815 18935 30821
rect 19334 30812 19340 30824
rect 19392 30852 19398 30864
rect 19978 30852 19984 30864
rect 19392 30824 19984 30852
rect 19392 30812 19398 30824
rect 19978 30812 19984 30824
rect 20036 30812 20042 30864
rect 18049 30787 18107 30793
rect 18049 30784 18061 30787
rect 17236 30756 18061 30784
rect 2041 30719 2099 30725
rect 2041 30685 2053 30719
rect 2087 30716 2099 30719
rect 2130 30716 2136 30728
rect 2087 30688 2136 30716
rect 2087 30685 2099 30688
rect 2041 30679 2099 30685
rect 2130 30676 2136 30688
rect 2188 30676 2194 30728
rect 17236 30725 17264 30756
rect 18049 30753 18061 30756
rect 18095 30753 18107 30787
rect 18049 30747 18107 30753
rect 18506 30744 18512 30796
rect 18564 30784 18570 30796
rect 19242 30784 19248 30796
rect 18564 30756 19248 30784
rect 18564 30744 18570 30756
rect 19242 30744 19248 30756
rect 19300 30784 19306 30796
rect 19521 30787 19579 30793
rect 19521 30784 19533 30787
rect 19300 30756 19533 30784
rect 19300 30744 19306 30756
rect 19521 30753 19533 30756
rect 19567 30753 19579 30787
rect 20346 30784 20352 30796
rect 20307 30756 20352 30784
rect 19521 30747 19579 30753
rect 20346 30744 20352 30756
rect 20404 30744 20410 30796
rect 17221 30719 17279 30725
rect 17221 30685 17233 30719
rect 17267 30685 17279 30719
rect 17770 30716 17776 30728
rect 17731 30688 17776 30716
rect 17221 30679 17279 30685
rect 17770 30676 17776 30688
rect 17828 30676 17834 30728
rect 17865 30719 17923 30725
rect 17865 30685 17877 30719
rect 17911 30716 17923 30719
rect 19058 30716 19064 30728
rect 17911 30688 19064 30716
rect 17911 30685 17923 30688
rect 17865 30679 17923 30685
rect 19058 30676 19064 30688
rect 19116 30676 19122 30728
rect 19426 30716 19432 30728
rect 19387 30688 19432 30716
rect 19426 30676 19432 30688
rect 19484 30676 19490 30728
rect 20616 30719 20674 30725
rect 20616 30685 20628 30719
rect 20662 30716 20674 30719
rect 21450 30716 21456 30728
rect 20662 30688 21456 30716
rect 20662 30685 20674 30688
rect 20616 30679 20674 30685
rect 21450 30676 21456 30688
rect 21508 30676 21514 30728
rect 21744 30716 21772 30883
rect 21910 30880 21916 30932
rect 21968 30920 21974 30932
rect 22189 30923 22247 30929
rect 22189 30920 22201 30923
rect 21968 30892 22201 30920
rect 21968 30880 21974 30892
rect 22189 30889 22201 30892
rect 22235 30889 22247 30923
rect 22189 30883 22247 30889
rect 22646 30880 22652 30932
rect 22704 30920 22710 30932
rect 24949 30923 25007 30929
rect 24949 30920 24961 30923
rect 22704 30892 24961 30920
rect 22704 30880 22710 30892
rect 24949 30889 24961 30892
rect 24995 30889 25007 30923
rect 24949 30883 25007 30889
rect 25130 30880 25136 30932
rect 25188 30920 25194 30932
rect 28902 30920 28908 30932
rect 25188 30892 28908 30920
rect 25188 30880 25194 30892
rect 28902 30880 28908 30892
rect 28960 30880 28966 30932
rect 29362 30880 29368 30932
rect 29420 30920 29426 30932
rect 29638 30920 29644 30932
rect 29420 30892 29644 30920
rect 29420 30880 29426 30892
rect 29638 30880 29644 30892
rect 29696 30880 29702 30932
rect 30193 30923 30251 30929
rect 30193 30889 30205 30923
rect 30239 30920 30251 30923
rect 31478 30920 31484 30932
rect 30239 30892 31484 30920
rect 30239 30889 30251 30892
rect 30193 30883 30251 30889
rect 31478 30880 31484 30892
rect 31536 30880 31542 30932
rect 32306 30920 32312 30932
rect 32048 30892 32312 30920
rect 23290 30812 23296 30864
rect 23348 30852 23354 30864
rect 23477 30855 23535 30861
rect 23477 30852 23489 30855
rect 23348 30824 23489 30852
rect 23348 30812 23354 30824
rect 23477 30821 23489 30824
rect 23523 30821 23535 30855
rect 23477 30815 23535 30821
rect 24029 30855 24087 30861
rect 24029 30821 24041 30855
rect 24075 30852 24087 30855
rect 29178 30852 29184 30864
rect 24075 30824 29184 30852
rect 24075 30821 24087 30824
rect 24029 30815 24087 30821
rect 29178 30812 29184 30824
rect 29236 30812 29242 30864
rect 31297 30855 31355 30861
rect 31297 30852 31309 30855
rect 30015 30824 31309 30852
rect 22373 30787 22431 30793
rect 22373 30753 22385 30787
rect 22419 30784 22431 30787
rect 22554 30784 22560 30796
rect 22419 30756 22560 30784
rect 22419 30753 22431 30756
rect 22373 30747 22431 30753
rect 22554 30744 22560 30756
rect 22612 30744 22618 30796
rect 24486 30784 24492 30796
rect 23676 30756 24492 30784
rect 22189 30719 22247 30725
rect 22189 30716 22201 30719
rect 21744 30688 22201 30716
rect 22189 30685 22201 30688
rect 22235 30685 22247 30719
rect 22189 30679 22247 30685
rect 22465 30719 22523 30725
rect 22465 30685 22477 30719
rect 22511 30716 22523 30719
rect 22922 30716 22928 30728
rect 22511 30688 22928 30716
rect 22511 30685 22523 30688
rect 22465 30679 22523 30685
rect 18506 30648 18512 30660
rect 18467 30620 18512 30648
rect 18506 30608 18512 30620
rect 18564 30608 18570 30660
rect 18725 30651 18783 30657
rect 18725 30617 18737 30651
rect 18771 30648 18783 30651
rect 19886 30648 19892 30660
rect 18771 30620 19892 30648
rect 18771 30617 18783 30620
rect 18725 30611 18783 30617
rect 19886 30608 19892 30620
rect 19944 30608 19950 30660
rect 21358 30608 21364 30660
rect 21416 30648 21422 30660
rect 22480 30648 22508 30679
rect 22922 30676 22928 30688
rect 22980 30676 22986 30728
rect 23676 30725 23704 30756
rect 24486 30744 24492 30756
rect 24544 30784 24550 30796
rect 24544 30756 24716 30784
rect 24544 30744 24550 30756
rect 24688 30728 24716 30756
rect 26418 30744 26424 30796
rect 26476 30784 26482 30796
rect 27154 30784 27160 30796
rect 26476 30756 27160 30784
rect 26476 30744 26482 30756
rect 27154 30744 27160 30756
rect 27212 30744 27218 30796
rect 29086 30784 29092 30796
rect 28368 30756 29092 30784
rect 23661 30719 23719 30725
rect 23661 30685 23673 30719
rect 23707 30685 23719 30719
rect 23661 30679 23719 30685
rect 23753 30719 23811 30725
rect 23753 30685 23765 30719
rect 23799 30716 23811 30719
rect 24026 30716 24032 30728
rect 23799 30688 24032 30716
rect 23799 30685 23811 30688
rect 23753 30679 23811 30685
rect 24026 30676 24032 30688
rect 24084 30676 24090 30728
rect 24670 30716 24676 30728
rect 24631 30688 24676 30716
rect 24670 30676 24676 30688
rect 24728 30676 24734 30728
rect 24765 30719 24823 30725
rect 24765 30685 24777 30719
rect 24811 30685 24823 30719
rect 28368 30716 28396 30756
rect 29086 30744 29092 30756
rect 29144 30744 29150 30796
rect 30015 30793 30043 30824
rect 31297 30821 31309 30824
rect 31343 30821 31355 30855
rect 31297 30815 31355 30821
rect 32048 30796 32076 30892
rect 32306 30880 32312 30892
rect 32364 30920 32370 30932
rect 32950 30920 32956 30932
rect 32364 30892 32956 30920
rect 32364 30880 32370 30892
rect 32950 30880 32956 30892
rect 33008 30880 33014 30932
rect 33410 30920 33416 30932
rect 33371 30892 33416 30920
rect 33410 30880 33416 30892
rect 33468 30880 33474 30932
rect 30009 30787 30067 30793
rect 30009 30753 30021 30787
rect 30055 30753 30067 30787
rect 30009 30747 30067 30753
rect 30742 30744 30748 30796
rect 30800 30784 30806 30796
rect 30837 30787 30895 30793
rect 30837 30784 30849 30787
rect 30800 30756 30849 30784
rect 30800 30744 30806 30756
rect 30837 30753 30849 30756
rect 30883 30784 30895 30787
rect 31754 30784 31760 30796
rect 30883 30756 31760 30784
rect 30883 30753 30895 30756
rect 30837 30747 30895 30753
rect 31754 30744 31760 30756
rect 31812 30744 31818 30796
rect 32030 30744 32036 30796
rect 32088 30784 32094 30796
rect 32088 30756 32181 30784
rect 32088 30744 32094 30756
rect 24765 30679 24823 30685
rect 24872 30688 28396 30716
rect 23842 30648 23848 30660
rect 21416 30620 22508 30648
rect 23803 30620 23848 30648
rect 21416 30608 21422 30620
rect 23842 30608 23848 30620
rect 23900 30608 23906 30660
rect 23934 30608 23940 30660
rect 23992 30648 23998 30660
rect 24780 30648 24808 30679
rect 23992 30620 24808 30648
rect 23992 30608 23998 30620
rect 17037 30583 17095 30589
rect 17037 30549 17049 30583
rect 17083 30580 17095 30583
rect 18966 30580 18972 30592
rect 17083 30552 18972 30580
rect 17083 30549 17095 30552
rect 17037 30543 17095 30549
rect 18966 30540 18972 30552
rect 19024 30540 19030 30592
rect 19794 30580 19800 30592
rect 19755 30552 19800 30580
rect 19794 30540 19800 30552
rect 19852 30540 19858 30592
rect 20162 30540 20168 30592
rect 20220 30580 20226 30592
rect 22649 30583 22707 30589
rect 22649 30580 22661 30583
rect 20220 30552 22661 30580
rect 20220 30540 20226 30552
rect 22649 30549 22661 30552
rect 22695 30549 22707 30583
rect 22649 30543 22707 30549
rect 23014 30540 23020 30592
rect 23072 30580 23078 30592
rect 24872 30580 24900 30688
rect 28442 30676 28448 30728
rect 28500 30716 28506 30728
rect 28721 30719 28779 30725
rect 28500 30688 28545 30716
rect 28500 30676 28506 30688
rect 28721 30685 28733 30719
rect 28767 30716 28779 30719
rect 28810 30716 28816 30728
rect 28767 30688 28816 30716
rect 28767 30685 28779 30688
rect 28721 30679 28779 30685
rect 28810 30676 28816 30688
rect 28868 30676 28874 30728
rect 29840 30725 29960 30726
rect 29840 30719 29975 30725
rect 29840 30698 29929 30719
rect 26053 30651 26111 30657
rect 26053 30617 26065 30651
rect 26099 30648 26111 30651
rect 28166 30648 28172 30660
rect 26099 30620 28172 30648
rect 26099 30617 26111 30620
rect 26053 30611 26111 30617
rect 28166 30608 28172 30620
rect 28224 30608 28230 30660
rect 28258 30608 28264 30660
rect 28316 30648 28322 30660
rect 28316 30620 28361 30648
rect 28316 30608 28322 30620
rect 28534 30608 28540 30660
rect 28592 30648 28598 30660
rect 29840 30648 29868 30698
rect 29917 30685 29929 30698
rect 29963 30685 29975 30719
rect 30926 30716 30932 30728
rect 30887 30688 30932 30716
rect 29917 30679 29975 30685
rect 30926 30676 30932 30688
rect 30984 30716 30990 30728
rect 31294 30716 31300 30728
rect 30984 30688 31300 30716
rect 30984 30676 30990 30688
rect 31294 30676 31300 30688
rect 31352 30676 31358 30728
rect 33410 30676 33416 30728
rect 33468 30716 33474 30728
rect 33873 30719 33931 30725
rect 33873 30716 33885 30719
rect 33468 30688 33885 30716
rect 33468 30676 33474 30688
rect 33873 30685 33885 30688
rect 33919 30685 33931 30719
rect 34054 30716 34060 30728
rect 34015 30688 34060 30716
rect 33873 30679 33931 30685
rect 34054 30676 34060 30688
rect 34112 30676 34118 30728
rect 28592 30620 28994 30648
rect 29840 30620 30972 30648
rect 28592 30608 28598 30620
rect 27338 30580 27344 30592
rect 23072 30552 24900 30580
rect 27299 30552 27344 30580
rect 23072 30540 23078 30552
rect 27338 30540 27344 30552
rect 27396 30540 27402 30592
rect 28074 30540 28080 30592
rect 28132 30580 28138 30592
rect 28552 30580 28580 30608
rect 28132 30552 28580 30580
rect 28629 30583 28687 30589
rect 28132 30540 28138 30552
rect 28629 30549 28641 30583
rect 28675 30580 28687 30583
rect 28718 30580 28724 30592
rect 28675 30552 28724 30580
rect 28675 30549 28687 30552
rect 28629 30543 28687 30549
rect 28718 30540 28724 30552
rect 28776 30540 28782 30592
rect 28966 30580 28994 30620
rect 30742 30580 30748 30592
rect 28966 30552 30748 30580
rect 30742 30540 30748 30552
rect 30800 30540 30806 30592
rect 30944 30580 30972 30620
rect 31018 30608 31024 30660
rect 31076 30648 31082 30660
rect 32278 30651 32336 30657
rect 32278 30648 32290 30651
rect 31076 30620 32290 30648
rect 31076 30608 31082 30620
rect 32278 30617 32290 30620
rect 32324 30617 32336 30651
rect 32278 30611 32336 30617
rect 32122 30580 32128 30592
rect 30944 30552 32128 30580
rect 32122 30540 32128 30552
rect 32180 30540 32186 30592
rect 34238 30580 34244 30592
rect 34199 30552 34244 30580
rect 34238 30540 34244 30552
rect 34296 30540 34302 30592
rect 1104 30490 35027 30512
rect 1104 30438 9390 30490
rect 9442 30438 9454 30490
rect 9506 30438 9518 30490
rect 9570 30438 9582 30490
rect 9634 30438 9646 30490
rect 9698 30438 17831 30490
rect 17883 30438 17895 30490
rect 17947 30438 17959 30490
rect 18011 30438 18023 30490
rect 18075 30438 18087 30490
rect 18139 30438 26272 30490
rect 26324 30438 26336 30490
rect 26388 30438 26400 30490
rect 26452 30438 26464 30490
rect 26516 30438 26528 30490
rect 26580 30438 34713 30490
rect 34765 30438 34777 30490
rect 34829 30438 34841 30490
rect 34893 30438 34905 30490
rect 34957 30438 34969 30490
rect 35021 30438 35027 30490
rect 1104 30416 35027 30438
rect 17497 30379 17555 30385
rect 17497 30345 17509 30379
rect 17543 30376 17555 30379
rect 21358 30376 21364 30388
rect 17543 30348 19334 30376
rect 21319 30348 21364 30376
rect 17543 30345 17555 30348
rect 17497 30339 17555 30345
rect 18397 30311 18455 30317
rect 18397 30277 18409 30311
rect 18443 30308 18455 30311
rect 18966 30308 18972 30320
rect 18443 30280 18972 30308
rect 18443 30277 18455 30280
rect 18397 30271 18455 30277
rect 18966 30268 18972 30280
rect 19024 30268 19030 30320
rect 19306 30308 19334 30348
rect 21358 30336 21364 30348
rect 21416 30336 21422 30388
rect 22646 30376 22652 30388
rect 21468 30348 22652 30376
rect 19610 30308 19616 30320
rect 19306 30280 19616 30308
rect 19610 30268 19616 30280
rect 19668 30268 19674 30320
rect 21468 30308 21496 30348
rect 22646 30336 22652 30348
rect 22704 30336 22710 30388
rect 23290 30336 23296 30388
rect 23348 30376 23354 30388
rect 23385 30379 23443 30385
rect 23385 30376 23397 30379
rect 23348 30348 23397 30376
rect 23348 30336 23354 30348
rect 23385 30345 23397 30348
rect 23431 30345 23443 30379
rect 23385 30339 23443 30345
rect 24854 30336 24860 30388
rect 24912 30376 24918 30388
rect 24912 30348 25452 30376
rect 24912 30336 24918 30348
rect 19812 30280 21496 30308
rect 17681 30243 17739 30249
rect 17681 30209 17693 30243
rect 17727 30209 17739 30243
rect 18138 30240 18144 30252
rect 18099 30212 18144 30240
rect 17681 30203 17739 30209
rect 17696 30172 17724 30203
rect 18138 30200 18144 30212
rect 18196 30200 18202 30252
rect 19812 30240 19840 30280
rect 21910 30268 21916 30320
rect 21968 30308 21974 30320
rect 22250 30311 22308 30317
rect 22250 30308 22262 30311
rect 21968 30280 22262 30308
rect 21968 30268 21974 30280
rect 22250 30277 22262 30280
rect 22296 30277 22308 30311
rect 22250 30271 22308 30277
rect 22462 30268 22468 30320
rect 22520 30308 22526 30320
rect 25032 30311 25090 30317
rect 22520 30280 24992 30308
rect 22520 30268 22526 30280
rect 18248 30212 19840 30240
rect 19904 30240 20116 30244
rect 20237 30243 20295 30249
rect 20237 30240 20249 30243
rect 19904 30216 20249 30240
rect 18248 30172 18276 30212
rect 17696 30144 18276 30172
rect 19242 30132 19248 30184
rect 19300 30172 19306 30184
rect 19904 30172 19932 30216
rect 20088 30212 20249 30216
rect 20237 30209 20249 30212
rect 20283 30209 20295 30243
rect 20237 30203 20295 30209
rect 22830 30200 22836 30252
rect 22888 30240 22894 30252
rect 24029 30243 24087 30249
rect 24029 30240 24041 30243
rect 22888 30212 24041 30240
rect 22888 30200 22894 30212
rect 24029 30209 24041 30212
rect 24075 30209 24087 30243
rect 24029 30203 24087 30209
rect 19300 30144 19932 30172
rect 19981 30175 20039 30181
rect 19300 30132 19306 30144
rect 19981 30141 19993 30175
rect 20027 30141 20039 30175
rect 19981 30135 20039 30141
rect 22005 30175 22063 30181
rect 22005 30141 22017 30175
rect 22051 30141 22063 30175
rect 23842 30172 23848 30184
rect 23803 30144 23848 30172
rect 22005 30135 22063 30141
rect 19150 30064 19156 30116
rect 19208 30104 19214 30116
rect 19996 30104 20024 30135
rect 19208 30076 20024 30104
rect 19208 30064 19214 30076
rect 17494 29996 17500 30048
rect 17552 30036 17558 30048
rect 18506 30036 18512 30048
rect 17552 30008 18512 30036
rect 17552 29996 17558 30008
rect 18506 29996 18512 30008
rect 18564 29996 18570 30048
rect 18782 29996 18788 30048
rect 18840 30036 18846 30048
rect 19242 30036 19248 30048
rect 18840 30008 19248 30036
rect 18840 29996 18846 30008
rect 19242 29996 19248 30008
rect 19300 29996 19306 30048
rect 19518 30036 19524 30048
rect 19479 30008 19524 30036
rect 19518 29996 19524 30008
rect 19576 29996 19582 30048
rect 19996 30036 20024 30076
rect 22020 30036 22048 30135
rect 23842 30132 23848 30144
rect 23900 30132 23906 30184
rect 24044 30172 24072 30203
rect 24578 30200 24584 30252
rect 24636 30240 24642 30252
rect 24765 30243 24823 30249
rect 24765 30240 24777 30243
rect 24636 30212 24777 30240
rect 24636 30200 24642 30212
rect 24765 30209 24777 30212
rect 24811 30209 24823 30243
rect 24765 30203 24823 30209
rect 24854 30200 24860 30252
rect 24912 30200 24918 30252
rect 24964 30240 24992 30280
rect 25032 30277 25044 30311
rect 25078 30308 25090 30311
rect 25314 30308 25320 30320
rect 25078 30280 25320 30308
rect 25078 30277 25090 30280
rect 25032 30271 25090 30277
rect 25314 30268 25320 30280
rect 25372 30268 25378 30320
rect 25424 30308 25452 30348
rect 25590 30336 25596 30388
rect 25648 30376 25654 30388
rect 25648 30348 25820 30376
rect 25648 30336 25654 30348
rect 25682 30308 25688 30320
rect 25424 30280 25688 30308
rect 25682 30268 25688 30280
rect 25740 30268 25746 30320
rect 25792 30308 25820 30348
rect 27982 30336 27988 30388
rect 28040 30376 28046 30388
rect 30374 30376 30380 30388
rect 28040 30348 30380 30376
rect 28040 30336 28046 30348
rect 30374 30336 30380 30348
rect 30432 30336 30438 30388
rect 30466 30336 30472 30388
rect 30524 30376 30530 30388
rect 31662 30376 31668 30388
rect 30524 30348 31668 30376
rect 30524 30336 30530 30348
rect 31662 30336 31668 30348
rect 31720 30336 31726 30388
rect 26050 30308 26056 30320
rect 25792 30280 26056 30308
rect 26050 30268 26056 30280
rect 26108 30268 26114 30320
rect 27792 30311 27850 30317
rect 27792 30277 27804 30311
rect 27838 30308 27850 30311
rect 28350 30308 28356 30320
rect 27838 30280 28356 30308
rect 27838 30277 27850 30280
rect 27792 30271 27850 30277
rect 28350 30268 28356 30280
rect 28408 30268 28414 30320
rect 29748 30280 30880 30308
rect 29748 30240 29776 30280
rect 24964 30212 29776 30240
rect 29825 30243 29883 30249
rect 29825 30209 29837 30243
rect 29871 30240 29883 30243
rect 30006 30240 30012 30252
rect 29871 30212 30012 30240
rect 29871 30209 29883 30212
rect 29825 30203 29883 30209
rect 30006 30200 30012 30212
rect 30064 30200 30070 30252
rect 30852 30249 30880 30280
rect 31570 30268 31576 30320
rect 31628 30308 31634 30320
rect 33226 30317 33232 30320
rect 32401 30311 32459 30317
rect 32401 30308 32413 30311
rect 31628 30280 32413 30308
rect 31628 30268 31634 30280
rect 32401 30277 32413 30280
rect 32447 30277 32459 30311
rect 33220 30308 33232 30317
rect 33187 30280 33232 30308
rect 32401 30271 32459 30277
rect 33220 30271 33232 30280
rect 33226 30268 33232 30271
rect 33284 30268 33290 30320
rect 30837 30243 30895 30249
rect 30837 30209 30849 30243
rect 30883 30240 30895 30243
rect 30883 30212 31616 30240
rect 30883 30209 30895 30212
rect 30837 30203 30895 30209
rect 24872 30172 24900 30200
rect 24044 30144 24900 30172
rect 26050 30132 26056 30184
rect 26108 30172 26114 30184
rect 27338 30172 27344 30184
rect 26108 30144 27344 30172
rect 26108 30132 26114 30144
rect 27338 30132 27344 30144
rect 27396 30172 27402 30184
rect 27525 30175 27583 30181
rect 27525 30172 27537 30175
rect 27396 30144 27537 30172
rect 27396 30132 27402 30144
rect 27525 30141 27537 30144
rect 27571 30141 27583 30175
rect 27525 30135 27583 30141
rect 28534 30132 28540 30184
rect 28592 30172 28598 30184
rect 29733 30175 29791 30181
rect 29733 30172 29745 30175
rect 28592 30144 29745 30172
rect 28592 30132 28598 30144
rect 29733 30141 29745 30144
rect 29779 30141 29791 30175
rect 29733 30135 29791 30141
rect 29914 30132 29920 30184
rect 29972 30172 29978 30184
rect 30193 30175 30251 30181
rect 30193 30172 30205 30175
rect 29972 30144 30205 30172
rect 29972 30132 29978 30144
rect 30193 30141 30205 30144
rect 30239 30172 30251 30175
rect 30466 30172 30472 30184
rect 30239 30144 30472 30172
rect 30239 30141 30251 30144
rect 30193 30135 30251 30141
rect 30466 30132 30472 30144
rect 30524 30132 30530 30184
rect 30926 30172 30932 30184
rect 30887 30144 30932 30172
rect 30926 30132 30932 30144
rect 30984 30132 30990 30184
rect 31588 30172 31616 30212
rect 31662 30200 31668 30252
rect 31720 30240 31726 30252
rect 32309 30243 32367 30249
rect 32309 30240 32321 30243
rect 31720 30212 32321 30240
rect 31720 30200 31726 30212
rect 32309 30209 32321 30212
rect 32355 30209 32367 30243
rect 32490 30240 32496 30252
rect 32451 30212 32496 30240
rect 32309 30203 32367 30209
rect 32490 30200 32496 30212
rect 32548 30200 32554 30252
rect 32950 30240 32956 30252
rect 32911 30212 32956 30240
rect 32950 30200 32956 30212
rect 33008 30200 33014 30252
rect 33042 30200 33048 30252
rect 33100 30200 33106 30252
rect 33060 30172 33088 30200
rect 31588 30144 33088 30172
rect 25774 30064 25780 30116
rect 25832 30104 25838 30116
rect 26145 30107 26203 30113
rect 26145 30104 26157 30107
rect 25832 30076 26157 30104
rect 25832 30064 25838 30076
rect 26145 30073 26157 30076
rect 26191 30073 26203 30107
rect 26145 30067 26203 30073
rect 28626 30064 28632 30116
rect 28684 30104 28690 30116
rect 28905 30107 28963 30113
rect 28905 30104 28917 30107
rect 28684 30076 28917 30104
rect 28684 30064 28690 30076
rect 28905 30073 28917 30076
rect 28951 30073 28963 30107
rect 28905 30067 28963 30073
rect 31386 30064 31392 30116
rect 31444 30104 31450 30116
rect 31444 30076 31616 30104
rect 31444 30064 31450 30076
rect 22738 30036 22744 30048
rect 19996 30008 22744 30036
rect 22738 29996 22744 30008
rect 22796 29996 22802 30048
rect 23014 29996 23020 30048
rect 23072 30036 23078 30048
rect 24213 30039 24271 30045
rect 24213 30036 24225 30039
rect 23072 30008 24225 30036
rect 23072 29996 23078 30008
rect 24213 30005 24225 30008
rect 24259 30005 24271 30039
rect 24213 29999 24271 30005
rect 27706 29996 27712 30048
rect 27764 30036 27770 30048
rect 28442 30036 28448 30048
rect 27764 30008 28448 30036
rect 27764 29996 27770 30008
rect 28442 29996 28448 30008
rect 28500 30036 28506 30048
rect 29086 30036 29092 30048
rect 28500 30008 29092 30036
rect 28500 29996 28506 30008
rect 29086 29996 29092 30008
rect 29144 29996 29150 30048
rect 31205 30039 31263 30045
rect 31205 30005 31217 30039
rect 31251 30036 31263 30039
rect 31478 30036 31484 30048
rect 31251 30008 31484 30036
rect 31251 30005 31263 30008
rect 31205 29999 31263 30005
rect 31478 29996 31484 30008
rect 31536 29996 31542 30048
rect 31588 30036 31616 30076
rect 32324 30076 32536 30104
rect 32324 30036 32352 30076
rect 31588 30008 32352 30036
rect 32508 30036 32536 30076
rect 34333 30039 34391 30045
rect 34333 30036 34345 30039
rect 32508 30008 34345 30036
rect 34333 30005 34345 30008
rect 34379 30005 34391 30039
rect 34333 29999 34391 30005
rect 1104 29946 34868 29968
rect 1104 29894 5170 29946
rect 5222 29894 5234 29946
rect 5286 29894 5298 29946
rect 5350 29894 5362 29946
rect 5414 29894 5426 29946
rect 5478 29894 13611 29946
rect 13663 29894 13675 29946
rect 13727 29894 13739 29946
rect 13791 29894 13803 29946
rect 13855 29894 13867 29946
rect 13919 29894 22052 29946
rect 22104 29894 22116 29946
rect 22168 29894 22180 29946
rect 22232 29894 22244 29946
rect 22296 29894 22308 29946
rect 22360 29894 30493 29946
rect 30545 29894 30557 29946
rect 30609 29894 30621 29946
rect 30673 29894 30685 29946
rect 30737 29894 30749 29946
rect 30801 29894 34868 29946
rect 1104 29872 34868 29894
rect 16206 29832 16212 29844
rect 16167 29804 16212 29832
rect 16206 29792 16212 29804
rect 16264 29792 16270 29844
rect 22922 29832 22928 29844
rect 16408 29804 22928 29832
rect 16408 29637 16436 29804
rect 22922 29792 22928 29804
rect 22980 29792 22986 29844
rect 23017 29835 23075 29841
rect 23017 29801 23029 29835
rect 23063 29832 23075 29835
rect 26142 29832 26148 29844
rect 23063 29804 26148 29832
rect 23063 29801 23075 29804
rect 23017 29795 23075 29801
rect 26142 29792 26148 29804
rect 26200 29792 26206 29844
rect 28626 29792 28632 29844
rect 28684 29832 28690 29844
rect 29270 29832 29276 29844
rect 28684 29804 29276 29832
rect 28684 29792 28690 29804
rect 29270 29792 29276 29804
rect 29328 29792 29334 29844
rect 29546 29792 29552 29844
rect 29604 29832 29610 29844
rect 29733 29835 29791 29841
rect 29733 29832 29745 29835
rect 29604 29804 29745 29832
rect 29604 29792 29610 29804
rect 29733 29801 29745 29804
rect 29779 29801 29791 29835
rect 34238 29832 34244 29844
rect 29733 29795 29791 29801
rect 29933 29804 34244 29832
rect 17494 29764 17500 29776
rect 17455 29736 17500 29764
rect 17494 29724 17500 29736
rect 17552 29724 17558 29776
rect 19610 29764 19616 29776
rect 17696 29736 19616 29764
rect 16393 29631 16451 29637
rect 16393 29597 16405 29631
rect 16439 29597 16451 29631
rect 16850 29628 16856 29640
rect 16811 29600 16856 29628
rect 16393 29591 16451 29597
rect 16850 29588 16856 29600
rect 16908 29588 16914 29640
rect 17221 29631 17279 29637
rect 17221 29597 17233 29631
rect 17267 29628 17279 29631
rect 17497 29631 17555 29637
rect 17497 29628 17509 29631
rect 17267 29600 17509 29628
rect 17267 29597 17279 29600
rect 17221 29591 17279 29597
rect 17497 29597 17509 29600
rect 17543 29628 17555 29631
rect 17696 29628 17724 29736
rect 19610 29724 19616 29736
rect 19668 29724 19674 29776
rect 19794 29724 19800 29776
rect 19852 29764 19858 29776
rect 20073 29767 20131 29773
rect 20073 29764 20085 29767
rect 19852 29736 20085 29764
rect 19852 29724 19858 29736
rect 20073 29733 20085 29736
rect 20119 29733 20131 29767
rect 20073 29727 20131 29733
rect 20162 29724 20168 29776
rect 20220 29764 20226 29776
rect 20220 29736 20265 29764
rect 20220 29724 20226 29736
rect 21818 29724 21824 29776
rect 21876 29764 21882 29776
rect 23845 29767 23903 29773
rect 23845 29764 23857 29767
rect 21876 29736 23857 29764
rect 21876 29724 21882 29736
rect 23845 29733 23857 29736
rect 23891 29733 23903 29767
rect 25958 29764 25964 29776
rect 25919 29736 25964 29764
rect 23845 29727 23903 29733
rect 25958 29724 25964 29736
rect 26016 29724 26022 29776
rect 27706 29764 27712 29776
rect 27667 29736 27712 29764
rect 27706 29724 27712 29736
rect 27764 29724 27770 29776
rect 18690 29696 18696 29708
rect 18524 29668 18696 29696
rect 17543 29600 17724 29628
rect 17773 29631 17831 29637
rect 17543 29597 17555 29600
rect 17497 29591 17555 29597
rect 17773 29597 17785 29631
rect 17819 29628 17831 29631
rect 17862 29628 17868 29640
rect 17819 29600 17868 29628
rect 17819 29597 17831 29600
rect 17773 29591 17831 29597
rect 17862 29588 17868 29600
rect 17920 29588 17926 29640
rect 18414 29628 18420 29640
rect 18375 29600 18420 29628
rect 18414 29588 18420 29600
rect 18472 29588 18478 29640
rect 18524 29637 18552 29668
rect 18690 29656 18696 29668
rect 18748 29656 18754 29708
rect 19518 29696 19524 29708
rect 18800 29668 19524 29696
rect 18509 29631 18567 29637
rect 18509 29597 18521 29631
rect 18555 29597 18567 29631
rect 18509 29591 18567 29597
rect 18601 29631 18659 29637
rect 18601 29597 18613 29631
rect 18647 29628 18659 29631
rect 18800 29628 18828 29668
rect 19518 29656 19524 29668
rect 19576 29656 19582 29708
rect 19803 29668 20300 29696
rect 18647 29600 18828 29628
rect 18877 29631 18935 29637
rect 18647 29597 18659 29600
rect 18601 29591 18659 29597
rect 18877 29597 18889 29631
rect 18923 29597 18935 29631
rect 18877 29591 18935 29597
rect 17586 29520 17592 29572
rect 17644 29560 17650 29572
rect 18233 29563 18291 29569
rect 18233 29560 18245 29563
rect 17644 29532 18245 29560
rect 17644 29520 17650 29532
rect 18233 29529 18245 29532
rect 18279 29529 18291 29563
rect 18233 29523 18291 29529
rect 18690 29520 18696 29572
rect 18748 29569 18754 29572
rect 18748 29563 18777 29569
rect 18765 29529 18777 29563
rect 18748 29523 18777 29529
rect 18748 29520 18754 29523
rect 16666 29492 16672 29504
rect 16627 29464 16672 29492
rect 16666 29452 16672 29464
rect 16724 29452 16730 29504
rect 17681 29495 17739 29501
rect 17681 29461 17693 29495
rect 17727 29492 17739 29495
rect 18598 29492 18604 29504
rect 17727 29464 18604 29492
rect 17727 29461 17739 29464
rect 17681 29455 17739 29461
rect 18598 29452 18604 29464
rect 18656 29452 18662 29504
rect 18892 29492 18920 29591
rect 18966 29588 18972 29640
rect 19024 29628 19030 29640
rect 19803 29628 19831 29668
rect 19024 29600 19831 29628
rect 19024 29588 19030 29600
rect 19978 29588 19984 29640
rect 20036 29628 20042 29640
rect 20272 29637 20300 29668
rect 23382 29656 23388 29708
rect 23440 29696 23446 29708
rect 24581 29699 24639 29705
rect 23440 29668 23704 29696
rect 23440 29656 23446 29668
rect 20257 29631 20315 29637
rect 20036 29600 20081 29628
rect 20036 29588 20042 29600
rect 20257 29597 20269 29631
rect 20303 29597 20315 29631
rect 20257 29591 20315 29597
rect 20809 29631 20867 29637
rect 20809 29597 20821 29631
rect 20855 29628 20867 29631
rect 20855 29600 22600 29628
rect 20855 29597 20867 29600
rect 20809 29591 20867 29597
rect 19242 29520 19248 29572
rect 19300 29560 19306 29572
rect 19797 29563 19855 29569
rect 19797 29560 19809 29563
rect 19300 29532 19809 29560
rect 19300 29520 19306 29532
rect 19797 29529 19809 29532
rect 19843 29529 19855 29563
rect 19797 29523 19855 29529
rect 21076 29563 21134 29569
rect 21076 29529 21088 29563
rect 21122 29560 21134 29563
rect 22278 29560 22284 29572
rect 21122 29532 22284 29560
rect 21122 29529 21134 29532
rect 21076 29523 21134 29529
rect 22278 29520 22284 29532
rect 22336 29520 22342 29572
rect 22572 29560 22600 29600
rect 22646 29588 22652 29640
rect 22704 29628 22710 29640
rect 22704 29600 22749 29628
rect 22704 29588 22710 29600
rect 22830 29588 22836 29640
rect 22888 29628 22894 29640
rect 23566 29628 23572 29640
rect 22888 29600 22933 29628
rect 23527 29600 23572 29628
rect 22888 29588 22894 29600
rect 23566 29588 23572 29600
rect 23624 29588 23630 29640
rect 23676 29637 23704 29668
rect 24581 29665 24593 29699
rect 24627 29696 24639 29699
rect 24854 29696 24860 29708
rect 24627 29668 24860 29696
rect 24627 29665 24639 29668
rect 24581 29659 24639 29665
rect 24854 29656 24860 29668
rect 24912 29656 24918 29708
rect 25038 29656 25044 29708
rect 25096 29696 25102 29708
rect 26053 29699 26111 29705
rect 26053 29696 26065 29699
rect 25096 29668 26065 29696
rect 25096 29656 25102 29668
rect 26053 29665 26065 29668
rect 26099 29665 26111 29699
rect 26053 29659 26111 29665
rect 27065 29699 27123 29705
rect 27065 29665 27077 29699
rect 27111 29696 27123 29699
rect 27430 29696 27436 29708
rect 27111 29668 27436 29696
rect 27111 29665 27123 29668
rect 27065 29659 27123 29665
rect 27430 29656 27436 29668
rect 27488 29656 27494 29708
rect 27982 29656 27988 29708
rect 28040 29696 28046 29708
rect 28718 29696 28724 29708
rect 28040 29668 28724 29696
rect 28040 29656 28046 29668
rect 28718 29656 28724 29668
rect 28776 29696 28782 29708
rect 28776 29668 28980 29696
rect 28776 29656 28782 29668
rect 23661 29631 23719 29637
rect 23661 29597 23673 29631
rect 23707 29597 23719 29631
rect 24762 29628 24768 29640
rect 24723 29600 24768 29628
rect 23661 29591 23719 29597
rect 24762 29588 24768 29600
rect 24820 29588 24826 29640
rect 24946 29628 24952 29640
rect 24907 29600 24952 29628
rect 24946 29588 24952 29600
rect 25004 29588 25010 29640
rect 25225 29631 25283 29637
rect 25225 29597 25237 29631
rect 25271 29628 25283 29631
rect 25590 29628 25596 29640
rect 25271 29600 25596 29628
rect 25271 29597 25283 29600
rect 25225 29591 25283 29597
rect 25590 29588 25596 29600
rect 25648 29588 25654 29640
rect 25866 29628 25872 29640
rect 25827 29600 25872 29628
rect 25866 29588 25872 29600
rect 25924 29588 25930 29640
rect 25958 29588 25964 29640
rect 26016 29628 26022 29640
rect 26145 29631 26203 29637
rect 26145 29628 26157 29631
rect 26016 29600 26157 29628
rect 26016 29588 26022 29600
rect 26145 29597 26157 29600
rect 26191 29597 26203 29631
rect 27338 29628 27344 29640
rect 27299 29600 27344 29628
rect 26145 29591 26203 29597
rect 27338 29588 27344 29600
rect 27396 29588 27402 29640
rect 27550 29631 27608 29637
rect 27550 29597 27562 29631
rect 27596 29628 27608 29631
rect 28534 29628 28540 29640
rect 27596 29600 28540 29628
rect 27596 29597 27608 29600
rect 27550 29591 27608 29597
rect 22738 29560 22744 29572
rect 22572 29532 22744 29560
rect 22738 29520 22744 29532
rect 22796 29560 22802 29572
rect 23198 29560 23204 29572
rect 22796 29532 23204 29560
rect 22796 29520 22802 29532
rect 23198 29520 23204 29532
rect 23256 29520 23262 29572
rect 24857 29563 24915 29569
rect 24857 29529 24869 29563
rect 24903 29529 24915 29563
rect 24857 29523 24915 29529
rect 25087 29563 25145 29569
rect 25087 29529 25099 29563
rect 25133 29560 25145 29563
rect 25685 29563 25743 29569
rect 25685 29560 25697 29563
rect 25133 29532 25697 29560
rect 25133 29529 25145 29532
rect 25087 29523 25145 29529
rect 25685 29529 25697 29532
rect 25731 29529 25743 29563
rect 25685 29523 25743 29529
rect 19334 29492 19340 29504
rect 18892 29464 19340 29492
rect 19334 29452 19340 29464
rect 19392 29492 19398 29504
rect 20254 29492 20260 29504
rect 19392 29464 20260 29492
rect 19392 29452 19398 29464
rect 20254 29452 20260 29464
rect 20312 29452 20318 29504
rect 22189 29495 22247 29501
rect 22189 29461 22201 29495
rect 22235 29492 22247 29495
rect 23842 29492 23848 29504
rect 22235 29464 23848 29492
rect 22235 29461 22247 29464
rect 22189 29455 22247 29461
rect 23842 29452 23848 29464
rect 23900 29452 23906 29504
rect 24872 29492 24900 29523
rect 26878 29520 26884 29572
rect 26936 29560 26942 29572
rect 27565 29560 27593 29591
rect 28534 29588 28540 29600
rect 28592 29588 28598 29640
rect 28952 29637 28980 29668
rect 28905 29631 28980 29637
rect 28813 29609 28871 29615
rect 28813 29575 28825 29609
rect 28859 29575 28871 29609
rect 28905 29597 28917 29631
rect 28951 29600 28980 29631
rect 29086 29628 29092 29640
rect 29047 29600 29092 29628
rect 28951 29597 28963 29600
rect 28905 29591 28963 29597
rect 29086 29588 29092 29600
rect 29144 29588 29150 29640
rect 29178 29588 29184 29640
rect 29236 29628 29242 29640
rect 29236 29600 29281 29628
rect 29236 29588 29242 29600
rect 29638 29588 29644 29640
rect 29696 29628 29702 29640
rect 29933 29637 29961 29804
rect 34238 29792 34244 29804
rect 34296 29792 34302 29844
rect 33226 29764 33232 29776
rect 33187 29736 33232 29764
rect 33226 29724 33232 29736
rect 33284 29724 33290 29776
rect 30098 29656 30104 29708
rect 30156 29696 30162 29708
rect 30193 29699 30251 29705
rect 30193 29696 30205 29699
rect 30156 29668 30205 29696
rect 30156 29656 30162 29668
rect 30193 29665 30205 29668
rect 30239 29665 30251 29699
rect 30193 29659 30251 29665
rect 32398 29656 32404 29708
rect 32456 29656 32462 29708
rect 32582 29656 32588 29708
rect 32640 29696 32646 29708
rect 33689 29699 33747 29705
rect 33689 29696 33701 29699
rect 32640 29668 33701 29696
rect 32640 29656 32646 29668
rect 33689 29665 33701 29668
rect 33735 29696 33747 29699
rect 34238 29696 34244 29708
rect 33735 29668 34244 29696
rect 33735 29665 33747 29668
rect 33689 29659 33747 29665
rect 34238 29656 34244 29668
rect 34296 29656 34302 29708
rect 29917 29631 29975 29637
rect 29917 29628 29929 29631
rect 29696 29600 29929 29628
rect 29696 29588 29702 29600
rect 29917 29597 29929 29600
rect 29963 29597 29975 29631
rect 29917 29591 29975 29597
rect 30009 29631 30067 29637
rect 30009 29597 30021 29631
rect 30055 29597 30067 29631
rect 30285 29631 30343 29637
rect 30285 29628 30297 29631
rect 30009 29591 30067 29597
rect 30116 29600 30297 29628
rect 28813 29572 28871 29575
rect 26936 29532 27593 29560
rect 26936 29520 26942 29532
rect 28810 29520 28816 29572
rect 28868 29560 28874 29572
rect 30024 29560 30052 29591
rect 28868 29532 30052 29560
rect 28868 29520 28874 29532
rect 25314 29492 25320 29504
rect 24872 29464 25320 29492
rect 25314 29452 25320 29464
rect 25372 29452 25378 29504
rect 25406 29452 25412 29504
rect 25464 29492 25470 29504
rect 25958 29492 25964 29504
rect 25464 29464 25964 29492
rect 25464 29452 25470 29464
rect 25958 29452 25964 29464
rect 26016 29452 26022 29504
rect 27433 29495 27491 29501
rect 27433 29461 27445 29495
rect 27479 29492 27491 29495
rect 27890 29492 27896 29504
rect 27479 29464 27896 29492
rect 27479 29461 27491 29464
rect 27433 29455 27491 29461
rect 27890 29452 27896 29464
rect 27948 29452 27954 29504
rect 28258 29452 28264 29504
rect 28316 29492 28322 29504
rect 28629 29495 28687 29501
rect 28629 29492 28641 29495
rect 28316 29464 28641 29492
rect 28316 29452 28322 29464
rect 28629 29461 28641 29464
rect 28675 29461 28687 29495
rect 28629 29455 28687 29461
rect 28718 29452 28724 29504
rect 28776 29492 28782 29504
rect 30116 29492 30144 29600
rect 30285 29597 30297 29600
rect 30331 29597 30343 29631
rect 30285 29591 30343 29597
rect 30374 29588 30380 29640
rect 30432 29628 30438 29640
rect 30929 29631 30987 29637
rect 30929 29628 30941 29631
rect 30432 29600 30941 29628
rect 30432 29588 30438 29600
rect 30929 29597 30941 29600
rect 30975 29597 30987 29631
rect 30929 29591 30987 29597
rect 31389 29631 31447 29637
rect 31389 29597 31401 29631
rect 31435 29628 31447 29631
rect 32030 29628 32036 29640
rect 31435 29600 32036 29628
rect 31435 29597 31447 29600
rect 31389 29591 31447 29597
rect 30190 29520 30196 29572
rect 30248 29560 30254 29572
rect 31404 29560 31432 29591
rect 32030 29588 32036 29600
rect 32088 29588 32094 29640
rect 32416 29628 32444 29656
rect 32140 29600 32444 29628
rect 31634 29563 31692 29569
rect 31634 29560 31646 29563
rect 30248 29532 31432 29560
rect 31496 29532 31646 29560
rect 30248 29520 30254 29532
rect 30742 29492 30748 29504
rect 28776 29464 30144 29492
rect 30703 29464 30748 29492
rect 28776 29452 28782 29464
rect 30742 29452 30748 29464
rect 30800 29452 30806 29504
rect 31110 29452 31116 29504
rect 31168 29492 31174 29504
rect 31496 29492 31524 29532
rect 31634 29529 31646 29532
rect 31680 29529 31692 29563
rect 31634 29523 31692 29529
rect 31168 29464 31524 29492
rect 31168 29452 31174 29464
rect 32030 29452 32036 29504
rect 32088 29492 32094 29504
rect 32140 29492 32168 29600
rect 33318 29588 33324 29640
rect 33376 29628 33382 29640
rect 33413 29631 33471 29637
rect 33413 29628 33425 29631
rect 33376 29600 33425 29628
rect 33376 29588 33382 29600
rect 33413 29597 33425 29600
rect 33459 29597 33471 29631
rect 33594 29628 33600 29640
rect 33555 29600 33600 29628
rect 33413 29591 33471 29597
rect 33594 29588 33600 29600
rect 33652 29588 33658 29640
rect 33778 29588 33784 29640
rect 33836 29628 33842 29640
rect 34054 29628 34060 29640
rect 33836 29600 34060 29628
rect 33836 29588 33842 29600
rect 34054 29588 34060 29600
rect 34112 29628 34118 29640
rect 34149 29631 34207 29637
rect 34149 29628 34161 29631
rect 34112 29600 34161 29628
rect 34112 29588 34118 29600
rect 34149 29597 34161 29600
rect 34195 29597 34207 29631
rect 34330 29628 34336 29640
rect 34291 29600 34336 29628
rect 34149 29591 34207 29597
rect 34330 29588 34336 29600
rect 34388 29588 34394 29640
rect 32214 29520 32220 29572
rect 32272 29560 32278 29572
rect 32272 29532 32536 29560
rect 32272 29520 32278 29532
rect 32088 29464 32168 29492
rect 32508 29492 32536 29532
rect 32766 29492 32772 29504
rect 32508 29464 32772 29492
rect 32088 29452 32094 29464
rect 32766 29452 32772 29464
rect 32824 29452 32830 29504
rect 33778 29452 33784 29504
rect 33836 29492 33842 29504
rect 34241 29495 34299 29501
rect 34241 29492 34253 29495
rect 33836 29464 34253 29492
rect 33836 29452 33842 29464
rect 34241 29461 34253 29464
rect 34287 29461 34299 29495
rect 34241 29455 34299 29461
rect 1104 29402 35027 29424
rect 1104 29350 9390 29402
rect 9442 29350 9454 29402
rect 9506 29350 9518 29402
rect 9570 29350 9582 29402
rect 9634 29350 9646 29402
rect 9698 29350 17831 29402
rect 17883 29350 17895 29402
rect 17947 29350 17959 29402
rect 18011 29350 18023 29402
rect 18075 29350 18087 29402
rect 18139 29350 26272 29402
rect 26324 29350 26336 29402
rect 26388 29350 26400 29402
rect 26452 29350 26464 29402
rect 26516 29350 26528 29402
rect 26580 29350 34713 29402
rect 34765 29350 34777 29402
rect 34829 29350 34841 29402
rect 34893 29350 34905 29402
rect 34957 29350 34969 29402
rect 35021 29350 35027 29402
rect 1104 29328 35027 29350
rect 16666 29248 16672 29300
rect 16724 29288 16730 29300
rect 20530 29288 20536 29300
rect 16724 29260 18828 29288
rect 20491 29260 20536 29288
rect 16724 29248 16730 29260
rect 18414 29220 18420 29232
rect 17328 29192 18420 29220
rect 17328 29161 17356 29192
rect 18414 29180 18420 29192
rect 18472 29180 18478 29232
rect 18800 29220 18828 29260
rect 20530 29248 20536 29260
rect 20588 29248 20594 29300
rect 20622 29248 20628 29300
rect 20680 29288 20686 29300
rect 21266 29288 21272 29300
rect 20680 29260 21272 29288
rect 20680 29248 20686 29260
rect 21266 29248 21272 29260
rect 21324 29288 21330 29300
rect 21361 29291 21419 29297
rect 21361 29288 21373 29291
rect 21324 29260 21373 29288
rect 21324 29248 21330 29260
rect 21361 29257 21373 29260
rect 21407 29257 21419 29291
rect 23566 29288 23572 29300
rect 21361 29251 21419 29257
rect 22112 29260 23572 29288
rect 19398 29223 19456 29229
rect 19398 29220 19410 29223
rect 18800 29192 19410 29220
rect 19398 29189 19410 29192
rect 19444 29189 19456 29223
rect 19398 29183 19456 29189
rect 20070 29180 20076 29232
rect 20128 29220 20134 29232
rect 20128 29192 20300 29220
rect 20128 29180 20134 29192
rect 17586 29161 17592 29164
rect 17313 29155 17371 29161
rect 17313 29121 17325 29155
rect 17359 29121 17371 29155
rect 17580 29152 17592 29161
rect 17547 29124 17592 29152
rect 17313 29115 17371 29121
rect 17580 29115 17592 29124
rect 17586 29112 17592 29115
rect 17644 29112 17650 29164
rect 18138 29112 18144 29164
rect 18196 29152 18202 29164
rect 19150 29152 19156 29164
rect 18196 29124 18368 29152
rect 19111 29124 19156 29152
rect 18196 29112 18202 29124
rect 18340 29016 18368 29124
rect 19150 29112 19156 29124
rect 19208 29112 19214 29164
rect 19242 29112 19248 29164
rect 19300 29152 19306 29164
rect 20272 29152 20300 29192
rect 20438 29180 20444 29232
rect 20496 29220 20502 29232
rect 21085 29223 21143 29229
rect 21085 29220 21097 29223
rect 20496 29192 21097 29220
rect 20496 29180 20502 29192
rect 21085 29189 21097 29192
rect 21131 29220 21143 29223
rect 21174 29220 21180 29232
rect 21131 29192 21180 29220
rect 21131 29189 21143 29192
rect 21085 29183 21143 29189
rect 21174 29180 21180 29192
rect 21232 29180 21238 29232
rect 22002 29152 22008 29164
rect 19300 29124 20208 29152
rect 20272 29124 22008 29152
rect 19300 29112 19306 29124
rect 18966 29044 18972 29096
rect 19024 29044 19030 29096
rect 20180 29084 20208 29124
rect 22002 29112 22008 29124
rect 22060 29112 22066 29164
rect 22112 29161 22140 29260
rect 23566 29248 23572 29260
rect 23624 29248 23630 29300
rect 24581 29291 24639 29297
rect 24581 29257 24593 29291
rect 24627 29288 24639 29291
rect 24670 29288 24676 29300
rect 24627 29260 24676 29288
rect 24627 29257 24639 29260
rect 24581 29251 24639 29257
rect 24670 29248 24676 29260
rect 24728 29248 24734 29300
rect 27430 29248 27436 29300
rect 27488 29248 27494 29300
rect 27706 29248 27712 29300
rect 27764 29288 27770 29300
rect 30742 29288 30748 29300
rect 27764 29260 30748 29288
rect 27764 29248 27770 29260
rect 30742 29248 30748 29260
rect 30800 29248 30806 29300
rect 31110 29288 31116 29300
rect 31071 29260 31116 29288
rect 31110 29248 31116 29260
rect 31168 29248 31174 29300
rect 31294 29248 31300 29300
rect 31352 29288 31358 29300
rect 31570 29288 31576 29300
rect 31352 29260 31576 29288
rect 31352 29248 31358 29260
rect 31570 29248 31576 29260
rect 31628 29248 31634 29300
rect 33134 29288 33140 29300
rect 31680 29260 33140 29288
rect 22373 29223 22431 29229
rect 22373 29189 22385 29223
rect 22419 29220 22431 29223
rect 24118 29220 24124 29232
rect 22419 29192 24124 29220
rect 22419 29189 22431 29192
rect 22373 29183 22431 29189
rect 24118 29180 24124 29192
rect 24176 29180 24182 29232
rect 25225 29223 25283 29229
rect 25225 29189 25237 29223
rect 25271 29220 25283 29223
rect 26418 29220 26424 29232
rect 25271 29192 26424 29220
rect 25271 29189 25283 29192
rect 25225 29183 25283 29189
rect 26418 29180 26424 29192
rect 26476 29220 26482 29232
rect 27448 29220 27476 29248
rect 26476 29192 27476 29220
rect 27632 29192 28111 29220
rect 26476 29180 26482 29192
rect 22097 29155 22155 29161
rect 22097 29121 22109 29155
rect 22143 29121 22155 29155
rect 22097 29115 22155 29121
rect 22189 29155 22247 29161
rect 22189 29121 22201 29155
rect 22235 29152 22247 29155
rect 22554 29152 22560 29164
rect 22235 29124 22560 29152
rect 22235 29121 22247 29124
rect 22189 29115 22247 29121
rect 22554 29112 22560 29124
rect 22612 29152 22618 29164
rect 22830 29152 22836 29164
rect 22612 29124 22836 29152
rect 22612 29112 22618 29124
rect 22830 29112 22836 29124
rect 22888 29112 22894 29164
rect 23474 29161 23480 29164
rect 23468 29152 23480 29161
rect 23435 29124 23480 29152
rect 23468 29115 23480 29124
rect 23474 29112 23480 29115
rect 23532 29112 23538 29164
rect 26145 29155 26203 29161
rect 26145 29121 26157 29155
rect 26191 29152 26203 29155
rect 26878 29152 26884 29164
rect 26191 29124 26884 29152
rect 26191 29121 26203 29124
rect 26145 29115 26203 29121
rect 23014 29084 23020 29096
rect 20180 29056 23020 29084
rect 23014 29044 23020 29056
rect 23072 29044 23078 29096
rect 23198 29084 23204 29096
rect 23159 29056 23204 29084
rect 23198 29044 23204 29056
rect 23256 29044 23262 29096
rect 26160 29084 26188 29115
rect 26878 29112 26884 29124
rect 26936 29112 26942 29164
rect 27246 29112 27252 29164
rect 27304 29152 27310 29164
rect 27632 29161 27660 29192
rect 27433 29155 27491 29161
rect 27433 29152 27445 29155
rect 27304 29124 27445 29152
rect 27304 29112 27310 29124
rect 27433 29121 27445 29124
rect 27479 29121 27491 29155
rect 27433 29115 27491 29121
rect 27617 29155 27675 29161
rect 27617 29121 27629 29155
rect 27663 29121 27675 29155
rect 27798 29152 27804 29164
rect 27759 29124 27804 29152
rect 27617 29115 27675 29121
rect 27798 29112 27804 29124
rect 27856 29112 27862 29164
rect 27890 29112 27896 29164
rect 27948 29152 27954 29164
rect 27985 29155 28043 29161
rect 27985 29152 27997 29155
rect 27948 29124 27997 29152
rect 27948 29112 27954 29124
rect 27985 29121 27997 29124
rect 28031 29121 28043 29155
rect 28083 29152 28111 29192
rect 28166 29180 28172 29232
rect 28224 29220 28230 29232
rect 28629 29223 28687 29229
rect 28629 29220 28641 29223
rect 28224 29192 28641 29220
rect 28224 29180 28230 29192
rect 28629 29189 28641 29192
rect 28675 29189 28687 29223
rect 28629 29183 28687 29189
rect 28810 29152 28816 29164
rect 28083 29124 28816 29152
rect 27985 29115 28043 29121
rect 28810 29112 28816 29124
rect 28868 29112 28874 29164
rect 29086 29112 29092 29164
rect 29144 29152 29150 29164
rect 30834 29152 30840 29164
rect 29144 29124 30840 29152
rect 29144 29112 29150 29124
rect 30834 29112 30840 29124
rect 30892 29152 30898 29164
rect 31110 29152 31116 29164
rect 30892 29124 31116 29152
rect 30892 29112 30898 29124
rect 31110 29112 31116 29124
rect 31168 29152 31174 29164
rect 31343 29155 31401 29161
rect 31475 29155 31481 29167
rect 31343 29152 31355 29155
rect 31168 29124 31355 29152
rect 31168 29112 31174 29124
rect 31343 29121 31355 29124
rect 31389 29121 31401 29155
rect 31436 29127 31481 29155
rect 31343 29115 31401 29121
rect 31475 29115 31481 29127
rect 31533 29115 31539 29167
rect 31573 29155 31631 29161
rect 31573 29121 31585 29155
rect 31619 29152 31631 29155
rect 31680 29152 31708 29260
rect 33134 29248 33140 29260
rect 33192 29248 33198 29300
rect 33689 29291 33747 29297
rect 33689 29257 33701 29291
rect 33735 29288 33747 29291
rect 33962 29288 33968 29300
rect 33735 29260 33968 29288
rect 33735 29257 33747 29260
rect 33689 29251 33747 29257
rect 33962 29248 33968 29260
rect 34020 29248 34026 29300
rect 31846 29180 31852 29232
rect 31904 29220 31910 29232
rect 32677 29223 32735 29229
rect 31904 29192 32628 29220
rect 31904 29180 31910 29192
rect 31619 29124 31708 29152
rect 31757 29155 31815 29161
rect 31619 29121 31631 29124
rect 31573 29115 31631 29121
rect 31757 29121 31769 29155
rect 31803 29121 31815 29155
rect 31757 29115 31815 29121
rect 27709 29087 27767 29093
rect 27709 29084 27721 29087
rect 25608 29056 26188 29084
rect 26344 29056 27721 29084
rect 18984 29016 19012 29044
rect 21818 29016 21824 29028
rect 18340 28988 19012 29016
rect 21192 28988 21824 29016
rect 18708 28957 18736 28988
rect 18693 28951 18751 28957
rect 18693 28917 18705 28951
rect 18739 28917 18751 28951
rect 18693 28911 18751 28917
rect 18966 28908 18972 28960
rect 19024 28948 19030 28960
rect 21192 28948 21220 28988
rect 21818 28976 21824 28988
rect 21876 28976 21882 29028
rect 25608 29025 25636 29056
rect 25593 29019 25651 29025
rect 25593 28985 25605 29019
rect 25639 28985 25651 29019
rect 25593 28979 25651 28985
rect 25685 29019 25743 29025
rect 25685 28985 25697 29019
rect 25731 29016 25743 29019
rect 26344 29016 26372 29056
rect 27709 29053 27721 29056
rect 27755 29084 27767 29087
rect 30098 29084 30104 29096
rect 27755 29056 30104 29084
rect 27755 29053 27767 29056
rect 27709 29047 27767 29053
rect 30098 29044 30104 29056
rect 30156 29044 30162 29096
rect 25731 28988 26372 29016
rect 25731 28985 25743 28988
rect 25685 28979 25743 28985
rect 26418 28976 26424 29028
rect 26476 29016 26482 29028
rect 26605 29019 26663 29025
rect 26476 28988 26521 29016
rect 26476 28976 26482 28988
rect 26605 28985 26617 29019
rect 26651 29016 26663 29019
rect 27890 29016 27896 29028
rect 26651 28988 27896 29016
rect 26651 28985 26663 28988
rect 26605 28979 26663 28985
rect 27890 28976 27896 28988
rect 27948 28976 27954 29028
rect 27982 28976 27988 29028
rect 28040 29016 28046 29028
rect 28169 29019 28227 29025
rect 28169 29016 28181 29019
rect 28040 28988 28181 29016
rect 28040 28976 28046 28988
rect 28169 28985 28181 28988
rect 28215 28985 28227 29019
rect 28169 28979 28227 28985
rect 29546 28976 29552 29028
rect 29604 29016 29610 29028
rect 30282 29016 30288 29028
rect 29604 28988 30288 29016
rect 29604 28976 29610 28988
rect 30282 28976 30288 28988
rect 30340 28976 30346 29028
rect 31662 28976 31668 29028
rect 31720 29016 31726 29028
rect 31772 29016 31800 29115
rect 31938 29112 31944 29164
rect 31996 29112 32002 29164
rect 32122 29112 32128 29164
rect 32180 29152 32186 29164
rect 32309 29155 32367 29161
rect 32309 29152 32321 29155
rect 32180 29124 32321 29152
rect 32180 29112 32186 29124
rect 32309 29121 32321 29124
rect 32355 29121 32367 29155
rect 32309 29115 32367 29121
rect 32398 29112 32404 29164
rect 32456 29158 32462 29164
rect 32493 29158 32551 29161
rect 32456 29155 32551 29158
rect 32456 29130 32505 29155
rect 32456 29112 32462 29130
rect 32493 29121 32505 29130
rect 32539 29121 32551 29155
rect 32600 29152 32628 29192
rect 32677 29189 32689 29223
rect 32723 29220 32735 29223
rect 32723 29192 32904 29220
rect 32723 29189 32735 29192
rect 32677 29183 32735 29189
rect 32769 29155 32827 29161
rect 32769 29152 32781 29155
rect 32600 29150 32711 29152
rect 32768 29150 32781 29152
rect 32600 29124 32781 29150
rect 32683 29122 32781 29124
rect 32493 29115 32551 29121
rect 32769 29121 32781 29122
rect 32815 29121 32827 29155
rect 32876 29152 32904 29192
rect 33042 29152 33048 29164
rect 32876 29124 33048 29152
rect 32769 29115 32827 29121
rect 33042 29112 33048 29124
rect 33100 29112 33106 29164
rect 33318 29112 33324 29164
rect 33376 29152 33382 29164
rect 33505 29155 33563 29161
rect 33505 29152 33517 29155
rect 33376 29124 33517 29152
rect 33376 29112 33382 29124
rect 33505 29121 33517 29124
rect 33551 29121 33563 29155
rect 33778 29152 33784 29164
rect 33739 29124 33784 29152
rect 33505 29115 33563 29121
rect 33778 29112 33784 29124
rect 33836 29112 33842 29164
rect 31956 29084 31984 29112
rect 31956 29056 32444 29084
rect 32416 29028 32444 29056
rect 31720 28988 31800 29016
rect 31720 28976 31726 28988
rect 32398 28976 32404 29028
rect 32456 28976 32462 29028
rect 33226 28976 33232 29028
rect 33284 29016 33290 29028
rect 33321 29019 33379 29025
rect 33321 29016 33333 29019
rect 33284 28988 33333 29016
rect 33284 28976 33290 28988
rect 33321 28985 33333 28988
rect 33367 28985 33379 29019
rect 34330 29016 34336 29028
rect 33321 28979 33379 28985
rect 33428 28988 34336 29016
rect 19024 28920 21220 28948
rect 19024 28908 19030 28920
rect 21266 28908 21272 28960
rect 21324 28948 21330 28960
rect 23382 28948 23388 28960
rect 21324 28920 23388 28948
rect 21324 28908 21330 28920
rect 23382 28908 23388 28920
rect 23440 28908 23446 28960
rect 23474 28908 23480 28960
rect 23532 28948 23538 28960
rect 28074 28948 28080 28960
rect 23532 28920 28080 28948
rect 23532 28908 23538 28920
rect 28074 28908 28080 28920
rect 28132 28908 28138 28960
rect 28442 28908 28448 28960
rect 28500 28948 28506 28960
rect 29178 28948 29184 28960
rect 28500 28920 29184 28948
rect 28500 28908 28506 28920
rect 29178 28908 29184 28920
rect 29236 28908 29242 28960
rect 29730 28908 29736 28960
rect 29788 28948 29794 28960
rect 29917 28951 29975 28957
rect 29917 28948 29929 28951
rect 29788 28920 29929 28948
rect 29788 28908 29794 28920
rect 29917 28917 29929 28920
rect 29963 28948 29975 28951
rect 30190 28948 30196 28960
rect 29963 28920 30196 28948
rect 29963 28917 29975 28920
rect 29917 28911 29975 28917
rect 30190 28908 30196 28920
rect 30248 28908 30254 28960
rect 31570 28908 31576 28960
rect 31628 28948 31634 28960
rect 33428 28948 33456 28988
rect 34330 28976 34336 28988
rect 34388 28976 34394 29028
rect 31628 28920 33456 28948
rect 31628 28908 31634 28920
rect 1104 28858 34868 28880
rect 1104 28806 5170 28858
rect 5222 28806 5234 28858
rect 5286 28806 5298 28858
rect 5350 28806 5362 28858
rect 5414 28806 5426 28858
rect 5478 28806 13611 28858
rect 13663 28806 13675 28858
rect 13727 28806 13739 28858
rect 13791 28806 13803 28858
rect 13855 28806 13867 28858
rect 13919 28806 22052 28858
rect 22104 28806 22116 28858
rect 22168 28806 22180 28858
rect 22232 28806 22244 28858
rect 22296 28806 22308 28858
rect 22360 28806 30493 28858
rect 30545 28806 30557 28858
rect 30609 28806 30621 28858
rect 30673 28806 30685 28858
rect 30737 28806 30749 28858
rect 30801 28806 34868 28858
rect 1104 28784 34868 28806
rect 16117 28747 16175 28753
rect 16117 28713 16129 28747
rect 16163 28744 16175 28747
rect 21266 28744 21272 28756
rect 16163 28716 21272 28744
rect 16163 28713 16175 28716
rect 16117 28707 16175 28713
rect 21266 28704 21272 28716
rect 21324 28704 21330 28756
rect 22281 28747 22339 28753
rect 22281 28713 22293 28747
rect 22327 28744 22339 28747
rect 22370 28744 22376 28756
rect 22327 28716 22376 28744
rect 22327 28713 22339 28716
rect 22281 28707 22339 28713
rect 22370 28704 22376 28716
rect 22428 28704 22434 28756
rect 25958 28744 25964 28756
rect 25919 28716 25964 28744
rect 25958 28704 25964 28716
rect 26016 28704 26022 28756
rect 27338 28704 27344 28756
rect 27396 28744 27402 28756
rect 27798 28744 27804 28756
rect 27396 28716 27804 28744
rect 27396 28704 27402 28716
rect 27798 28704 27804 28716
rect 27856 28704 27862 28756
rect 28994 28704 29000 28756
rect 29052 28744 29058 28756
rect 31938 28744 31944 28756
rect 29052 28716 31944 28744
rect 29052 28704 29058 28716
rect 31938 28704 31944 28716
rect 31996 28704 32002 28756
rect 32122 28704 32128 28756
rect 32180 28744 32186 28756
rect 32858 28744 32864 28756
rect 32180 28716 32864 28744
rect 32180 28704 32186 28716
rect 32858 28704 32864 28716
rect 32916 28704 32922 28756
rect 33870 28744 33876 28756
rect 33831 28716 33876 28744
rect 33870 28704 33876 28716
rect 33928 28704 33934 28756
rect 17405 28679 17463 28685
rect 17405 28645 17417 28679
rect 17451 28676 17463 28679
rect 18782 28676 18788 28688
rect 17451 28648 18788 28676
rect 17451 28645 17463 28648
rect 17405 28639 17463 28645
rect 18782 28636 18788 28648
rect 18840 28636 18846 28688
rect 22738 28636 22744 28688
rect 22796 28676 22802 28688
rect 23845 28679 23903 28685
rect 23845 28676 23857 28679
rect 22796 28648 23857 28676
rect 22796 28636 22802 28648
rect 23845 28645 23857 28648
rect 23891 28645 23903 28679
rect 23845 28639 23903 28645
rect 28828 28648 29592 28676
rect 19242 28608 19248 28620
rect 16960 28580 19248 28608
rect 16298 28540 16304 28552
rect 16259 28512 16304 28540
rect 16298 28500 16304 28512
rect 16356 28500 16362 28552
rect 16960 28549 16988 28580
rect 19242 28568 19248 28580
rect 19300 28568 19306 28620
rect 19797 28611 19855 28617
rect 19797 28608 19809 28611
rect 19352 28580 19809 28608
rect 16945 28543 17003 28549
rect 16945 28509 16957 28543
rect 16991 28509 17003 28543
rect 17586 28540 17592 28552
rect 17547 28512 17592 28540
rect 16945 28503 17003 28509
rect 17586 28500 17592 28512
rect 17644 28500 17650 28552
rect 18138 28540 18144 28552
rect 18099 28512 18144 28540
rect 18138 28500 18144 28512
rect 18196 28500 18202 28552
rect 18233 28543 18291 28549
rect 18233 28509 18245 28543
rect 18279 28540 18291 28543
rect 18279 28512 18644 28540
rect 18279 28509 18291 28512
rect 18233 28503 18291 28509
rect 17126 28432 17132 28484
rect 17184 28472 17190 28484
rect 18417 28475 18475 28481
rect 18417 28472 18429 28475
rect 17184 28444 18429 28472
rect 17184 28432 17190 28444
rect 18417 28441 18429 28444
rect 18463 28441 18475 28475
rect 18417 28435 18475 28441
rect 18616 28416 18644 28512
rect 18966 28500 18972 28552
rect 19024 28540 19030 28552
rect 19352 28540 19380 28580
rect 19797 28577 19809 28580
rect 19843 28577 19855 28611
rect 19797 28571 19855 28577
rect 23198 28568 23204 28620
rect 23256 28608 23262 28620
rect 28828 28617 28856 28648
rect 28813 28611 28871 28617
rect 23256 28580 24624 28608
rect 23256 28568 23262 28580
rect 24596 28552 24624 28580
rect 28813 28577 28825 28611
rect 28859 28577 28871 28611
rect 28813 28571 28871 28577
rect 28994 28568 29000 28620
rect 29052 28608 29058 28620
rect 29564 28608 29592 28648
rect 31110 28636 31116 28688
rect 31168 28676 31174 28688
rect 33318 28676 33324 28688
rect 31168 28648 33324 28676
rect 31168 28636 31174 28648
rect 33318 28636 33324 28648
rect 33376 28636 33382 28688
rect 29052 28580 29097 28608
rect 29564 28580 29868 28608
rect 29052 28568 29058 28580
rect 29840 28552 29868 28580
rect 31846 28568 31852 28620
rect 31904 28608 31910 28620
rect 32769 28611 32827 28617
rect 32769 28608 32781 28611
rect 31904 28580 32781 28608
rect 31904 28568 31910 28580
rect 32769 28577 32781 28580
rect 32815 28577 32827 28611
rect 32769 28571 32827 28577
rect 32953 28611 33011 28617
rect 32953 28577 32965 28611
rect 32999 28608 33011 28611
rect 33505 28611 33563 28617
rect 33505 28608 33517 28611
rect 32999 28580 33517 28608
rect 32999 28577 33011 28580
rect 32953 28571 33011 28577
rect 33505 28577 33517 28580
rect 33551 28577 33563 28611
rect 33505 28571 33563 28577
rect 19518 28540 19524 28552
rect 19024 28512 19380 28540
rect 19479 28512 19524 28540
rect 19024 28500 19030 28512
rect 19518 28500 19524 28512
rect 19576 28500 19582 28552
rect 19613 28543 19671 28549
rect 19613 28509 19625 28543
rect 19659 28540 19671 28543
rect 24026 28540 24032 28552
rect 19659 28512 19748 28540
rect 23987 28512 24032 28540
rect 19659 28509 19671 28512
rect 19613 28503 19671 28509
rect 16758 28404 16764 28416
rect 16719 28376 16764 28404
rect 16758 28364 16764 28376
rect 16816 28364 16822 28416
rect 18598 28364 18604 28416
rect 18656 28364 18662 28416
rect 19058 28364 19064 28416
rect 19116 28404 19122 28416
rect 19720 28404 19748 28512
rect 24026 28500 24032 28512
rect 24084 28500 24090 28552
rect 24578 28540 24584 28552
rect 24539 28512 24584 28540
rect 24578 28500 24584 28512
rect 24636 28500 24642 28552
rect 24854 28549 24860 28552
rect 24848 28540 24860 28549
rect 24815 28512 24860 28540
rect 24848 28503 24860 28512
rect 24854 28500 24860 28503
rect 24912 28500 24918 28552
rect 26050 28500 26056 28552
rect 26108 28540 26114 28552
rect 26694 28549 26700 28552
rect 26421 28543 26479 28549
rect 26421 28540 26433 28543
rect 26108 28512 26433 28540
rect 26108 28500 26114 28512
rect 26421 28509 26433 28512
rect 26467 28509 26479 28543
rect 26421 28503 26479 28509
rect 26688 28503 26700 28549
rect 26752 28540 26758 28552
rect 28905 28543 28963 28549
rect 26752 28512 26788 28540
rect 26694 28500 26700 28503
rect 26752 28500 26758 28512
rect 28905 28509 28917 28543
rect 28951 28509 28963 28543
rect 29086 28540 29092 28552
rect 29047 28512 29092 28540
rect 28905 28503 28963 28509
rect 20806 28472 20812 28484
rect 20767 28444 20812 28472
rect 20806 28432 20812 28444
rect 20864 28432 20870 28484
rect 22094 28432 22100 28484
rect 22152 28472 22158 28484
rect 22554 28472 22560 28484
rect 22152 28444 22560 28472
rect 22152 28432 22158 28444
rect 22554 28432 22560 28444
rect 22612 28432 22618 28484
rect 23017 28475 23075 28481
rect 23017 28441 23029 28475
rect 23063 28472 23075 28475
rect 23106 28472 23112 28484
rect 23063 28444 23112 28472
rect 23063 28441 23075 28444
rect 23017 28435 23075 28441
rect 23106 28432 23112 28444
rect 23164 28432 23170 28484
rect 23201 28475 23259 28481
rect 23201 28441 23213 28475
rect 23247 28472 23259 28475
rect 24394 28472 24400 28484
rect 23247 28444 24400 28472
rect 23247 28441 23259 28444
rect 23201 28435 23259 28441
rect 24394 28432 24400 28444
rect 24452 28432 24458 28484
rect 28920 28472 28948 28503
rect 29086 28500 29092 28512
rect 29144 28500 29150 28552
rect 29730 28540 29736 28552
rect 29691 28512 29736 28540
rect 29730 28500 29736 28512
rect 29788 28500 29794 28552
rect 29822 28500 29828 28552
rect 29880 28500 29886 28552
rect 30282 28500 30288 28552
rect 30340 28540 30346 28552
rect 31573 28543 31631 28549
rect 31573 28540 31585 28543
rect 30340 28512 31585 28540
rect 30340 28500 30346 28512
rect 31573 28509 31585 28512
rect 31619 28509 31631 28543
rect 32677 28543 32735 28549
rect 32677 28540 32689 28543
rect 31573 28503 31631 28509
rect 32232 28512 32689 28540
rect 29178 28472 29184 28484
rect 28920 28444 29184 28472
rect 29178 28432 29184 28444
rect 29236 28472 29242 28484
rect 29638 28472 29644 28484
rect 29236 28444 29644 28472
rect 29236 28432 29242 28444
rect 29638 28432 29644 28444
rect 29696 28432 29702 28484
rect 30006 28481 30012 28484
rect 30000 28435 30012 28481
rect 30064 28472 30070 28484
rect 30064 28444 30100 28472
rect 30006 28432 30012 28435
rect 30064 28432 30070 28444
rect 31478 28432 31484 28484
rect 31536 28472 31542 28484
rect 32232 28472 32260 28512
rect 32677 28509 32689 28512
rect 32723 28509 32735 28543
rect 32677 28503 32735 28509
rect 32858 28500 32864 28552
rect 32916 28540 32922 28552
rect 33597 28543 33655 28549
rect 33597 28540 33609 28543
rect 32916 28512 33609 28540
rect 32916 28500 32922 28512
rect 33597 28509 33609 28512
rect 33643 28509 33655 28543
rect 33597 28503 33655 28509
rect 31536 28444 32260 28472
rect 31536 28432 31542 28444
rect 19116 28376 19748 28404
rect 19116 28364 19122 28376
rect 21174 28364 21180 28416
rect 21232 28404 21238 28416
rect 22922 28404 22928 28416
rect 21232 28376 22928 28404
rect 21232 28364 21238 28376
rect 22922 28364 22928 28376
rect 22980 28364 22986 28416
rect 23385 28407 23443 28413
rect 23385 28373 23397 28407
rect 23431 28404 23443 28407
rect 23474 28404 23480 28416
rect 23431 28376 23480 28404
rect 23431 28373 23443 28376
rect 23385 28367 23443 28373
rect 23474 28364 23480 28376
rect 23532 28364 23538 28416
rect 24486 28364 24492 28416
rect 24544 28404 24550 28416
rect 27246 28404 27252 28416
rect 24544 28376 27252 28404
rect 24544 28364 24550 28376
rect 27246 28364 27252 28376
rect 27304 28404 27310 28416
rect 28442 28404 28448 28416
rect 27304 28376 28448 28404
rect 27304 28364 27310 28376
rect 28442 28364 28448 28376
rect 28500 28364 28506 28416
rect 28629 28407 28687 28413
rect 28629 28373 28641 28407
rect 28675 28404 28687 28407
rect 29546 28404 29552 28416
rect 28675 28376 29552 28404
rect 28675 28373 28687 28376
rect 28629 28367 28687 28373
rect 29546 28364 29552 28376
rect 29604 28364 29610 28416
rect 29822 28364 29828 28416
rect 29880 28404 29886 28416
rect 30098 28404 30104 28416
rect 29880 28376 30104 28404
rect 29880 28364 29886 28376
rect 30098 28364 30104 28376
rect 30156 28404 30162 28416
rect 30834 28404 30840 28416
rect 30156 28376 30840 28404
rect 30156 28364 30162 28376
rect 30834 28364 30840 28376
rect 30892 28404 30898 28416
rect 31113 28407 31171 28413
rect 31113 28404 31125 28407
rect 30892 28376 31125 28404
rect 30892 28364 30898 28376
rect 31113 28373 31125 28376
rect 31159 28373 31171 28407
rect 31113 28367 31171 28373
rect 31757 28407 31815 28413
rect 31757 28373 31769 28407
rect 31803 28404 31815 28407
rect 32122 28404 32128 28416
rect 31803 28376 32128 28404
rect 31803 28373 31815 28376
rect 31757 28367 31815 28373
rect 32122 28364 32128 28376
rect 32180 28364 32186 28416
rect 32232 28404 32260 28444
rect 32309 28475 32367 28481
rect 32309 28441 32321 28475
rect 32355 28472 32367 28475
rect 33778 28472 33784 28484
rect 32355 28444 33784 28472
rect 32355 28441 32367 28444
rect 32309 28435 32367 28441
rect 33778 28432 33784 28444
rect 33836 28432 33842 28484
rect 33594 28404 33600 28416
rect 32232 28376 33600 28404
rect 33594 28364 33600 28376
rect 33652 28364 33658 28416
rect 1104 28314 35027 28336
rect 1104 28262 9390 28314
rect 9442 28262 9454 28314
rect 9506 28262 9518 28314
rect 9570 28262 9582 28314
rect 9634 28262 9646 28314
rect 9698 28262 17831 28314
rect 17883 28262 17895 28314
rect 17947 28262 17959 28314
rect 18011 28262 18023 28314
rect 18075 28262 18087 28314
rect 18139 28262 26272 28314
rect 26324 28262 26336 28314
rect 26388 28262 26400 28314
rect 26452 28262 26464 28314
rect 26516 28262 26528 28314
rect 26580 28262 34713 28314
rect 34765 28262 34777 28314
rect 34829 28262 34841 28314
rect 34893 28262 34905 28314
rect 34957 28262 34969 28314
rect 35021 28262 35027 28314
rect 1104 28240 35027 28262
rect 16758 28160 16764 28212
rect 16816 28200 16822 28212
rect 20162 28200 20168 28212
rect 16816 28172 20168 28200
rect 16816 28160 16822 28172
rect 20162 28160 20168 28172
rect 20220 28160 20226 28212
rect 20622 28200 20628 28212
rect 20272 28172 20628 28200
rect 17589 28135 17647 28141
rect 17589 28101 17601 28135
rect 17635 28132 17647 28135
rect 17678 28132 17684 28144
rect 17635 28104 17684 28132
rect 17635 28101 17647 28104
rect 17589 28095 17647 28101
rect 17678 28092 17684 28104
rect 17736 28092 17742 28144
rect 18414 28092 18420 28144
rect 18472 28132 18478 28144
rect 19150 28132 19156 28144
rect 18472 28104 19156 28132
rect 18472 28092 18478 28104
rect 16114 28064 16120 28076
rect 16075 28036 16120 28064
rect 16114 28024 16120 28036
rect 16172 28024 16178 28076
rect 16301 28067 16359 28073
rect 16301 28033 16313 28067
rect 16347 28064 16359 28067
rect 17034 28064 17040 28076
rect 16347 28036 17040 28064
rect 16347 28033 16359 28036
rect 16301 28027 16359 28033
rect 17034 28024 17040 28036
rect 17092 28024 17098 28076
rect 17126 28024 17132 28076
rect 17184 28064 17190 28076
rect 18524 28073 18552 28104
rect 19150 28092 19156 28104
rect 19208 28092 19214 28144
rect 20272 28132 20300 28172
rect 20622 28160 20628 28172
rect 20680 28160 20686 28212
rect 23290 28200 23296 28212
rect 21284 28172 23296 28200
rect 20438 28132 20444 28144
rect 19260 28104 20300 28132
rect 20399 28104 20444 28132
rect 18509 28067 18567 28073
rect 17184 28036 17229 28064
rect 17184 28024 17190 28036
rect 18509 28033 18521 28067
rect 18555 28033 18567 28067
rect 18765 28067 18823 28073
rect 18765 28064 18777 28067
rect 18509 28027 18567 28033
rect 18616 28036 18777 28064
rect 18616 27996 18644 28036
rect 18765 28033 18777 28036
rect 18811 28033 18823 28067
rect 18765 28027 18823 28033
rect 19058 28024 19064 28076
rect 19116 28064 19122 28076
rect 19260 28064 19288 28104
rect 20438 28092 20444 28104
rect 20496 28092 20502 28144
rect 21284 28132 21312 28172
rect 23290 28160 23296 28172
rect 23348 28160 23354 28212
rect 23477 28203 23535 28209
rect 23477 28169 23489 28203
rect 23523 28200 23535 28203
rect 23566 28200 23572 28212
rect 23523 28172 23572 28200
rect 23523 28169 23535 28172
rect 23477 28163 23535 28169
rect 23566 28160 23572 28172
rect 23624 28160 23630 28212
rect 26050 28200 26056 28212
rect 24596 28172 26056 28200
rect 22462 28132 22468 28144
rect 21192 28104 21312 28132
rect 22112 28104 22468 28132
rect 21192 28073 21220 28104
rect 19116 28036 19288 28064
rect 21177 28067 21235 28073
rect 19116 28024 19122 28036
rect 21177 28033 21189 28067
rect 21223 28033 21235 28067
rect 21177 28027 21235 28033
rect 21269 28067 21327 28073
rect 21269 28033 21281 28067
rect 21315 28064 21327 28067
rect 22002 28064 22008 28076
rect 21315 28036 22008 28064
rect 21315 28033 21327 28036
rect 21269 28027 21327 28033
rect 17788 27968 18644 27996
rect 20625 27999 20683 28005
rect 16945 27931 17003 27937
rect 16945 27897 16957 27931
rect 16991 27928 17003 27931
rect 17788 27928 17816 27968
rect 20625 27965 20637 27999
rect 20671 27996 20683 27999
rect 21284 27996 21312 28027
rect 22002 28024 22008 28036
rect 22060 28024 22066 28076
rect 22112 28073 22140 28104
rect 22462 28092 22468 28104
rect 22520 28132 22526 28144
rect 23198 28132 23204 28144
rect 22520 28104 23204 28132
rect 22520 28092 22526 28104
rect 23198 28092 23204 28104
rect 23256 28092 23262 28144
rect 22097 28067 22155 28073
rect 22097 28033 22109 28067
rect 22143 28033 22155 28067
rect 22353 28067 22411 28073
rect 22353 28064 22365 28067
rect 22097 28027 22155 28033
rect 22204 28036 22365 28064
rect 22204 27996 22232 28036
rect 22353 28033 22365 28036
rect 22399 28033 22411 28067
rect 24118 28064 24124 28076
rect 24079 28036 24124 28064
rect 22353 28027 22411 28033
rect 24118 28024 24124 28036
rect 24176 28024 24182 28076
rect 24596 28073 24624 28172
rect 26050 28160 26056 28172
rect 26108 28160 26114 28212
rect 27062 28160 27068 28212
rect 27120 28200 27126 28212
rect 27525 28203 27583 28209
rect 27525 28200 27537 28203
rect 27120 28172 27537 28200
rect 27120 28160 27126 28172
rect 27525 28169 27537 28172
rect 27571 28169 27583 28203
rect 27525 28163 27583 28169
rect 30926 28160 30932 28212
rect 30984 28200 30990 28212
rect 31205 28203 31263 28209
rect 31205 28200 31217 28203
rect 30984 28172 31217 28200
rect 30984 28160 30990 28172
rect 31205 28169 31217 28172
rect 31251 28169 31263 28203
rect 31205 28163 31263 28169
rect 31662 28160 31668 28212
rect 31720 28200 31726 28212
rect 34054 28200 34060 28212
rect 31720 28172 34060 28200
rect 31720 28160 31726 28172
rect 34054 28160 34060 28172
rect 34112 28160 34118 28212
rect 25038 28092 25044 28144
rect 25096 28132 25102 28144
rect 28810 28132 28816 28144
rect 25096 28104 28816 28132
rect 25096 28092 25102 28104
rect 28810 28092 28816 28104
rect 28868 28092 28874 28144
rect 29638 28132 29644 28144
rect 29472 28104 29644 28132
rect 24581 28067 24639 28073
rect 24581 28033 24593 28067
rect 24627 28033 24639 28067
rect 24837 28067 24895 28073
rect 24837 28064 24849 28067
rect 24581 28027 24639 28033
rect 24688 28036 24849 28064
rect 20671 27968 21312 27996
rect 21376 27968 22232 27996
rect 20671 27965 20683 27968
rect 20625 27959 20683 27965
rect 16991 27900 17816 27928
rect 17957 27931 18015 27937
rect 16991 27897 17003 27900
rect 16945 27891 17003 27897
rect 17957 27897 17969 27931
rect 18003 27928 18015 27931
rect 18230 27928 18236 27940
rect 18003 27900 18236 27928
rect 18003 27897 18015 27900
rect 17957 27891 18015 27897
rect 16117 27863 16175 27869
rect 16117 27829 16129 27863
rect 16163 27860 16175 27863
rect 16298 27860 16304 27872
rect 16163 27832 16304 27860
rect 16163 27829 16175 27832
rect 16117 27823 16175 27829
rect 16298 27820 16304 27832
rect 16356 27820 16362 27872
rect 17402 27820 17408 27872
rect 17460 27860 17466 27872
rect 17972 27860 18000 27891
rect 18230 27888 18236 27900
rect 18288 27888 18294 27940
rect 20162 27888 20168 27940
rect 20220 27928 20226 27940
rect 21376 27928 21404 27968
rect 23382 27956 23388 28008
rect 23440 27996 23446 28008
rect 24688 27996 24716 28036
rect 24837 28033 24849 28036
rect 24883 28033 24895 28067
rect 24837 28027 24895 28033
rect 26142 28024 26148 28076
rect 26200 28064 26206 28076
rect 26605 28067 26663 28073
rect 26605 28064 26617 28067
rect 26200 28036 26617 28064
rect 26200 28024 26206 28036
rect 26605 28033 26617 28036
rect 26651 28033 26663 28067
rect 26605 28027 26663 28033
rect 27341 28067 27399 28073
rect 27341 28033 27353 28067
rect 27387 28064 27399 28067
rect 27522 28064 27528 28076
rect 27387 28036 27528 28064
rect 27387 28033 27399 28036
rect 27341 28027 27399 28033
rect 27522 28024 27528 28036
rect 27580 28024 27586 28076
rect 28445 28067 28503 28073
rect 28445 28033 28457 28067
rect 28491 28033 28503 28067
rect 28445 28027 28503 28033
rect 27154 27996 27160 28008
rect 23440 27968 24716 27996
rect 27115 27968 27160 27996
rect 23440 27956 23446 27968
rect 27154 27956 27160 27968
rect 27212 27956 27218 28008
rect 28350 27996 28356 28008
rect 28311 27968 28356 27996
rect 28350 27956 28356 27968
rect 28408 27956 28414 28008
rect 24486 27928 24492 27940
rect 20220 27900 21404 27928
rect 23492 27900 24492 27928
rect 20220 27888 20226 27900
rect 17460 27832 18000 27860
rect 18049 27863 18107 27869
rect 17460 27820 17466 27832
rect 18049 27829 18061 27863
rect 18095 27860 18107 27863
rect 18414 27860 18420 27872
rect 18095 27832 18420 27860
rect 18095 27829 18107 27832
rect 18049 27823 18107 27829
rect 18414 27820 18420 27832
rect 18472 27820 18478 27872
rect 18506 27820 18512 27872
rect 18564 27860 18570 27872
rect 19889 27863 19947 27869
rect 19889 27860 19901 27863
rect 18564 27832 19901 27860
rect 18564 27820 18570 27832
rect 19889 27829 19901 27832
rect 19935 27829 19947 27863
rect 19889 27823 19947 27829
rect 21453 27863 21511 27869
rect 21453 27829 21465 27863
rect 21499 27860 21511 27863
rect 22370 27860 22376 27872
rect 21499 27832 22376 27860
rect 21499 27829 21511 27832
rect 21453 27823 21511 27829
rect 22370 27820 22376 27832
rect 22428 27820 22434 27872
rect 22830 27820 22836 27872
rect 22888 27860 22894 27872
rect 23492 27860 23520 27900
rect 24486 27888 24492 27900
rect 24544 27888 24550 27940
rect 25590 27888 25596 27940
rect 25648 27928 25654 27940
rect 26421 27931 26479 27937
rect 25648 27900 26096 27928
rect 25648 27888 25654 27900
rect 22888 27832 23520 27860
rect 22888 27820 22894 27832
rect 23566 27820 23572 27872
rect 23624 27860 23630 27872
rect 23937 27863 23995 27869
rect 23937 27860 23949 27863
rect 23624 27832 23949 27860
rect 23624 27820 23630 27832
rect 23937 27829 23949 27832
rect 23983 27829 23995 27863
rect 23937 27823 23995 27829
rect 24946 27820 24952 27872
rect 25004 27860 25010 27872
rect 25961 27863 26019 27869
rect 25961 27860 25973 27863
rect 25004 27832 25973 27860
rect 25004 27820 25010 27832
rect 25961 27829 25973 27832
rect 26007 27829 26019 27863
rect 26068 27860 26096 27900
rect 26421 27897 26433 27931
rect 26467 27928 26479 27931
rect 26878 27928 26884 27940
rect 26467 27900 26884 27928
rect 26467 27897 26479 27900
rect 26421 27891 26479 27897
rect 26878 27888 26884 27900
rect 26936 27888 26942 27940
rect 28074 27860 28080 27872
rect 26068 27832 28080 27860
rect 25961 27823 26019 27829
rect 28074 27820 28080 27832
rect 28132 27820 28138 27872
rect 28460 27860 28488 28027
rect 28994 28024 29000 28076
rect 29052 28064 29058 28076
rect 29273 28067 29331 28073
rect 29472 28071 29500 28104
rect 29638 28092 29644 28104
rect 29696 28092 29702 28144
rect 30006 28092 30012 28144
rect 30064 28132 30070 28144
rect 31018 28132 31024 28144
rect 30064 28104 30109 28132
rect 30484 28104 31024 28132
rect 30064 28092 30070 28104
rect 29273 28064 29285 28067
rect 29052 28036 29285 28064
rect 29052 28024 29058 28036
rect 29273 28033 29285 28036
rect 29319 28033 29331 28067
rect 29273 28027 29331 28033
rect 29457 28065 29515 28071
rect 29457 28031 29469 28065
rect 29503 28031 29515 28065
rect 29457 28025 29515 28031
rect 29543 28067 29601 28073
rect 29543 28033 29555 28067
rect 29589 28033 29601 28067
rect 29543 28027 29601 28033
rect 28813 27999 28871 28005
rect 28813 27965 28825 27999
rect 28859 27996 28871 27999
rect 29086 27996 29092 28008
rect 28859 27968 29092 27996
rect 28859 27965 28871 27968
rect 28813 27959 28871 27965
rect 29086 27956 29092 27968
rect 29144 27956 29150 28008
rect 29564 27872 29592 28027
rect 29822 28024 29828 28076
rect 29880 28073 29886 28076
rect 30484 28073 30512 28104
rect 31018 28092 31024 28104
rect 31076 28092 31082 28144
rect 29880 28067 29894 28073
rect 29882 28064 29894 28067
rect 30469 28067 30527 28073
rect 29882 28036 29925 28064
rect 29882 28033 29894 28036
rect 29880 28027 29894 28033
rect 30469 28033 30481 28067
rect 30515 28033 30527 28067
rect 30469 28027 30527 28033
rect 30653 28067 30711 28073
rect 30653 28033 30665 28067
rect 30699 28033 30711 28067
rect 30653 28027 30711 28033
rect 30745 28067 30803 28073
rect 30745 28033 30757 28067
rect 30791 28064 30803 28067
rect 31110 28064 31116 28076
rect 30791 28036 31116 28064
rect 30791 28033 30803 28036
rect 30745 28027 30803 28033
rect 29880 28024 29886 28027
rect 29638 27956 29644 28008
rect 29696 27996 29702 28008
rect 30668 27996 30696 28027
rect 31110 28024 31116 28036
rect 31168 28024 31174 28076
rect 31481 28067 31539 28073
rect 31481 28033 31493 28067
rect 31527 28064 31539 28067
rect 31680 28064 31708 28160
rect 32674 28132 32680 28144
rect 32635 28104 32680 28132
rect 32674 28092 32680 28104
rect 32732 28092 32738 28144
rect 32490 28064 32496 28076
rect 31527 28036 31708 28064
rect 32451 28036 32496 28064
rect 31527 28033 31539 28036
rect 31481 28027 31539 28033
rect 32490 28024 32496 28036
rect 32548 28024 32554 28076
rect 30926 27996 30932 28008
rect 29696 27968 29741 27996
rect 30668 27968 30932 27996
rect 29696 27956 29702 27968
rect 30926 27956 30932 27968
rect 30984 27956 30990 28008
rect 31389 27999 31447 28005
rect 31389 27965 31401 27999
rect 31435 27965 31447 27999
rect 31570 27996 31576 28008
rect 31531 27968 31576 27996
rect 31389 27959 31447 27965
rect 31404 27928 31432 27959
rect 31570 27956 31576 27968
rect 31628 27956 31634 28008
rect 31665 27999 31723 28005
rect 31665 27965 31677 27999
rect 31711 27996 31723 27999
rect 32398 27996 32404 28008
rect 31711 27968 32404 27996
rect 31711 27965 31723 27968
rect 31665 27959 31723 27965
rect 32398 27956 32404 27968
rect 32456 27956 32462 28008
rect 34330 27996 34336 28008
rect 34291 27968 34336 27996
rect 34330 27956 34336 27968
rect 34388 27956 34394 28008
rect 32858 27928 32864 27940
rect 31404 27900 32864 27928
rect 32858 27888 32864 27900
rect 32916 27888 32922 27940
rect 29362 27860 29368 27872
rect 28460 27832 29368 27860
rect 29362 27820 29368 27832
rect 29420 27820 29426 27872
rect 29546 27820 29552 27872
rect 29604 27820 29610 27872
rect 30374 27820 30380 27872
rect 30432 27860 30438 27872
rect 30469 27863 30527 27869
rect 30469 27860 30481 27863
rect 30432 27832 30481 27860
rect 30432 27820 30438 27832
rect 30469 27829 30481 27832
rect 30515 27829 30527 27863
rect 30469 27823 30527 27829
rect 31294 27820 31300 27872
rect 31352 27860 31358 27872
rect 31846 27860 31852 27872
rect 31352 27832 31852 27860
rect 31352 27820 31358 27832
rect 31846 27820 31852 27832
rect 31904 27860 31910 27872
rect 32398 27860 32404 27872
rect 31904 27832 32404 27860
rect 31904 27820 31910 27832
rect 32398 27820 32404 27832
rect 32456 27820 32462 27872
rect 1104 27770 34868 27792
rect 1104 27718 5170 27770
rect 5222 27718 5234 27770
rect 5286 27718 5298 27770
rect 5350 27718 5362 27770
rect 5414 27718 5426 27770
rect 5478 27718 13611 27770
rect 13663 27718 13675 27770
rect 13727 27718 13739 27770
rect 13791 27718 13803 27770
rect 13855 27718 13867 27770
rect 13919 27718 22052 27770
rect 22104 27718 22116 27770
rect 22168 27718 22180 27770
rect 22232 27718 22244 27770
rect 22296 27718 22308 27770
rect 22360 27718 30493 27770
rect 30545 27718 30557 27770
rect 30609 27718 30621 27770
rect 30673 27718 30685 27770
rect 30737 27718 30749 27770
rect 30801 27718 34868 27770
rect 1104 27696 34868 27718
rect 17034 27616 17040 27668
rect 17092 27656 17098 27668
rect 22830 27656 22836 27668
rect 17092 27628 22836 27656
rect 17092 27616 17098 27628
rect 22830 27616 22836 27628
rect 22888 27616 22894 27668
rect 22922 27616 22928 27668
rect 22980 27656 22986 27668
rect 24765 27659 24823 27665
rect 24765 27656 24777 27659
rect 22980 27628 24777 27656
rect 22980 27616 22986 27628
rect 24765 27625 24777 27628
rect 24811 27656 24823 27659
rect 25866 27656 25872 27668
rect 24811 27628 25872 27656
rect 24811 27625 24823 27628
rect 24765 27619 24823 27625
rect 25866 27616 25872 27628
rect 25924 27656 25930 27668
rect 27522 27656 27528 27668
rect 25924 27628 27528 27656
rect 25924 27616 25930 27628
rect 27522 27616 27528 27628
rect 27580 27616 27586 27668
rect 30006 27656 30012 27668
rect 29656 27628 30012 27656
rect 16853 27591 16911 27597
rect 16853 27557 16865 27591
rect 16899 27588 16911 27591
rect 17586 27588 17592 27600
rect 16899 27560 17592 27588
rect 16899 27557 16911 27560
rect 16853 27551 16911 27557
rect 17586 27548 17592 27560
rect 17644 27548 17650 27600
rect 18506 27588 18512 27600
rect 17696 27560 18512 27588
rect 6457 27523 6515 27529
rect 6457 27489 6469 27523
rect 6503 27520 6515 27523
rect 7650 27520 7656 27532
rect 6503 27492 7656 27520
rect 6503 27489 6515 27492
rect 6457 27483 6515 27489
rect 7650 27480 7656 27492
rect 7708 27480 7714 27532
rect 7837 27523 7895 27529
rect 7837 27489 7849 27523
rect 7883 27489 7895 27523
rect 7837 27483 7895 27489
rect 6638 27384 6644 27396
rect 6599 27356 6644 27384
rect 6638 27344 6644 27356
rect 6696 27344 6702 27396
rect 3510 27276 3516 27328
rect 3568 27316 3574 27328
rect 7852 27316 7880 27483
rect 17034 27480 17040 27532
rect 17092 27520 17098 27532
rect 17696 27529 17724 27560
rect 18506 27548 18512 27560
rect 18564 27548 18570 27600
rect 22646 27548 22652 27600
rect 22704 27588 22710 27600
rect 23109 27591 23167 27597
rect 23109 27588 23121 27591
rect 22704 27560 23121 27588
rect 22704 27548 22710 27560
rect 23109 27557 23121 27560
rect 23155 27557 23167 27591
rect 23109 27551 23167 27557
rect 25498 27548 25504 27600
rect 25556 27588 25562 27600
rect 25961 27591 26019 27597
rect 25961 27588 25973 27591
rect 25556 27560 25973 27588
rect 25556 27548 25562 27560
rect 25961 27557 25973 27560
rect 26007 27557 26019 27591
rect 25961 27551 26019 27557
rect 26697 27591 26755 27597
rect 26697 27557 26709 27591
rect 26743 27557 26755 27591
rect 26697 27551 26755 27557
rect 27801 27591 27859 27597
rect 27801 27557 27813 27591
rect 27847 27588 27859 27591
rect 29454 27588 29460 27600
rect 27847 27560 29460 27588
rect 27847 27557 27859 27560
rect 27801 27551 27859 27557
rect 17681 27523 17739 27529
rect 17681 27520 17693 27523
rect 17092 27492 17693 27520
rect 17092 27480 17098 27492
rect 17681 27489 17693 27492
rect 17727 27489 17739 27523
rect 17681 27483 17739 27489
rect 17862 27480 17868 27532
rect 17920 27529 17926 27532
rect 17920 27523 17948 27529
rect 17936 27489 17948 27523
rect 19058 27520 19064 27532
rect 17920 27483 17948 27489
rect 18616 27492 19064 27520
rect 17920 27480 17926 27483
rect 18616 27464 18644 27492
rect 19058 27480 19064 27492
rect 19116 27480 19122 27532
rect 16022 27452 16028 27464
rect 15983 27424 16028 27452
rect 16022 27412 16028 27424
rect 16080 27412 16086 27464
rect 16485 27455 16543 27461
rect 16485 27421 16497 27455
rect 16531 27452 16543 27455
rect 17402 27452 17408 27464
rect 16531 27424 17408 27452
rect 16531 27421 16543 27424
rect 16485 27415 16543 27421
rect 17402 27412 17408 27424
rect 17460 27412 17466 27464
rect 17773 27455 17831 27461
rect 17773 27421 17785 27455
rect 17819 27452 17831 27455
rect 18322 27452 18328 27464
rect 17819 27424 18328 27452
rect 17819 27421 17831 27424
rect 17773 27415 17831 27421
rect 18322 27412 18328 27424
rect 18380 27412 18386 27464
rect 18598 27452 18604 27464
rect 18559 27424 18604 27452
rect 18598 27412 18604 27424
rect 18656 27412 18662 27464
rect 18693 27455 18751 27461
rect 18693 27421 18705 27455
rect 18739 27452 18751 27455
rect 19150 27452 19156 27464
rect 18739 27424 19156 27452
rect 18739 27421 18751 27424
rect 18693 27415 18751 27421
rect 19150 27412 19156 27424
rect 19208 27412 19214 27464
rect 19426 27452 19432 27464
rect 19339 27424 19432 27452
rect 19426 27412 19432 27424
rect 19484 27452 19490 27464
rect 21269 27455 21327 27461
rect 21269 27452 21281 27455
rect 19484 27424 21281 27452
rect 19484 27412 19490 27424
rect 21269 27421 21281 27424
rect 21315 27452 21327 27455
rect 22462 27452 22468 27464
rect 21315 27424 22468 27452
rect 21315 27421 21327 27424
rect 21269 27415 21327 27421
rect 22462 27412 22468 27424
rect 22520 27412 22526 27464
rect 16868 27356 17816 27384
rect 3568 27288 7880 27316
rect 15841 27319 15899 27325
rect 3568 27276 3574 27288
rect 15841 27285 15853 27319
rect 15887 27316 15899 27319
rect 16868 27316 16896 27356
rect 15887 27288 16896 27316
rect 16945 27319 17003 27325
rect 15887 27285 15899 27288
rect 15841 27279 15899 27285
rect 16945 27285 16957 27319
rect 16991 27316 17003 27319
rect 17402 27316 17408 27328
rect 16991 27288 17408 27316
rect 16991 27285 17003 27288
rect 16945 27279 17003 27285
rect 17402 27276 17408 27288
rect 17460 27276 17466 27328
rect 17788 27316 17816 27356
rect 17972 27356 19472 27384
rect 17972 27316 18000 27356
rect 17788 27288 18000 27316
rect 18049 27319 18107 27325
rect 18049 27285 18061 27319
rect 18095 27316 18107 27319
rect 18230 27316 18236 27328
rect 18095 27288 18236 27316
rect 18095 27285 18107 27288
rect 18049 27279 18107 27285
rect 18230 27276 18236 27288
rect 18288 27276 18294 27328
rect 18877 27319 18935 27325
rect 18877 27285 18889 27319
rect 18923 27316 18935 27319
rect 19334 27316 19340 27328
rect 18923 27288 19340 27316
rect 18923 27285 18935 27288
rect 18877 27279 18935 27285
rect 19334 27276 19340 27288
rect 19392 27276 19398 27328
rect 19444 27316 19472 27356
rect 19518 27344 19524 27396
rect 19576 27384 19582 27396
rect 19674 27387 19732 27393
rect 19674 27384 19686 27387
rect 19576 27356 19686 27384
rect 19576 27344 19582 27356
rect 19674 27353 19686 27356
rect 19720 27353 19732 27387
rect 19674 27347 19732 27353
rect 21536 27387 21594 27393
rect 21536 27353 21548 27387
rect 21582 27384 21594 27387
rect 21910 27384 21916 27396
rect 21582 27356 21916 27384
rect 21582 27353 21594 27356
rect 21536 27347 21594 27353
rect 21910 27344 21916 27356
rect 21968 27344 21974 27396
rect 22664 27384 22692 27548
rect 23842 27520 23848 27532
rect 22066 27356 22692 27384
rect 23032 27492 23848 27520
rect 20438 27316 20444 27328
rect 19444 27288 20444 27316
rect 20438 27276 20444 27288
rect 20496 27276 20502 27328
rect 20809 27319 20867 27325
rect 20809 27285 20821 27319
rect 20855 27316 20867 27319
rect 22066 27316 22094 27356
rect 20855 27288 22094 27316
rect 22649 27319 22707 27325
rect 20855 27285 20867 27288
rect 20809 27279 20867 27285
rect 22649 27285 22661 27319
rect 22695 27316 22707 27319
rect 22830 27316 22836 27328
rect 22695 27288 22836 27316
rect 22695 27285 22707 27288
rect 22649 27279 22707 27285
rect 22830 27276 22836 27288
rect 22888 27276 22894 27328
rect 23032 27316 23060 27492
rect 23842 27480 23848 27492
rect 23900 27520 23906 27532
rect 24118 27520 24124 27532
rect 23900 27492 24124 27520
rect 23900 27480 23906 27492
rect 24118 27480 24124 27492
rect 24176 27480 24182 27532
rect 26050 27480 26056 27532
rect 26108 27520 26114 27532
rect 26712 27520 26740 27551
rect 29454 27548 29460 27560
rect 29512 27588 29518 27600
rect 29656 27588 29684 27628
rect 30006 27616 30012 27628
rect 30064 27616 30070 27668
rect 34238 27616 34244 27668
rect 34296 27656 34302 27668
rect 34333 27659 34391 27665
rect 34333 27656 34345 27659
rect 34296 27628 34345 27656
rect 34296 27616 34302 27628
rect 34333 27625 34345 27628
rect 34379 27625 34391 27659
rect 34333 27619 34391 27625
rect 29512 27560 29684 27588
rect 29512 27548 29518 27560
rect 29730 27548 29736 27600
rect 29788 27588 29794 27600
rect 29788 27560 32996 27588
rect 29788 27548 29794 27560
rect 26108 27492 26740 27520
rect 26108 27480 26114 27492
rect 29086 27480 29092 27532
rect 29144 27520 29150 27532
rect 29914 27520 29920 27532
rect 29144 27492 29500 27520
rect 29875 27492 29920 27520
rect 29144 27480 29150 27492
rect 23290 27412 23296 27464
rect 23348 27452 23354 27464
rect 23477 27455 23535 27461
rect 23477 27452 23489 27455
rect 23348 27424 23489 27452
rect 23348 27412 23354 27424
rect 23477 27421 23489 27424
rect 23523 27421 23535 27455
rect 24670 27452 24676 27464
rect 24631 27424 24676 27452
rect 23477 27415 23535 27421
rect 24670 27412 24676 27424
rect 24728 27412 24734 27464
rect 24762 27412 24768 27464
rect 24820 27452 24826 27464
rect 25317 27455 25375 27461
rect 25317 27452 25329 27455
rect 24820 27424 25329 27452
rect 24820 27412 24826 27424
rect 25317 27421 25329 27424
rect 25363 27452 25375 27455
rect 26421 27455 26479 27461
rect 26421 27452 26433 27455
rect 25363 27424 26433 27452
rect 25363 27421 25375 27424
rect 25317 27415 25375 27421
rect 26421 27421 26433 27424
rect 26467 27452 26479 27455
rect 27154 27452 27160 27464
rect 26467 27424 27160 27452
rect 26467 27421 26479 27424
rect 26421 27415 26479 27421
rect 27154 27412 27160 27424
rect 27212 27412 27218 27464
rect 27982 27452 27988 27464
rect 27943 27424 27988 27452
rect 27982 27412 27988 27424
rect 28040 27412 28046 27464
rect 28258 27452 28264 27464
rect 28219 27424 28264 27452
rect 28258 27412 28264 27424
rect 28316 27412 28322 27464
rect 28902 27452 28908 27464
rect 28863 27424 28908 27452
rect 28902 27412 28908 27424
rect 28960 27412 28966 27464
rect 29178 27452 29184 27464
rect 29139 27424 29184 27452
rect 29178 27412 29184 27424
rect 29236 27412 29242 27464
rect 29472 27452 29500 27492
rect 29914 27480 29920 27492
rect 29972 27480 29978 27532
rect 30190 27520 30196 27532
rect 30151 27492 30196 27520
rect 30190 27480 30196 27492
rect 30248 27480 30254 27532
rect 30282 27480 30288 27532
rect 30340 27520 30346 27532
rect 31294 27520 31300 27532
rect 30340 27492 31300 27520
rect 30340 27480 30346 27492
rect 31294 27480 31300 27492
rect 31352 27480 31358 27532
rect 31662 27480 31668 27532
rect 31720 27520 31726 27532
rect 31757 27523 31815 27529
rect 31757 27520 31769 27523
rect 31720 27492 31769 27520
rect 31720 27480 31726 27492
rect 31757 27489 31769 27492
rect 31803 27489 31815 27523
rect 31757 27483 31815 27489
rect 32214 27480 32220 27532
rect 32272 27520 32278 27532
rect 32968 27529 32996 27560
rect 32309 27523 32367 27529
rect 32309 27520 32321 27523
rect 32272 27492 32321 27520
rect 32272 27480 32278 27492
rect 32309 27489 32321 27492
rect 32355 27489 32367 27523
rect 32309 27483 32367 27489
rect 32953 27523 33011 27529
rect 32953 27489 32965 27523
rect 32999 27489 33011 27523
rect 32953 27483 33011 27489
rect 29822 27452 29828 27464
rect 29472 27424 29828 27452
rect 29822 27412 29828 27424
rect 29880 27452 29886 27464
rect 30009 27455 30067 27461
rect 30009 27452 30021 27455
rect 29880 27424 30021 27452
rect 29880 27412 29886 27424
rect 30009 27421 30021 27424
rect 30055 27421 30067 27455
rect 30009 27415 30067 27421
rect 30098 27412 30104 27464
rect 30156 27452 30162 27464
rect 30156 27424 30201 27452
rect 30156 27412 30162 27424
rect 31110 27412 31116 27464
rect 31168 27452 31174 27464
rect 31389 27455 31447 27461
rect 31389 27452 31401 27455
rect 31168 27424 31401 27452
rect 31168 27412 31174 27424
rect 31389 27421 31401 27424
rect 31435 27452 31447 27455
rect 31478 27452 31484 27464
rect 31435 27424 31484 27452
rect 31435 27421 31447 27424
rect 31389 27415 31447 27421
rect 31478 27412 31484 27424
rect 31536 27412 31542 27464
rect 32030 27452 32036 27464
rect 31991 27424 32036 27452
rect 32030 27412 32036 27424
rect 32088 27412 32094 27464
rect 32125 27455 32183 27461
rect 32125 27421 32137 27455
rect 32171 27452 32183 27455
rect 32490 27452 32496 27464
rect 32171 27424 32496 27452
rect 32171 27421 32183 27424
rect 32125 27415 32183 27421
rect 23198 27344 23204 27396
rect 23256 27384 23262 27396
rect 23661 27387 23719 27393
rect 23661 27384 23673 27387
rect 23256 27356 23673 27384
rect 23256 27344 23262 27356
rect 23661 27353 23673 27356
rect 23707 27353 23719 27387
rect 23661 27347 23719 27353
rect 24854 27344 24860 27396
rect 24912 27384 24918 27396
rect 25802 27387 25860 27393
rect 25802 27384 25814 27387
rect 24912 27356 25814 27384
rect 24912 27344 24918 27356
rect 25802 27353 25814 27356
rect 25848 27384 25860 27387
rect 25958 27384 25964 27396
rect 25848 27356 25964 27384
rect 25848 27353 25860 27356
rect 25802 27347 25860 27353
rect 25958 27344 25964 27356
rect 26016 27344 26022 27396
rect 27062 27384 27068 27396
rect 26068 27356 27068 27384
rect 23293 27319 23351 27325
rect 23293 27316 23305 27319
rect 23032 27288 23305 27316
rect 23293 27285 23305 27288
rect 23339 27285 23351 27319
rect 23293 27279 23351 27285
rect 23385 27319 23443 27325
rect 23385 27285 23397 27319
rect 23431 27316 23443 27319
rect 23750 27316 23756 27328
rect 23431 27288 23756 27316
rect 23431 27285 23443 27288
rect 23385 27279 23443 27285
rect 23750 27276 23756 27288
rect 23808 27276 23814 27328
rect 25590 27316 25596 27328
rect 25551 27288 25596 27316
rect 25590 27276 25596 27288
rect 25648 27276 25654 27328
rect 25685 27319 25743 27325
rect 25685 27285 25697 27319
rect 25731 27316 25743 27319
rect 26068 27316 26096 27356
rect 27062 27344 27068 27356
rect 27120 27344 27126 27396
rect 28074 27344 28080 27396
rect 28132 27384 28138 27396
rect 28920 27384 28948 27412
rect 31570 27384 31576 27396
rect 28132 27356 28948 27384
rect 29748 27356 31576 27384
rect 28132 27344 28138 27356
rect 25731 27288 26096 27316
rect 25731 27285 25743 27288
rect 25685 27279 25743 27285
rect 26142 27276 26148 27328
rect 26200 27316 26206 27328
rect 26881 27319 26939 27325
rect 26881 27316 26893 27319
rect 26200 27288 26893 27316
rect 26200 27276 26206 27288
rect 26881 27285 26893 27288
rect 26927 27285 26939 27319
rect 26881 27279 26939 27285
rect 27614 27276 27620 27328
rect 27672 27316 27678 27328
rect 28169 27319 28227 27325
rect 28169 27316 28181 27319
rect 27672 27288 28181 27316
rect 27672 27276 27678 27288
rect 28169 27285 28181 27288
rect 28215 27285 28227 27319
rect 28718 27316 28724 27328
rect 28679 27288 28724 27316
rect 28169 27279 28227 27285
rect 28718 27276 28724 27288
rect 28776 27276 28782 27328
rect 29089 27319 29147 27325
rect 29089 27285 29101 27319
rect 29135 27316 29147 27319
rect 29454 27316 29460 27328
rect 29135 27288 29460 27316
rect 29135 27285 29147 27288
rect 29089 27279 29147 27285
rect 29454 27276 29460 27288
rect 29512 27276 29518 27328
rect 29748 27325 29776 27356
rect 31570 27344 31576 27356
rect 31628 27344 31634 27396
rect 31662 27344 31668 27396
rect 31720 27384 31726 27396
rect 32140 27384 32168 27415
rect 32490 27412 32496 27424
rect 32548 27412 32554 27464
rect 33198 27387 33256 27393
rect 33198 27384 33210 27387
rect 31720 27356 32168 27384
rect 32600 27356 33210 27384
rect 31720 27344 31726 27356
rect 32600 27328 32628 27356
rect 33198 27353 33210 27356
rect 33244 27353 33256 27387
rect 33198 27347 33256 27353
rect 29733 27319 29791 27325
rect 29733 27285 29745 27319
rect 29779 27285 29791 27319
rect 29733 27279 29791 27285
rect 30098 27276 30104 27328
rect 30156 27316 30162 27328
rect 32309 27319 32367 27325
rect 32309 27316 32321 27319
rect 30156 27288 32321 27316
rect 30156 27276 30162 27288
rect 32309 27285 32321 27288
rect 32355 27285 32367 27319
rect 32582 27316 32588 27328
rect 32543 27288 32588 27316
rect 32309 27279 32367 27285
rect 32582 27276 32588 27288
rect 32640 27276 32646 27328
rect 1104 27226 35027 27248
rect 1104 27174 9390 27226
rect 9442 27174 9454 27226
rect 9506 27174 9518 27226
rect 9570 27174 9582 27226
rect 9634 27174 9646 27226
rect 9698 27174 17831 27226
rect 17883 27174 17895 27226
rect 17947 27174 17959 27226
rect 18011 27174 18023 27226
rect 18075 27174 18087 27226
rect 18139 27174 26272 27226
rect 26324 27174 26336 27226
rect 26388 27174 26400 27226
rect 26452 27174 26464 27226
rect 26516 27174 26528 27226
rect 26580 27174 34713 27226
rect 34765 27174 34777 27226
rect 34829 27174 34841 27226
rect 34893 27174 34905 27226
rect 34957 27174 34969 27226
rect 35021 27174 35027 27226
rect 1104 27152 35027 27174
rect 6638 27112 6644 27124
rect 6599 27084 6644 27112
rect 6638 27072 6644 27084
rect 6696 27072 6702 27124
rect 7650 27072 7656 27124
rect 7708 27112 7714 27124
rect 8757 27115 8815 27121
rect 8757 27112 8769 27115
rect 7708 27084 8769 27112
rect 7708 27072 7714 27084
rect 8757 27081 8769 27084
rect 8803 27081 8815 27115
rect 18322 27112 18328 27124
rect 8757 27075 8815 27081
rect 16684 27084 18328 27112
rect 2130 26936 2136 26988
rect 2188 26976 2194 26988
rect 6546 26976 6552 26988
rect 2188 26948 6552 26976
rect 2188 26936 2194 26948
rect 6546 26936 6552 26948
rect 6604 26936 6610 26988
rect 8938 26976 8944 26988
rect 8899 26948 8944 26976
rect 8938 26936 8944 26948
rect 8996 26936 9002 26988
rect 16117 26979 16175 26985
rect 16117 26945 16129 26979
rect 16163 26945 16175 26979
rect 16298 26976 16304 26988
rect 16259 26948 16304 26976
rect 16117 26939 16175 26945
rect 16132 26908 16160 26939
rect 16298 26936 16304 26948
rect 16356 26936 16362 26988
rect 16684 26976 16712 27084
rect 18322 27072 18328 27084
rect 18380 27112 18386 27124
rect 20809 27115 20867 27121
rect 20809 27112 20821 27115
rect 18380 27084 20821 27112
rect 18380 27072 18386 27084
rect 16758 27004 16764 27056
rect 16816 27044 16822 27056
rect 18230 27044 18236 27056
rect 16816 27016 18236 27044
rect 16816 27004 16822 27016
rect 16853 26979 16911 26985
rect 16853 26976 16865 26979
rect 16684 26948 16865 26976
rect 16853 26945 16865 26948
rect 16899 26945 16911 26979
rect 17034 26976 17040 26988
rect 16995 26948 17040 26976
rect 16853 26939 16911 26945
rect 17034 26936 17040 26948
rect 17092 26936 17098 26988
rect 17972 26985 18000 27016
rect 18230 27004 18236 27016
rect 18288 27004 18294 27056
rect 17681 26979 17739 26985
rect 17681 26945 17693 26979
rect 17727 26945 17739 26979
rect 17681 26939 17739 26945
rect 17773 26979 17831 26985
rect 17773 26945 17785 26979
rect 17819 26945 17831 26979
rect 17773 26939 17831 26945
rect 17957 26979 18015 26985
rect 17957 26945 17969 26979
rect 18003 26945 18015 26979
rect 17957 26939 18015 26945
rect 16942 26908 16948 26920
rect 16132 26880 16948 26908
rect 16942 26868 16948 26880
rect 17000 26868 17006 26920
rect 17696 26908 17724 26939
rect 17052 26880 17724 26908
rect 17788 26908 17816 26939
rect 18046 26936 18052 26988
rect 18104 26976 18110 26988
rect 18506 26976 18512 26988
rect 18104 26948 18149 26976
rect 18467 26948 18512 26976
rect 18104 26936 18110 26948
rect 18506 26936 18512 26948
rect 18564 26936 18570 26988
rect 18708 26985 18736 27084
rect 20809 27081 20821 27084
rect 20855 27081 20867 27115
rect 20809 27075 20867 27081
rect 20916 27084 26924 27112
rect 18782 27004 18788 27056
rect 18840 27044 18846 27056
rect 19702 27053 19708 27056
rect 19696 27044 19708 27053
rect 18840 27016 19564 27044
rect 19663 27016 19708 27044
rect 18840 27004 18846 27016
rect 18693 26979 18751 26985
rect 18693 26945 18705 26979
rect 18739 26945 18751 26979
rect 19426 26976 19432 26988
rect 19387 26948 19432 26976
rect 18693 26939 18751 26945
rect 19426 26936 19432 26948
rect 19484 26936 19490 26988
rect 19536 26976 19564 27016
rect 19696 27007 19708 27016
rect 19702 27004 19708 27007
rect 19760 27004 19766 27056
rect 20916 26976 20944 27084
rect 22462 27044 22468 27056
rect 22020 27016 22468 27044
rect 21450 26976 21456 26988
rect 19536 26948 20944 26976
rect 21411 26948 21456 26976
rect 21450 26936 21456 26948
rect 21508 26936 21514 26988
rect 22020 26985 22048 27016
rect 22462 27004 22468 27016
rect 22520 27004 22526 27056
rect 22646 27004 22652 27056
rect 22704 27044 22710 27056
rect 23014 27044 23020 27056
rect 22704 27016 23020 27044
rect 22704 27004 22710 27016
rect 23014 27004 23020 27016
rect 23072 27004 23078 27056
rect 23290 27004 23296 27056
rect 23348 27044 23354 27056
rect 23937 27047 23995 27053
rect 23937 27044 23949 27047
rect 23348 27016 23949 27044
rect 23348 27004 23354 27016
rect 23937 27013 23949 27016
rect 23983 27013 23995 27047
rect 26896 27044 26924 27084
rect 28166 27072 28172 27124
rect 28224 27112 28230 27124
rect 28445 27115 28503 27121
rect 28445 27112 28457 27115
rect 28224 27084 28457 27112
rect 28224 27072 28230 27084
rect 28445 27081 28457 27084
rect 28491 27112 28503 27115
rect 28534 27112 28540 27124
rect 28491 27084 28540 27112
rect 28491 27081 28503 27084
rect 28445 27075 28503 27081
rect 28534 27072 28540 27084
rect 28592 27072 28598 27124
rect 32582 27112 32588 27124
rect 28644 27084 32588 27112
rect 28644 27044 28672 27084
rect 32582 27072 32588 27084
rect 32640 27072 32646 27124
rect 26896 27016 28672 27044
rect 23937 27007 23995 27013
rect 28718 27004 28724 27056
rect 28776 27044 28782 27056
rect 32950 27044 32956 27056
rect 28776 27016 29868 27044
rect 28776 27004 28782 27016
rect 22005 26979 22063 26985
rect 22005 26945 22017 26979
rect 22051 26945 22063 26979
rect 22005 26939 22063 26945
rect 22272 26979 22330 26985
rect 22272 26945 22284 26979
rect 22318 26976 22330 26979
rect 23566 26976 23572 26988
rect 22318 26948 23572 26976
rect 22318 26945 22330 26948
rect 22272 26939 22330 26945
rect 23566 26936 23572 26948
rect 23624 26936 23630 26988
rect 24213 26979 24271 26985
rect 24213 26976 24225 26979
rect 23676 26948 24225 26976
rect 18138 26908 18144 26920
rect 17788 26880 18144 26908
rect 17052 26784 17080 26880
rect 18138 26868 18144 26880
rect 18196 26908 18202 26920
rect 18414 26908 18420 26920
rect 18196 26880 18420 26908
rect 18196 26868 18202 26880
rect 18414 26868 18420 26880
rect 18472 26868 18478 26920
rect 23014 26868 23020 26920
rect 23072 26908 23078 26920
rect 23676 26908 23704 26948
rect 24213 26945 24225 26948
rect 24259 26945 24271 26979
rect 24213 26939 24271 26945
rect 24578 26936 24584 26988
rect 24636 26976 24642 26988
rect 25225 26979 25283 26985
rect 25225 26976 25237 26979
rect 24636 26948 25237 26976
rect 24636 26936 24642 26948
rect 25225 26945 25237 26948
rect 25271 26945 25283 26979
rect 25481 26979 25539 26985
rect 25481 26976 25493 26979
rect 25225 26939 25283 26945
rect 25332 26948 25493 26976
rect 23072 26880 23704 26908
rect 23072 26868 23078 26880
rect 23750 26868 23756 26920
rect 23808 26908 23814 26920
rect 24029 26911 24087 26917
rect 24029 26908 24041 26911
rect 23808 26880 24041 26908
rect 23808 26868 23814 26880
rect 24029 26877 24041 26880
rect 24075 26877 24087 26911
rect 25332 26908 25360 26948
rect 25481 26945 25493 26948
rect 25527 26945 25539 26979
rect 27154 26976 27160 26988
rect 27115 26948 27160 26976
rect 25481 26939 25539 26945
rect 27154 26936 27160 26948
rect 27212 26936 27218 26988
rect 29362 26936 29368 26988
rect 29420 26976 29426 26988
rect 29638 26976 29644 26988
rect 29420 26948 29644 26976
rect 29420 26936 29426 26948
rect 29638 26936 29644 26948
rect 29696 26936 29702 26988
rect 29840 26985 29868 27016
rect 29932 27016 30696 27044
rect 29733 26979 29791 26985
rect 29733 26945 29745 26979
rect 29779 26945 29791 26979
rect 29733 26939 29791 26945
rect 29825 26979 29883 26985
rect 29825 26945 29837 26979
rect 29871 26945 29883 26979
rect 29825 26939 29883 26945
rect 29178 26908 29184 26920
rect 24029 26871 24087 26877
rect 24136 26880 25360 26908
rect 26252 26880 29184 26908
rect 17497 26843 17555 26849
rect 17497 26809 17509 26843
rect 17543 26840 17555 26843
rect 18230 26840 18236 26852
rect 17543 26812 18236 26840
rect 17543 26809 17555 26812
rect 17497 26803 17555 26809
rect 18230 26800 18236 26812
rect 18288 26800 18294 26852
rect 20438 26800 20444 26852
rect 20496 26840 20502 26852
rect 24136 26840 24164 26880
rect 24394 26840 24400 26852
rect 20496 26812 21404 26840
rect 20496 26800 20502 26812
rect 16114 26772 16120 26784
rect 16075 26744 16120 26772
rect 16114 26732 16120 26744
rect 16172 26732 16178 26784
rect 16853 26775 16911 26781
rect 16853 26741 16865 26775
rect 16899 26772 16911 26775
rect 17034 26772 17040 26784
rect 16899 26744 17040 26772
rect 16899 26741 16911 26744
rect 16853 26735 16911 26741
rect 17034 26732 17040 26744
rect 17092 26732 17098 26784
rect 17862 26732 17868 26784
rect 17920 26772 17926 26784
rect 18877 26775 18935 26781
rect 18877 26772 18889 26775
rect 17920 26744 18889 26772
rect 17920 26732 17926 26744
rect 18877 26741 18889 26744
rect 18923 26741 18935 26775
rect 21266 26772 21272 26784
rect 21227 26744 21272 26772
rect 18877 26735 18935 26741
rect 21266 26732 21272 26744
rect 21324 26732 21330 26784
rect 21376 26772 21404 26812
rect 23308 26812 24164 26840
rect 24355 26812 24400 26840
rect 23308 26772 23336 26812
rect 24394 26800 24400 26812
rect 24452 26800 24458 26852
rect 21376 26744 23336 26772
rect 23382 26732 23388 26784
rect 23440 26772 23446 26784
rect 24118 26772 24124 26784
rect 23440 26744 23485 26772
rect 24079 26744 24124 26772
rect 23440 26732 23446 26744
rect 24118 26732 24124 26744
rect 24176 26732 24182 26784
rect 24578 26732 24584 26784
rect 24636 26772 24642 26784
rect 26252 26772 26280 26880
rect 29178 26868 29184 26880
rect 29236 26868 29242 26920
rect 29546 26868 29552 26920
rect 29604 26908 29610 26920
rect 29748 26908 29776 26939
rect 29932 26908 29960 27016
rect 30009 26979 30067 26985
rect 30009 26945 30021 26979
rect 30055 26945 30067 26979
rect 30009 26939 30067 26945
rect 29604 26880 29960 26908
rect 29604 26868 29610 26880
rect 26326 26800 26332 26852
rect 26384 26840 26390 26852
rect 27982 26840 27988 26852
rect 26384 26812 27988 26840
rect 26384 26800 26390 26812
rect 27982 26800 27988 26812
rect 28040 26800 28046 26852
rect 28166 26800 28172 26852
rect 28224 26840 28230 26852
rect 30024 26840 30052 26939
rect 30668 26908 30696 27016
rect 31588 27016 32956 27044
rect 31110 26936 31116 26988
rect 31168 26976 31174 26988
rect 31389 26979 31447 26985
rect 31389 26976 31401 26979
rect 31168 26948 31401 26976
rect 31168 26936 31174 26948
rect 31389 26945 31401 26948
rect 31435 26945 31447 26979
rect 31389 26939 31447 26945
rect 31478 26982 31536 26988
rect 31588 26985 31616 27016
rect 32950 27004 32956 27016
rect 33008 27004 33014 27056
rect 33594 27044 33600 27056
rect 33244 27016 33600 27044
rect 31478 26948 31490 26982
rect 31524 26948 31536 26982
rect 31478 26942 31536 26948
rect 31573 26979 31631 26985
rect 31573 26945 31585 26979
rect 31619 26945 31631 26979
rect 31754 26976 31760 26988
rect 31715 26948 31760 26976
rect 31493 26908 31521 26942
rect 31573 26939 31631 26945
rect 31754 26936 31760 26948
rect 31812 26936 31818 26988
rect 32493 26979 32551 26985
rect 32493 26945 32505 26979
rect 32539 26976 32551 26979
rect 33244 26976 33272 27016
rect 33594 27004 33600 27016
rect 33652 27044 33658 27056
rect 34238 27044 34244 27056
rect 33652 27016 34244 27044
rect 33652 27004 33658 27016
rect 34238 27004 34244 27016
rect 34296 27004 34302 27056
rect 33502 26976 33508 26988
rect 32539 26948 33272 26976
rect 33463 26948 33508 26976
rect 32539 26945 32551 26948
rect 32493 26939 32551 26945
rect 33502 26936 33508 26948
rect 33560 26936 33566 26988
rect 33686 26976 33692 26988
rect 33647 26948 33692 26976
rect 33686 26936 33692 26948
rect 33744 26936 33750 26988
rect 33781 26979 33839 26985
rect 33781 26945 33793 26979
rect 33827 26945 33839 26979
rect 33781 26939 33839 26945
rect 32122 26908 32128 26920
rect 30668 26880 32128 26908
rect 32122 26868 32128 26880
rect 32180 26868 32186 26920
rect 32398 26908 32404 26920
rect 32359 26880 32404 26908
rect 32398 26868 32404 26880
rect 32456 26868 32462 26920
rect 32858 26908 32864 26920
rect 32819 26880 32864 26908
rect 32858 26868 32864 26880
rect 32916 26868 32922 26920
rect 33042 26868 33048 26920
rect 33100 26908 33106 26920
rect 33796 26908 33824 26939
rect 33100 26880 33824 26908
rect 33100 26868 33106 26880
rect 28224 26812 30052 26840
rect 28224 26800 28230 26812
rect 30926 26800 30932 26852
rect 30984 26840 30990 26852
rect 34238 26840 34244 26852
rect 30984 26812 34244 26840
rect 30984 26800 30990 26812
rect 34238 26800 34244 26812
rect 34296 26800 34302 26852
rect 24636 26744 26280 26772
rect 26605 26775 26663 26781
rect 24636 26732 24642 26744
rect 26605 26741 26617 26775
rect 26651 26772 26663 26775
rect 27062 26772 27068 26784
rect 26651 26744 27068 26772
rect 26651 26741 26663 26744
rect 26605 26735 26663 26741
rect 27062 26732 27068 26744
rect 27120 26732 27126 26784
rect 29362 26772 29368 26784
rect 29323 26744 29368 26772
rect 29362 26732 29368 26744
rect 29420 26732 29426 26784
rect 29638 26732 29644 26784
rect 29696 26772 29702 26784
rect 29914 26772 29920 26784
rect 29696 26744 29920 26772
rect 29696 26732 29702 26744
rect 29914 26732 29920 26744
rect 29972 26732 29978 26784
rect 31113 26775 31171 26781
rect 31113 26741 31125 26775
rect 31159 26772 31171 26775
rect 32398 26772 32404 26784
rect 31159 26744 32404 26772
rect 31159 26741 31171 26744
rect 31113 26735 31171 26741
rect 32398 26732 32404 26744
rect 32456 26732 32462 26784
rect 33318 26772 33324 26784
rect 33279 26744 33324 26772
rect 33318 26732 33324 26744
rect 33376 26732 33382 26784
rect 1104 26682 34868 26704
rect 1104 26630 5170 26682
rect 5222 26630 5234 26682
rect 5286 26630 5298 26682
rect 5350 26630 5362 26682
rect 5414 26630 5426 26682
rect 5478 26630 13611 26682
rect 13663 26630 13675 26682
rect 13727 26630 13739 26682
rect 13791 26630 13803 26682
rect 13855 26630 13867 26682
rect 13919 26630 22052 26682
rect 22104 26630 22116 26682
rect 22168 26630 22180 26682
rect 22232 26630 22244 26682
rect 22296 26630 22308 26682
rect 22360 26630 30493 26682
rect 30545 26630 30557 26682
rect 30609 26630 30621 26682
rect 30673 26630 30685 26682
rect 30737 26630 30749 26682
rect 30801 26630 34868 26682
rect 1104 26608 34868 26630
rect 16942 26528 16948 26580
rect 17000 26568 17006 26580
rect 19058 26568 19064 26580
rect 17000 26540 19064 26568
rect 17000 26528 17006 26540
rect 19058 26528 19064 26540
rect 19116 26528 19122 26580
rect 26142 26568 26148 26580
rect 26103 26540 26148 26568
rect 26142 26528 26148 26540
rect 26200 26528 26206 26580
rect 28997 26571 29055 26577
rect 28997 26568 29009 26571
rect 26252 26540 29009 26568
rect 16114 26460 16120 26512
rect 16172 26500 16178 26512
rect 18966 26500 18972 26512
rect 16172 26472 18972 26500
rect 16172 26460 16178 26472
rect 18966 26460 18972 26472
rect 19024 26460 19030 26512
rect 19426 26460 19432 26512
rect 19484 26500 19490 26512
rect 19484 26472 19529 26500
rect 19484 26460 19490 26472
rect 24394 26460 24400 26512
rect 24452 26500 24458 26512
rect 24762 26500 24768 26512
rect 24452 26472 24768 26500
rect 24452 26460 24458 26472
rect 24762 26460 24768 26472
rect 24820 26500 24826 26512
rect 24949 26503 25007 26509
rect 24949 26500 24961 26503
rect 24820 26472 24961 26500
rect 24820 26460 24826 26472
rect 24949 26469 24961 26472
rect 24995 26469 25007 26503
rect 24949 26463 25007 26469
rect 25038 26460 25044 26512
rect 25096 26500 25102 26512
rect 26252 26500 26280 26540
rect 28997 26537 29009 26540
rect 29043 26537 29055 26571
rect 28997 26531 29055 26537
rect 29178 26528 29184 26580
rect 29236 26568 29242 26580
rect 30101 26571 30159 26577
rect 29236 26540 29868 26568
rect 29236 26528 29242 26540
rect 25096 26472 26280 26500
rect 25096 26460 25102 26472
rect 28258 26460 28264 26512
rect 28316 26500 28322 26512
rect 28442 26500 28448 26512
rect 28316 26472 28448 26500
rect 28316 26460 28322 26472
rect 28442 26460 28448 26472
rect 28500 26500 28506 26512
rect 28537 26503 28595 26509
rect 28537 26500 28549 26503
rect 28500 26472 28549 26500
rect 28500 26460 28506 26472
rect 28537 26469 28549 26472
rect 28583 26500 28595 26503
rect 29638 26500 29644 26512
rect 28583 26472 29644 26500
rect 28583 26469 28595 26472
rect 28537 26463 28595 26469
rect 29638 26460 29644 26472
rect 29696 26460 29702 26512
rect 17862 26432 17868 26444
rect 17052 26404 17724 26432
rect 17823 26404 17868 26432
rect 17052 26376 17080 26404
rect 17696 26376 17724 26404
rect 17862 26392 17868 26404
rect 17920 26392 17926 26444
rect 18782 26392 18788 26444
rect 18840 26432 18846 26444
rect 22462 26432 22468 26444
rect 18840 26404 20208 26432
rect 22423 26404 22468 26432
rect 18840 26392 18846 26404
rect 16758 26364 16764 26376
rect 16719 26336 16764 26364
rect 16758 26324 16764 26336
rect 16816 26324 16822 26376
rect 17034 26364 17040 26376
rect 16995 26336 17040 26364
rect 17034 26324 17040 26336
rect 17092 26324 17098 26376
rect 17310 26324 17316 26376
rect 17368 26364 17374 26376
rect 17494 26364 17500 26376
rect 17368 26336 17500 26364
rect 17368 26324 17374 26336
rect 17494 26324 17500 26336
rect 17552 26324 17558 26376
rect 17678 26364 17684 26376
rect 17591 26336 17684 26364
rect 17678 26324 17684 26336
rect 17736 26324 17742 26376
rect 17773 26367 17831 26373
rect 17773 26333 17785 26367
rect 17819 26333 17831 26367
rect 17773 26327 17831 26333
rect 18049 26367 18107 26373
rect 18049 26333 18061 26367
rect 18095 26364 18107 26367
rect 18138 26364 18144 26376
rect 18095 26336 18144 26364
rect 18095 26333 18107 26336
rect 18049 26327 18107 26333
rect 16022 26256 16028 26308
rect 16080 26296 16086 26308
rect 16577 26299 16635 26305
rect 16577 26296 16589 26299
rect 16080 26268 16589 26296
rect 16080 26256 16086 26268
rect 16577 26265 16589 26268
rect 16623 26265 16635 26299
rect 16577 26259 16635 26265
rect 16945 26299 17003 26305
rect 16945 26265 16957 26299
rect 16991 26296 17003 26299
rect 16991 26268 17356 26296
rect 16991 26265 17003 26268
rect 16945 26259 17003 26265
rect 17328 26228 17356 26268
rect 17402 26256 17408 26308
rect 17460 26296 17466 26308
rect 17788 26296 17816 26327
rect 18138 26324 18144 26336
rect 18196 26324 18202 26376
rect 18233 26367 18291 26373
rect 18233 26333 18245 26367
rect 18279 26364 18291 26367
rect 18598 26364 18604 26376
rect 18279 26336 18604 26364
rect 18279 26333 18291 26336
rect 18233 26327 18291 26333
rect 18598 26324 18604 26336
rect 18656 26364 18662 26376
rect 18693 26367 18751 26373
rect 18693 26364 18705 26367
rect 18656 26336 18705 26364
rect 18656 26324 18662 26336
rect 18693 26333 18705 26336
rect 18739 26333 18751 26367
rect 18874 26364 18880 26376
rect 18835 26336 18880 26364
rect 18693 26327 18751 26333
rect 18874 26324 18880 26336
rect 18932 26324 18938 26376
rect 19334 26324 19340 26376
rect 19392 26364 19398 26376
rect 20180 26373 20208 26404
rect 22462 26392 22468 26404
rect 22520 26392 22526 26444
rect 23661 26435 23719 26441
rect 23661 26401 23673 26435
rect 23707 26432 23719 26435
rect 23842 26432 23848 26444
rect 23707 26404 23848 26432
rect 23707 26401 23719 26404
rect 23661 26395 23719 26401
rect 23842 26392 23848 26404
rect 23900 26392 23906 26444
rect 24673 26435 24731 26441
rect 24673 26401 24685 26435
rect 24719 26432 24731 26435
rect 24854 26432 24860 26444
rect 24719 26404 24860 26432
rect 24719 26401 24731 26404
rect 24673 26395 24731 26401
rect 24854 26392 24860 26404
rect 24912 26392 24918 26444
rect 25133 26435 25191 26441
rect 25133 26401 25145 26435
rect 25179 26432 25191 26435
rect 26237 26435 26295 26441
rect 26237 26432 26249 26435
rect 25179 26404 26249 26432
rect 25179 26401 25191 26404
rect 25133 26395 25191 26401
rect 26237 26401 26249 26404
rect 26283 26432 26295 26435
rect 26602 26432 26608 26444
rect 26283 26404 26608 26432
rect 26283 26401 26295 26404
rect 26237 26395 26295 26401
rect 26602 26392 26608 26404
rect 26660 26392 26666 26444
rect 29730 26432 29736 26444
rect 28920 26404 29736 26432
rect 19613 26367 19671 26373
rect 19613 26364 19625 26367
rect 19392 26336 19625 26364
rect 19392 26324 19398 26336
rect 19613 26333 19625 26336
rect 19659 26333 19671 26367
rect 19613 26327 19671 26333
rect 20165 26367 20223 26373
rect 20165 26333 20177 26367
rect 20211 26333 20223 26367
rect 20806 26364 20812 26376
rect 20767 26336 20812 26364
rect 20165 26327 20223 26333
rect 20806 26324 20812 26336
rect 20864 26324 20870 26376
rect 23198 26364 23204 26376
rect 23159 26336 23204 26364
rect 23198 26324 23204 26336
rect 23256 26324 23262 26376
rect 23474 26324 23480 26376
rect 23532 26373 23538 26376
rect 23532 26367 23561 26373
rect 23549 26333 23561 26367
rect 23532 26327 23561 26333
rect 25869 26367 25927 26373
rect 25869 26333 25881 26367
rect 25915 26333 25927 26367
rect 25869 26327 25927 26333
rect 25961 26367 26019 26373
rect 25961 26333 25973 26367
rect 26007 26364 26019 26367
rect 26786 26364 26792 26376
rect 26007 26336 26792 26364
rect 26007 26333 26019 26336
rect 25961 26327 26019 26333
rect 23532 26324 23538 26327
rect 17460 26268 17816 26296
rect 18156 26296 18184 26324
rect 18322 26296 18328 26308
rect 18156 26268 18328 26296
rect 17460 26256 17466 26268
rect 18156 26228 18184 26268
rect 18322 26256 18328 26268
rect 18380 26256 18386 26308
rect 20257 26299 20315 26305
rect 20257 26265 20269 26299
rect 20303 26296 20315 26299
rect 20530 26296 20536 26308
rect 20303 26268 20536 26296
rect 20303 26265 20315 26268
rect 20257 26259 20315 26265
rect 20530 26256 20536 26268
rect 20588 26256 20594 26308
rect 23290 26296 23296 26308
rect 23251 26268 23296 26296
rect 23290 26256 23296 26268
rect 23348 26256 23354 26308
rect 23382 26256 23388 26308
rect 23440 26296 23446 26308
rect 25406 26296 25412 26308
rect 23440 26268 25412 26296
rect 23440 26256 23446 26268
rect 25406 26256 25412 26268
rect 25464 26256 25470 26308
rect 25884 26296 25912 26327
rect 26786 26324 26792 26336
rect 26844 26324 26850 26376
rect 27157 26367 27215 26373
rect 27157 26333 27169 26367
rect 27203 26364 27215 26367
rect 28920 26364 28948 26404
rect 29730 26392 29736 26404
rect 29788 26392 29794 26444
rect 29840 26432 29868 26540
rect 30101 26537 30113 26571
rect 30147 26568 30159 26571
rect 30190 26568 30196 26580
rect 30147 26540 30196 26568
rect 30147 26537 30159 26540
rect 30101 26531 30159 26537
rect 30190 26528 30196 26540
rect 30248 26528 30254 26580
rect 31573 26571 31631 26577
rect 31573 26537 31585 26571
rect 31619 26568 31631 26571
rect 33686 26568 33692 26580
rect 31619 26540 33692 26568
rect 31619 26537 31631 26540
rect 31573 26531 31631 26537
rect 33686 26528 33692 26540
rect 33744 26528 33750 26580
rect 29914 26460 29920 26512
rect 29972 26500 29978 26512
rect 30469 26503 30527 26509
rect 30469 26500 30481 26503
rect 29972 26472 30481 26500
rect 29972 26460 29978 26472
rect 30469 26469 30481 26472
rect 30515 26469 30527 26503
rect 32033 26503 32091 26509
rect 30469 26463 30527 26469
rect 30852 26472 31892 26500
rect 30852 26444 30880 26472
rect 30561 26435 30619 26441
rect 29840 26404 30420 26432
rect 27203 26336 28948 26364
rect 28997 26367 29055 26373
rect 27203 26333 27215 26336
rect 27157 26327 27215 26333
rect 28997 26333 29009 26367
rect 29043 26333 29055 26367
rect 28997 26327 29055 26333
rect 29181 26367 29239 26373
rect 29181 26333 29193 26367
rect 29227 26333 29239 26367
rect 30282 26364 30288 26376
rect 30243 26336 30288 26364
rect 29181 26327 29239 26333
rect 26050 26296 26056 26308
rect 25884 26268 26056 26296
rect 26050 26256 26056 26268
rect 26108 26256 26114 26308
rect 27424 26299 27482 26305
rect 27424 26265 27436 26299
rect 27470 26296 27482 26299
rect 27522 26296 27528 26308
rect 27470 26268 27528 26296
rect 27470 26265 27482 26268
rect 27424 26259 27482 26265
rect 27522 26256 27528 26268
rect 27580 26256 27586 26308
rect 29012 26296 29040 26327
rect 27632 26268 29040 26296
rect 29196 26296 29224 26327
rect 30282 26324 30288 26336
rect 30340 26324 30346 26376
rect 30392 26364 30420 26404
rect 30561 26401 30573 26435
rect 30607 26432 30619 26435
rect 30834 26432 30840 26444
rect 30607 26404 30840 26432
rect 30607 26401 30619 26404
rect 30561 26395 30619 26401
rect 30834 26392 30840 26404
rect 30892 26392 30898 26444
rect 31570 26364 31576 26376
rect 30392 26336 31576 26364
rect 31570 26324 31576 26336
rect 31628 26324 31634 26376
rect 31754 26364 31760 26376
rect 31715 26336 31760 26364
rect 31754 26324 31760 26336
rect 31812 26324 31818 26376
rect 31864 26373 31892 26472
rect 32033 26469 32045 26503
rect 32079 26500 32091 26503
rect 32674 26500 32680 26512
rect 32079 26472 32680 26500
rect 32079 26469 32091 26472
rect 32033 26463 32091 26469
rect 32674 26460 32680 26472
rect 32732 26460 32738 26512
rect 32398 26392 32404 26444
rect 32456 26432 32462 26444
rect 32456 26404 32904 26432
rect 32456 26392 32462 26404
rect 31849 26367 31907 26373
rect 31849 26333 31861 26367
rect 31895 26333 31907 26367
rect 32122 26364 32128 26376
rect 32083 26336 32128 26364
rect 31849 26327 31907 26333
rect 30926 26296 30932 26308
rect 29196 26268 30932 26296
rect 17328 26200 18184 26228
rect 18414 26188 18420 26240
rect 18472 26228 18478 26240
rect 18785 26231 18843 26237
rect 18785 26228 18797 26231
rect 18472 26200 18797 26228
rect 18472 26188 18478 26200
rect 18785 26197 18797 26200
rect 18831 26197 18843 26231
rect 23014 26228 23020 26240
rect 22975 26200 23020 26228
rect 18785 26191 18843 26197
rect 23014 26188 23020 26200
rect 23072 26188 23078 26240
rect 25590 26188 25596 26240
rect 25648 26228 25654 26240
rect 25685 26231 25743 26237
rect 25685 26228 25697 26231
rect 25648 26200 25697 26228
rect 25648 26188 25654 26200
rect 25685 26197 25697 26200
rect 25731 26197 25743 26231
rect 25685 26191 25743 26197
rect 26878 26188 26884 26240
rect 26936 26228 26942 26240
rect 27632 26228 27660 26268
rect 30926 26256 30932 26268
rect 30984 26256 30990 26308
rect 31864 26296 31892 26327
rect 32122 26324 32128 26336
rect 32180 26324 32186 26376
rect 32306 26324 32312 26376
rect 32364 26364 32370 26376
rect 32769 26367 32827 26373
rect 32769 26364 32781 26367
rect 32364 26336 32781 26364
rect 32364 26324 32370 26336
rect 32769 26333 32781 26336
rect 32815 26333 32827 26367
rect 32876 26364 32904 26404
rect 33025 26367 33083 26373
rect 33025 26364 33037 26367
rect 32876 26336 33037 26364
rect 32769 26327 32827 26333
rect 33025 26333 33037 26336
rect 33071 26333 33083 26367
rect 33025 26327 33083 26333
rect 32398 26296 32404 26308
rect 31864 26268 32404 26296
rect 32398 26256 32404 26268
rect 32456 26256 32462 26308
rect 32674 26256 32680 26308
rect 32732 26296 32738 26308
rect 33410 26296 33416 26308
rect 32732 26268 33416 26296
rect 32732 26256 32738 26268
rect 33410 26256 33416 26268
rect 33468 26256 33474 26308
rect 26936 26200 27660 26228
rect 26936 26188 26942 26200
rect 27798 26188 27804 26240
rect 27856 26228 27862 26240
rect 28258 26228 28264 26240
rect 27856 26200 28264 26228
rect 27856 26188 27862 26200
rect 28258 26188 28264 26200
rect 28316 26188 28322 26240
rect 28718 26188 28724 26240
rect 28776 26228 28782 26240
rect 29546 26228 29552 26240
rect 28776 26200 29552 26228
rect 28776 26188 28782 26200
rect 29546 26188 29552 26200
rect 29604 26188 29610 26240
rect 29730 26188 29736 26240
rect 29788 26228 29794 26240
rect 31018 26228 31024 26240
rect 29788 26200 31024 26228
rect 29788 26188 29794 26200
rect 31018 26188 31024 26200
rect 31076 26188 31082 26240
rect 31478 26188 31484 26240
rect 31536 26228 31542 26240
rect 32122 26228 32128 26240
rect 31536 26200 32128 26228
rect 31536 26188 31542 26200
rect 32122 26188 32128 26200
rect 32180 26228 32186 26240
rect 33226 26228 33232 26240
rect 32180 26200 33232 26228
rect 32180 26188 32186 26200
rect 33226 26188 33232 26200
rect 33284 26228 33290 26240
rect 34149 26231 34207 26237
rect 34149 26228 34161 26231
rect 33284 26200 34161 26228
rect 33284 26188 33290 26200
rect 34149 26197 34161 26200
rect 34195 26197 34207 26231
rect 34149 26191 34207 26197
rect 1104 26138 35027 26160
rect 1104 26086 9390 26138
rect 9442 26086 9454 26138
rect 9506 26086 9518 26138
rect 9570 26086 9582 26138
rect 9634 26086 9646 26138
rect 9698 26086 17831 26138
rect 17883 26086 17895 26138
rect 17947 26086 17959 26138
rect 18011 26086 18023 26138
rect 18075 26086 18087 26138
rect 18139 26086 26272 26138
rect 26324 26086 26336 26138
rect 26388 26086 26400 26138
rect 26452 26086 26464 26138
rect 26516 26086 26528 26138
rect 26580 26086 34713 26138
rect 34765 26086 34777 26138
rect 34829 26086 34841 26138
rect 34893 26086 34905 26138
rect 34957 26086 34969 26138
rect 35021 26086 35027 26138
rect 1104 26064 35027 26086
rect 25774 26024 25780 26036
rect 15672 25996 25780 26024
rect 15672 25897 15700 25996
rect 25774 25984 25780 25996
rect 25832 25984 25838 26036
rect 26513 26027 26571 26033
rect 26513 25993 26525 26027
rect 26559 25993 26571 26027
rect 26513 25987 26571 25993
rect 17405 25959 17463 25965
rect 17405 25925 17417 25959
rect 17451 25956 17463 25959
rect 18138 25956 18144 25968
rect 17451 25928 18144 25956
rect 17451 25925 17463 25928
rect 17405 25919 17463 25925
rect 18138 25916 18144 25928
rect 18196 25916 18202 25968
rect 18230 25916 18236 25968
rect 18288 25956 18294 25968
rect 20714 25956 20720 25968
rect 18288 25928 18920 25956
rect 18288 25916 18294 25928
rect 15657 25891 15715 25897
rect 15657 25857 15669 25891
rect 15703 25857 15715 25891
rect 17586 25888 17592 25900
rect 17547 25860 17592 25888
rect 15657 25851 15715 25857
rect 17586 25848 17592 25860
rect 17644 25848 17650 25900
rect 17678 25848 17684 25900
rect 17736 25888 17742 25900
rect 17957 25891 18015 25897
rect 17736 25860 17781 25888
rect 17736 25848 17742 25860
rect 17957 25857 17969 25891
rect 18003 25888 18015 25891
rect 18322 25888 18328 25900
rect 18003 25860 18328 25888
rect 18003 25857 18015 25860
rect 17957 25851 18015 25857
rect 18322 25848 18328 25860
rect 18380 25848 18386 25900
rect 18598 25888 18604 25900
rect 18559 25860 18604 25888
rect 18598 25848 18604 25860
rect 18656 25848 18662 25900
rect 18782 25888 18788 25900
rect 18743 25860 18788 25888
rect 18782 25848 18788 25860
rect 18840 25848 18846 25900
rect 18892 25897 18920 25928
rect 19352 25928 20720 25956
rect 19352 25897 19380 25928
rect 20714 25916 20720 25928
rect 20772 25916 20778 25968
rect 22916 25959 22974 25965
rect 21468 25928 22876 25956
rect 18877 25891 18935 25897
rect 18877 25857 18889 25891
rect 18923 25857 18935 25891
rect 18877 25851 18935 25857
rect 19337 25891 19395 25897
rect 19337 25857 19349 25891
rect 19383 25857 19395 25891
rect 19337 25851 19395 25857
rect 19426 25848 19432 25900
rect 19484 25888 19490 25900
rect 21468 25897 21496 25928
rect 19593 25891 19651 25897
rect 19593 25888 19605 25891
rect 19484 25860 19605 25888
rect 19484 25848 19490 25860
rect 19593 25857 19605 25860
rect 19639 25857 19651 25891
rect 19593 25851 19651 25857
rect 21177 25891 21235 25897
rect 21177 25857 21189 25891
rect 21223 25857 21235 25891
rect 21177 25851 21235 25857
rect 21361 25891 21419 25897
rect 21361 25857 21373 25891
rect 21407 25857 21419 25891
rect 21361 25851 21419 25857
rect 21453 25891 21511 25897
rect 21453 25857 21465 25891
rect 21499 25857 21511 25891
rect 21453 25851 21511 25857
rect 22189 25891 22247 25897
rect 22189 25857 22201 25891
rect 22235 25888 22247 25891
rect 22370 25888 22376 25900
rect 22235 25860 22376 25888
rect 22235 25857 22247 25860
rect 22189 25851 22247 25857
rect 17402 25780 17408 25832
rect 17460 25820 17466 25832
rect 17865 25823 17923 25829
rect 17865 25820 17877 25823
rect 17460 25792 17877 25820
rect 17460 25780 17466 25792
rect 17865 25789 17877 25792
rect 17911 25789 17923 25823
rect 17865 25783 17923 25789
rect 16301 25755 16359 25761
rect 16301 25721 16313 25755
rect 16347 25752 16359 25755
rect 19334 25752 19340 25764
rect 16347 25724 19340 25752
rect 16347 25721 16359 25724
rect 16301 25715 16359 25721
rect 19334 25712 19340 25724
rect 19392 25712 19398 25764
rect 20438 25712 20444 25764
rect 20496 25752 20502 25764
rect 21192 25752 21220 25851
rect 20496 25724 21220 25752
rect 20496 25712 20502 25724
rect 1578 25644 1584 25696
rect 1636 25684 1642 25696
rect 2041 25687 2099 25693
rect 2041 25684 2053 25687
rect 1636 25656 2053 25684
rect 1636 25644 1642 25656
rect 2041 25653 2053 25656
rect 2087 25653 2099 25687
rect 2041 25647 2099 25653
rect 17402 25644 17408 25696
rect 17460 25684 17466 25696
rect 18417 25687 18475 25693
rect 18417 25684 18429 25687
rect 17460 25656 18429 25684
rect 17460 25644 17466 25656
rect 18417 25653 18429 25656
rect 18463 25653 18475 25687
rect 18417 25647 18475 25653
rect 19610 25644 19616 25696
rect 19668 25684 19674 25696
rect 20717 25687 20775 25693
rect 20717 25684 20729 25687
rect 19668 25656 20729 25684
rect 19668 25644 19674 25656
rect 20717 25653 20729 25656
rect 20763 25684 20775 25687
rect 20898 25684 20904 25696
rect 20763 25656 20904 25684
rect 20763 25653 20775 25656
rect 20717 25647 20775 25653
rect 20898 25644 20904 25656
rect 20956 25644 20962 25696
rect 21174 25684 21180 25696
rect 21135 25656 21180 25684
rect 21174 25644 21180 25656
rect 21232 25644 21238 25696
rect 21376 25684 21404 25851
rect 22370 25848 22376 25860
rect 22428 25848 22434 25900
rect 22462 25848 22468 25900
rect 22520 25888 22526 25900
rect 22649 25891 22707 25897
rect 22649 25888 22661 25891
rect 22520 25860 22661 25888
rect 22520 25848 22526 25860
rect 22649 25857 22661 25860
rect 22695 25857 22707 25891
rect 22848 25888 22876 25928
rect 22916 25925 22928 25959
rect 22962 25956 22974 25959
rect 23014 25956 23020 25968
rect 22962 25928 23020 25956
rect 22962 25925 22974 25928
rect 22916 25919 22974 25925
rect 23014 25916 23020 25928
rect 23072 25916 23078 25968
rect 23842 25916 23848 25968
rect 23900 25956 23906 25968
rect 24734 25959 24792 25965
rect 24734 25956 24746 25959
rect 23900 25928 24746 25956
rect 23900 25916 23906 25928
rect 24734 25925 24746 25928
rect 24780 25925 24792 25959
rect 24734 25919 24792 25925
rect 25406 25916 25412 25968
rect 25464 25956 25470 25968
rect 26528 25956 26556 25987
rect 27430 25984 27436 26036
rect 27488 26024 27494 26036
rect 27488 25996 32536 26024
rect 27488 25984 27494 25996
rect 27522 25956 27528 25968
rect 25464 25928 26556 25956
rect 27483 25928 27528 25956
rect 25464 25916 25470 25928
rect 24578 25888 24584 25900
rect 22848 25860 24584 25888
rect 22649 25851 22707 25857
rect 24578 25848 24584 25860
rect 24636 25848 24642 25900
rect 25866 25848 25872 25900
rect 25924 25888 25930 25900
rect 26329 25891 26387 25897
rect 26329 25888 26341 25891
rect 25924 25860 26341 25888
rect 25924 25848 25930 25860
rect 26329 25857 26341 25860
rect 26375 25857 26387 25891
rect 26329 25851 26387 25857
rect 24302 25780 24308 25832
rect 24360 25820 24366 25832
rect 24489 25823 24547 25829
rect 24489 25820 24501 25823
rect 24360 25792 24501 25820
rect 24360 25780 24366 25792
rect 24489 25789 24501 25792
rect 24535 25789 24547 25823
rect 26528 25820 26556 25928
rect 27522 25916 27528 25928
rect 27580 25916 27586 25968
rect 29086 25956 29092 25968
rect 27908 25928 28580 25956
rect 27908 25900 27936 25928
rect 27338 25848 27344 25900
rect 27396 25888 27402 25900
rect 27614 25888 27620 25900
rect 27396 25860 27620 25888
rect 27396 25848 27402 25860
rect 27614 25848 27620 25860
rect 27672 25848 27678 25900
rect 27798 25888 27804 25900
rect 27759 25860 27804 25888
rect 27798 25848 27804 25860
rect 27856 25848 27862 25900
rect 27893 25894 27951 25900
rect 27893 25860 27905 25894
rect 27939 25860 27951 25894
rect 27893 25854 27951 25860
rect 27982 25848 27988 25900
rect 28040 25888 28046 25900
rect 28040 25860 28085 25888
rect 28040 25848 28046 25860
rect 28166 25848 28172 25900
rect 28224 25888 28230 25900
rect 28224 25860 28269 25888
rect 28224 25848 28230 25860
rect 28552 25820 28580 25928
rect 28644 25928 29092 25956
rect 28644 25897 28672 25928
rect 29086 25916 29092 25928
rect 29144 25916 29150 25968
rect 31297 25959 31355 25965
rect 31297 25925 31309 25959
rect 31343 25956 31355 25959
rect 31754 25956 31760 25968
rect 31343 25928 31760 25956
rect 31343 25925 31355 25928
rect 31297 25919 31355 25925
rect 31754 25916 31760 25928
rect 31812 25916 31818 25968
rect 28629 25891 28687 25897
rect 28629 25857 28641 25891
rect 28675 25857 28687 25891
rect 28629 25851 28687 25857
rect 28718 25848 28724 25900
rect 28776 25848 28782 25900
rect 28896 25891 28954 25897
rect 28896 25857 28908 25891
rect 28942 25888 28954 25891
rect 29362 25888 29368 25900
rect 28942 25860 29368 25888
rect 28942 25857 28954 25860
rect 28896 25851 28954 25857
rect 29362 25848 29368 25860
rect 29420 25848 29426 25900
rect 31018 25888 31024 25900
rect 30979 25860 31024 25888
rect 31018 25848 31024 25860
rect 31076 25848 31082 25900
rect 31169 25891 31227 25897
rect 31169 25857 31181 25891
rect 31215 25888 31227 25891
rect 31386 25888 31392 25900
rect 31215 25857 31248 25888
rect 31347 25860 31392 25888
rect 31169 25851 31248 25857
rect 28736 25820 28764 25848
rect 26528 25792 27936 25820
rect 24489 25783 24547 25789
rect 27908 25764 27936 25792
rect 28552 25792 28764 25820
rect 31220 25820 31248 25851
rect 31386 25848 31392 25860
rect 31444 25848 31450 25900
rect 31478 25848 31484 25900
rect 31536 25897 31542 25900
rect 32508 25897 32536 25996
rect 31536 25888 31544 25897
rect 32493 25891 32551 25897
rect 31536 25860 31581 25888
rect 31536 25851 31544 25860
rect 32493 25857 32505 25891
rect 32539 25857 32551 25891
rect 34330 25888 34336 25900
rect 34291 25860 34336 25888
rect 32493 25851 32551 25857
rect 31536 25848 31542 25851
rect 34330 25848 34336 25860
rect 34388 25848 34394 25900
rect 31938 25820 31944 25832
rect 31220 25792 31944 25820
rect 22002 25752 22008 25764
rect 21963 25724 22008 25752
rect 22002 25712 22008 25724
rect 22060 25712 22066 25764
rect 24029 25755 24087 25761
rect 24029 25721 24041 25755
rect 24075 25752 24087 25755
rect 24394 25752 24400 25764
rect 24075 25724 24400 25752
rect 24075 25721 24087 25724
rect 24029 25715 24087 25721
rect 24394 25712 24400 25724
rect 24452 25712 24458 25764
rect 25682 25712 25688 25764
rect 25740 25752 25746 25764
rect 25869 25755 25927 25761
rect 25869 25752 25881 25755
rect 25740 25724 25881 25752
rect 25740 25712 25746 25724
rect 25869 25721 25881 25724
rect 25915 25752 25927 25755
rect 26970 25752 26976 25764
rect 25915 25724 26976 25752
rect 25915 25721 25927 25724
rect 25869 25715 25927 25721
rect 26970 25712 26976 25724
rect 27028 25752 27034 25764
rect 27246 25752 27252 25764
rect 27028 25724 27252 25752
rect 27028 25712 27034 25724
rect 27246 25712 27252 25724
rect 27304 25712 27310 25764
rect 27890 25712 27896 25764
rect 27948 25712 27954 25764
rect 28166 25712 28172 25764
rect 28224 25752 28230 25764
rect 28552 25752 28580 25792
rect 31938 25780 31944 25792
rect 31996 25780 32002 25832
rect 32677 25823 32735 25829
rect 32677 25789 32689 25823
rect 32723 25789 32735 25823
rect 32677 25783 32735 25789
rect 32692 25752 32720 25783
rect 28224 25724 28580 25752
rect 29564 25724 32720 25752
rect 28224 25712 28230 25724
rect 24486 25684 24492 25696
rect 21376 25656 24492 25684
rect 24486 25644 24492 25656
rect 24544 25644 24550 25696
rect 26418 25644 26424 25696
rect 26476 25684 26482 25696
rect 29564 25684 29592 25724
rect 26476 25656 29592 25684
rect 26476 25644 26482 25656
rect 29914 25644 29920 25696
rect 29972 25684 29978 25696
rect 30009 25687 30067 25693
rect 30009 25684 30021 25687
rect 29972 25656 30021 25684
rect 29972 25644 29978 25656
rect 30009 25653 30021 25656
rect 30055 25684 30067 25687
rect 31202 25684 31208 25696
rect 30055 25656 31208 25684
rect 30055 25653 30067 25656
rect 30009 25647 30067 25653
rect 31202 25644 31208 25656
rect 31260 25644 31266 25696
rect 31662 25684 31668 25696
rect 31623 25656 31668 25684
rect 31662 25644 31668 25656
rect 31720 25644 31726 25696
rect 1104 25594 34868 25616
rect 1104 25542 5170 25594
rect 5222 25542 5234 25594
rect 5286 25542 5298 25594
rect 5350 25542 5362 25594
rect 5414 25542 5426 25594
rect 5478 25542 13611 25594
rect 13663 25542 13675 25594
rect 13727 25542 13739 25594
rect 13791 25542 13803 25594
rect 13855 25542 13867 25594
rect 13919 25542 22052 25594
rect 22104 25542 22116 25594
rect 22168 25542 22180 25594
rect 22232 25542 22244 25594
rect 22296 25542 22308 25594
rect 22360 25542 30493 25594
rect 30545 25542 30557 25594
rect 30609 25542 30621 25594
rect 30673 25542 30685 25594
rect 30737 25542 30749 25594
rect 30801 25542 34868 25594
rect 1104 25520 34868 25542
rect 16577 25483 16635 25489
rect 16577 25449 16589 25483
rect 16623 25480 16635 25483
rect 18874 25480 18880 25492
rect 16623 25452 18880 25480
rect 16623 25449 16635 25452
rect 16577 25443 16635 25449
rect 18874 25440 18880 25452
rect 18932 25440 18938 25492
rect 19426 25480 19432 25492
rect 19387 25452 19432 25480
rect 19426 25440 19432 25452
rect 19484 25440 19490 25492
rect 23290 25440 23296 25492
rect 23348 25480 23354 25492
rect 23385 25483 23443 25489
rect 23385 25480 23397 25483
rect 23348 25452 23397 25480
rect 23348 25440 23354 25452
rect 23385 25449 23397 25452
rect 23431 25449 23443 25483
rect 24946 25480 24952 25492
rect 24907 25452 24952 25480
rect 23385 25443 23443 25449
rect 24946 25440 24952 25452
rect 25004 25440 25010 25492
rect 27893 25483 27951 25489
rect 27893 25449 27905 25483
rect 27939 25480 27951 25483
rect 27982 25480 27988 25492
rect 27939 25452 27988 25480
rect 27939 25449 27951 25452
rect 27893 25443 27951 25449
rect 27982 25440 27988 25452
rect 28040 25440 28046 25492
rect 28350 25440 28356 25492
rect 28408 25480 28414 25492
rect 29270 25480 29276 25492
rect 28408 25452 29276 25480
rect 28408 25440 28414 25452
rect 29270 25440 29276 25452
rect 29328 25440 29334 25492
rect 31018 25440 31024 25492
rect 31076 25480 31082 25492
rect 32033 25483 32091 25489
rect 32033 25480 32045 25483
rect 31076 25452 32045 25480
rect 31076 25440 31082 25452
rect 32033 25449 32045 25452
rect 32079 25449 32091 25483
rect 32033 25443 32091 25449
rect 20622 25412 20628 25424
rect 15948 25384 20628 25412
rect 1578 25344 1584 25356
rect 1539 25316 1584 25344
rect 1578 25304 1584 25316
rect 1636 25304 1642 25356
rect 2774 25344 2780 25356
rect 2735 25316 2780 25344
rect 2774 25304 2780 25316
rect 2832 25304 2838 25356
rect 15286 25276 15292 25288
rect 15247 25248 15292 25276
rect 15286 25236 15292 25248
rect 15344 25236 15350 25288
rect 15948 25285 15976 25384
rect 20622 25372 20628 25384
rect 20680 25372 20686 25424
rect 26050 25372 26056 25424
rect 26108 25412 26114 25424
rect 26108 25384 27384 25412
rect 26108 25372 26114 25384
rect 16025 25347 16083 25353
rect 16025 25313 16037 25347
rect 16071 25344 16083 25347
rect 18414 25344 18420 25356
rect 16071 25316 18296 25344
rect 18375 25316 18420 25344
rect 16071 25313 16083 25316
rect 16025 25307 16083 25313
rect 15933 25279 15991 25285
rect 15933 25245 15945 25279
rect 15979 25245 15991 25279
rect 16574 25276 16580 25288
rect 16535 25248 16580 25276
rect 15933 25239 15991 25245
rect 16574 25236 16580 25248
rect 16632 25236 16638 25288
rect 16761 25279 16819 25285
rect 16761 25245 16773 25279
rect 16807 25276 16819 25279
rect 17034 25276 17040 25288
rect 16807 25248 17040 25276
rect 16807 25245 16819 25248
rect 16761 25239 16819 25245
rect 17034 25236 17040 25248
rect 17092 25236 17098 25288
rect 17126 25236 17132 25288
rect 17184 25276 17190 25288
rect 17402 25276 17408 25288
rect 17184 25248 17408 25276
rect 17184 25236 17190 25248
rect 17402 25236 17408 25248
rect 17460 25236 17466 25288
rect 1762 25208 1768 25220
rect 1723 25180 1768 25208
rect 1762 25168 1768 25180
rect 1820 25168 1826 25220
rect 16850 25168 16856 25220
rect 16908 25208 16914 25220
rect 17221 25211 17279 25217
rect 17221 25208 17233 25211
rect 16908 25180 17233 25208
rect 16908 25168 16914 25180
rect 17221 25177 17233 25180
rect 17267 25177 17279 25211
rect 18046 25208 18052 25220
rect 17221 25171 17279 25177
rect 17420 25180 18052 25208
rect 15381 25143 15439 25149
rect 15381 25109 15393 25143
rect 15427 25140 15439 25143
rect 17420 25140 17448 25180
rect 18046 25168 18052 25180
rect 18104 25168 18110 25220
rect 18268 25208 18296 25316
rect 18414 25304 18420 25316
rect 18472 25304 18478 25356
rect 22462 25304 22468 25356
rect 22520 25344 22526 25356
rect 22830 25344 22836 25356
rect 22520 25316 22836 25344
rect 22520 25304 22526 25316
rect 22830 25304 22836 25316
rect 22888 25304 22894 25356
rect 25961 25347 26019 25353
rect 25961 25313 25973 25347
rect 26007 25344 26019 25347
rect 26142 25344 26148 25356
rect 26007 25316 26148 25344
rect 26007 25313 26019 25316
rect 25961 25307 26019 25313
rect 26142 25304 26148 25316
rect 26200 25304 26206 25356
rect 26326 25304 26332 25356
rect 26384 25344 26390 25356
rect 26421 25347 26479 25353
rect 26421 25344 26433 25347
rect 26384 25316 26433 25344
rect 26384 25304 26390 25316
rect 26421 25313 26433 25316
rect 26467 25344 26479 25347
rect 26510 25344 26516 25356
rect 26467 25316 26516 25344
rect 26467 25313 26479 25316
rect 26421 25307 26479 25313
rect 26510 25304 26516 25316
rect 26568 25304 26574 25356
rect 26694 25304 26700 25356
rect 26752 25344 26758 25356
rect 27356 25344 27384 25384
rect 27522 25372 27528 25424
rect 27580 25412 27586 25424
rect 28995 25412 29001 25424
rect 27580 25384 29001 25412
rect 27580 25372 27586 25384
rect 28995 25372 29001 25384
rect 29053 25372 29059 25424
rect 29181 25415 29239 25421
rect 29181 25381 29193 25415
rect 29227 25381 29239 25415
rect 29181 25375 29239 25381
rect 29196 25344 29224 25375
rect 31570 25344 31576 25356
rect 26752 25316 27292 25344
rect 27356 25316 29224 25344
rect 31531 25316 31576 25344
rect 26752 25304 26758 25316
rect 18325 25279 18383 25285
rect 18325 25245 18337 25279
rect 18371 25276 18383 25279
rect 18782 25276 18788 25288
rect 18371 25248 18788 25276
rect 18371 25245 18383 25248
rect 18325 25239 18383 25245
rect 18782 25236 18788 25248
rect 18840 25236 18846 25288
rect 19610 25236 19616 25288
rect 19668 25276 19674 25288
rect 19705 25279 19763 25285
rect 19705 25276 19717 25279
rect 19668 25248 19717 25276
rect 19668 25236 19674 25248
rect 19705 25245 19717 25248
rect 19751 25245 19763 25279
rect 19705 25239 19763 25245
rect 19797 25279 19855 25285
rect 19797 25245 19809 25279
rect 19843 25245 19855 25279
rect 19797 25239 19855 25245
rect 18598 25208 18604 25220
rect 18268 25180 18604 25208
rect 18598 25168 18604 25180
rect 18656 25168 18662 25220
rect 19058 25168 19064 25220
rect 19116 25208 19122 25220
rect 19812 25208 19840 25239
rect 19886 25236 19892 25288
rect 19944 25285 19950 25288
rect 19944 25276 19952 25285
rect 19944 25248 19989 25276
rect 19944 25239 19952 25248
rect 19944 25236 19950 25239
rect 20070 25236 20076 25288
rect 20128 25276 20134 25288
rect 20128 25248 20173 25276
rect 20128 25236 20134 25248
rect 20714 25236 20720 25288
rect 20772 25276 20778 25288
rect 20809 25279 20867 25285
rect 20809 25276 20821 25279
rect 20772 25248 20821 25276
rect 20772 25236 20778 25248
rect 20809 25245 20821 25248
rect 20855 25276 20867 25279
rect 21910 25276 21916 25288
rect 20855 25248 21916 25276
rect 20855 25245 20867 25248
rect 20809 25239 20867 25245
rect 21910 25236 21916 25248
rect 21968 25236 21974 25288
rect 23014 25236 23020 25288
rect 23072 25276 23078 25288
rect 23109 25279 23167 25285
rect 23109 25276 23121 25279
rect 23072 25248 23121 25276
rect 23072 25236 23078 25248
rect 23109 25245 23121 25248
rect 23155 25245 23167 25279
rect 23109 25239 23167 25245
rect 23382 25236 23388 25288
rect 23440 25276 23446 25288
rect 23845 25279 23903 25285
rect 23845 25276 23857 25279
rect 23440 25248 23857 25276
rect 23440 25236 23446 25248
rect 23845 25245 23857 25248
rect 23891 25245 23903 25279
rect 23845 25239 23903 25245
rect 24210 25236 24216 25288
rect 24268 25276 24274 25288
rect 25682 25276 25688 25288
rect 24268 25248 24624 25276
rect 25643 25248 25688 25276
rect 24268 25236 24274 25248
rect 24596 25220 24624 25248
rect 25682 25236 25688 25248
rect 25740 25236 25746 25288
rect 25869 25279 25927 25285
rect 25869 25245 25881 25279
rect 25915 25245 25927 25279
rect 26050 25276 26056 25288
rect 26011 25248 26056 25276
rect 25869 25239 25927 25245
rect 19116 25180 19840 25208
rect 21076 25211 21134 25217
rect 19116 25168 19122 25180
rect 21076 25177 21088 25211
rect 21122 25208 21134 25211
rect 21266 25208 21272 25220
rect 21122 25180 21272 25208
rect 21122 25177 21134 25180
rect 21076 25171 21134 25177
rect 21266 25168 21272 25180
rect 21324 25168 21330 25220
rect 23201 25211 23259 25217
rect 23201 25177 23213 25211
rect 23247 25208 23259 25211
rect 23290 25208 23296 25220
rect 23247 25180 23296 25208
rect 23247 25177 23259 25180
rect 23201 25171 23259 25177
rect 23290 25168 23296 25180
rect 23348 25168 23354 25220
rect 24578 25168 24584 25220
rect 24636 25208 24642 25220
rect 24673 25211 24731 25217
rect 24673 25208 24685 25211
rect 24636 25180 24685 25208
rect 24636 25168 24642 25180
rect 24673 25177 24685 25180
rect 24719 25208 24731 25211
rect 25406 25208 25412 25220
rect 24719 25180 25412 25208
rect 24719 25177 24731 25180
rect 24673 25171 24731 25177
rect 25406 25168 25412 25180
rect 25464 25168 25470 25220
rect 25884 25208 25912 25239
rect 26050 25236 26056 25248
rect 26108 25236 26114 25288
rect 26237 25279 26295 25285
rect 26237 25245 26249 25279
rect 26283 25276 26295 25279
rect 26602 25276 26608 25288
rect 26283 25248 26608 25276
rect 26283 25245 26295 25248
rect 26237 25239 26295 25245
rect 26602 25236 26608 25248
rect 26660 25236 26666 25288
rect 26786 25276 26792 25288
rect 26712 25248 26792 25276
rect 25884 25180 26556 25208
rect 17586 25140 17592 25152
rect 15427 25112 17448 25140
rect 17547 25112 17592 25140
rect 15427 25109 15439 25112
rect 15381 25103 15439 25109
rect 17586 25100 17592 25112
rect 17644 25100 17650 25152
rect 18693 25143 18751 25149
rect 18693 25109 18705 25143
rect 18739 25140 18751 25143
rect 18874 25140 18880 25152
rect 18739 25112 18880 25140
rect 18739 25109 18751 25112
rect 18693 25103 18751 25109
rect 18874 25100 18880 25112
rect 18932 25100 18938 25152
rect 22189 25143 22247 25149
rect 22189 25109 22201 25143
rect 22235 25140 22247 25143
rect 22922 25140 22928 25152
rect 22235 25112 22928 25140
rect 22235 25109 22247 25112
rect 22189 25103 22247 25109
rect 22922 25100 22928 25112
rect 22980 25140 22986 25152
rect 23017 25143 23075 25149
rect 23017 25140 23029 25143
rect 22980 25112 23029 25140
rect 22980 25100 22986 25112
rect 23017 25109 23029 25112
rect 23063 25109 23075 25143
rect 23017 25103 23075 25109
rect 23566 25100 23572 25152
rect 23624 25140 23630 25152
rect 23937 25143 23995 25149
rect 23937 25140 23949 25143
rect 23624 25112 23949 25140
rect 23624 25100 23630 25112
rect 23937 25109 23949 25112
rect 23983 25109 23995 25143
rect 26528 25140 26556 25180
rect 26712 25140 26740 25248
rect 26786 25236 26792 25248
rect 26844 25276 26850 25288
rect 27065 25279 27123 25285
rect 27065 25276 27077 25279
rect 26844 25248 27077 25276
rect 26844 25236 26850 25248
rect 27065 25245 27077 25248
rect 27111 25245 27123 25279
rect 27065 25239 27123 25245
rect 27157 25279 27215 25285
rect 27157 25245 27169 25279
rect 27203 25245 27215 25279
rect 27264 25276 27292 25316
rect 31570 25304 31576 25316
rect 31628 25304 31634 25356
rect 31665 25347 31723 25353
rect 31665 25313 31677 25347
rect 31711 25344 31723 25347
rect 31754 25344 31760 25356
rect 31711 25316 31760 25344
rect 31711 25313 31723 25316
rect 31665 25307 31723 25313
rect 31754 25304 31760 25316
rect 31812 25304 31818 25356
rect 32030 25304 32036 25356
rect 32088 25344 32094 25356
rect 32493 25347 32551 25353
rect 32493 25344 32505 25347
rect 32088 25316 32505 25344
rect 32088 25304 32094 25316
rect 32493 25313 32505 25316
rect 32539 25313 32551 25347
rect 32493 25307 32551 25313
rect 32677 25347 32735 25353
rect 32677 25313 32689 25347
rect 32723 25344 32735 25347
rect 32858 25344 32864 25356
rect 32723 25316 32864 25344
rect 32723 25313 32735 25316
rect 32677 25307 32735 25313
rect 32858 25304 32864 25316
rect 32916 25304 32922 25356
rect 27341 25279 27399 25285
rect 27341 25276 27353 25279
rect 27264 25248 27353 25276
rect 27157 25239 27215 25245
rect 27341 25245 27353 25248
rect 27387 25245 27399 25279
rect 27341 25239 27399 25245
rect 26970 25168 26976 25220
rect 27028 25208 27034 25220
rect 27172 25208 27200 25239
rect 27430 25236 27436 25288
rect 27488 25276 27494 25288
rect 28074 25276 28080 25288
rect 27488 25248 27533 25276
rect 28035 25248 28080 25276
rect 27488 25236 27494 25248
rect 28074 25236 28080 25248
rect 28132 25236 28138 25288
rect 28350 25276 28356 25288
rect 28311 25248 28356 25276
rect 28350 25236 28356 25248
rect 28408 25236 28414 25288
rect 28813 25279 28871 25285
rect 28813 25245 28825 25279
rect 28859 25274 28871 25279
rect 28997 25279 29055 25285
rect 28859 25245 28872 25274
rect 28813 25239 28872 25245
rect 28997 25245 29009 25279
rect 29043 25245 29055 25279
rect 28997 25239 29055 25245
rect 27028 25180 27200 25208
rect 27028 25168 27034 25180
rect 27246 25168 27252 25220
rect 27304 25208 27310 25220
rect 28844 25208 28872 25239
rect 27304 25180 28872 25208
rect 27304 25168 27310 25180
rect 26878 25140 26884 25152
rect 26528 25112 26740 25140
rect 26839 25112 26884 25140
rect 23937 25103 23995 25109
rect 26878 25100 26884 25112
rect 26936 25100 26942 25152
rect 28261 25143 28319 25149
rect 28261 25109 28273 25143
rect 28307 25140 28319 25143
rect 28350 25140 28356 25152
rect 28307 25112 28356 25140
rect 28307 25109 28319 25112
rect 28261 25103 28319 25109
rect 28350 25100 28356 25112
rect 28408 25100 28414 25152
rect 28442 25100 28448 25152
rect 28500 25140 28506 25152
rect 29012 25140 29040 25239
rect 30098 25236 30104 25288
rect 30156 25276 30162 25288
rect 30285 25279 30343 25285
rect 30285 25276 30297 25279
rect 30156 25248 30297 25276
rect 30156 25236 30162 25248
rect 30285 25245 30297 25248
rect 30331 25245 30343 25279
rect 30650 25276 30656 25288
rect 30611 25248 30656 25276
rect 30285 25239 30343 25245
rect 30650 25236 30656 25248
rect 30708 25236 30714 25288
rect 31110 25236 31116 25288
rect 31168 25276 31174 25288
rect 31297 25279 31355 25285
rect 31297 25276 31309 25279
rect 31168 25248 31309 25276
rect 31168 25236 31174 25248
rect 31297 25245 31309 25248
rect 31343 25245 31355 25279
rect 31297 25239 31355 25245
rect 31481 25279 31539 25285
rect 31481 25245 31493 25279
rect 31527 25245 31539 25279
rect 31481 25239 31539 25245
rect 31849 25279 31907 25285
rect 31849 25245 31861 25279
rect 31895 25276 31907 25279
rect 31938 25276 31944 25288
rect 31895 25248 31944 25276
rect 31895 25245 31907 25248
rect 31849 25239 31907 25245
rect 30374 25168 30380 25220
rect 30432 25208 30438 25220
rect 30469 25211 30527 25217
rect 30469 25208 30481 25211
rect 30432 25180 30481 25208
rect 30432 25168 30438 25180
rect 30469 25177 30481 25180
rect 30515 25177 30527 25211
rect 30469 25171 30527 25177
rect 30561 25211 30619 25217
rect 30561 25177 30573 25211
rect 30607 25208 30619 25211
rect 30742 25208 30748 25220
rect 30607 25180 30748 25208
rect 30607 25177 30619 25180
rect 30561 25171 30619 25177
rect 28500 25112 29040 25140
rect 28500 25100 28506 25112
rect 29638 25100 29644 25152
rect 29696 25140 29702 25152
rect 30576 25140 30604 25171
rect 30742 25168 30748 25180
rect 30800 25168 30806 25220
rect 31496 25208 31524 25239
rect 31938 25236 31944 25248
rect 31996 25236 32002 25288
rect 34054 25208 34060 25220
rect 31496 25180 34060 25208
rect 34054 25168 34060 25180
rect 34112 25168 34118 25220
rect 34330 25208 34336 25220
rect 34291 25180 34336 25208
rect 34330 25168 34336 25180
rect 34388 25168 34394 25220
rect 29696 25112 30604 25140
rect 30837 25143 30895 25149
rect 29696 25100 29702 25112
rect 30837 25109 30849 25143
rect 30883 25140 30895 25143
rect 31570 25140 31576 25152
rect 30883 25112 31576 25140
rect 30883 25109 30895 25112
rect 30837 25103 30895 25109
rect 31570 25100 31576 25112
rect 31628 25100 31634 25152
rect 1104 25050 35027 25072
rect 1104 24998 9390 25050
rect 9442 24998 9454 25050
rect 9506 24998 9518 25050
rect 9570 24998 9582 25050
rect 9634 24998 9646 25050
rect 9698 24998 17831 25050
rect 17883 24998 17895 25050
rect 17947 24998 17959 25050
rect 18011 24998 18023 25050
rect 18075 24998 18087 25050
rect 18139 24998 26272 25050
rect 26324 24998 26336 25050
rect 26388 24998 26400 25050
rect 26452 24998 26464 25050
rect 26516 24998 26528 25050
rect 26580 24998 34713 25050
rect 34765 24998 34777 25050
rect 34829 24998 34841 25050
rect 34893 24998 34905 25050
rect 34957 24998 34969 25050
rect 35021 24998 35027 25050
rect 1104 24976 35027 24998
rect 1762 24896 1768 24948
rect 1820 24936 1826 24948
rect 2133 24939 2191 24945
rect 2133 24936 2145 24939
rect 1820 24908 2145 24936
rect 1820 24896 1826 24908
rect 2133 24905 2145 24908
rect 2179 24905 2191 24939
rect 2133 24899 2191 24905
rect 16209 24939 16267 24945
rect 16209 24905 16221 24939
rect 16255 24936 16267 24939
rect 16574 24936 16580 24948
rect 16255 24908 16580 24936
rect 16255 24905 16267 24908
rect 16209 24899 16267 24905
rect 16574 24896 16580 24908
rect 16632 24896 16638 24948
rect 17310 24896 17316 24948
rect 17368 24936 17374 24948
rect 19610 24936 19616 24948
rect 17368 24908 19616 24936
rect 17368 24896 17374 24908
rect 19610 24896 19616 24908
rect 19668 24896 19674 24948
rect 23014 24896 23020 24948
rect 23072 24936 23078 24948
rect 23198 24936 23204 24948
rect 23072 24908 23204 24936
rect 23072 24896 23078 24908
rect 23198 24896 23204 24908
rect 23256 24936 23262 24948
rect 25685 24939 25743 24945
rect 25685 24936 25697 24939
rect 23256 24908 25697 24936
rect 23256 24896 23262 24908
rect 25685 24905 25697 24908
rect 25731 24905 25743 24939
rect 25685 24899 25743 24905
rect 26513 24939 26571 24945
rect 26513 24905 26525 24939
rect 26559 24936 26571 24939
rect 26602 24936 26608 24948
rect 26559 24908 26608 24936
rect 26559 24905 26571 24908
rect 26513 24899 26571 24905
rect 26602 24896 26608 24908
rect 26660 24936 26666 24948
rect 26970 24936 26976 24948
rect 26660 24908 26976 24936
rect 26660 24896 26666 24908
rect 26970 24896 26976 24908
rect 27028 24896 27034 24948
rect 27614 24896 27620 24948
rect 27672 24936 27678 24948
rect 27893 24939 27951 24945
rect 27893 24936 27905 24939
rect 27672 24908 27905 24936
rect 27672 24896 27678 24908
rect 27893 24905 27905 24908
rect 27939 24905 27951 24939
rect 27893 24899 27951 24905
rect 28350 24896 28356 24948
rect 28408 24936 28414 24948
rect 31938 24936 31944 24948
rect 28408 24908 31944 24936
rect 28408 24896 28414 24908
rect 31938 24896 31944 24908
rect 31996 24896 32002 24948
rect 17402 24868 17408 24880
rect 17363 24840 17408 24868
rect 17402 24828 17408 24840
rect 17460 24828 17466 24880
rect 17494 24828 17500 24880
rect 17552 24868 17558 24880
rect 17605 24871 17663 24877
rect 17605 24868 17617 24871
rect 17552 24840 17617 24868
rect 17552 24828 17558 24840
rect 17605 24837 17617 24840
rect 17651 24837 17663 24871
rect 17605 24831 17663 24837
rect 18969 24871 19027 24877
rect 18969 24837 18981 24871
rect 19015 24868 19027 24871
rect 19886 24868 19892 24880
rect 19015 24840 19892 24868
rect 19015 24837 19027 24840
rect 18969 24831 19027 24837
rect 19886 24828 19892 24840
rect 19944 24828 19950 24880
rect 20714 24868 20720 24880
rect 20272 24840 20720 24868
rect 2038 24800 2044 24812
rect 1999 24772 2044 24800
rect 2038 24760 2044 24772
rect 2096 24800 2102 24812
rect 3050 24800 3056 24812
rect 2096 24772 3056 24800
rect 2096 24760 2102 24772
rect 3050 24760 3056 24772
rect 3108 24760 3114 24812
rect 16022 24800 16028 24812
rect 15983 24772 16028 24800
rect 16022 24760 16028 24772
rect 16080 24760 16086 24812
rect 17218 24760 17224 24812
rect 17276 24800 17282 24812
rect 18233 24803 18291 24809
rect 18233 24800 18245 24803
rect 17276 24772 18245 24800
rect 17276 24760 17282 24772
rect 18233 24769 18245 24772
rect 18279 24769 18291 24803
rect 18233 24763 18291 24769
rect 18322 24760 18328 24812
rect 18380 24800 18386 24812
rect 18417 24803 18475 24809
rect 18417 24800 18429 24803
rect 18380 24772 18429 24800
rect 18380 24760 18386 24772
rect 18417 24769 18429 24772
rect 18463 24769 18475 24803
rect 18874 24800 18880 24812
rect 18835 24772 18880 24800
rect 18417 24763 18475 24769
rect 18874 24760 18880 24772
rect 18932 24760 18938 24812
rect 19058 24800 19064 24812
rect 19019 24772 19064 24800
rect 19058 24760 19064 24772
rect 19116 24760 19122 24812
rect 19705 24803 19763 24809
rect 19705 24769 19717 24803
rect 19751 24800 19763 24803
rect 20272 24800 20300 24840
rect 20714 24828 20720 24840
rect 20772 24828 20778 24880
rect 22554 24868 22560 24880
rect 21284 24840 22560 24868
rect 19751 24772 20300 24800
rect 20349 24803 20407 24809
rect 19751 24769 19763 24772
rect 19705 24763 19763 24769
rect 20349 24769 20361 24803
rect 20395 24769 20407 24803
rect 20349 24763 20407 24769
rect 20441 24803 20499 24809
rect 20441 24769 20453 24803
rect 20487 24800 20499 24803
rect 21174 24800 21180 24812
rect 20487 24772 21180 24800
rect 20487 24769 20499 24772
rect 20441 24763 20499 24769
rect 18598 24692 18604 24744
rect 18656 24732 18662 24744
rect 19076 24732 19104 24760
rect 18656 24704 19104 24732
rect 20364 24732 20392 24763
rect 21174 24760 21180 24772
rect 21232 24760 21238 24812
rect 21284 24809 21312 24840
rect 22554 24828 22560 24840
rect 22612 24828 22618 24880
rect 22664 24840 22968 24868
rect 21269 24803 21327 24809
rect 21269 24769 21281 24803
rect 21315 24769 21327 24803
rect 21450 24800 21456 24812
rect 21411 24772 21456 24800
rect 21269 24763 21327 24769
rect 21450 24760 21456 24772
rect 21508 24760 21514 24812
rect 21910 24760 21916 24812
rect 21968 24800 21974 24812
rect 22465 24803 22523 24809
rect 22465 24800 22477 24803
rect 21968 24772 22477 24800
rect 21968 24760 21974 24772
rect 22465 24769 22477 24772
rect 22511 24800 22523 24803
rect 22664 24800 22692 24840
rect 22738 24809 22744 24812
rect 22511 24772 22692 24800
rect 22511 24769 22523 24772
rect 22465 24763 22523 24769
rect 22732 24763 22744 24809
rect 22796 24800 22802 24812
rect 22940 24800 22968 24840
rect 24670 24828 24676 24880
rect 24728 24828 24734 24880
rect 25498 24828 25504 24880
rect 25556 24868 25562 24880
rect 26694 24868 26700 24880
rect 25556 24840 26700 24868
rect 25556 24828 25562 24840
rect 24302 24800 24308 24812
rect 22796 24772 22832 24800
rect 22940 24772 24308 24800
rect 22738 24760 22744 24763
rect 22796 24760 22802 24772
rect 24302 24760 24308 24772
rect 24360 24760 24366 24812
rect 24561 24803 24619 24809
rect 24561 24800 24573 24803
rect 24412 24772 24573 24800
rect 20530 24732 20536 24744
rect 20364 24704 20536 24732
rect 18656 24692 18662 24704
rect 20530 24692 20536 24704
rect 20588 24692 20594 24744
rect 20625 24735 20683 24741
rect 20625 24701 20637 24735
rect 20671 24732 20683 24735
rect 20990 24732 20996 24744
rect 20671 24704 20996 24732
rect 20671 24701 20683 24704
rect 20625 24695 20683 24701
rect 20990 24692 20996 24704
rect 21048 24692 21054 24744
rect 21085 24735 21143 24741
rect 21085 24701 21097 24735
rect 21131 24732 21143 24735
rect 22370 24732 22376 24744
rect 21131 24704 22376 24732
rect 21131 24701 21143 24704
rect 21085 24695 21143 24701
rect 22370 24692 22376 24704
rect 22428 24692 22434 24744
rect 24412 24732 24440 24772
rect 24561 24769 24573 24772
rect 24607 24769 24619 24803
rect 24688 24800 24716 24828
rect 26344 24809 26372 24840
rect 26694 24828 26700 24840
rect 26752 24828 26758 24880
rect 27062 24828 27068 24880
rect 27120 24868 27126 24880
rect 28442 24868 28448 24880
rect 27120 24840 28448 24868
rect 27120 24828 27126 24840
rect 28442 24828 28448 24840
rect 28500 24828 28506 24880
rect 29730 24868 29736 24880
rect 28644 24840 29736 24868
rect 26329 24803 26387 24809
rect 24688 24772 26280 24800
rect 24561 24763 24619 24769
rect 23492 24704 24440 24732
rect 26252 24732 26280 24772
rect 26329 24769 26341 24803
rect 26375 24769 26387 24803
rect 26329 24763 26387 24769
rect 26605 24803 26663 24809
rect 26605 24769 26617 24803
rect 26651 24800 26663 24803
rect 26786 24800 26792 24812
rect 26651 24772 26792 24800
rect 26651 24769 26663 24772
rect 26605 24763 26663 24769
rect 26786 24760 26792 24772
rect 26844 24760 26850 24812
rect 27709 24803 27767 24809
rect 27709 24800 27721 24803
rect 26896 24772 27721 24800
rect 26896 24732 26924 24772
rect 27709 24769 27721 24772
rect 27755 24769 27767 24803
rect 27709 24763 27767 24769
rect 27985 24803 28043 24809
rect 27985 24769 27997 24803
rect 28031 24800 28043 24803
rect 28166 24800 28172 24812
rect 28031 24772 28172 24800
rect 28031 24769 28043 24772
rect 27985 24763 28043 24769
rect 28166 24760 28172 24772
rect 28224 24760 28230 24812
rect 28644 24800 28672 24840
rect 29730 24828 29736 24840
rect 29788 24828 29794 24880
rect 30558 24868 30564 24880
rect 30116 24840 30564 24868
rect 28368 24772 28672 24800
rect 28712 24803 28770 24809
rect 26252 24704 26924 24732
rect 27525 24735 27583 24741
rect 19521 24667 19579 24673
rect 19521 24633 19533 24667
rect 19567 24664 19579 24667
rect 19567 24636 22094 24664
rect 19567 24633 19579 24636
rect 19521 24627 19579 24633
rect 17310 24556 17316 24608
rect 17368 24596 17374 24608
rect 17589 24599 17647 24605
rect 17589 24596 17601 24599
rect 17368 24568 17601 24596
rect 17368 24556 17374 24568
rect 17589 24565 17601 24568
rect 17635 24565 17647 24599
rect 17589 24559 17647 24565
rect 17678 24556 17684 24608
rect 17736 24596 17742 24608
rect 17773 24599 17831 24605
rect 17773 24596 17785 24599
rect 17736 24568 17785 24596
rect 17736 24556 17742 24568
rect 17773 24565 17785 24568
rect 17819 24565 17831 24599
rect 18322 24596 18328 24608
rect 18283 24568 18328 24596
rect 17773 24559 17831 24565
rect 18322 24556 18328 24568
rect 18380 24556 18386 24608
rect 20533 24599 20591 24605
rect 20533 24565 20545 24599
rect 20579 24596 20591 24599
rect 20622 24596 20628 24608
rect 20579 24568 20628 24596
rect 20579 24565 20591 24568
rect 20533 24559 20591 24565
rect 20622 24556 20628 24568
rect 20680 24556 20686 24608
rect 22066 24596 22094 24636
rect 23492 24596 23520 24704
rect 27525 24701 27537 24735
rect 27571 24732 27583 24735
rect 28368 24732 28396 24772
rect 28712 24769 28724 24803
rect 28758 24800 28770 24803
rect 30116 24800 30144 24840
rect 30558 24828 30564 24840
rect 30616 24828 30622 24880
rect 30650 24828 30656 24880
rect 30708 24868 30714 24880
rect 31570 24868 31576 24880
rect 30708 24840 31576 24868
rect 30708 24828 30714 24840
rect 28758 24772 30144 24800
rect 28758 24769 28770 24772
rect 28712 24763 28770 24769
rect 30190 24760 30196 24812
rect 30248 24800 30254 24812
rect 30285 24803 30343 24809
rect 30285 24800 30297 24803
rect 30248 24772 30297 24800
rect 30248 24760 30254 24772
rect 30285 24769 30297 24772
rect 30331 24769 30343 24803
rect 30285 24763 30343 24769
rect 30469 24803 30527 24809
rect 30469 24769 30481 24803
rect 30515 24800 30527 24803
rect 31018 24800 31024 24812
rect 30515 24772 31024 24800
rect 30515 24769 30527 24772
rect 30469 24763 30527 24769
rect 27571 24704 28396 24732
rect 28445 24735 28503 24741
rect 27571 24701 27583 24704
rect 27525 24695 27583 24701
rect 28445 24701 28457 24735
rect 28491 24701 28503 24735
rect 28445 24695 28503 24701
rect 23842 24596 23848 24608
rect 22066 24568 23520 24596
rect 23803 24568 23848 24596
rect 23842 24556 23848 24568
rect 23900 24556 23906 24608
rect 26145 24599 26203 24605
rect 26145 24565 26157 24599
rect 26191 24596 26203 24599
rect 27062 24596 27068 24608
rect 26191 24568 27068 24596
rect 26191 24565 26203 24568
rect 26145 24559 26203 24565
rect 27062 24556 27068 24568
rect 27120 24556 27126 24608
rect 28460 24596 28488 24695
rect 29546 24692 29552 24744
rect 29604 24732 29610 24744
rect 30484 24732 30512 24763
rect 31018 24760 31024 24772
rect 31076 24760 31082 24812
rect 31312 24809 31340 24840
rect 31570 24828 31576 24840
rect 31628 24828 31634 24880
rect 31846 24828 31852 24880
rect 31904 24868 31910 24880
rect 33594 24868 33600 24880
rect 31904 24840 32720 24868
rect 33555 24840 33600 24868
rect 31904 24828 31910 24840
rect 32692 24812 32720 24840
rect 33594 24828 33600 24840
rect 33652 24828 33658 24880
rect 31297 24803 31355 24809
rect 31297 24769 31309 24803
rect 31343 24769 31355 24803
rect 31297 24763 31355 24769
rect 31389 24803 31447 24809
rect 31389 24769 31401 24803
rect 31435 24800 31447 24803
rect 31478 24800 31484 24812
rect 31435 24772 31484 24800
rect 31435 24769 31447 24772
rect 31389 24763 31447 24769
rect 31478 24760 31484 24772
rect 31536 24760 31542 24812
rect 31665 24803 31723 24809
rect 31665 24769 31677 24803
rect 31711 24800 31723 24803
rect 32309 24803 32367 24809
rect 32309 24800 32321 24803
rect 31711 24772 32321 24800
rect 31711 24769 31723 24772
rect 31665 24763 31723 24769
rect 32309 24769 32321 24772
rect 32355 24769 32367 24803
rect 32309 24763 32367 24769
rect 32493 24803 32551 24809
rect 32493 24769 32505 24803
rect 32539 24769 32551 24803
rect 32493 24763 32551 24769
rect 32585 24803 32643 24809
rect 32585 24769 32597 24803
rect 32631 24769 32643 24803
rect 32585 24763 32643 24769
rect 29604 24704 30512 24732
rect 29604 24692 29610 24704
rect 31202 24692 31208 24744
rect 31260 24732 31266 24744
rect 31680 24732 31708 24763
rect 32508 24732 32536 24763
rect 31260 24704 31708 24732
rect 32140 24704 32536 24732
rect 31260 24692 31266 24704
rect 32140 24676 32168 24704
rect 30742 24624 30748 24676
rect 30800 24664 30806 24676
rect 31478 24664 31484 24676
rect 30800 24636 31484 24664
rect 30800 24624 30806 24636
rect 31478 24624 31484 24636
rect 31536 24624 31542 24676
rect 31573 24667 31631 24673
rect 31573 24633 31585 24667
rect 31619 24664 31631 24667
rect 32122 24664 32128 24676
rect 31619 24636 32128 24664
rect 31619 24633 31631 24636
rect 31573 24627 31631 24633
rect 32122 24624 32128 24636
rect 32180 24624 32186 24676
rect 32398 24624 32404 24676
rect 32456 24664 32462 24676
rect 32600 24664 32628 24763
rect 32674 24760 32680 24812
rect 32732 24800 32738 24812
rect 32732 24772 32777 24800
rect 32732 24760 32738 24772
rect 33226 24760 33232 24812
rect 33284 24800 33290 24812
rect 33321 24803 33379 24809
rect 33321 24800 33333 24803
rect 33284 24772 33333 24800
rect 33284 24760 33290 24772
rect 33321 24769 33333 24772
rect 33367 24769 33379 24803
rect 33321 24763 33379 24769
rect 33410 24760 33416 24812
rect 33468 24800 33474 24812
rect 33505 24803 33563 24809
rect 33505 24800 33517 24803
rect 33468 24772 33517 24800
rect 33468 24760 33474 24772
rect 33505 24769 33517 24772
rect 33551 24769 33563 24803
rect 33505 24763 33563 24769
rect 33689 24803 33747 24809
rect 33689 24769 33701 24803
rect 33735 24800 33747 24803
rect 34054 24800 34060 24812
rect 33735 24772 34060 24800
rect 33735 24769 33747 24772
rect 33689 24763 33747 24769
rect 34054 24760 34060 24772
rect 34112 24760 34118 24812
rect 32456 24636 32628 24664
rect 32456 24624 32462 24636
rect 33502 24624 33508 24676
rect 33560 24664 33566 24676
rect 33873 24667 33931 24673
rect 33873 24664 33885 24667
rect 33560 24636 33885 24664
rect 33560 24624 33566 24636
rect 33873 24633 33885 24636
rect 33919 24633 33931 24667
rect 33873 24627 33931 24633
rect 29086 24596 29092 24608
rect 28460 24568 29092 24596
rect 29086 24556 29092 24568
rect 29144 24556 29150 24608
rect 29730 24556 29736 24608
rect 29788 24596 29794 24608
rect 29825 24599 29883 24605
rect 29825 24596 29837 24599
rect 29788 24568 29837 24596
rect 29788 24556 29794 24568
rect 29825 24565 29837 24568
rect 29871 24565 29883 24599
rect 29825 24559 29883 24565
rect 29914 24556 29920 24608
rect 29972 24596 29978 24608
rect 30653 24599 30711 24605
rect 30653 24596 30665 24599
rect 29972 24568 30665 24596
rect 29972 24556 29978 24568
rect 30653 24565 30665 24568
rect 30699 24565 30711 24599
rect 31110 24596 31116 24608
rect 31071 24568 31116 24596
rect 30653 24559 30711 24565
rect 31110 24556 31116 24568
rect 31168 24556 31174 24608
rect 31846 24556 31852 24608
rect 31904 24596 31910 24608
rect 32861 24599 32919 24605
rect 32861 24596 32873 24599
rect 31904 24568 32873 24596
rect 31904 24556 31910 24568
rect 32861 24565 32873 24568
rect 32907 24565 32919 24599
rect 32861 24559 32919 24565
rect 1104 24506 34868 24528
rect 1104 24454 5170 24506
rect 5222 24454 5234 24506
rect 5286 24454 5298 24506
rect 5350 24454 5362 24506
rect 5414 24454 5426 24506
rect 5478 24454 13611 24506
rect 13663 24454 13675 24506
rect 13727 24454 13739 24506
rect 13791 24454 13803 24506
rect 13855 24454 13867 24506
rect 13919 24454 22052 24506
rect 22104 24454 22116 24506
rect 22168 24454 22180 24506
rect 22232 24454 22244 24506
rect 22296 24454 22308 24506
rect 22360 24454 30493 24506
rect 30545 24454 30557 24506
rect 30609 24454 30621 24506
rect 30673 24454 30685 24506
rect 30737 24454 30749 24506
rect 30801 24454 34868 24506
rect 1104 24432 34868 24454
rect 16761 24395 16819 24401
rect 16761 24361 16773 24395
rect 16807 24392 16819 24395
rect 16850 24392 16856 24404
rect 16807 24364 16856 24392
rect 16807 24361 16819 24364
rect 16761 24355 16819 24361
rect 16776 24324 16804 24355
rect 16850 24352 16856 24364
rect 16908 24352 16914 24404
rect 17218 24392 17224 24404
rect 17179 24364 17224 24392
rect 17218 24352 17224 24364
rect 17276 24352 17282 24404
rect 18414 24352 18420 24404
rect 18472 24392 18478 24404
rect 20070 24392 20076 24404
rect 18472 24364 18736 24392
rect 18472 24352 18478 24364
rect 15672 24296 16804 24324
rect 15565 24191 15623 24197
rect 15565 24157 15577 24191
rect 15611 24188 15623 24191
rect 15672 24188 15700 24296
rect 16022 24216 16028 24268
rect 16080 24256 16086 24268
rect 16301 24259 16359 24265
rect 16301 24256 16313 24259
rect 16080 24228 16313 24256
rect 16080 24216 16086 24228
rect 16301 24225 16313 24228
rect 16347 24225 16359 24259
rect 16758 24256 16764 24268
rect 16301 24219 16359 24225
rect 16439 24228 16764 24256
rect 15611 24160 15700 24188
rect 15611 24157 15623 24160
rect 15565 24151 15623 24157
rect 15746 24148 15752 24200
rect 15804 24188 15810 24200
rect 16439 24197 16467 24228
rect 16758 24216 16764 24228
rect 16816 24256 16822 24268
rect 16816 24228 18184 24256
rect 16816 24216 16822 24228
rect 16393 24191 16467 24197
rect 15804 24160 15849 24188
rect 15804 24148 15810 24160
rect 16393 24157 16405 24191
rect 16439 24157 16467 24191
rect 17405 24191 17463 24197
rect 17405 24157 17417 24191
rect 17451 24188 17463 24191
rect 17494 24188 17500 24200
rect 17451 24160 17500 24188
rect 17451 24157 17463 24160
rect 16393 24151 16451 24157
rect 17405 24151 17463 24157
rect 17494 24148 17500 24160
rect 17552 24148 17558 24200
rect 17681 24191 17739 24197
rect 17681 24157 17693 24191
rect 17727 24157 17739 24191
rect 17681 24151 17739 24157
rect 18156 24188 18184 24228
rect 18463 24191 18521 24197
rect 18463 24188 18475 24191
rect 18156 24160 18475 24188
rect 15657 24123 15715 24129
rect 15657 24089 15669 24123
rect 15703 24120 15715 24123
rect 17310 24120 17316 24132
rect 15703 24092 17316 24120
rect 15703 24089 15715 24092
rect 15657 24083 15715 24089
rect 17310 24080 17316 24092
rect 17368 24120 17374 24132
rect 17696 24120 17724 24151
rect 17368 24092 17724 24120
rect 17368 24080 17374 24092
rect 16666 24012 16672 24064
rect 16724 24052 16730 24064
rect 17402 24052 17408 24064
rect 16724 24024 17408 24052
rect 16724 24012 16730 24024
rect 17402 24012 17408 24024
rect 17460 24052 17466 24064
rect 17589 24055 17647 24061
rect 17589 24052 17601 24055
rect 17460 24024 17601 24052
rect 17460 24012 17466 24024
rect 17589 24021 17601 24024
rect 17635 24021 17647 24055
rect 18156 24052 18184 24160
rect 18463 24157 18475 24160
rect 18509 24157 18521 24191
rect 18598 24188 18604 24200
rect 18559 24160 18604 24188
rect 18463 24151 18521 24157
rect 18598 24148 18604 24160
rect 18656 24148 18662 24200
rect 18708 24197 18736 24364
rect 18892 24364 20076 24392
rect 18892 24200 18920 24364
rect 20070 24352 20076 24364
rect 20128 24352 20134 24404
rect 20990 24352 20996 24404
rect 21048 24392 21054 24404
rect 22005 24395 22063 24401
rect 22005 24392 22017 24395
rect 21048 24364 22017 24392
rect 21048 24352 21054 24364
rect 22005 24361 22017 24364
rect 22051 24392 22063 24395
rect 22370 24392 22376 24404
rect 22051 24364 22376 24392
rect 22051 24361 22063 24364
rect 22005 24355 22063 24361
rect 22370 24352 22376 24364
rect 22428 24352 22434 24404
rect 22462 24352 22468 24404
rect 22520 24392 22526 24404
rect 22922 24392 22928 24404
rect 22520 24364 22784 24392
rect 22883 24364 22928 24392
rect 22520 24352 22526 24364
rect 22756 24324 22784 24364
rect 22922 24352 22928 24364
rect 22980 24352 22986 24404
rect 23106 24392 23112 24404
rect 23067 24364 23112 24392
rect 23106 24352 23112 24364
rect 23164 24352 23170 24404
rect 23937 24395 23995 24401
rect 23937 24361 23949 24395
rect 23983 24392 23995 24395
rect 24026 24392 24032 24404
rect 23983 24364 24032 24392
rect 23983 24361 23995 24364
rect 23937 24355 23995 24361
rect 24026 24352 24032 24364
rect 24084 24352 24090 24404
rect 26970 24352 26976 24404
rect 27028 24392 27034 24404
rect 27430 24392 27436 24404
rect 27028 24364 27436 24392
rect 27028 24352 27034 24364
rect 27430 24352 27436 24364
rect 27488 24392 27494 24404
rect 30101 24395 30159 24401
rect 30101 24392 30113 24395
rect 27488 24364 30113 24392
rect 27488 24352 27494 24364
rect 30101 24361 30113 24364
rect 30147 24361 30159 24395
rect 30101 24355 30159 24361
rect 30929 24395 30987 24401
rect 30929 24361 30941 24395
rect 30975 24392 30987 24395
rect 31386 24392 31392 24404
rect 30975 24364 31392 24392
rect 30975 24361 30987 24364
rect 30929 24355 30987 24361
rect 31386 24352 31392 24364
rect 31444 24352 31450 24404
rect 31573 24395 31631 24401
rect 31573 24361 31585 24395
rect 31619 24392 31631 24395
rect 33042 24392 33048 24404
rect 31619 24364 33048 24392
rect 31619 24361 31631 24364
rect 31573 24355 31631 24361
rect 33042 24352 33048 24364
rect 33100 24352 33106 24404
rect 22756 24296 22961 24324
rect 21174 24216 21180 24268
rect 21232 24256 21238 24268
rect 22462 24256 22468 24268
rect 21232 24228 22468 24256
rect 21232 24216 21238 24228
rect 22462 24216 22468 24228
rect 22520 24216 22526 24268
rect 18708 24191 18772 24197
rect 18708 24160 18726 24191
rect 18714 24157 18726 24160
rect 18760 24157 18772 24191
rect 18714 24151 18772 24157
rect 18874 24148 18880 24200
rect 18932 24188 18938 24200
rect 18932 24160 19025 24188
rect 18932 24148 18938 24160
rect 19058 24148 19064 24200
rect 19116 24188 19122 24200
rect 19429 24191 19487 24197
rect 19429 24188 19441 24191
rect 19116 24160 19441 24188
rect 19116 24148 19122 24160
rect 19429 24157 19441 24160
rect 19475 24188 19487 24191
rect 21726 24188 21732 24200
rect 19475 24160 21732 24188
rect 19475 24157 19487 24160
rect 19429 24151 19487 24157
rect 21726 24148 21732 24160
rect 21784 24148 21790 24200
rect 22278 24188 22284 24200
rect 21836 24160 22284 24188
rect 21836 24129 21864 24160
rect 22278 24148 22284 24160
rect 22336 24148 22342 24200
rect 22933 24197 22961 24296
rect 24394 24284 24400 24336
rect 24452 24324 24458 24336
rect 32398 24324 32404 24336
rect 24452 24296 32404 24324
rect 24452 24284 24458 24296
rect 32398 24284 32404 24296
rect 32456 24284 32462 24336
rect 23106 24216 23112 24268
rect 23164 24256 23170 24268
rect 23569 24259 23627 24265
rect 23569 24256 23581 24259
rect 23164 24228 23581 24256
rect 23164 24216 23170 24228
rect 23569 24225 23581 24228
rect 23615 24225 23627 24259
rect 24946 24256 24952 24268
rect 24907 24228 24952 24256
rect 23569 24219 23627 24225
rect 24946 24216 24952 24228
rect 25004 24216 25010 24268
rect 27062 24256 27068 24268
rect 25056 24228 26096 24256
rect 27023 24228 27068 24256
rect 25056 24200 25084 24228
rect 22833 24191 22891 24197
rect 22833 24157 22845 24191
rect 22879 24157 22891 24191
rect 22833 24151 22891 24157
rect 22925 24191 22983 24197
rect 22925 24157 22937 24191
rect 22971 24157 22983 24191
rect 22925 24151 22983 24157
rect 23753 24191 23811 24197
rect 23753 24157 23765 24191
rect 23799 24157 23811 24191
rect 23753 24151 23811 24157
rect 24857 24191 24915 24197
rect 24857 24157 24869 24191
rect 24903 24188 24915 24191
rect 25038 24188 25044 24200
rect 24903 24160 25044 24188
rect 24903 24157 24915 24160
rect 24857 24151 24915 24157
rect 18233 24123 18291 24129
rect 18233 24089 18245 24123
rect 18279 24120 18291 24123
rect 19674 24123 19732 24129
rect 19674 24120 19686 24123
rect 18279 24092 19686 24120
rect 18279 24089 18291 24092
rect 18233 24083 18291 24089
rect 19674 24089 19686 24092
rect 19720 24089 19732 24123
rect 19674 24083 19732 24089
rect 21821 24123 21879 24129
rect 21821 24089 21833 24123
rect 21867 24089 21879 24123
rect 21821 24083 21879 24089
rect 22037 24123 22095 24129
rect 22037 24089 22049 24123
rect 22083 24120 22095 24123
rect 22554 24120 22560 24132
rect 22083 24092 22560 24120
rect 22083 24089 22095 24092
rect 22037 24083 22095 24089
rect 22554 24080 22560 24092
rect 22612 24080 22618 24132
rect 22646 24080 22652 24132
rect 22704 24120 22710 24132
rect 22848 24120 22876 24151
rect 23198 24120 23204 24132
rect 22704 24092 22749 24120
rect 22848 24092 23204 24120
rect 22704 24080 22710 24092
rect 23198 24080 23204 24092
rect 23256 24080 23262 24132
rect 20809 24055 20867 24061
rect 20809 24052 20821 24055
rect 18156 24024 20821 24052
rect 17589 24015 17647 24021
rect 20809 24021 20821 24024
rect 20855 24052 20867 24055
rect 21174 24052 21180 24064
rect 20855 24024 21180 24052
rect 20855 24021 20867 24024
rect 20809 24015 20867 24021
rect 21174 24012 21180 24024
rect 21232 24012 21238 24064
rect 22186 24052 22192 24064
rect 22147 24024 22192 24052
rect 22186 24012 22192 24024
rect 22244 24012 22250 24064
rect 22278 24012 22284 24064
rect 22336 24052 22342 24064
rect 22738 24052 22744 24064
rect 22336 24024 22744 24052
rect 22336 24012 22342 24024
rect 22738 24012 22744 24024
rect 22796 24052 22802 24064
rect 23768 24052 23796 24151
rect 25038 24148 25044 24160
rect 25096 24148 25102 24200
rect 25869 24191 25927 24197
rect 25869 24157 25881 24191
rect 25915 24188 25927 24191
rect 25958 24188 25964 24200
rect 25915 24160 25964 24188
rect 25915 24157 25927 24160
rect 25869 24151 25927 24157
rect 25958 24148 25964 24160
rect 26016 24148 26022 24200
rect 26068 24197 26096 24228
rect 27062 24216 27068 24228
rect 27120 24216 27126 24268
rect 27341 24259 27399 24265
rect 27341 24225 27353 24259
rect 27387 24256 27399 24259
rect 28442 24256 28448 24268
rect 27387 24228 28448 24256
rect 27387 24225 27399 24228
rect 27341 24219 27399 24225
rect 28442 24216 28448 24228
rect 28500 24216 28506 24268
rect 28537 24259 28595 24265
rect 28537 24225 28549 24259
rect 28583 24256 28595 24259
rect 28718 24256 28724 24268
rect 28583 24228 28724 24256
rect 28583 24225 28595 24228
rect 28537 24219 28595 24225
rect 28718 24216 28724 24228
rect 28776 24256 28782 24268
rect 29546 24256 29552 24268
rect 28776 24228 29552 24256
rect 28776 24216 28782 24228
rect 29546 24216 29552 24228
rect 29604 24216 29610 24268
rect 30193 24259 30251 24265
rect 30193 24225 30205 24259
rect 30239 24256 30251 24259
rect 30926 24256 30932 24268
rect 30239 24228 30932 24256
rect 30239 24225 30251 24228
rect 30193 24219 30251 24225
rect 30926 24216 30932 24228
rect 30984 24216 30990 24268
rect 31018 24216 31024 24268
rect 31076 24256 31082 24268
rect 34146 24256 34152 24268
rect 31076 24228 34152 24256
rect 31076 24216 31082 24228
rect 34146 24216 34152 24228
rect 34204 24216 34210 24268
rect 26053 24191 26111 24197
rect 26053 24157 26065 24191
rect 26099 24157 26111 24191
rect 26053 24151 26111 24157
rect 26145 24191 26203 24197
rect 26145 24157 26157 24191
rect 26191 24188 26203 24191
rect 26878 24188 26884 24200
rect 26191 24160 26884 24188
rect 26191 24157 26203 24160
rect 26145 24151 26203 24157
rect 26878 24148 26884 24160
rect 26936 24148 26942 24200
rect 26970 24148 26976 24200
rect 27028 24188 27034 24200
rect 28350 24188 28356 24200
rect 27028 24160 27073 24188
rect 28311 24160 28356 24188
rect 27028 24148 27034 24160
rect 28350 24148 28356 24160
rect 28408 24148 28414 24200
rect 28629 24191 28687 24197
rect 28629 24157 28641 24191
rect 28675 24188 28687 24191
rect 29733 24191 29791 24197
rect 29733 24188 29745 24191
rect 28675 24160 29745 24188
rect 28675 24157 28687 24160
rect 28629 24151 28687 24157
rect 29733 24157 29745 24160
rect 29779 24157 29791 24191
rect 29733 24151 29791 24157
rect 29917 24191 29975 24197
rect 29917 24157 29929 24191
rect 29963 24188 29975 24191
rect 30282 24188 30288 24200
rect 29963 24160 30288 24188
rect 29963 24157 29975 24160
rect 29917 24151 29975 24157
rect 30282 24148 30288 24160
rect 30340 24148 30346 24200
rect 30650 24188 30656 24200
rect 30611 24160 30656 24188
rect 30650 24148 30656 24160
rect 30708 24148 30714 24200
rect 31110 24148 31116 24200
rect 31168 24148 31174 24200
rect 31757 24191 31815 24197
rect 31757 24157 31769 24191
rect 31803 24188 31815 24191
rect 31846 24188 31852 24200
rect 31803 24160 31852 24188
rect 31803 24157 31815 24160
rect 31757 24151 31815 24157
rect 31846 24148 31852 24160
rect 31904 24148 31910 24200
rect 32030 24188 32036 24200
rect 31991 24160 32036 24188
rect 32030 24148 32036 24160
rect 32088 24148 32094 24200
rect 32490 24188 32496 24200
rect 32451 24160 32496 24188
rect 32490 24148 32496 24160
rect 32548 24148 32554 24200
rect 26694 24120 26700 24132
rect 25240 24092 26700 24120
rect 25240 24061 25268 24092
rect 26694 24080 26700 24092
rect 26752 24080 26758 24132
rect 28718 24120 28724 24132
rect 27586 24092 28724 24120
rect 22796 24024 23796 24052
rect 25225 24055 25283 24061
rect 22796 24012 22802 24024
rect 25225 24021 25237 24055
rect 25271 24021 25283 24055
rect 25225 24015 25283 24021
rect 25685 24055 25743 24061
rect 25685 24021 25697 24055
rect 25731 24052 25743 24055
rect 27586 24052 27614 24092
rect 28718 24080 28724 24092
rect 28776 24080 28782 24132
rect 31128 24120 31156 24148
rect 31941 24123 31999 24129
rect 31941 24120 31953 24123
rect 31128 24092 31953 24120
rect 31941 24089 31953 24092
rect 31987 24089 31999 24123
rect 32674 24120 32680 24132
rect 32635 24092 32680 24120
rect 31941 24083 31999 24089
rect 32674 24080 32680 24092
rect 32732 24080 32738 24132
rect 34330 24120 34336 24132
rect 34291 24092 34336 24120
rect 34330 24080 34336 24092
rect 34388 24080 34394 24132
rect 28166 24052 28172 24064
rect 25731 24024 27614 24052
rect 28127 24024 28172 24052
rect 25731 24021 25743 24024
rect 25685 24015 25743 24021
rect 28166 24012 28172 24024
rect 28224 24012 28230 24064
rect 28442 24012 28448 24064
rect 28500 24052 28506 24064
rect 30190 24052 30196 24064
rect 28500 24024 30196 24052
rect 28500 24012 28506 24024
rect 30190 24012 30196 24024
rect 30248 24012 30254 24064
rect 31113 24055 31171 24061
rect 31113 24021 31125 24055
rect 31159 24052 31171 24055
rect 31846 24052 31852 24064
rect 31159 24024 31852 24052
rect 31159 24021 31171 24024
rect 31113 24015 31171 24021
rect 31846 24012 31852 24024
rect 31904 24052 31910 24064
rect 32214 24052 32220 24064
rect 31904 24024 32220 24052
rect 31904 24012 31910 24024
rect 32214 24012 32220 24024
rect 32272 24012 32278 24064
rect 1104 23962 35027 23984
rect 1104 23910 9390 23962
rect 9442 23910 9454 23962
rect 9506 23910 9518 23962
rect 9570 23910 9582 23962
rect 9634 23910 9646 23962
rect 9698 23910 17831 23962
rect 17883 23910 17895 23962
rect 17947 23910 17959 23962
rect 18011 23910 18023 23962
rect 18075 23910 18087 23962
rect 18139 23910 26272 23962
rect 26324 23910 26336 23962
rect 26388 23910 26400 23962
rect 26452 23910 26464 23962
rect 26516 23910 26528 23962
rect 26580 23910 34713 23962
rect 34765 23910 34777 23962
rect 34829 23910 34841 23962
rect 34893 23910 34905 23962
rect 34957 23910 34969 23962
rect 35021 23910 35027 23962
rect 1104 23888 35027 23910
rect 8938 23808 8944 23860
rect 8996 23848 9002 23860
rect 22186 23848 22192 23860
rect 8996 23820 22192 23848
rect 8996 23808 9002 23820
rect 22186 23808 22192 23820
rect 22244 23808 22250 23860
rect 22370 23808 22376 23860
rect 22428 23848 22434 23860
rect 22465 23851 22523 23857
rect 22465 23848 22477 23851
rect 22428 23820 22477 23848
rect 22428 23808 22434 23820
rect 22465 23817 22477 23820
rect 22511 23817 22523 23851
rect 22465 23811 22523 23817
rect 22646 23808 22652 23860
rect 22704 23848 22710 23860
rect 23290 23848 23296 23860
rect 22704 23820 23296 23848
rect 22704 23808 22710 23820
rect 23290 23808 23296 23820
rect 23348 23848 23354 23860
rect 23842 23848 23848 23860
rect 23348 23820 23848 23848
rect 23348 23808 23354 23820
rect 23842 23808 23848 23820
rect 23900 23808 23906 23860
rect 27614 23808 27620 23860
rect 27672 23848 27678 23860
rect 29730 23848 29736 23860
rect 27672 23820 29736 23848
rect 27672 23808 27678 23820
rect 29730 23808 29736 23820
rect 29788 23808 29794 23860
rect 31754 23808 31760 23860
rect 31812 23848 31818 23860
rect 32398 23848 32404 23860
rect 31812 23820 32404 23848
rect 31812 23808 31818 23820
rect 32398 23808 32404 23820
rect 32456 23808 32462 23860
rect 17494 23780 17500 23792
rect 17052 23752 17500 23780
rect 17052 23721 17080 23752
rect 17494 23740 17500 23752
rect 17552 23740 17558 23792
rect 17678 23740 17684 23792
rect 17736 23780 17742 23792
rect 18601 23783 18659 23789
rect 17736 23752 18092 23780
rect 17736 23740 17742 23752
rect 15933 23715 15991 23721
rect 15933 23681 15945 23715
rect 15979 23712 15991 23715
rect 17037 23715 17095 23721
rect 17037 23712 17049 23715
rect 15979 23684 16252 23712
rect 15979 23681 15991 23684
rect 15933 23675 15991 23681
rect 16022 23644 16028 23656
rect 15983 23616 16028 23644
rect 16022 23604 16028 23616
rect 16080 23604 16086 23656
rect 16224 23576 16252 23684
rect 16316 23684 17049 23712
rect 16316 23653 16344 23684
rect 17037 23681 17049 23684
rect 17083 23681 17095 23715
rect 17218 23712 17224 23724
rect 17179 23684 17224 23712
rect 17037 23675 17095 23681
rect 17218 23672 17224 23684
rect 17276 23672 17282 23724
rect 17865 23715 17923 23721
rect 17865 23681 17877 23715
rect 17911 23712 17923 23715
rect 17954 23712 17960 23724
rect 17911 23684 17960 23712
rect 17911 23681 17923 23684
rect 17865 23675 17923 23681
rect 17954 23672 17960 23684
rect 18012 23672 18018 23724
rect 18064 23721 18092 23752
rect 18601 23749 18613 23783
rect 18647 23780 18659 23783
rect 19306 23783 19364 23789
rect 19306 23780 19318 23783
rect 18647 23752 19318 23780
rect 18647 23749 18659 23752
rect 18601 23743 18659 23749
rect 19306 23749 19318 23752
rect 19352 23749 19364 23783
rect 22278 23780 22284 23792
rect 19306 23743 19364 23749
rect 21284 23752 22284 23780
rect 18049 23715 18107 23721
rect 18049 23681 18061 23715
rect 18095 23681 18107 23715
rect 18049 23675 18107 23681
rect 18141 23715 18199 23721
rect 18141 23681 18153 23715
rect 18187 23712 18199 23715
rect 18322 23712 18328 23724
rect 18187 23684 18328 23712
rect 18187 23681 18199 23684
rect 18141 23675 18199 23681
rect 18322 23672 18328 23684
rect 18380 23672 18386 23724
rect 18417 23715 18475 23721
rect 18417 23681 18429 23715
rect 18463 23712 18475 23715
rect 19058 23712 19064 23724
rect 18463 23684 18920 23712
rect 19019 23684 19064 23712
rect 18463 23681 18475 23684
rect 18417 23675 18475 23681
rect 16301 23647 16359 23653
rect 16301 23613 16313 23647
rect 16347 23613 16359 23647
rect 16301 23607 16359 23613
rect 16850 23604 16856 23656
rect 16908 23644 16914 23656
rect 17129 23647 17187 23653
rect 17129 23644 17141 23647
rect 16908 23616 17141 23644
rect 16908 23604 16914 23616
rect 17129 23613 17141 23616
rect 17175 23613 17187 23647
rect 17129 23607 17187 23613
rect 17310 23604 17316 23656
rect 17368 23644 17374 23656
rect 18233 23647 18291 23653
rect 17368 23616 17413 23644
rect 17368 23604 17374 23616
rect 18233 23613 18245 23647
rect 18279 23644 18291 23647
rect 18598 23644 18604 23656
rect 18279 23616 18604 23644
rect 18279 23613 18291 23616
rect 18233 23607 18291 23613
rect 18598 23604 18604 23616
rect 18656 23604 18662 23656
rect 17494 23576 17500 23588
rect 16224 23548 17500 23576
rect 17494 23536 17500 23548
rect 17552 23576 17558 23588
rect 18892 23576 18920 23684
rect 19058 23672 19064 23684
rect 19116 23672 19122 23724
rect 21284 23721 21312 23752
rect 22278 23740 22284 23752
rect 22336 23740 22342 23792
rect 23382 23780 23388 23792
rect 22388 23752 23388 23780
rect 21269 23715 21327 23721
rect 21269 23681 21281 23715
rect 21315 23681 21327 23715
rect 21269 23675 21327 23681
rect 22005 23715 22063 23721
rect 22005 23681 22017 23715
rect 22051 23712 22063 23715
rect 22388 23712 22416 23752
rect 23382 23740 23388 23752
rect 23440 23740 23446 23792
rect 24302 23780 24308 23792
rect 23584 23752 24308 23780
rect 22051 23684 22416 23712
rect 22051 23681 22063 23684
rect 22005 23675 22063 23681
rect 22462 23672 22468 23724
rect 22520 23712 22526 23724
rect 23584 23721 23612 23752
rect 24302 23740 24308 23752
rect 24360 23740 24366 23792
rect 26878 23780 26884 23792
rect 25700 23752 26884 23780
rect 25700 23724 25728 23752
rect 26878 23740 26884 23752
rect 26936 23740 26942 23792
rect 28534 23740 28540 23792
rect 28592 23780 28598 23792
rect 28629 23783 28687 23789
rect 28629 23780 28641 23783
rect 28592 23752 28641 23780
rect 28592 23740 28598 23752
rect 28629 23749 28641 23752
rect 28675 23749 28687 23783
rect 29748 23780 29776 23808
rect 34333 23783 34391 23789
rect 29748 23752 31754 23780
rect 28629 23743 28687 23749
rect 22925 23715 22983 23721
rect 22925 23712 22937 23715
rect 22520 23684 22937 23712
rect 22520 23672 22526 23684
rect 22925 23681 22937 23684
rect 22971 23681 22983 23715
rect 22925 23675 22983 23681
rect 23109 23715 23167 23721
rect 23109 23681 23121 23715
rect 23155 23681 23167 23715
rect 23109 23675 23167 23681
rect 23569 23715 23627 23721
rect 23569 23681 23581 23715
rect 23615 23681 23627 23715
rect 23569 23675 23627 23681
rect 23836 23715 23894 23721
rect 23836 23681 23848 23715
rect 23882 23712 23894 23715
rect 24394 23712 24400 23724
rect 23882 23684 24400 23712
rect 23882 23681 23894 23684
rect 23836 23675 23894 23681
rect 21085 23647 21143 23653
rect 21085 23613 21097 23647
rect 21131 23644 21143 23647
rect 22646 23644 22652 23656
rect 21131 23616 22652 23644
rect 21131 23613 21143 23616
rect 21085 23607 21143 23613
rect 22646 23604 22652 23616
rect 22704 23604 22710 23656
rect 17552 23548 18920 23576
rect 17552 23536 17558 23548
rect 16114 23468 16120 23520
rect 16172 23508 16178 23520
rect 16853 23511 16911 23517
rect 16853 23508 16865 23511
rect 16172 23480 16865 23508
rect 16172 23468 16178 23480
rect 16853 23477 16865 23480
rect 16899 23477 16911 23511
rect 18892 23508 18920 23548
rect 20714 23536 20720 23588
rect 20772 23576 20778 23588
rect 21453 23579 21511 23585
rect 21453 23576 21465 23579
rect 20772 23548 21465 23576
rect 20772 23536 20778 23548
rect 21453 23545 21465 23548
rect 21499 23545 21511 23579
rect 23124 23576 23152 23675
rect 24394 23672 24400 23684
rect 24452 23672 24458 23724
rect 25682 23712 25688 23724
rect 25643 23684 25688 23712
rect 25682 23672 25688 23684
rect 25740 23672 25746 23724
rect 25777 23715 25835 23721
rect 25777 23681 25789 23715
rect 25823 23681 25835 23715
rect 25777 23675 25835 23681
rect 25869 23715 25927 23721
rect 25869 23681 25881 23715
rect 25915 23681 25927 23715
rect 25869 23675 25927 23681
rect 21453 23539 21511 23545
rect 21551 23548 23152 23576
rect 25792 23576 25820 23675
rect 25884 23644 25912 23675
rect 25958 23672 25964 23724
rect 26016 23712 26022 23724
rect 26053 23715 26111 23721
rect 26053 23712 26065 23715
rect 26016 23684 26065 23712
rect 26016 23672 26022 23684
rect 26053 23681 26065 23684
rect 26099 23681 26111 23715
rect 26053 23675 26111 23681
rect 26970 23672 26976 23724
rect 27028 23712 27034 23724
rect 27341 23715 27399 23721
rect 27341 23712 27353 23715
rect 27028 23684 27353 23712
rect 27028 23672 27034 23684
rect 27341 23681 27353 23684
rect 27387 23712 27399 23715
rect 28994 23712 29000 23724
rect 27387 23684 29000 23712
rect 27387 23681 27399 23684
rect 27341 23675 27399 23681
rect 28994 23672 29000 23684
rect 29052 23672 29058 23724
rect 31021 23715 31079 23721
rect 31021 23681 31033 23715
rect 31067 23712 31079 23715
rect 31478 23712 31484 23724
rect 31067 23684 31484 23712
rect 31067 23681 31079 23684
rect 31021 23675 31079 23681
rect 31478 23672 31484 23684
rect 31536 23672 31542 23724
rect 26602 23644 26608 23656
rect 25884 23616 26608 23644
rect 26602 23604 26608 23616
rect 26660 23604 26666 23656
rect 27062 23604 27068 23656
rect 27120 23644 27126 23656
rect 27249 23647 27307 23653
rect 27249 23644 27261 23647
rect 27120 23616 27261 23644
rect 27120 23604 27126 23616
rect 27249 23613 27261 23616
rect 27295 23613 27307 23647
rect 27249 23607 27307 23613
rect 28442 23604 28448 23656
rect 28500 23644 28506 23656
rect 28810 23644 28816 23656
rect 28500 23616 28816 23644
rect 28500 23604 28506 23616
rect 28810 23604 28816 23616
rect 28868 23604 28874 23656
rect 29086 23604 29092 23656
rect 29144 23644 29150 23656
rect 30098 23644 30104 23656
rect 29144 23616 30104 23644
rect 29144 23604 29150 23616
rect 30098 23604 30104 23616
rect 30156 23644 30162 23656
rect 30377 23647 30435 23653
rect 30377 23644 30389 23647
rect 30156 23616 30389 23644
rect 30156 23604 30162 23616
rect 30377 23613 30389 23616
rect 30423 23613 30435 23647
rect 30377 23607 30435 23613
rect 27522 23576 27528 23588
rect 25792 23548 27528 23576
rect 20254 23508 20260 23520
rect 18892 23480 20260 23508
rect 16853 23471 16911 23477
rect 20254 23468 20260 23480
rect 20312 23508 20318 23520
rect 20441 23511 20499 23517
rect 20441 23508 20453 23511
rect 20312 23480 20453 23508
rect 20312 23468 20318 23480
rect 20441 23477 20453 23480
rect 20487 23477 20499 23511
rect 20441 23471 20499 23477
rect 20530 23468 20536 23520
rect 20588 23508 20594 23520
rect 21551 23508 21579 23548
rect 27522 23536 27528 23548
rect 27580 23536 27586 23588
rect 28626 23536 28632 23588
rect 28684 23576 28690 23588
rect 30282 23576 30288 23588
rect 28684 23548 30288 23576
rect 28684 23536 28690 23548
rect 30282 23536 30288 23548
rect 30340 23536 30346 23588
rect 30392 23576 30420 23607
rect 30650 23604 30656 23656
rect 30708 23644 30714 23656
rect 31297 23647 31355 23653
rect 31297 23644 31309 23647
rect 30708 23616 31309 23644
rect 30708 23604 30714 23616
rect 31297 23613 31309 23616
rect 31343 23644 31355 23647
rect 31386 23644 31392 23656
rect 31343 23616 31392 23644
rect 31343 23613 31355 23616
rect 31297 23607 31355 23613
rect 31386 23604 31392 23616
rect 31444 23604 31450 23656
rect 31726 23576 31754 23752
rect 34333 23749 34345 23783
rect 34379 23780 34391 23783
rect 34422 23780 34428 23792
rect 34379 23752 34428 23780
rect 34379 23749 34391 23752
rect 34333 23743 34391 23749
rect 34422 23740 34428 23752
rect 34480 23740 34486 23792
rect 32490 23644 32496 23656
rect 32451 23616 32496 23644
rect 32490 23604 32496 23616
rect 32548 23604 32554 23656
rect 32674 23644 32680 23656
rect 32635 23616 32680 23644
rect 32674 23604 32680 23616
rect 32732 23604 32738 23656
rect 32030 23576 32036 23588
rect 30392 23548 31340 23576
rect 31726 23548 32036 23576
rect 20588 23480 21579 23508
rect 22281 23511 22339 23517
rect 20588 23468 20594 23480
rect 22281 23477 22293 23511
rect 22327 23508 22339 23511
rect 22370 23508 22376 23520
rect 22327 23480 22376 23508
rect 22327 23477 22339 23480
rect 22281 23471 22339 23477
rect 22370 23468 22376 23480
rect 22428 23468 22434 23520
rect 23014 23508 23020 23520
rect 22975 23480 23020 23508
rect 23014 23468 23020 23480
rect 23072 23468 23078 23520
rect 24949 23511 25007 23517
rect 24949 23477 24961 23511
rect 24995 23508 25007 23511
rect 25038 23508 25044 23520
rect 24995 23480 25044 23508
rect 24995 23477 25007 23480
rect 24949 23471 25007 23477
rect 25038 23468 25044 23480
rect 25096 23468 25102 23520
rect 25406 23508 25412 23520
rect 25367 23480 25412 23508
rect 25406 23468 25412 23480
rect 25464 23468 25470 23520
rect 27709 23511 27767 23517
rect 27709 23477 27721 23511
rect 27755 23508 27767 23511
rect 28350 23508 28356 23520
rect 27755 23480 28356 23508
rect 27755 23477 27767 23480
rect 27709 23471 27767 23477
rect 28350 23468 28356 23480
rect 28408 23508 28414 23520
rect 28902 23508 28908 23520
rect 28408 23480 28908 23508
rect 28408 23468 28414 23480
rect 28902 23468 28908 23480
rect 28960 23468 28966 23520
rect 30834 23508 30840 23520
rect 30795 23480 30840 23508
rect 30834 23468 30840 23480
rect 30892 23468 30898 23520
rect 30926 23468 30932 23520
rect 30984 23508 30990 23520
rect 31205 23511 31263 23517
rect 31205 23508 31217 23511
rect 30984 23480 31217 23508
rect 30984 23468 30990 23480
rect 31205 23477 31217 23480
rect 31251 23477 31263 23511
rect 31312 23508 31340 23548
rect 32030 23536 32036 23548
rect 32088 23576 32094 23588
rect 32858 23576 32864 23588
rect 32088 23548 32864 23576
rect 32088 23536 32094 23548
rect 32858 23536 32864 23548
rect 32916 23536 32922 23588
rect 32306 23508 32312 23520
rect 31312 23480 32312 23508
rect 31205 23471 31263 23477
rect 32306 23468 32312 23480
rect 32364 23468 32370 23520
rect 1104 23418 34868 23440
rect 1104 23366 5170 23418
rect 5222 23366 5234 23418
rect 5286 23366 5298 23418
rect 5350 23366 5362 23418
rect 5414 23366 5426 23418
rect 5478 23366 13611 23418
rect 13663 23366 13675 23418
rect 13727 23366 13739 23418
rect 13791 23366 13803 23418
rect 13855 23366 13867 23418
rect 13919 23366 22052 23418
rect 22104 23366 22116 23418
rect 22168 23366 22180 23418
rect 22232 23366 22244 23418
rect 22296 23366 22308 23418
rect 22360 23366 30493 23418
rect 30545 23366 30557 23418
rect 30609 23366 30621 23418
rect 30673 23366 30685 23418
rect 30737 23366 30749 23418
rect 30801 23366 34868 23418
rect 1104 23344 34868 23366
rect 16666 23304 16672 23316
rect 16627 23276 16672 23304
rect 16666 23264 16672 23276
rect 16724 23264 16730 23316
rect 17865 23307 17923 23313
rect 17865 23273 17877 23307
rect 17911 23304 17923 23307
rect 18414 23304 18420 23316
rect 17911 23276 18420 23304
rect 17911 23273 17923 23276
rect 17865 23267 17923 23273
rect 18414 23264 18420 23276
rect 18472 23264 18478 23316
rect 18690 23264 18696 23316
rect 18748 23304 18754 23316
rect 19797 23307 19855 23313
rect 19797 23304 19809 23307
rect 18748 23276 19809 23304
rect 18748 23264 18754 23276
rect 19797 23273 19809 23276
rect 19843 23273 19855 23307
rect 19797 23267 19855 23273
rect 21910 23264 21916 23316
rect 21968 23304 21974 23316
rect 22097 23307 22155 23313
rect 22097 23304 22109 23307
rect 21968 23276 22109 23304
rect 21968 23264 21974 23276
rect 22097 23273 22109 23276
rect 22143 23273 22155 23307
rect 28258 23304 28264 23316
rect 22097 23267 22155 23273
rect 25148 23276 28264 23304
rect 18601 23239 18659 23245
rect 18601 23205 18613 23239
rect 18647 23205 18659 23239
rect 18601 23199 18659 23205
rect 17586 23168 17592 23180
rect 17547 23140 17592 23168
rect 17586 23128 17592 23140
rect 17644 23128 17650 23180
rect 18616 23168 18644 23199
rect 18782 23196 18788 23248
rect 18840 23236 18846 23248
rect 18840 23208 19717 23236
rect 18840 23196 18846 23208
rect 19689 23180 19717 23208
rect 22370 23196 22376 23248
rect 22428 23236 22434 23248
rect 22554 23236 22560 23248
rect 22428 23208 22560 23236
rect 22428 23196 22434 23208
rect 22554 23196 22560 23208
rect 22612 23196 22618 23248
rect 18616 23140 19656 23168
rect 19689 23140 19708 23180
rect 16574 23100 16580 23112
rect 16535 23072 16580 23100
rect 16574 23060 16580 23072
rect 16632 23060 16638 23112
rect 16758 23100 16764 23112
rect 16719 23072 16764 23100
rect 16758 23060 16764 23072
rect 16816 23060 16822 23112
rect 17402 23060 17408 23112
rect 17460 23100 17466 23112
rect 19628 23109 19656 23140
rect 19702 23128 19708 23140
rect 19760 23168 19766 23180
rect 19889 23171 19947 23177
rect 19889 23168 19901 23171
rect 19760 23140 19901 23168
rect 19760 23128 19766 23140
rect 19889 23137 19901 23140
rect 19935 23137 19947 23171
rect 19889 23131 19947 23137
rect 20070 23128 20076 23180
rect 20128 23168 20134 23180
rect 25148 23168 25176 23276
rect 28258 23264 28264 23276
rect 28316 23264 28322 23316
rect 29086 23304 29092 23316
rect 28368 23276 29092 23304
rect 26878 23236 26884 23248
rect 26839 23208 26884 23236
rect 26878 23196 26884 23208
rect 26936 23196 26942 23248
rect 20128 23140 25176 23168
rect 20128 23128 20134 23140
rect 17681 23103 17739 23109
rect 17681 23100 17693 23103
rect 17460 23072 17693 23100
rect 17460 23060 17466 23072
rect 17681 23069 17693 23072
rect 17727 23069 17739 23103
rect 18877 23103 18935 23109
rect 18877 23100 18889 23103
rect 17681 23063 17739 23069
rect 18248 23072 18889 23100
rect 18248 23044 18276 23072
rect 18877 23069 18889 23072
rect 18923 23069 18935 23103
rect 18877 23063 18935 23069
rect 19613 23103 19671 23109
rect 19613 23069 19625 23103
rect 19659 23069 19671 23103
rect 19978 23100 19984 23112
rect 19891 23072 19984 23100
rect 19613 23063 19671 23069
rect 17221 23035 17279 23041
rect 17221 23001 17233 23035
rect 17267 23032 17279 23035
rect 18230 23032 18236 23044
rect 17267 23004 18236 23032
rect 17267 23001 17279 23004
rect 17221 22995 17279 23001
rect 18230 22992 18236 23004
rect 18288 22992 18294 23044
rect 18601 23035 18659 23041
rect 18601 23001 18613 23035
rect 18647 23032 18659 23035
rect 19904 23032 19932 23072
rect 19978 23060 19984 23072
rect 20036 23100 20042 23112
rect 20438 23100 20444 23112
rect 20036 23072 20444 23100
rect 20036 23060 20042 23072
rect 20438 23060 20444 23072
rect 20496 23060 20502 23112
rect 20806 23100 20812 23112
rect 20767 23072 20812 23100
rect 20806 23060 20812 23072
rect 20864 23060 20870 23112
rect 23198 23100 23204 23112
rect 23159 23072 23204 23100
rect 23198 23060 23204 23072
rect 23256 23060 23262 23112
rect 23474 23100 23480 23112
rect 23435 23072 23480 23100
rect 23474 23060 23480 23072
rect 23532 23060 23538 23112
rect 24765 23103 24823 23109
rect 24765 23069 24777 23103
rect 24811 23069 24823 23103
rect 24946 23100 24952 23112
rect 24907 23072 24952 23100
rect 24765 23063 24823 23069
rect 18647 23004 19932 23032
rect 18647 23001 18659 23004
rect 18601 22995 18659 23001
rect 20346 22992 20352 23044
rect 20404 23032 20410 23044
rect 23385 23035 23443 23041
rect 23385 23032 23397 23035
rect 20404 23004 23397 23032
rect 20404 22992 20410 23004
rect 23385 23001 23397 23004
rect 23431 23001 23443 23035
rect 24780 23032 24808 23063
rect 24946 23060 24952 23072
rect 25004 23060 25010 23112
rect 25041 23103 25099 23109
rect 25041 23069 25053 23103
rect 25087 23100 25099 23103
rect 25222 23100 25228 23112
rect 25087 23072 25228 23100
rect 25087 23069 25099 23072
rect 25041 23063 25099 23069
rect 25222 23060 25228 23072
rect 25280 23060 25286 23112
rect 25501 23103 25559 23109
rect 25501 23069 25513 23103
rect 25547 23100 25559 23103
rect 28368 23100 28396 23276
rect 29086 23264 29092 23276
rect 29144 23264 29150 23316
rect 31938 23264 31944 23316
rect 31996 23304 32002 23316
rect 32033 23307 32091 23313
rect 32033 23304 32045 23307
rect 31996 23276 32045 23304
rect 31996 23264 32002 23276
rect 32033 23273 32045 23276
rect 32079 23273 32091 23307
rect 32033 23267 32091 23273
rect 29362 23236 29368 23248
rect 28745 23208 29368 23236
rect 28745 23177 28773 23208
rect 29362 23196 29368 23208
rect 29420 23196 29426 23248
rect 31294 23236 31300 23248
rect 31255 23208 31300 23236
rect 31294 23196 31300 23208
rect 31352 23196 31358 23248
rect 28721 23171 28779 23177
rect 28721 23137 28733 23171
rect 28767 23137 28779 23171
rect 28721 23131 28779 23137
rect 28810 23128 28816 23180
rect 28868 23168 28874 23180
rect 28868 23140 28913 23168
rect 29488 23140 29776 23168
rect 28868 23128 28874 23140
rect 25547 23072 28396 23100
rect 25547 23069 25559 23072
rect 25501 23063 25559 23069
rect 28442 23060 28448 23112
rect 28500 23100 28506 23112
rect 28629 23103 28687 23109
rect 28500 23072 28545 23100
rect 28500 23060 28506 23072
rect 28629 23069 28641 23103
rect 28675 23069 28687 23103
rect 28629 23063 28687 23069
rect 25314 23032 25320 23044
rect 24780 23004 25320 23032
rect 23385 22995 23443 23001
rect 25314 22992 25320 23004
rect 25372 22992 25378 23044
rect 25406 22992 25412 23044
rect 25464 23032 25470 23044
rect 25746 23035 25804 23041
rect 25746 23032 25758 23035
rect 25464 23004 25758 23032
rect 25464 22992 25470 23004
rect 25746 23001 25758 23004
rect 25792 23001 25804 23035
rect 25746 22995 25804 23001
rect 27062 22992 27068 23044
rect 27120 23032 27126 23044
rect 27433 23035 27491 23041
rect 27433 23032 27445 23035
rect 27120 23004 27445 23032
rect 27120 22992 27126 23004
rect 27433 23001 27445 23004
rect 27479 23001 27491 23035
rect 27433 22995 27491 23001
rect 27522 22992 27528 23044
rect 27580 23032 27586 23044
rect 27614 23032 27620 23044
rect 27580 23004 27620 23032
rect 27580 22992 27586 23004
rect 27614 22992 27620 23004
rect 27672 22992 27678 23044
rect 28350 22992 28356 23044
rect 28408 23032 28414 23044
rect 28644 23032 28672 23063
rect 28994 23060 29000 23112
rect 29052 23109 29058 23112
rect 29052 23103 29066 23109
rect 29054 23100 29066 23103
rect 29488 23100 29516 23140
rect 29054 23072 29516 23100
rect 29641 23103 29699 23109
rect 29054 23069 29066 23072
rect 29052 23063 29066 23069
rect 29641 23069 29653 23103
rect 29687 23069 29699 23103
rect 29748 23100 29776 23140
rect 31018 23100 31024 23112
rect 29748 23072 31024 23100
rect 29641 23063 29699 23069
rect 29052 23060 29058 23063
rect 28408 23004 28672 23032
rect 28408 22992 28414 23004
rect 18782 22964 18788 22976
rect 18743 22936 18788 22964
rect 18782 22924 18788 22936
rect 18840 22924 18846 22976
rect 19426 22964 19432 22976
rect 19387 22936 19432 22964
rect 19426 22924 19432 22936
rect 19484 22924 19490 22976
rect 22738 22924 22744 22976
rect 22796 22964 22802 22976
rect 23017 22967 23075 22973
rect 23017 22964 23029 22967
rect 22796 22936 23029 22964
rect 22796 22924 22802 22936
rect 23017 22933 23029 22936
rect 23063 22933 23075 22967
rect 24578 22964 24584 22976
rect 24539 22936 24584 22964
rect 23017 22927 23075 22933
rect 24578 22924 24584 22936
rect 24636 22924 24642 22976
rect 27709 22967 27767 22973
rect 27709 22933 27721 22967
rect 27755 22964 27767 22967
rect 28626 22964 28632 22976
rect 27755 22936 28632 22964
rect 27755 22933 27767 22936
rect 27709 22927 27767 22933
rect 28626 22924 28632 22936
rect 28684 22924 28690 22976
rect 29178 22964 29184 22976
rect 29139 22936 29184 22964
rect 29178 22924 29184 22936
rect 29236 22924 29242 22976
rect 29656 22964 29684 23063
rect 31018 23060 31024 23072
rect 31076 23060 31082 23112
rect 31312 23100 31340 23196
rect 34330 23168 34336 23180
rect 34291 23140 34336 23168
rect 34330 23128 34336 23140
rect 34388 23128 34394 23180
rect 31665 23103 31723 23109
rect 31665 23100 31677 23103
rect 31312 23072 31677 23100
rect 31665 23069 31677 23072
rect 31711 23069 31723 23103
rect 31665 23063 31723 23069
rect 31849 23103 31907 23109
rect 31849 23069 31861 23103
rect 31895 23100 31907 23103
rect 32030 23100 32036 23112
rect 31895 23072 32036 23100
rect 31895 23069 31907 23072
rect 31849 23063 31907 23069
rect 32030 23060 32036 23072
rect 32088 23060 32094 23112
rect 32490 23100 32496 23112
rect 32451 23072 32496 23100
rect 32490 23060 32496 23072
rect 32548 23060 32554 23112
rect 29908 23035 29966 23041
rect 29908 23001 29920 23035
rect 29954 23032 29966 23035
rect 32674 23032 32680 23044
rect 29954 23004 31432 23032
rect 32635 23004 32680 23032
rect 29954 23001 29966 23004
rect 29908 22995 29966 23001
rect 30098 22964 30104 22976
rect 29656 22936 30104 22964
rect 30098 22924 30104 22936
rect 30156 22924 30162 22976
rect 30282 22924 30288 22976
rect 30340 22964 30346 22976
rect 30466 22964 30472 22976
rect 30340 22936 30472 22964
rect 30340 22924 30346 22936
rect 30466 22924 30472 22936
rect 30524 22924 30530 22976
rect 31021 22967 31079 22973
rect 31021 22933 31033 22967
rect 31067 22964 31079 22967
rect 31110 22964 31116 22976
rect 31067 22936 31116 22964
rect 31067 22933 31079 22936
rect 31021 22927 31079 22933
rect 31110 22924 31116 22936
rect 31168 22924 31174 22976
rect 31404 22964 31432 23004
rect 32674 22992 32680 23004
rect 32732 22992 32738 23044
rect 34514 22964 34520 22976
rect 31404 22936 34520 22964
rect 34514 22924 34520 22936
rect 34572 22924 34578 22976
rect 1104 22874 35027 22896
rect 1104 22822 9390 22874
rect 9442 22822 9454 22874
rect 9506 22822 9518 22874
rect 9570 22822 9582 22874
rect 9634 22822 9646 22874
rect 9698 22822 17831 22874
rect 17883 22822 17895 22874
rect 17947 22822 17959 22874
rect 18011 22822 18023 22874
rect 18075 22822 18087 22874
rect 18139 22822 26272 22874
rect 26324 22822 26336 22874
rect 26388 22822 26400 22874
rect 26452 22822 26464 22874
rect 26516 22822 26528 22874
rect 26580 22822 34713 22874
rect 34765 22822 34777 22874
rect 34829 22822 34841 22874
rect 34893 22822 34905 22874
rect 34957 22822 34969 22874
rect 35021 22822 35027 22874
rect 1104 22800 35027 22822
rect 17037 22763 17095 22769
rect 17037 22729 17049 22763
rect 17083 22760 17095 22763
rect 17310 22760 17316 22772
rect 17083 22732 17316 22760
rect 17083 22729 17095 22732
rect 17037 22723 17095 22729
rect 17310 22720 17316 22732
rect 17368 22720 17374 22772
rect 19702 22720 19708 22772
rect 19760 22760 19766 22772
rect 19797 22763 19855 22769
rect 19797 22760 19809 22763
rect 19760 22732 19809 22760
rect 19760 22720 19766 22732
rect 19797 22729 19809 22732
rect 19843 22729 19855 22763
rect 19797 22723 19855 22729
rect 21177 22763 21235 22769
rect 21177 22729 21189 22763
rect 21223 22760 21235 22763
rect 23474 22760 23480 22772
rect 21223 22732 23480 22760
rect 21223 22729 21235 22732
rect 21177 22723 21235 22729
rect 23474 22720 23480 22732
rect 23532 22720 23538 22772
rect 25222 22760 25228 22772
rect 24872 22732 25228 22760
rect 19058 22692 19064 22704
rect 18432 22664 19064 22692
rect 16574 22584 16580 22636
rect 16632 22624 16638 22636
rect 17221 22627 17279 22633
rect 17221 22624 17233 22627
rect 16632 22596 17233 22624
rect 16632 22584 16638 22596
rect 17221 22593 17233 22596
rect 17267 22624 17279 22627
rect 17586 22624 17592 22636
rect 17267 22596 17592 22624
rect 17267 22593 17279 22596
rect 17221 22587 17279 22593
rect 17586 22584 17592 22596
rect 17644 22584 17650 22636
rect 18432 22633 18460 22664
rect 19058 22652 19064 22664
rect 19116 22652 19122 22704
rect 20809 22695 20867 22701
rect 20809 22661 20821 22695
rect 20855 22692 20867 22695
rect 22272 22695 22330 22701
rect 20855 22664 22094 22692
rect 20855 22661 20867 22664
rect 20809 22655 20867 22661
rect 18417 22627 18475 22633
rect 18417 22593 18429 22627
rect 18463 22593 18475 22627
rect 18417 22587 18475 22593
rect 18684 22627 18742 22633
rect 18684 22593 18696 22627
rect 18730 22624 18742 22627
rect 19426 22624 19432 22636
rect 18730 22596 19432 22624
rect 18730 22593 18742 22596
rect 18684 22587 18742 22593
rect 19426 22584 19432 22596
rect 19484 22584 19490 22636
rect 20622 22624 20628 22636
rect 20583 22596 20628 22624
rect 20622 22584 20628 22596
rect 20680 22584 20686 22636
rect 20714 22584 20720 22636
rect 20772 22624 20778 22636
rect 20898 22624 20904 22636
rect 20772 22596 20904 22624
rect 20772 22584 20778 22596
rect 20898 22584 20904 22596
rect 20956 22584 20962 22636
rect 20990 22584 20996 22636
rect 21048 22624 21054 22636
rect 22066 22624 22094 22664
rect 22272 22661 22284 22695
rect 22318 22692 22330 22695
rect 24578 22692 24584 22704
rect 22318 22664 24584 22692
rect 22318 22661 22330 22664
rect 22272 22655 22330 22661
rect 24578 22652 24584 22664
rect 24636 22652 24642 22704
rect 23014 22624 23020 22636
rect 21048 22596 21093 22624
rect 22066 22596 23020 22624
rect 21048 22584 21054 22596
rect 23014 22584 23020 22596
rect 23072 22584 23078 22636
rect 24118 22633 24124 22636
rect 24112 22587 24124 22633
rect 24176 22624 24182 22636
rect 24176 22596 24212 22624
rect 24118 22584 24124 22587
rect 24176 22584 24182 22596
rect 17494 22556 17500 22568
rect 17455 22528 17500 22556
rect 17494 22516 17500 22528
rect 17552 22516 17558 22568
rect 21910 22516 21916 22568
rect 21968 22556 21974 22568
rect 22005 22559 22063 22565
rect 22005 22556 22017 22559
rect 21968 22528 22017 22556
rect 21968 22516 21974 22528
rect 22005 22525 22017 22528
rect 22051 22525 22063 22559
rect 22005 22519 22063 22525
rect 23474 22516 23480 22568
rect 23532 22556 23538 22568
rect 23845 22559 23903 22565
rect 23845 22556 23857 22559
rect 23532 22528 23857 22556
rect 23532 22516 23538 22528
rect 23845 22525 23857 22528
rect 23891 22525 23903 22559
rect 23845 22519 23903 22525
rect 16758 22448 16764 22500
rect 16816 22488 16822 22500
rect 17405 22491 17463 22497
rect 17405 22488 17417 22491
rect 16816 22460 17417 22488
rect 16816 22448 16822 22460
rect 17405 22457 17417 22460
rect 17451 22457 17463 22491
rect 17405 22451 17463 22457
rect 16390 22380 16396 22432
rect 16448 22420 16454 22432
rect 20070 22420 20076 22432
rect 16448 22392 20076 22420
rect 16448 22380 16454 22392
rect 20070 22380 20076 22392
rect 20128 22380 20134 22432
rect 23382 22420 23388 22432
rect 23295 22392 23388 22420
rect 23382 22380 23388 22392
rect 23440 22420 23446 22432
rect 24872 22420 24900 22732
rect 25222 22720 25228 22732
rect 25280 22760 25286 22772
rect 25869 22763 25927 22769
rect 25869 22760 25881 22763
rect 25280 22732 25881 22760
rect 25280 22720 25286 22732
rect 25869 22729 25881 22732
rect 25915 22729 25927 22763
rect 26602 22760 26608 22772
rect 26563 22732 26608 22760
rect 25869 22723 25927 22729
rect 26602 22720 26608 22732
rect 26660 22720 26666 22772
rect 26878 22720 26884 22772
rect 26936 22760 26942 22772
rect 29089 22763 29147 22769
rect 26936 22732 28948 22760
rect 26936 22720 26942 22732
rect 24946 22652 24952 22704
rect 25004 22692 25010 22704
rect 25130 22692 25136 22704
rect 25004 22664 25136 22692
rect 25004 22652 25010 22664
rect 25130 22652 25136 22664
rect 25188 22692 25194 22704
rect 26694 22692 26700 22704
rect 25188 22664 26004 22692
rect 25188 22652 25194 22664
rect 25406 22584 25412 22636
rect 25464 22624 25470 22636
rect 25976 22633 26004 22664
rect 26436 22664 26700 22692
rect 26436 22633 26464 22664
rect 26694 22652 26700 22664
rect 26752 22652 26758 22704
rect 28920 22692 28948 22732
rect 29089 22729 29101 22763
rect 29135 22729 29147 22763
rect 29089 22723 29147 22729
rect 28994 22692 29000 22704
rect 28920 22664 29000 22692
rect 28994 22652 29000 22664
rect 29052 22652 29058 22704
rect 29104 22692 29132 22723
rect 30466 22720 30472 22772
rect 30524 22760 30530 22772
rect 31386 22760 31392 22772
rect 30524 22732 30972 22760
rect 31347 22732 31392 22760
rect 30524 22720 30530 22732
rect 29270 22692 29276 22704
rect 29104 22664 29276 22692
rect 29270 22652 29276 22664
rect 29328 22652 29334 22704
rect 30276 22695 30334 22701
rect 30276 22661 30288 22695
rect 30322 22692 30334 22695
rect 30834 22692 30840 22704
rect 30322 22664 30840 22692
rect 30322 22661 30334 22664
rect 30276 22655 30334 22661
rect 30834 22652 30840 22664
rect 30892 22652 30898 22704
rect 30944 22692 30972 22732
rect 31386 22720 31392 22732
rect 31444 22720 31450 22772
rect 31496 22732 34192 22760
rect 31496 22692 31524 22732
rect 30944 22664 31524 22692
rect 25685 22627 25743 22633
rect 25685 22624 25697 22627
rect 25464 22596 25697 22624
rect 25464 22584 25470 22596
rect 25685 22593 25697 22596
rect 25731 22593 25743 22627
rect 25685 22587 25743 22593
rect 25961 22627 26019 22633
rect 25961 22593 25973 22627
rect 26007 22593 26019 22627
rect 25961 22587 26019 22593
rect 26421 22627 26479 22633
rect 26421 22593 26433 22627
rect 26467 22593 26479 22627
rect 26421 22587 26479 22593
rect 26605 22627 26663 22633
rect 26605 22593 26617 22627
rect 26651 22624 26663 22627
rect 27246 22624 27252 22636
rect 26651 22596 27252 22624
rect 26651 22593 26663 22596
rect 26605 22587 26663 22593
rect 27246 22584 27252 22596
rect 27304 22624 27310 22636
rect 27522 22624 27528 22636
rect 27304 22596 27528 22624
rect 27304 22584 27310 22596
rect 27522 22584 27528 22596
rect 27580 22584 27586 22636
rect 28902 22624 28908 22636
rect 28863 22596 28908 22624
rect 28902 22584 28908 22596
rect 28960 22584 28966 22636
rect 29181 22627 29239 22633
rect 29181 22593 29193 22627
rect 29227 22624 29239 22627
rect 30009 22627 30067 22633
rect 29227 22596 29261 22624
rect 29227 22593 29239 22596
rect 29181 22587 29239 22593
rect 30009 22593 30021 22627
rect 30055 22624 30067 22627
rect 30098 22624 30104 22636
rect 30055 22596 30104 22624
rect 30055 22593 30067 22596
rect 30009 22587 30067 22593
rect 25590 22516 25596 22568
rect 25648 22556 25654 22568
rect 27617 22559 27675 22565
rect 27617 22556 27629 22559
rect 25648 22528 27629 22556
rect 25648 22516 25654 22528
rect 27617 22525 27629 22528
rect 27663 22525 27675 22559
rect 27617 22519 27675 22525
rect 27985 22559 28043 22565
rect 27985 22525 27997 22559
rect 28031 22525 28043 22559
rect 27985 22519 28043 22525
rect 28077 22559 28135 22565
rect 28077 22525 28089 22559
rect 28123 22556 28135 22559
rect 29196 22556 29224 22587
rect 30098 22584 30104 22596
rect 30156 22584 30162 22636
rect 32306 22624 32312 22636
rect 32267 22596 32312 22624
rect 32306 22584 32312 22596
rect 32364 22584 32370 22636
rect 32576 22627 32634 22633
rect 32576 22593 32588 22627
rect 32622 22624 32634 22627
rect 33134 22624 33140 22636
rect 32622 22596 33140 22624
rect 32622 22593 32634 22596
rect 32576 22587 32634 22593
rect 33134 22584 33140 22596
rect 33192 22584 33198 22636
rect 34164 22633 34192 22732
rect 34238 22720 34244 22772
rect 34296 22760 34302 22772
rect 34296 22732 34341 22760
rect 34296 22720 34302 22732
rect 34149 22627 34207 22633
rect 34149 22593 34161 22627
rect 34195 22593 34207 22627
rect 34330 22624 34336 22636
rect 34291 22596 34336 22624
rect 34149 22587 34207 22593
rect 34330 22584 34336 22596
rect 34388 22584 34394 22636
rect 29730 22556 29736 22568
rect 28123 22528 29736 22556
rect 28123 22525 28135 22528
rect 28077 22519 28135 22525
rect 25314 22448 25320 22500
rect 25372 22488 25378 22500
rect 25685 22491 25743 22497
rect 25685 22488 25697 22491
rect 25372 22460 25697 22488
rect 25372 22448 25378 22460
rect 25685 22457 25697 22460
rect 25731 22457 25743 22491
rect 28000 22488 28028 22519
rect 29730 22516 29736 22528
rect 29788 22516 29794 22568
rect 29914 22488 29920 22500
rect 28000 22460 29920 22488
rect 25685 22451 25743 22457
rect 29914 22448 29920 22460
rect 29972 22448 29978 22500
rect 31294 22448 31300 22500
rect 31352 22488 31358 22500
rect 31352 22460 31754 22488
rect 31352 22448 31358 22460
rect 25222 22420 25228 22432
rect 23440 22392 24900 22420
rect 25183 22392 25228 22420
rect 23440 22380 23446 22392
rect 25222 22380 25228 22392
rect 25280 22380 25286 22432
rect 27798 22380 27804 22432
rect 27856 22420 27862 22432
rect 28261 22423 28319 22429
rect 28261 22420 28273 22423
rect 27856 22392 28273 22420
rect 27856 22380 27862 22392
rect 28261 22389 28273 22392
rect 28307 22389 28319 22423
rect 28718 22420 28724 22432
rect 28679 22392 28724 22420
rect 28261 22383 28319 22389
rect 28718 22380 28724 22392
rect 28776 22380 28782 22432
rect 31726 22420 31754 22460
rect 33689 22423 33747 22429
rect 33689 22420 33701 22423
rect 31726 22392 33701 22420
rect 33689 22389 33701 22392
rect 33735 22389 33747 22423
rect 33689 22383 33747 22389
rect 1104 22330 34868 22352
rect 1104 22278 5170 22330
rect 5222 22278 5234 22330
rect 5286 22278 5298 22330
rect 5350 22278 5362 22330
rect 5414 22278 5426 22330
rect 5478 22278 13611 22330
rect 13663 22278 13675 22330
rect 13727 22278 13739 22330
rect 13791 22278 13803 22330
rect 13855 22278 13867 22330
rect 13919 22278 22052 22330
rect 22104 22278 22116 22330
rect 22168 22278 22180 22330
rect 22232 22278 22244 22330
rect 22296 22278 22308 22330
rect 22360 22278 30493 22330
rect 30545 22278 30557 22330
rect 30609 22278 30621 22330
rect 30673 22278 30685 22330
rect 30737 22278 30749 22330
rect 30801 22278 34868 22330
rect 1104 22256 34868 22278
rect 19705 22219 19763 22225
rect 19705 22185 19717 22219
rect 19751 22216 19763 22219
rect 21818 22216 21824 22228
rect 19751 22188 21824 22216
rect 19751 22185 19763 22188
rect 19705 22179 19763 22185
rect 21818 22176 21824 22188
rect 21876 22176 21882 22228
rect 24394 22176 24400 22228
rect 24452 22216 24458 22228
rect 24581 22219 24639 22225
rect 24581 22216 24593 22219
rect 24452 22188 24593 22216
rect 24452 22176 24458 22188
rect 24581 22185 24593 22188
rect 24627 22185 24639 22219
rect 28810 22216 28816 22228
rect 28771 22188 28816 22216
rect 24581 22179 24639 22185
rect 28810 22176 28816 22188
rect 28868 22176 28874 22228
rect 30098 22216 30104 22228
rect 29748 22188 30104 22216
rect 16574 22148 16580 22160
rect 16224 22120 16580 22148
rect 16224 22089 16252 22120
rect 16574 22108 16580 22120
rect 16632 22108 16638 22160
rect 17589 22151 17647 22157
rect 17589 22117 17601 22151
rect 17635 22148 17647 22151
rect 18690 22148 18696 22160
rect 17635 22120 18460 22148
rect 18651 22120 18696 22148
rect 17635 22117 17647 22120
rect 17589 22111 17647 22117
rect 16209 22083 16267 22089
rect 16209 22049 16221 22083
rect 16255 22049 16267 22083
rect 16482 22080 16488 22092
rect 16443 22052 16488 22080
rect 16209 22043 16267 22049
rect 16482 22040 16488 22052
rect 16540 22040 16546 22092
rect 17310 22080 17316 22092
rect 17271 22052 17316 22080
rect 17310 22040 17316 22052
rect 17368 22040 17374 22092
rect 16117 22015 16175 22021
rect 16117 21981 16129 22015
rect 16163 21981 16175 22015
rect 16117 21975 16175 21981
rect 16132 21944 16160 21975
rect 16666 21972 16672 22024
rect 16724 22012 16730 22024
rect 18432 22021 18460 22120
rect 18690 22108 18696 22120
rect 18748 22108 18754 22160
rect 23106 22148 23112 22160
rect 20640 22120 23112 22148
rect 20346 22080 20352 22092
rect 20307 22052 20352 22080
rect 20346 22040 20352 22052
rect 20404 22040 20410 22092
rect 20640 22080 20668 22120
rect 23106 22108 23112 22120
rect 23164 22148 23170 22160
rect 23845 22151 23903 22157
rect 23164 22120 23704 22148
rect 23164 22108 23170 22120
rect 20456 22052 20668 22080
rect 20809 22083 20867 22089
rect 17221 22015 17279 22021
rect 17221 22012 17233 22015
rect 16724 21984 17233 22012
rect 16724 21972 16730 21984
rect 17221 21981 17233 21984
rect 17267 21981 17279 22015
rect 17221 21975 17279 21981
rect 18417 22015 18475 22021
rect 18417 21981 18429 22015
rect 18463 21981 18475 22015
rect 18598 22012 18604 22024
rect 18559 21984 18604 22012
rect 18417 21975 18475 21981
rect 18598 21972 18604 21984
rect 18656 21972 18662 22024
rect 18785 22015 18843 22021
rect 18785 21981 18797 22015
rect 18831 22012 18843 22015
rect 19058 22012 19064 22024
rect 18831 21984 19064 22012
rect 18831 21981 18843 21984
rect 18785 21975 18843 21981
rect 19058 21972 19064 21984
rect 19116 21972 19122 22024
rect 17494 21944 17500 21956
rect 16132 21916 17500 21944
rect 17494 21904 17500 21916
rect 17552 21904 17558 21956
rect 18877 21947 18935 21953
rect 18877 21913 18889 21947
rect 18923 21944 18935 21947
rect 18966 21944 18972 21956
rect 18923 21916 18972 21944
rect 18923 21913 18935 21916
rect 18877 21907 18935 21913
rect 18966 21904 18972 21916
rect 19024 21904 19030 21956
rect 19521 21947 19579 21953
rect 19521 21913 19533 21947
rect 19567 21944 19579 21947
rect 20456 21944 20484 22052
rect 20809 22049 20821 22083
rect 20855 22080 20867 22083
rect 21082 22080 21088 22092
rect 20855 22052 21088 22080
rect 20855 22049 20867 22052
rect 20809 22043 20867 22049
rect 21082 22040 21088 22052
rect 21140 22080 21146 22092
rect 22002 22080 22008 22092
rect 21140 22052 22008 22080
rect 21140 22040 21146 22052
rect 22002 22040 22008 22052
rect 22060 22040 22066 22092
rect 23566 22080 23572 22092
rect 22572 22052 23572 22080
rect 20533 22015 20591 22021
rect 20533 21981 20545 22015
rect 20579 21981 20591 22015
rect 20533 21975 20591 21981
rect 20625 22015 20683 22021
rect 20625 21981 20637 22015
rect 20671 22012 20683 22015
rect 20714 22012 20720 22024
rect 20671 21984 20720 22012
rect 20671 21981 20683 21984
rect 20625 21975 20683 21981
rect 19567 21916 20484 21944
rect 20548 21944 20576 21975
rect 20714 21972 20720 21984
rect 20772 21972 20778 22024
rect 20901 22015 20959 22021
rect 20901 21981 20913 22015
rect 20947 22012 20959 22015
rect 21174 22012 21180 22024
rect 20947 21984 21180 22012
rect 20947 21981 20959 21984
rect 20901 21975 20959 21981
rect 21174 21972 21180 21984
rect 21232 22012 21238 22024
rect 21358 22012 21364 22024
rect 21232 21984 21364 22012
rect 21232 21972 21238 21984
rect 21358 21972 21364 21984
rect 21416 21972 21422 22024
rect 21450 21972 21456 22024
rect 21508 22012 21514 22024
rect 21637 22015 21695 22021
rect 21637 22012 21649 22015
rect 21508 21984 21649 22012
rect 21508 21972 21514 21984
rect 21637 21981 21649 21984
rect 21683 21981 21695 22015
rect 21637 21975 21695 21981
rect 21730 22015 21788 22021
rect 21730 21981 21742 22015
rect 21776 21981 21788 22015
rect 21730 21975 21788 21981
rect 22143 22015 22201 22021
rect 22143 21981 22155 22015
rect 22189 22012 22201 22015
rect 22572 22012 22600 22052
rect 23566 22040 23572 22052
rect 23624 22040 23630 22092
rect 23676 22080 23704 22120
rect 23845 22117 23857 22151
rect 23891 22148 23903 22151
rect 23934 22148 23940 22160
rect 23891 22120 23940 22148
rect 23891 22117 23903 22120
rect 23845 22111 23903 22117
rect 23934 22108 23940 22120
rect 23992 22108 23998 22160
rect 27246 22148 27252 22160
rect 25976 22120 27252 22148
rect 24026 22080 24032 22092
rect 23676 22052 23796 22080
rect 23987 22052 24032 22080
rect 22738 22012 22744 22024
rect 22189 21984 22600 22012
rect 22699 21984 22744 22012
rect 22189 21981 22201 21984
rect 22143 21975 22201 21981
rect 20806 21944 20812 21956
rect 20548 21916 20812 21944
rect 19567 21913 19579 21916
rect 19521 21907 19579 21913
rect 20806 21904 20812 21916
rect 20864 21944 20870 21956
rect 20990 21944 20996 21956
rect 20864 21916 20996 21944
rect 20864 21904 20870 21916
rect 20990 21904 20996 21916
rect 21048 21904 21054 21956
rect 21744 21944 21772 21975
rect 22738 21972 22744 21984
rect 22796 21972 22802 22024
rect 22830 21972 22836 22024
rect 22888 22012 22894 22024
rect 23768 22021 23796 22052
rect 24026 22040 24032 22052
rect 24084 22080 24090 22092
rect 24394 22080 24400 22092
rect 24084 22052 24400 22080
rect 24084 22040 24090 22052
rect 24394 22040 24400 22052
rect 24452 22040 24458 22092
rect 24949 22083 25007 22089
rect 24949 22049 24961 22083
rect 24995 22080 25007 22083
rect 25976 22080 26004 22120
rect 27246 22108 27252 22120
rect 27304 22108 27310 22160
rect 28350 22108 28356 22160
rect 28408 22148 28414 22160
rect 29638 22148 29644 22160
rect 28408 22120 29644 22148
rect 28408 22108 28414 22120
rect 29638 22108 29644 22120
rect 29696 22108 29702 22160
rect 28442 22080 28448 22092
rect 24995 22052 26004 22080
rect 26068 22052 28448 22080
rect 24995 22049 25007 22052
rect 24949 22043 25007 22049
rect 23109 22015 23167 22021
rect 23109 22012 23121 22015
rect 22888 21984 23121 22012
rect 22888 21972 22894 21984
rect 23109 21981 23121 21984
rect 23155 21981 23167 22015
rect 23109 21975 23167 21981
rect 23753 22015 23811 22021
rect 23753 21981 23765 22015
rect 23799 21981 23811 22015
rect 24762 22012 24768 22024
rect 24723 21984 24768 22012
rect 23753 21975 23811 21981
rect 24762 21972 24768 21984
rect 24820 21972 24826 22024
rect 25038 22012 25044 22024
rect 24999 21984 25044 22012
rect 25038 21972 25044 21984
rect 25096 21972 25102 22024
rect 26068 22021 26096 22052
rect 28442 22040 28448 22052
rect 28500 22040 28506 22092
rect 29748 22089 29776 22188
rect 30098 22176 30104 22188
rect 30156 22176 30162 22228
rect 31018 22176 31024 22228
rect 31076 22216 31082 22228
rect 31113 22219 31171 22225
rect 31113 22216 31125 22219
rect 31076 22188 31125 22216
rect 31076 22176 31082 22188
rect 31113 22185 31125 22188
rect 31159 22185 31171 22219
rect 31113 22179 31171 22185
rect 29733 22083 29791 22089
rect 29733 22049 29745 22083
rect 29779 22049 29791 22083
rect 32582 22080 32588 22092
rect 29733 22043 29791 22049
rect 31956 22052 32588 22080
rect 31956 22024 31984 22052
rect 32582 22040 32588 22052
rect 32640 22040 32646 22092
rect 26053 22015 26111 22021
rect 26053 21981 26065 22015
rect 26099 21981 26111 22015
rect 26053 21975 26111 21981
rect 26421 22015 26479 22021
rect 26421 21981 26433 22015
rect 26467 22012 26479 22015
rect 27062 22012 27068 22024
rect 26467 21984 27068 22012
rect 26467 21981 26479 21984
rect 26421 21975 26479 21981
rect 27062 21972 27068 21984
rect 27120 21972 27126 22024
rect 27430 21972 27436 22024
rect 27488 22012 27494 22024
rect 27617 22015 27675 22021
rect 27617 22012 27629 22015
rect 27488 21984 27629 22012
rect 27488 21972 27494 21984
rect 27617 21981 27629 21984
rect 27663 21981 27675 22015
rect 27617 21975 27675 21981
rect 27709 22015 27767 22021
rect 27709 21981 27721 22015
rect 27755 21981 27767 22015
rect 27709 21975 27767 21981
rect 21192 21916 21772 21944
rect 21913 21947 21971 21953
rect 21192 21888 21220 21916
rect 21913 21913 21925 21947
rect 21959 21913 21971 21947
rect 21913 21907 21971 21913
rect 22005 21947 22063 21953
rect 22005 21913 22017 21947
rect 22051 21944 22063 21947
rect 22462 21944 22468 21956
rect 22051 21916 22468 21944
rect 22051 21913 22063 21916
rect 22005 21907 22063 21913
rect 19702 21836 19708 21888
rect 19760 21885 19766 21888
rect 19760 21879 19779 21885
rect 19767 21845 19779 21879
rect 19760 21839 19779 21845
rect 19889 21879 19947 21885
rect 19889 21845 19901 21879
rect 19935 21876 19947 21879
rect 20530 21876 20536 21888
rect 19935 21848 20536 21876
rect 19935 21845 19947 21848
rect 19889 21839 19947 21845
rect 19760 21836 19766 21839
rect 20530 21836 20536 21848
rect 20588 21836 20594 21888
rect 21174 21836 21180 21888
rect 21232 21836 21238 21888
rect 21726 21836 21732 21888
rect 21784 21876 21790 21888
rect 21928 21876 21956 21907
rect 22204 21888 22232 21916
rect 22462 21904 22468 21916
rect 22520 21904 22526 21956
rect 22554 21904 22560 21956
rect 22612 21944 22618 21956
rect 22925 21947 22983 21953
rect 22925 21944 22937 21947
rect 22612 21916 22937 21944
rect 22612 21904 22618 21916
rect 22925 21913 22937 21916
rect 22971 21913 22983 21947
rect 22925 21907 22983 21913
rect 23014 21904 23020 21956
rect 23072 21944 23078 21956
rect 23072 21916 23117 21944
rect 23072 21904 23078 21916
rect 25682 21904 25688 21956
rect 25740 21944 25746 21956
rect 26237 21947 26295 21953
rect 26237 21944 26249 21947
rect 25740 21916 26249 21944
rect 25740 21904 25746 21916
rect 26237 21913 26249 21916
rect 26283 21913 26295 21947
rect 26237 21907 26295 21913
rect 26329 21947 26387 21953
rect 26329 21913 26341 21947
rect 26375 21944 26387 21947
rect 26878 21944 26884 21956
rect 26375 21916 26884 21944
rect 26375 21913 26387 21916
rect 26329 21907 26387 21913
rect 26878 21904 26884 21916
rect 26936 21904 26942 21956
rect 27246 21904 27252 21956
rect 27304 21944 27310 21956
rect 27724 21944 27752 21975
rect 27798 21972 27804 22024
rect 27856 22012 27862 22024
rect 27985 22015 28043 22021
rect 27856 21984 27901 22012
rect 27856 21972 27862 21984
rect 27985 21981 27997 22015
rect 28031 22012 28043 22015
rect 28074 22012 28080 22024
rect 28031 21984 28080 22012
rect 28031 21981 28043 21984
rect 27985 21975 28043 21981
rect 28074 21972 28080 21984
rect 28132 21972 28138 22024
rect 29178 21972 29184 22024
rect 29236 22012 29242 22024
rect 29989 22015 30047 22021
rect 29989 22012 30001 22015
rect 29236 21984 30001 22012
rect 29236 21972 29242 21984
rect 29989 21981 30001 21984
rect 30035 21981 30047 22015
rect 29989 21975 30047 21981
rect 31754 21972 31760 22024
rect 31812 22012 31818 22024
rect 31938 22012 31944 22024
rect 31812 21984 31857 22012
rect 31899 21984 31944 22012
rect 31812 21972 31818 21984
rect 31938 21972 31944 21984
rect 31996 21972 32002 22024
rect 32033 22015 32091 22021
rect 32033 21981 32045 22015
rect 32079 22012 32091 22015
rect 32398 22012 32404 22024
rect 32079 21984 32404 22012
rect 32079 21981 32091 21984
rect 32033 21975 32091 21981
rect 32398 21972 32404 21984
rect 32456 21972 32462 22024
rect 32766 22012 32772 22024
rect 32727 21984 32772 22012
rect 32766 21972 32772 21984
rect 32824 21972 32830 22024
rect 27304 21916 27752 21944
rect 27304 21904 27310 21916
rect 27890 21904 27896 21956
rect 27948 21944 27954 21956
rect 28629 21947 28687 21953
rect 28629 21944 28641 21947
rect 27948 21916 28641 21944
rect 27948 21904 27954 21916
rect 28629 21913 28641 21916
rect 28675 21944 28687 21947
rect 31573 21947 31631 21953
rect 28675 21916 29132 21944
rect 28675 21913 28687 21916
rect 28629 21907 28687 21913
rect 21784 21848 21956 21876
rect 21784 21836 21790 21848
rect 22186 21836 22192 21888
rect 22244 21836 22250 21888
rect 22281 21879 22339 21885
rect 22281 21845 22293 21879
rect 22327 21876 22339 21879
rect 22370 21876 22376 21888
rect 22327 21848 22376 21876
rect 22327 21845 22339 21848
rect 22281 21839 22339 21845
rect 22370 21836 22376 21848
rect 22428 21836 22434 21888
rect 23290 21876 23296 21888
rect 23251 21848 23296 21876
rect 23290 21836 23296 21848
rect 23348 21836 23354 21888
rect 24026 21876 24032 21888
rect 23987 21848 24032 21876
rect 24026 21836 24032 21848
rect 24084 21836 24090 21888
rect 25774 21836 25780 21888
rect 25832 21876 25838 21888
rect 26605 21879 26663 21885
rect 26605 21876 26617 21879
rect 25832 21848 26617 21876
rect 25832 21836 25838 21848
rect 26605 21845 26617 21848
rect 26651 21845 26663 21879
rect 27338 21876 27344 21888
rect 27299 21848 27344 21876
rect 26605 21839 26663 21845
rect 27338 21836 27344 21848
rect 27396 21836 27402 21888
rect 27982 21836 27988 21888
rect 28040 21876 28046 21888
rect 28829 21879 28887 21885
rect 28829 21876 28841 21879
rect 28040 21848 28841 21876
rect 28040 21836 28046 21848
rect 28829 21845 28841 21848
rect 28875 21845 28887 21879
rect 28994 21876 29000 21888
rect 28955 21848 29000 21876
rect 28829 21839 28887 21845
rect 28994 21836 29000 21848
rect 29052 21836 29058 21888
rect 29104 21876 29132 21916
rect 31573 21913 31585 21947
rect 31619 21944 31631 21947
rect 33014 21947 33072 21953
rect 33014 21944 33026 21947
rect 31619 21916 33026 21944
rect 31619 21913 31631 21916
rect 31573 21907 31631 21913
rect 33014 21913 33026 21916
rect 33060 21913 33072 21947
rect 33014 21907 33072 21913
rect 30282 21876 30288 21888
rect 29104 21848 30288 21876
rect 30282 21836 30288 21848
rect 30340 21836 30346 21888
rect 32398 21836 32404 21888
rect 32456 21876 32462 21888
rect 34149 21879 34207 21885
rect 34149 21876 34161 21879
rect 32456 21848 34161 21876
rect 32456 21836 32462 21848
rect 34149 21845 34161 21848
rect 34195 21845 34207 21879
rect 34149 21839 34207 21845
rect 1104 21786 35027 21808
rect 1104 21734 9390 21786
rect 9442 21734 9454 21786
rect 9506 21734 9518 21786
rect 9570 21734 9582 21786
rect 9634 21734 9646 21786
rect 9698 21734 17831 21786
rect 17883 21734 17895 21786
rect 17947 21734 17959 21786
rect 18011 21734 18023 21786
rect 18075 21734 18087 21786
rect 18139 21734 26272 21786
rect 26324 21734 26336 21786
rect 26388 21734 26400 21786
rect 26452 21734 26464 21786
rect 26516 21734 26528 21786
rect 26580 21734 34713 21786
rect 34765 21734 34777 21786
rect 34829 21734 34841 21786
rect 34893 21734 34905 21786
rect 34957 21734 34969 21786
rect 35021 21734 35027 21786
rect 1104 21712 35027 21734
rect 15289 21675 15347 21681
rect 15289 21641 15301 21675
rect 15335 21672 15347 21675
rect 17126 21672 17132 21684
rect 15335 21644 17132 21672
rect 15335 21641 15347 21644
rect 15289 21635 15347 21641
rect 17126 21632 17132 21644
rect 17184 21632 17190 21684
rect 17310 21632 17316 21684
rect 17368 21672 17374 21684
rect 17773 21675 17831 21681
rect 17773 21672 17785 21675
rect 17368 21644 17785 21672
rect 17368 21632 17374 21644
rect 17773 21641 17785 21644
rect 17819 21641 17831 21675
rect 17773 21635 17831 21641
rect 19794 21632 19800 21684
rect 19852 21672 19858 21684
rect 21174 21672 21180 21684
rect 19852 21644 21180 21672
rect 19852 21632 19858 21644
rect 21174 21632 21180 21644
rect 21232 21632 21238 21684
rect 21450 21672 21456 21684
rect 21411 21644 21456 21672
rect 21450 21632 21456 21644
rect 21508 21632 21514 21684
rect 22557 21675 22615 21681
rect 22557 21641 22569 21675
rect 22603 21672 22615 21675
rect 23198 21672 23204 21684
rect 22603 21644 23204 21672
rect 22603 21641 22615 21644
rect 22557 21635 22615 21641
rect 23198 21632 23204 21644
rect 23256 21632 23262 21684
rect 27154 21632 27160 21684
rect 27212 21672 27218 21684
rect 33042 21672 33048 21684
rect 27212 21644 33048 21672
rect 27212 21632 27218 21644
rect 33042 21632 33048 21644
rect 33100 21632 33106 21684
rect 16114 21604 16120 21616
rect 15304 21576 16120 21604
rect 15304 21545 15332 21576
rect 16114 21564 16120 21576
rect 16172 21564 16178 21616
rect 20254 21564 20260 21616
rect 20312 21604 20318 21616
rect 21542 21604 21548 21616
rect 20312 21576 21548 21604
rect 20312 21564 20318 21576
rect 21542 21564 21548 21576
rect 21600 21604 21606 21616
rect 22281 21607 22339 21613
rect 22281 21604 22293 21607
rect 21600 21576 22293 21604
rect 21600 21564 21606 21576
rect 22281 21573 22293 21576
rect 22327 21573 22339 21607
rect 22281 21567 22339 21573
rect 25038 21564 25044 21616
rect 25096 21604 25102 21616
rect 25501 21607 25559 21613
rect 25501 21604 25513 21607
rect 25096 21576 25513 21604
rect 25096 21564 25102 21576
rect 25501 21573 25513 21576
rect 25547 21573 25559 21607
rect 26878 21604 26884 21616
rect 25501 21567 25559 21573
rect 26344 21576 26884 21604
rect 15105 21539 15163 21545
rect 15105 21505 15117 21539
rect 15151 21505 15163 21539
rect 15105 21499 15163 21505
rect 15289 21539 15347 21545
rect 15289 21505 15301 21539
rect 15335 21505 15347 21539
rect 16022 21536 16028 21548
rect 15983 21508 16028 21536
rect 15289 21499 15347 21505
rect 15120 21400 15148 21499
rect 16022 21496 16028 21508
rect 16080 21496 16086 21548
rect 17586 21536 17592 21548
rect 17547 21508 17592 21536
rect 17586 21496 17592 21508
rect 17644 21496 17650 21548
rect 18966 21545 18972 21548
rect 18960 21536 18972 21545
rect 18927 21508 18972 21536
rect 18960 21499 18972 21508
rect 18966 21496 18972 21499
rect 19024 21496 19030 21548
rect 20717 21539 20775 21545
rect 20717 21505 20729 21539
rect 20763 21505 20775 21539
rect 20717 21499 20775 21505
rect 20901 21539 20959 21545
rect 20901 21505 20913 21539
rect 20947 21505 20959 21539
rect 20901 21499 20959 21505
rect 15930 21468 15936 21480
rect 15891 21440 15936 21468
rect 15930 21428 15936 21440
rect 15988 21428 15994 21480
rect 16114 21468 16120 21480
rect 16075 21440 16120 21468
rect 16114 21428 16120 21440
rect 16172 21428 16178 21480
rect 16209 21471 16267 21477
rect 16209 21437 16221 21471
rect 16255 21468 16267 21471
rect 16850 21468 16856 21480
rect 16255 21440 16856 21468
rect 16255 21437 16267 21440
rect 16209 21431 16267 21437
rect 16850 21428 16856 21440
rect 16908 21428 16914 21480
rect 17494 21468 17500 21480
rect 17455 21440 17500 21468
rect 17494 21428 17500 21440
rect 17552 21428 17558 21480
rect 18693 21471 18751 21477
rect 18693 21437 18705 21471
rect 18739 21437 18751 21471
rect 18693 21431 18751 21437
rect 16022 21400 16028 21412
rect 15120 21372 16028 21400
rect 16022 21360 16028 21372
rect 16080 21400 16086 21412
rect 16482 21400 16488 21412
rect 16080 21372 16488 21400
rect 16080 21360 16086 21372
rect 16482 21360 16488 21372
rect 16540 21400 16546 21412
rect 17586 21400 17592 21412
rect 16540 21372 17592 21400
rect 16540 21360 16546 21372
rect 17586 21360 17592 21372
rect 17644 21360 17650 21412
rect 15749 21335 15807 21341
rect 15749 21301 15761 21335
rect 15795 21332 15807 21335
rect 16942 21332 16948 21344
rect 15795 21304 16948 21332
rect 15795 21301 15807 21304
rect 15749 21295 15807 21301
rect 16942 21292 16948 21304
rect 17000 21292 17006 21344
rect 18708 21332 18736 21431
rect 19426 21332 19432 21344
rect 18708 21304 19432 21332
rect 19426 21292 19432 21304
rect 19484 21292 19490 21344
rect 20070 21332 20076 21344
rect 20031 21304 20076 21332
rect 20070 21292 20076 21304
rect 20128 21292 20134 21344
rect 20732 21332 20760 21499
rect 20916 21400 20944 21499
rect 20990 21496 20996 21548
rect 21048 21536 21054 21548
rect 21048 21508 21093 21536
rect 21048 21496 21054 21508
rect 21174 21496 21180 21548
rect 21232 21536 21238 21548
rect 21269 21539 21327 21545
rect 21269 21536 21281 21539
rect 21232 21508 21281 21536
rect 21232 21496 21238 21508
rect 21269 21505 21281 21508
rect 21315 21505 21327 21539
rect 21269 21499 21327 21505
rect 21358 21496 21364 21548
rect 21416 21536 21422 21548
rect 22005 21539 22063 21545
rect 22005 21536 22017 21539
rect 21416 21508 22017 21536
rect 21416 21496 21422 21508
rect 22005 21505 22017 21508
rect 22051 21505 22063 21539
rect 22005 21499 22063 21505
rect 22094 21496 22100 21548
rect 22152 21536 22158 21548
rect 22189 21539 22247 21545
rect 22189 21536 22201 21539
rect 22152 21508 22201 21536
rect 22152 21496 22158 21508
rect 22189 21505 22201 21508
rect 22235 21505 22247 21539
rect 22189 21499 22247 21505
rect 22373 21539 22431 21545
rect 22373 21505 22385 21539
rect 22419 21536 22431 21539
rect 22419 21508 23152 21536
rect 22419 21505 22431 21508
rect 22373 21499 22431 21505
rect 21085 21471 21143 21477
rect 21085 21437 21097 21471
rect 21131 21468 21143 21471
rect 21450 21468 21456 21480
rect 21131 21440 21456 21468
rect 21131 21437 21143 21440
rect 21085 21431 21143 21437
rect 21450 21428 21456 21440
rect 21508 21428 21514 21480
rect 22462 21400 22468 21412
rect 20916 21372 22468 21400
rect 22462 21360 22468 21372
rect 22520 21360 22526 21412
rect 23124 21400 23152 21508
rect 23566 21496 23572 21548
rect 23624 21536 23630 21548
rect 23733 21539 23791 21545
rect 23733 21536 23745 21539
rect 23624 21508 23745 21536
rect 23624 21496 23630 21508
rect 23733 21505 23745 21508
rect 23779 21505 23791 21539
rect 23733 21499 23791 21505
rect 25317 21539 25375 21545
rect 25317 21505 25329 21539
rect 25363 21536 25375 21539
rect 25406 21536 25412 21548
rect 25363 21508 25412 21536
rect 25363 21505 25375 21508
rect 25317 21499 25375 21505
rect 25406 21496 25412 21508
rect 25464 21496 25470 21548
rect 25590 21536 25596 21548
rect 25551 21508 25596 21536
rect 25590 21496 25596 21508
rect 25648 21496 25654 21548
rect 26344 21545 26372 21576
rect 26878 21564 26884 21576
rect 26936 21564 26942 21616
rect 27338 21564 27344 21616
rect 27396 21604 27402 21616
rect 27678 21607 27736 21613
rect 27678 21604 27690 21607
rect 27396 21576 27690 21604
rect 27396 21564 27402 21576
rect 27678 21573 27690 21576
rect 27724 21573 27736 21607
rect 27678 21567 27736 21573
rect 27890 21564 27896 21616
rect 27948 21604 27954 21616
rect 28074 21604 28080 21616
rect 27948 21576 28080 21604
rect 27948 21564 27954 21576
rect 28074 21564 28080 21576
rect 28132 21564 28138 21616
rect 29270 21604 29276 21616
rect 29231 21576 29276 21604
rect 29270 21564 29276 21576
rect 29328 21564 29334 21616
rect 29473 21607 29531 21613
rect 29473 21604 29485 21607
rect 29380 21576 29485 21604
rect 26237 21539 26295 21545
rect 26237 21505 26249 21539
rect 26283 21505 26295 21539
rect 26237 21499 26295 21505
rect 26329 21539 26387 21545
rect 26329 21505 26341 21539
rect 26375 21505 26387 21539
rect 26329 21499 26387 21505
rect 26605 21539 26663 21545
rect 26605 21505 26617 21539
rect 26651 21536 26663 21539
rect 27433 21539 27491 21545
rect 26651 21508 27200 21536
rect 26651 21505 26663 21508
rect 26605 21499 26663 21505
rect 23474 21468 23480 21480
rect 23435 21440 23480 21468
rect 23474 21428 23480 21440
rect 23532 21428 23538 21480
rect 26252 21468 26280 21499
rect 27062 21468 27068 21480
rect 26252 21440 27068 21468
rect 27062 21428 27068 21440
rect 27120 21428 27126 21480
rect 23124 21372 23520 21400
rect 23382 21332 23388 21344
rect 20732 21304 23388 21332
rect 23382 21292 23388 21304
rect 23440 21292 23446 21344
rect 23492 21332 23520 21372
rect 24762 21360 24768 21412
rect 24820 21400 24826 21412
rect 25317 21403 25375 21409
rect 25317 21400 25329 21403
rect 24820 21372 25329 21400
rect 24820 21360 24826 21372
rect 25317 21369 25329 21372
rect 25363 21369 25375 21403
rect 25317 21363 25375 21369
rect 23658 21332 23664 21344
rect 23492 21304 23664 21332
rect 23658 21292 23664 21304
rect 23716 21292 23722 21344
rect 24857 21335 24915 21341
rect 24857 21301 24869 21335
rect 24903 21332 24915 21335
rect 25130 21332 25136 21344
rect 24903 21304 25136 21332
rect 24903 21301 24915 21304
rect 24857 21295 24915 21301
rect 25130 21292 25136 21304
rect 25188 21292 25194 21344
rect 26050 21332 26056 21344
rect 26011 21304 26056 21332
rect 26050 21292 26056 21304
rect 26108 21292 26114 21344
rect 26510 21332 26516 21344
rect 26471 21304 26516 21332
rect 26510 21292 26516 21304
rect 26568 21292 26574 21344
rect 26878 21292 26884 21344
rect 26936 21332 26942 21344
rect 27172 21332 27200 21508
rect 27433 21505 27445 21539
rect 27479 21536 27491 21539
rect 27522 21536 27528 21548
rect 27479 21508 27528 21536
rect 27479 21505 27491 21508
rect 27433 21499 27491 21505
rect 27522 21496 27528 21508
rect 27580 21496 27586 21548
rect 28258 21496 28264 21548
rect 28316 21536 28322 21548
rect 28316 21508 28856 21536
rect 28316 21496 28322 21508
rect 28828 21468 28856 21508
rect 28902 21496 28908 21548
rect 28960 21536 28966 21548
rect 29380 21536 29408 21576
rect 29473 21573 29485 21576
rect 29519 21573 29531 21607
rect 30282 21604 30288 21616
rect 30243 21576 30288 21604
rect 29473 21567 29531 21573
rect 30282 21564 30288 21576
rect 30340 21564 30346 21616
rect 30501 21607 30559 21613
rect 30501 21573 30513 21607
rect 30547 21604 30559 21607
rect 31662 21604 31668 21616
rect 30547 21576 31668 21604
rect 30547 21573 30559 21576
rect 30501 21567 30559 21573
rect 31662 21564 31668 21576
rect 31720 21564 31726 21616
rect 28960 21508 29408 21536
rect 31297 21539 31355 21545
rect 28960 21496 28966 21508
rect 31297 21505 31309 21539
rect 31343 21536 31355 21539
rect 31754 21536 31760 21548
rect 31343 21508 31760 21536
rect 31343 21505 31355 21508
rect 31297 21499 31355 21505
rect 31754 21496 31760 21508
rect 31812 21496 31818 21548
rect 32766 21496 32772 21548
rect 32824 21536 32830 21548
rect 33134 21545 33140 21548
rect 32861 21539 32919 21545
rect 32861 21536 32873 21539
rect 32824 21508 32873 21536
rect 32824 21496 32830 21508
rect 32861 21505 32873 21508
rect 32907 21505 32919 21539
rect 32861 21499 32919 21505
rect 33128 21499 33140 21545
rect 33192 21536 33198 21548
rect 33192 21508 33228 21536
rect 33134 21496 33140 21499
rect 33192 21496 33198 21508
rect 28828 21440 29776 21468
rect 29638 21400 29644 21412
rect 29599 21372 29644 21400
rect 29638 21360 29644 21372
rect 29696 21360 29702 21412
rect 29748 21400 29776 21440
rect 30926 21428 30932 21480
rect 30984 21468 30990 21480
rect 31110 21468 31116 21480
rect 30984 21440 31116 21468
rect 30984 21428 30990 21440
rect 31110 21428 31116 21440
rect 31168 21428 31174 21480
rect 30653 21403 30711 21409
rect 30653 21400 30665 21403
rect 29748 21372 30665 21400
rect 30653 21369 30665 21372
rect 30699 21369 30711 21403
rect 31846 21400 31852 21412
rect 30653 21363 30711 21369
rect 30760 21372 31852 21400
rect 27430 21332 27436 21344
rect 26936 21304 27436 21332
rect 26936 21292 26942 21304
rect 27430 21292 27436 21304
rect 27488 21332 27494 21344
rect 28813 21335 28871 21341
rect 28813 21332 28825 21335
rect 27488 21304 28825 21332
rect 27488 21292 27494 21304
rect 28813 21301 28825 21304
rect 28859 21301 28871 21335
rect 28813 21295 28871 21301
rect 29457 21335 29515 21341
rect 29457 21301 29469 21335
rect 29503 21332 29515 21335
rect 29730 21332 29736 21344
rect 29503 21304 29736 21332
rect 29503 21301 29515 21304
rect 29457 21295 29515 21301
rect 29730 21292 29736 21304
rect 29788 21292 29794 21344
rect 30469 21335 30527 21341
rect 30469 21301 30481 21335
rect 30515 21332 30527 21335
rect 30760 21332 30788 21372
rect 31846 21360 31852 21372
rect 31904 21360 31910 21412
rect 30515 21304 30788 21332
rect 30515 21301 30527 21304
rect 30469 21295 30527 21301
rect 30834 21292 30840 21344
rect 30892 21332 30898 21344
rect 31110 21332 31116 21344
rect 30892 21304 31116 21332
rect 30892 21292 30898 21304
rect 31110 21292 31116 21304
rect 31168 21332 31174 21344
rect 31481 21335 31539 21341
rect 31481 21332 31493 21335
rect 31168 21304 31493 21332
rect 31168 21292 31174 21304
rect 31481 21301 31493 21304
rect 31527 21301 31539 21335
rect 31481 21295 31539 21301
rect 31570 21292 31576 21344
rect 31628 21332 31634 21344
rect 33594 21332 33600 21344
rect 31628 21304 33600 21332
rect 31628 21292 31634 21304
rect 33594 21292 33600 21304
rect 33652 21332 33658 21344
rect 34241 21335 34299 21341
rect 34241 21332 34253 21335
rect 33652 21304 34253 21332
rect 33652 21292 33658 21304
rect 34241 21301 34253 21304
rect 34287 21301 34299 21335
rect 34241 21295 34299 21301
rect 1104 21242 34868 21264
rect 1104 21190 5170 21242
rect 5222 21190 5234 21242
rect 5286 21190 5298 21242
rect 5350 21190 5362 21242
rect 5414 21190 5426 21242
rect 5478 21190 13611 21242
rect 13663 21190 13675 21242
rect 13727 21190 13739 21242
rect 13791 21190 13803 21242
rect 13855 21190 13867 21242
rect 13919 21190 22052 21242
rect 22104 21190 22116 21242
rect 22168 21190 22180 21242
rect 22232 21190 22244 21242
rect 22296 21190 22308 21242
rect 22360 21190 30493 21242
rect 30545 21190 30557 21242
rect 30609 21190 30621 21242
rect 30673 21190 30685 21242
rect 30737 21190 30749 21242
rect 30801 21190 34868 21242
rect 1104 21168 34868 21190
rect 15930 21088 15936 21140
rect 15988 21128 15994 21140
rect 16666 21128 16672 21140
rect 15988 21100 16672 21128
rect 15988 21088 15994 21100
rect 16666 21088 16672 21100
rect 16724 21088 16730 21140
rect 19702 21088 19708 21140
rect 19760 21128 19766 21140
rect 22646 21128 22652 21140
rect 19760 21100 22652 21128
rect 19760 21088 19766 21100
rect 22646 21088 22652 21100
rect 22704 21088 22710 21140
rect 23566 21128 23572 21140
rect 23527 21100 23572 21128
rect 23566 21088 23572 21100
rect 23624 21088 23630 21140
rect 25130 21128 25136 21140
rect 24136 21100 25136 21128
rect 17773 21063 17831 21069
rect 17773 21029 17785 21063
rect 17819 21060 17831 21063
rect 20073 21063 20131 21069
rect 17819 21032 18757 21060
rect 17819 21029 17831 21032
rect 17773 21023 17831 21029
rect 16393 20995 16451 21001
rect 16393 20961 16405 20995
rect 16439 20992 16451 20995
rect 16574 20992 16580 21004
rect 16439 20964 16580 20992
rect 16439 20961 16451 20964
rect 16393 20955 16451 20961
rect 16574 20952 16580 20964
rect 16632 20952 16638 21004
rect 17497 20995 17555 21001
rect 17497 20961 17509 20995
rect 17543 20992 17555 20995
rect 18230 20992 18236 21004
rect 17543 20964 18236 20992
rect 17543 20961 17555 20964
rect 17497 20955 17555 20961
rect 18230 20952 18236 20964
rect 18288 20952 18294 21004
rect 16301 20927 16359 20933
rect 16301 20893 16313 20927
rect 16347 20924 16359 20927
rect 16666 20924 16672 20936
rect 16347 20896 16672 20924
rect 16347 20893 16359 20896
rect 16301 20887 16359 20893
rect 16666 20884 16672 20896
rect 16724 20884 16730 20936
rect 17126 20884 17132 20936
rect 17184 20924 17190 20936
rect 17589 20927 17647 20933
rect 17589 20924 17601 20927
rect 17184 20896 17601 20924
rect 17184 20884 17190 20896
rect 17589 20893 17601 20896
rect 17635 20893 17647 20927
rect 17589 20887 17647 20893
rect 18414 20884 18420 20936
rect 18472 20934 18478 20936
rect 18472 20933 18506 20934
rect 18729 20933 18757 21032
rect 20073 21029 20085 21063
rect 20119 21060 20131 21063
rect 24136 21060 24164 21100
rect 25130 21088 25136 21100
rect 25188 21088 25194 21140
rect 29454 21088 29460 21140
rect 29512 21128 29518 21140
rect 30101 21131 30159 21137
rect 30101 21128 30113 21131
rect 29512 21100 30113 21128
rect 29512 21088 29518 21100
rect 30101 21097 30113 21100
rect 30147 21097 30159 21131
rect 31570 21128 31576 21140
rect 30101 21091 30159 21097
rect 30668 21100 31576 21128
rect 20119 21032 23796 21060
rect 20119 21029 20131 21032
rect 20073 21023 20131 21029
rect 20272 20964 22094 20992
rect 18472 20927 18521 20933
rect 18714 20927 18772 20933
rect 18472 20893 18475 20927
rect 18509 20893 18521 20927
rect 18614 20921 18672 20927
rect 18614 20914 18626 20921
rect 18472 20887 18521 20893
rect 18472 20884 18478 20887
rect 18598 20862 18604 20914
rect 18660 20887 18672 20921
rect 18714 20893 18726 20927
rect 18760 20893 18772 20927
rect 18874 20924 18880 20936
rect 18835 20896 18880 20924
rect 18714 20887 18772 20893
rect 18656 20881 18672 20887
rect 18874 20884 18880 20896
rect 18932 20884 18938 20936
rect 20272 20933 20300 20964
rect 19429 20927 19487 20933
rect 19429 20893 19441 20927
rect 19475 20924 19487 20927
rect 20257 20927 20315 20933
rect 19475 20896 19932 20924
rect 19475 20893 19487 20896
rect 19429 20887 19487 20893
rect 18656 20862 18662 20881
rect 17129 20791 17187 20797
rect 17129 20757 17141 20791
rect 17175 20788 17187 20791
rect 18138 20788 18144 20800
rect 17175 20760 18144 20788
rect 17175 20757 17187 20760
rect 17129 20751 17187 20757
rect 18138 20748 18144 20760
rect 18196 20748 18202 20800
rect 18233 20791 18291 20797
rect 18233 20757 18245 20791
rect 18279 20788 18291 20791
rect 19334 20788 19340 20800
rect 18279 20760 19340 20788
rect 18279 20757 18291 20760
rect 18233 20751 18291 20757
rect 19334 20748 19340 20760
rect 19392 20748 19398 20800
rect 19518 20788 19524 20800
rect 19479 20760 19524 20788
rect 19518 20748 19524 20760
rect 19576 20748 19582 20800
rect 19904 20788 19932 20896
rect 20257 20893 20269 20927
rect 20303 20893 20315 20927
rect 20257 20887 20315 20893
rect 20346 20884 20352 20936
rect 20404 20924 20410 20936
rect 20809 20927 20867 20933
rect 20404 20896 20449 20924
rect 20404 20884 20410 20896
rect 20809 20893 20821 20927
rect 20855 20924 20867 20927
rect 20898 20924 20904 20936
rect 20855 20896 20904 20924
rect 20855 20893 20867 20896
rect 20809 20887 20867 20893
rect 20898 20884 20904 20896
rect 20956 20884 20962 20936
rect 21450 20884 21456 20936
rect 21508 20924 21514 20936
rect 21726 20924 21732 20936
rect 21508 20896 21732 20924
rect 21508 20884 21514 20896
rect 21726 20884 21732 20896
rect 21784 20884 21790 20936
rect 22066 20924 22094 20964
rect 23768 20933 23796 21032
rect 23952 21032 24164 21060
rect 23952 20992 23980 21032
rect 23860 20964 23980 20992
rect 23753 20927 23811 20933
rect 22204 20924 22324 20926
rect 22066 20898 23612 20924
rect 22066 20896 22232 20898
rect 22296 20896 23612 20898
rect 19978 20816 19984 20868
rect 20036 20856 20042 20868
rect 20073 20859 20131 20865
rect 20073 20856 20085 20859
rect 20036 20828 20085 20856
rect 20036 20816 20042 20828
rect 20073 20825 20085 20828
rect 20119 20825 20131 20859
rect 20916 20856 20944 20884
rect 22094 20856 22100 20868
rect 20916 20828 22100 20856
rect 20073 20819 20131 20825
rect 22094 20816 22100 20828
rect 22152 20816 22158 20868
rect 22557 20859 22615 20865
rect 22557 20825 22569 20859
rect 22603 20856 22615 20859
rect 23474 20856 23480 20868
rect 22603 20828 23480 20856
rect 22603 20825 22615 20828
rect 22557 20819 22615 20825
rect 23474 20816 23480 20828
rect 23532 20816 23538 20868
rect 23584 20856 23612 20896
rect 23753 20893 23765 20927
rect 23799 20893 23811 20927
rect 23753 20887 23811 20893
rect 23860 20856 23888 20964
rect 23937 20927 23995 20933
rect 23937 20893 23949 20927
rect 23983 20893 23995 20927
rect 23937 20887 23995 20893
rect 24029 20927 24087 20933
rect 24029 20893 24041 20927
rect 24075 20924 24087 20927
rect 24136 20924 24164 21032
rect 24486 21020 24492 21072
rect 24544 21060 24550 21072
rect 24544 21032 29132 21060
rect 24544 21020 24550 21032
rect 24210 20952 24216 21004
rect 24268 20992 24274 21004
rect 24268 20964 26096 20992
rect 24268 20952 24274 20964
rect 25038 20924 25044 20936
rect 24075 20896 24164 20924
rect 24596 20896 25044 20924
rect 24075 20893 24087 20896
rect 24029 20887 24087 20893
rect 23584 20828 23888 20856
rect 23952 20856 23980 20887
rect 24486 20856 24492 20868
rect 23952 20828 24492 20856
rect 24486 20816 24492 20828
rect 24544 20816 24550 20868
rect 24596 20788 24624 20896
rect 25038 20884 25044 20896
rect 25096 20884 25102 20936
rect 26068 20933 26096 20964
rect 28350 20952 28356 21004
rect 28408 20992 28414 21004
rect 28718 20992 28724 21004
rect 28408 20964 28724 20992
rect 28408 20952 28414 20964
rect 28718 20952 28724 20964
rect 28776 20952 28782 21004
rect 28994 20992 29000 21004
rect 28955 20964 29000 20992
rect 28994 20952 29000 20964
rect 29052 20952 29058 21004
rect 29104 20992 29132 21032
rect 29270 21020 29276 21072
rect 29328 21060 29334 21072
rect 29914 21060 29920 21072
rect 29328 21032 29920 21060
rect 29328 21020 29334 21032
rect 29914 21020 29920 21032
rect 29972 21020 29978 21072
rect 30466 20992 30472 21004
rect 29104 20964 30472 20992
rect 30466 20952 30472 20964
rect 30524 20952 30530 21004
rect 30561 20995 30619 21001
rect 30561 20961 30573 20995
rect 30607 20992 30619 20995
rect 30668 20992 30696 21100
rect 31570 21088 31576 21100
rect 31628 21088 31634 21140
rect 31849 21131 31907 21137
rect 31849 21097 31861 21131
rect 31895 21128 31907 21131
rect 31895 21100 32260 21128
rect 31895 21097 31907 21100
rect 31849 21091 31907 21097
rect 32122 21060 32128 21072
rect 30607 20964 30696 20992
rect 30760 21032 32128 21060
rect 30607 20961 30619 20964
rect 30561 20955 30619 20961
rect 26053 20927 26111 20933
rect 26053 20893 26065 20927
rect 26099 20924 26111 20927
rect 28534 20924 28540 20936
rect 26099 20896 28540 20924
rect 26099 20893 26111 20896
rect 26053 20887 26111 20893
rect 28534 20884 28540 20896
rect 28592 20884 28598 20936
rect 28629 20927 28687 20933
rect 28629 20893 28641 20927
rect 28675 20924 28687 20927
rect 29086 20924 29092 20936
rect 28675 20896 29092 20924
rect 28675 20893 28687 20896
rect 28629 20887 28687 20893
rect 29086 20884 29092 20896
rect 29144 20884 29150 20936
rect 29733 20927 29791 20933
rect 29733 20893 29745 20927
rect 29779 20924 29791 20927
rect 29822 20924 29828 20936
rect 29779 20896 29828 20924
rect 29779 20893 29791 20896
rect 29733 20887 29791 20893
rect 29822 20884 29828 20896
rect 29880 20884 29886 20936
rect 29917 20927 29975 20933
rect 29917 20893 29929 20927
rect 29963 20924 29975 20927
rect 30098 20924 30104 20936
rect 29963 20896 30104 20924
rect 29963 20893 29975 20896
rect 29917 20887 29975 20893
rect 30098 20884 30104 20896
rect 30156 20884 30162 20936
rect 30760 20933 30788 21032
rect 32122 21020 32128 21032
rect 32180 21020 32186 21072
rect 30834 20952 30840 21004
rect 30892 20992 30898 21004
rect 31386 20992 31392 21004
rect 30892 20964 31392 20992
rect 30892 20952 30898 20964
rect 31386 20952 31392 20964
rect 31444 20952 31450 21004
rect 31570 20952 31576 21004
rect 31628 20992 31634 21004
rect 32232 20992 32260 21100
rect 32398 20992 32404 21004
rect 31628 20964 32404 20992
rect 31628 20952 31634 20964
rect 32398 20952 32404 20964
rect 32456 20952 32462 21004
rect 30745 20927 30803 20933
rect 30745 20893 30757 20927
rect 30791 20893 30803 20927
rect 30745 20887 30803 20893
rect 31294 20884 31300 20936
rect 31352 20924 31358 20936
rect 32490 20924 32496 20936
rect 31352 20896 31708 20924
rect 32451 20896 32496 20924
rect 31352 20884 31358 20896
rect 24670 20816 24676 20868
rect 24728 20856 24734 20868
rect 24728 20828 24773 20856
rect 24728 20816 24734 20828
rect 26510 20816 26516 20868
rect 26568 20856 26574 20868
rect 27430 20856 27436 20868
rect 26568 20828 27436 20856
rect 26568 20816 26574 20828
rect 27430 20816 27436 20828
rect 27488 20816 27494 20868
rect 30006 20816 30012 20868
rect 30064 20856 30070 20868
rect 31680 20865 31708 20896
rect 32490 20884 32496 20896
rect 32548 20884 32554 20936
rect 31665 20859 31723 20865
rect 30064 20828 31524 20856
rect 30064 20816 30070 20828
rect 19904 20760 24624 20788
rect 24949 20791 25007 20797
rect 24949 20757 24961 20791
rect 24995 20788 25007 20791
rect 25406 20788 25412 20800
rect 24995 20760 25412 20788
rect 24995 20757 25007 20760
rect 24949 20751 25007 20757
rect 25406 20748 25412 20760
rect 25464 20748 25470 20800
rect 25958 20748 25964 20800
rect 26016 20788 26022 20800
rect 26878 20788 26884 20800
rect 26016 20760 26884 20788
rect 26016 20748 26022 20760
rect 26878 20748 26884 20760
rect 26936 20748 26942 20800
rect 27522 20788 27528 20800
rect 27483 20760 27528 20788
rect 27522 20748 27528 20760
rect 27580 20748 27586 20800
rect 30929 20791 30987 20797
rect 30929 20757 30941 20791
rect 30975 20788 30987 20791
rect 31386 20788 31392 20800
rect 30975 20760 31392 20788
rect 30975 20757 30987 20760
rect 30929 20751 30987 20757
rect 31386 20748 31392 20760
rect 31444 20748 31450 20800
rect 31496 20788 31524 20828
rect 31665 20825 31677 20859
rect 31711 20825 31723 20859
rect 32677 20859 32735 20865
rect 32677 20856 32689 20859
rect 31665 20819 31723 20825
rect 31772 20828 32689 20856
rect 31772 20788 31800 20828
rect 32677 20825 32689 20828
rect 32723 20825 32735 20859
rect 34330 20856 34336 20868
rect 34291 20828 34336 20856
rect 32677 20819 32735 20825
rect 34330 20816 34336 20828
rect 34388 20816 34394 20868
rect 31496 20760 31800 20788
rect 31846 20748 31852 20800
rect 31904 20797 31910 20800
rect 31904 20791 31923 20797
rect 31911 20757 31923 20791
rect 31904 20751 31923 20757
rect 32033 20791 32091 20797
rect 32033 20757 32045 20791
rect 32079 20788 32091 20791
rect 32122 20788 32128 20800
rect 32079 20760 32128 20788
rect 32079 20757 32091 20760
rect 32033 20751 32091 20757
rect 31904 20748 31910 20751
rect 32122 20748 32128 20760
rect 32180 20788 32186 20800
rect 32950 20788 32956 20800
rect 32180 20760 32956 20788
rect 32180 20748 32186 20760
rect 32950 20748 32956 20760
rect 33008 20748 33014 20800
rect 1104 20698 35027 20720
rect 1104 20646 9390 20698
rect 9442 20646 9454 20698
rect 9506 20646 9518 20698
rect 9570 20646 9582 20698
rect 9634 20646 9646 20698
rect 9698 20646 17831 20698
rect 17883 20646 17895 20698
rect 17947 20646 17959 20698
rect 18011 20646 18023 20698
rect 18075 20646 18087 20698
rect 18139 20646 26272 20698
rect 26324 20646 26336 20698
rect 26388 20646 26400 20698
rect 26452 20646 26464 20698
rect 26516 20646 26528 20698
rect 26580 20646 34713 20698
rect 34765 20646 34777 20698
rect 34829 20646 34841 20698
rect 34893 20646 34905 20698
rect 34957 20646 34969 20698
rect 35021 20646 35027 20698
rect 1104 20624 35027 20646
rect 16850 20544 16856 20596
rect 16908 20584 16914 20596
rect 17129 20587 17187 20593
rect 17129 20584 17141 20587
rect 16908 20556 17141 20584
rect 16908 20544 16914 20556
rect 17129 20553 17141 20556
rect 17175 20553 17187 20587
rect 17129 20547 17187 20553
rect 18230 20544 18236 20596
rect 18288 20584 18294 20596
rect 18417 20587 18475 20593
rect 18417 20584 18429 20587
rect 18288 20556 18429 20584
rect 18288 20544 18294 20556
rect 18417 20553 18429 20556
rect 18463 20553 18475 20587
rect 18417 20547 18475 20553
rect 20806 20544 20812 20596
rect 20864 20584 20870 20596
rect 21361 20587 21419 20593
rect 21361 20584 21373 20587
rect 20864 20556 21373 20584
rect 20864 20544 20870 20556
rect 21361 20553 21373 20556
rect 21407 20553 21419 20587
rect 21361 20547 21419 20553
rect 21634 20544 21640 20596
rect 21692 20584 21698 20596
rect 23014 20584 23020 20596
rect 21692 20556 23020 20584
rect 21692 20544 21698 20556
rect 23014 20544 23020 20556
rect 23072 20544 23078 20596
rect 23382 20544 23388 20596
rect 23440 20584 23446 20596
rect 24305 20587 24363 20593
rect 24305 20584 24317 20587
rect 23440 20556 24317 20584
rect 23440 20544 23446 20556
rect 24305 20553 24317 20556
rect 24351 20553 24363 20587
rect 24305 20547 24363 20553
rect 24486 20544 24492 20596
rect 24544 20584 24550 20596
rect 25038 20584 25044 20596
rect 24544 20556 25044 20584
rect 24544 20544 24550 20556
rect 25038 20544 25044 20556
rect 25096 20584 25102 20596
rect 25222 20584 25228 20596
rect 25096 20556 25228 20584
rect 25096 20544 25102 20556
rect 25222 20544 25228 20556
rect 25280 20544 25286 20596
rect 25501 20587 25559 20593
rect 25501 20553 25513 20587
rect 25547 20584 25559 20587
rect 26050 20584 26056 20596
rect 25547 20556 26056 20584
rect 25547 20553 25559 20556
rect 25501 20547 25559 20553
rect 26050 20544 26056 20556
rect 26108 20544 26114 20596
rect 26326 20544 26332 20596
rect 26384 20584 26390 20596
rect 26970 20584 26976 20596
rect 26384 20556 26976 20584
rect 26384 20544 26390 20556
rect 26970 20544 26976 20556
rect 27028 20544 27034 20596
rect 30190 20544 30196 20596
rect 30248 20584 30254 20596
rect 30248 20556 34192 20584
rect 30248 20544 30254 20556
rect 16114 20476 16120 20528
rect 16172 20516 16178 20528
rect 16172 20488 17448 20516
rect 16172 20476 16178 20488
rect 16022 20448 16028 20460
rect 15983 20420 16028 20448
rect 16022 20408 16028 20420
rect 16080 20408 16086 20460
rect 16206 20448 16212 20460
rect 16167 20420 16212 20448
rect 16206 20408 16212 20420
rect 16264 20408 16270 20460
rect 16574 20408 16580 20460
rect 16632 20448 16638 20460
rect 17313 20451 17371 20457
rect 17313 20448 17325 20451
rect 16632 20420 17325 20448
rect 16632 20408 16638 20420
rect 17313 20417 17325 20420
rect 17359 20417 17371 20451
rect 17420 20448 17448 20488
rect 17586 20476 17592 20528
rect 17644 20516 17650 20528
rect 18049 20519 18107 20525
rect 18049 20516 18061 20519
rect 17644 20488 18061 20516
rect 17644 20476 17650 20488
rect 18049 20485 18061 20488
rect 18095 20485 18107 20519
rect 18049 20479 18107 20485
rect 19334 20476 19340 20528
rect 19392 20516 19398 20528
rect 19674 20519 19732 20525
rect 19674 20516 19686 20519
rect 19392 20488 19686 20516
rect 19392 20476 19398 20488
rect 19674 20485 19686 20488
rect 19720 20485 19732 20519
rect 19674 20479 19732 20485
rect 22370 20476 22376 20528
rect 22428 20516 22434 20528
rect 22830 20516 22836 20528
rect 22428 20488 22836 20516
rect 22428 20476 22434 20488
rect 22830 20476 22836 20488
rect 22888 20476 22894 20528
rect 26237 20519 26295 20525
rect 26237 20485 26249 20519
rect 26283 20516 26295 20519
rect 26602 20516 26608 20528
rect 26283 20488 26608 20516
rect 26283 20485 26295 20488
rect 26237 20479 26295 20485
rect 26602 20476 26608 20488
rect 26660 20476 26666 20528
rect 27522 20516 27528 20528
rect 27172 20488 27528 20516
rect 18233 20451 18291 20457
rect 18233 20448 18245 20451
rect 17420 20420 18245 20448
rect 17313 20411 17371 20417
rect 18233 20417 18245 20420
rect 18279 20417 18291 20451
rect 19426 20448 19432 20460
rect 19387 20420 19432 20448
rect 18233 20411 18291 20417
rect 19426 20408 19432 20420
rect 19484 20408 19490 20460
rect 19536 20420 20484 20448
rect 16666 20340 16672 20392
rect 16724 20380 16730 20392
rect 17589 20383 17647 20389
rect 17589 20380 17601 20383
rect 16724 20352 17601 20380
rect 16724 20340 16730 20352
rect 17589 20349 17601 20352
rect 17635 20380 17647 20383
rect 19334 20380 19340 20392
rect 17635 20352 19340 20380
rect 17635 20349 17647 20352
rect 17589 20343 17647 20349
rect 19334 20340 19340 20352
rect 19392 20340 19398 20392
rect 19536 20380 19564 20420
rect 19444 20352 19564 20380
rect 16758 20272 16764 20324
rect 16816 20312 16822 20324
rect 17494 20312 17500 20324
rect 16816 20284 17172 20312
rect 17407 20284 17500 20312
rect 16816 20272 16822 20284
rect 16025 20247 16083 20253
rect 16025 20213 16037 20247
rect 16071 20244 16083 20247
rect 17034 20244 17040 20256
rect 16071 20216 17040 20244
rect 16071 20213 16083 20216
rect 16025 20207 16083 20213
rect 17034 20204 17040 20216
rect 17092 20204 17098 20256
rect 17144 20244 17172 20284
rect 17494 20272 17500 20284
rect 17552 20312 17558 20324
rect 18506 20312 18512 20324
rect 17552 20284 18512 20312
rect 17552 20272 17558 20284
rect 18506 20272 18512 20284
rect 18564 20312 18570 20324
rect 19444 20312 19472 20352
rect 18564 20284 19472 20312
rect 20456 20312 20484 20420
rect 20806 20408 20812 20460
rect 20864 20448 20870 20460
rect 21269 20451 21327 20457
rect 21269 20448 21281 20451
rect 20864 20420 21281 20448
rect 20864 20408 20870 20420
rect 21269 20417 21281 20420
rect 21315 20417 21327 20451
rect 21269 20411 21327 20417
rect 21910 20408 21916 20460
rect 21968 20448 21974 20460
rect 22005 20451 22063 20457
rect 22005 20448 22017 20451
rect 21968 20420 22017 20448
rect 21968 20408 21974 20420
rect 22005 20417 22017 20420
rect 22051 20417 22063 20451
rect 22005 20411 22063 20417
rect 22272 20451 22330 20457
rect 22272 20417 22284 20451
rect 22318 20448 22330 20451
rect 22738 20448 22744 20460
rect 22318 20420 22744 20448
rect 22318 20417 22330 20420
rect 22272 20411 22330 20417
rect 22738 20408 22744 20420
rect 22796 20408 22802 20460
rect 23750 20408 23756 20460
rect 23808 20448 23814 20460
rect 23845 20451 23903 20457
rect 23845 20448 23857 20451
rect 23808 20420 23857 20448
rect 23808 20408 23814 20420
rect 23845 20417 23857 20420
rect 23891 20417 23903 20451
rect 23845 20411 23903 20417
rect 25317 20451 25375 20457
rect 25317 20417 25329 20451
rect 25363 20417 25375 20451
rect 25317 20411 25375 20417
rect 25593 20451 25651 20457
rect 25593 20417 25605 20451
rect 25639 20448 25651 20451
rect 25774 20448 25780 20460
rect 25639 20420 25780 20448
rect 25639 20417 25651 20420
rect 25593 20411 25651 20417
rect 25332 20380 25360 20411
rect 25774 20408 25780 20420
rect 25832 20408 25838 20460
rect 25958 20408 25964 20460
rect 26016 20448 26022 20460
rect 26053 20451 26111 20457
rect 26053 20448 26065 20451
rect 26016 20420 26065 20448
rect 26016 20408 26022 20420
rect 26053 20417 26065 20420
rect 26099 20417 26111 20451
rect 26326 20448 26332 20460
rect 26287 20420 26332 20448
rect 26053 20411 26111 20417
rect 26326 20408 26332 20420
rect 26384 20408 26390 20460
rect 26418 20408 26424 20460
rect 26476 20448 26482 20460
rect 27172 20457 27200 20488
rect 27522 20476 27528 20488
rect 27580 20516 27586 20528
rect 29822 20516 29828 20528
rect 27580 20488 29828 20516
rect 27580 20476 27586 20488
rect 29822 20476 29828 20488
rect 29880 20476 29886 20528
rect 32766 20516 32772 20528
rect 32324 20488 32772 20516
rect 32324 20460 32352 20488
rect 32766 20476 32772 20488
rect 32824 20476 32830 20528
rect 27157 20451 27215 20457
rect 26476 20420 26521 20448
rect 26476 20408 26482 20420
rect 27157 20417 27169 20451
rect 27203 20417 27215 20451
rect 27157 20411 27215 20417
rect 27246 20408 27252 20460
rect 27304 20448 27310 20460
rect 27413 20451 27471 20457
rect 27413 20448 27425 20451
rect 27304 20420 27425 20448
rect 27304 20408 27310 20420
rect 27413 20417 27425 20420
rect 27459 20417 27471 20451
rect 27413 20411 27471 20417
rect 28166 20408 28172 20460
rect 28224 20448 28230 20460
rect 28902 20448 28908 20460
rect 28224 20420 28908 20448
rect 28224 20408 28230 20420
rect 28902 20408 28908 20420
rect 28960 20408 28966 20460
rect 28994 20408 29000 20460
rect 29052 20448 29058 20460
rect 29181 20451 29239 20457
rect 29181 20448 29193 20451
rect 29052 20420 29193 20448
rect 29052 20408 29058 20420
rect 29181 20417 29193 20420
rect 29227 20448 29239 20451
rect 30193 20451 30251 20457
rect 30193 20448 30205 20451
rect 29227 20420 30205 20448
rect 29227 20417 29239 20420
rect 29181 20411 29239 20417
rect 30193 20417 30205 20420
rect 30239 20417 30251 20451
rect 31202 20448 31208 20460
rect 31163 20420 31208 20448
rect 30193 20411 30251 20417
rect 31202 20408 31208 20420
rect 31260 20408 31266 20460
rect 31386 20448 31392 20460
rect 31347 20420 31392 20448
rect 31386 20408 31392 20420
rect 31444 20408 31450 20460
rect 32306 20408 32312 20460
rect 32364 20448 32370 20460
rect 32576 20451 32634 20457
rect 32364 20420 32457 20448
rect 32364 20408 32370 20420
rect 32576 20417 32588 20451
rect 32622 20448 32634 20451
rect 33686 20448 33692 20460
rect 32622 20420 33692 20448
rect 32622 20417 32634 20420
rect 32576 20411 32634 20417
rect 33686 20408 33692 20420
rect 33744 20408 33750 20460
rect 34164 20457 34192 20556
rect 34238 20544 34244 20596
rect 34296 20584 34302 20596
rect 34296 20556 34341 20584
rect 34296 20544 34302 20556
rect 34149 20451 34207 20457
rect 34149 20417 34161 20451
rect 34195 20417 34207 20451
rect 34149 20411 34207 20417
rect 34238 20408 34244 20460
rect 34296 20448 34302 20460
rect 34333 20451 34391 20457
rect 34333 20448 34345 20451
rect 34296 20420 34345 20448
rect 34296 20408 34302 20420
rect 34333 20417 34345 20420
rect 34379 20417 34391 20451
rect 34333 20411 34391 20417
rect 25332 20352 26648 20380
rect 20809 20315 20867 20321
rect 20809 20312 20821 20315
rect 20456 20284 20821 20312
rect 18564 20272 18570 20284
rect 20809 20281 20821 20284
rect 20855 20312 20867 20315
rect 21634 20312 21640 20324
rect 20855 20284 21640 20312
rect 20855 20281 20867 20284
rect 20809 20275 20867 20281
rect 21634 20272 21640 20284
rect 21692 20272 21698 20324
rect 23014 20272 23020 20324
rect 23072 20312 23078 20324
rect 23072 20284 23980 20312
rect 23072 20272 23078 20284
rect 21358 20244 21364 20256
rect 17144 20216 21364 20244
rect 21358 20204 21364 20216
rect 21416 20204 21422 20256
rect 23106 20204 23112 20256
rect 23164 20244 23170 20256
rect 23382 20244 23388 20256
rect 23164 20216 23388 20244
rect 23164 20204 23170 20216
rect 23382 20204 23388 20216
rect 23440 20204 23446 20256
rect 23952 20253 23980 20284
rect 26050 20272 26056 20324
rect 26108 20312 26114 20324
rect 26418 20312 26424 20324
rect 26108 20284 26424 20312
rect 26108 20272 26114 20284
rect 26418 20272 26424 20284
rect 26476 20272 26482 20324
rect 26620 20321 26648 20352
rect 28810 20340 28816 20392
rect 28868 20380 28874 20392
rect 29273 20383 29331 20389
rect 29273 20380 29285 20383
rect 28868 20352 29285 20380
rect 28868 20340 28874 20352
rect 29273 20349 29285 20352
rect 29319 20349 29331 20383
rect 29273 20343 29331 20349
rect 29365 20383 29423 20389
rect 29365 20349 29377 20383
rect 29411 20349 29423 20383
rect 29365 20343 29423 20349
rect 26605 20315 26663 20321
rect 26605 20281 26617 20315
rect 26651 20281 26663 20315
rect 26605 20275 26663 20281
rect 28537 20315 28595 20321
rect 28537 20281 28549 20315
rect 28583 20312 28595 20315
rect 28718 20312 28724 20324
rect 28583 20284 28724 20312
rect 28583 20281 28595 20284
rect 28537 20275 28595 20281
rect 28718 20272 28724 20284
rect 28776 20272 28782 20324
rect 28902 20272 28908 20324
rect 28960 20312 28966 20324
rect 29380 20312 29408 20343
rect 29454 20340 29460 20392
rect 29512 20380 29518 20392
rect 30098 20380 30104 20392
rect 29512 20352 29557 20380
rect 30059 20352 30104 20380
rect 29512 20340 29518 20352
rect 30098 20340 30104 20352
rect 30156 20340 30162 20392
rect 31481 20383 31539 20389
rect 31481 20349 31493 20383
rect 31527 20380 31539 20383
rect 31846 20380 31852 20392
rect 31527 20352 31852 20380
rect 31527 20349 31539 20352
rect 31481 20343 31539 20349
rect 31846 20340 31852 20352
rect 31904 20340 31910 20392
rect 28960 20284 29408 20312
rect 30561 20315 30619 20321
rect 28960 20272 28966 20284
rect 30561 20281 30573 20315
rect 30607 20312 30619 20315
rect 31938 20312 31944 20324
rect 30607 20284 31944 20312
rect 30607 20281 30619 20284
rect 30561 20275 30619 20281
rect 31938 20272 31944 20284
rect 31996 20272 32002 20324
rect 23937 20247 23995 20253
rect 23937 20213 23949 20247
rect 23983 20213 23995 20247
rect 23937 20207 23995 20213
rect 25133 20247 25191 20253
rect 25133 20213 25145 20247
rect 25179 20244 25191 20247
rect 26510 20244 26516 20256
rect 25179 20216 26516 20244
rect 25179 20213 25191 20216
rect 25133 20207 25191 20213
rect 26510 20204 26516 20216
rect 26568 20204 26574 20256
rect 28626 20204 28632 20256
rect 28684 20244 28690 20256
rect 28997 20247 29055 20253
rect 28997 20244 29009 20247
rect 28684 20216 29009 20244
rect 28684 20204 28690 20216
rect 28997 20213 29009 20216
rect 29043 20213 29055 20247
rect 31018 20244 31024 20256
rect 30979 20216 31024 20244
rect 28997 20207 29055 20213
rect 31018 20204 31024 20216
rect 31076 20204 31082 20256
rect 33689 20247 33747 20253
rect 33689 20213 33701 20247
rect 33735 20244 33747 20247
rect 33778 20244 33784 20256
rect 33735 20216 33784 20244
rect 33735 20213 33747 20216
rect 33689 20207 33747 20213
rect 33778 20204 33784 20216
rect 33836 20204 33842 20256
rect 1104 20154 34868 20176
rect 1104 20102 5170 20154
rect 5222 20102 5234 20154
rect 5286 20102 5298 20154
rect 5350 20102 5362 20154
rect 5414 20102 5426 20154
rect 5478 20102 13611 20154
rect 13663 20102 13675 20154
rect 13727 20102 13739 20154
rect 13791 20102 13803 20154
rect 13855 20102 13867 20154
rect 13919 20102 22052 20154
rect 22104 20102 22116 20154
rect 22168 20102 22180 20154
rect 22232 20102 22244 20154
rect 22296 20102 22308 20154
rect 22360 20102 30493 20154
rect 30545 20102 30557 20154
rect 30609 20102 30621 20154
rect 30673 20102 30685 20154
rect 30737 20102 30749 20154
rect 30801 20102 34868 20154
rect 1104 20080 34868 20102
rect 18414 20040 18420 20052
rect 15948 20012 18420 20040
rect 1946 19796 1952 19848
rect 2004 19836 2010 19848
rect 2041 19839 2099 19845
rect 2041 19836 2053 19839
rect 2004 19808 2053 19836
rect 2004 19796 2010 19808
rect 2041 19805 2053 19808
rect 2087 19836 2099 19839
rect 2498 19836 2504 19848
rect 2087 19808 2504 19836
rect 2087 19805 2099 19808
rect 2041 19799 2099 19805
rect 2498 19796 2504 19808
rect 2556 19796 2562 19848
rect 15948 19836 15976 20012
rect 18414 20000 18420 20012
rect 18472 20000 18478 20052
rect 21082 20040 21088 20052
rect 19444 20012 21088 20040
rect 16022 19932 16028 19984
rect 16080 19932 16086 19984
rect 17773 19975 17831 19981
rect 17773 19941 17785 19975
rect 17819 19972 17831 19975
rect 19444 19972 19472 20012
rect 21082 20000 21088 20012
rect 21140 20000 21146 20052
rect 21269 20043 21327 20049
rect 21269 20009 21281 20043
rect 21315 20040 21327 20043
rect 22554 20040 22560 20052
rect 21315 20012 22560 20040
rect 21315 20009 21327 20012
rect 21269 20003 21327 20009
rect 22554 20000 22560 20012
rect 22612 20000 22618 20052
rect 26513 20043 26571 20049
rect 26513 20009 26525 20043
rect 26559 20040 26571 20043
rect 27246 20040 27252 20052
rect 26559 20012 27252 20040
rect 26559 20009 26571 20012
rect 26513 20003 26571 20009
rect 27246 20000 27252 20012
rect 27304 20000 27310 20052
rect 31757 20043 31815 20049
rect 31757 20009 31769 20043
rect 31803 20040 31815 20043
rect 31846 20040 31852 20052
rect 31803 20012 31852 20040
rect 31803 20009 31815 20012
rect 31757 20003 31815 20009
rect 31846 20000 31852 20012
rect 31904 20000 31910 20052
rect 31938 20000 31944 20052
rect 31996 20040 32002 20052
rect 33226 20040 33232 20052
rect 31996 20012 33232 20040
rect 31996 20000 32002 20012
rect 33226 20000 33232 20012
rect 33284 20000 33290 20052
rect 17819 19944 19472 19972
rect 20809 19975 20867 19981
rect 17819 19941 17831 19944
rect 17773 19935 17831 19941
rect 20809 19941 20821 19975
rect 20855 19972 20867 19975
rect 21358 19972 21364 19984
rect 20855 19944 21364 19972
rect 20855 19941 20867 19944
rect 20809 19935 20867 19941
rect 21358 19932 21364 19944
rect 21416 19932 21422 19984
rect 21729 19975 21787 19981
rect 21729 19972 21741 19975
rect 21468 19944 21741 19972
rect 16040 19904 16068 19932
rect 16040 19876 16896 19904
rect 16025 19839 16083 19845
rect 16025 19836 16037 19839
rect 15948 19808 16037 19836
rect 16025 19805 16037 19808
rect 16071 19805 16083 19839
rect 16025 19799 16083 19805
rect 16209 19839 16267 19845
rect 16209 19805 16221 19839
rect 16255 19836 16267 19839
rect 16758 19836 16764 19848
rect 16255 19808 16764 19836
rect 16255 19805 16267 19808
rect 16209 19799 16267 19805
rect 16758 19796 16764 19808
rect 16816 19796 16822 19848
rect 16868 19845 16896 19876
rect 16942 19864 16948 19916
rect 17000 19904 17006 19916
rect 19426 19904 19432 19916
rect 17000 19876 17172 19904
rect 17000 19864 17006 19876
rect 17144 19848 17172 19876
rect 17696 19876 19288 19904
rect 19387 19876 19432 19904
rect 16853 19839 16911 19845
rect 16853 19805 16865 19839
rect 16899 19805 16911 19839
rect 17034 19836 17040 19848
rect 16995 19808 17040 19836
rect 16853 19799 16911 19805
rect 17034 19796 17040 19808
rect 17092 19796 17098 19848
rect 17126 19796 17132 19848
rect 17184 19836 17190 19848
rect 17696 19845 17724 19876
rect 17681 19839 17739 19845
rect 17184 19808 17277 19836
rect 17184 19796 17190 19808
rect 17681 19805 17693 19839
rect 17727 19805 17739 19839
rect 18601 19839 18659 19845
rect 18601 19836 18613 19839
rect 17681 19799 17739 19805
rect 17788 19808 18613 19836
rect 16117 19771 16175 19777
rect 16117 19737 16129 19771
rect 16163 19768 16175 19771
rect 17788 19768 17816 19808
rect 18601 19805 18613 19808
rect 18647 19805 18659 19839
rect 18601 19799 18659 19805
rect 18693 19839 18751 19845
rect 18693 19805 18705 19839
rect 18739 19836 18751 19839
rect 19058 19836 19064 19848
rect 18739 19808 19064 19836
rect 18739 19805 18751 19808
rect 18693 19799 18751 19805
rect 19058 19796 19064 19808
rect 19116 19796 19122 19848
rect 19260 19836 19288 19876
rect 19426 19864 19432 19876
rect 19484 19864 19490 19916
rect 20438 19864 20444 19916
rect 20496 19904 20502 19916
rect 21468 19904 21496 19944
rect 21729 19941 21741 19944
rect 21775 19972 21787 19975
rect 22370 19972 22376 19984
rect 21775 19944 22376 19972
rect 21775 19941 21787 19944
rect 21729 19935 21787 19941
rect 22370 19932 22376 19944
rect 22428 19932 22434 19984
rect 29730 19972 29736 19984
rect 27586 19944 29736 19972
rect 20496 19876 21496 19904
rect 20496 19864 20502 19876
rect 21634 19864 21640 19916
rect 21692 19904 21698 19916
rect 27338 19904 27344 19916
rect 21692 19876 21864 19904
rect 21692 19864 21698 19876
rect 20714 19836 20720 19848
rect 19260 19808 20720 19836
rect 20714 19796 20720 19808
rect 20772 19836 20778 19848
rect 21082 19836 21088 19848
rect 20772 19808 21088 19836
rect 20772 19796 20778 19808
rect 21082 19796 21088 19808
rect 21140 19796 21146 19848
rect 21450 19836 21456 19848
rect 21411 19808 21456 19836
rect 21450 19796 21456 19808
rect 21508 19796 21514 19848
rect 21542 19796 21548 19848
rect 21600 19836 21606 19848
rect 21836 19845 21864 19876
rect 26896 19876 27344 19904
rect 21821 19839 21879 19845
rect 21600 19808 21645 19836
rect 21600 19796 21606 19808
rect 21821 19805 21833 19839
rect 21867 19805 21879 19839
rect 21821 19799 21879 19805
rect 21910 19796 21916 19848
rect 21968 19836 21974 19848
rect 22373 19839 22431 19845
rect 22373 19836 22385 19839
rect 21968 19808 22385 19836
rect 21968 19796 21974 19808
rect 22373 19805 22385 19808
rect 22419 19836 22431 19839
rect 23474 19836 23480 19848
rect 22419 19808 23480 19836
rect 22419 19805 22431 19808
rect 22373 19799 22431 19805
rect 23474 19796 23480 19808
rect 23532 19836 23538 19848
rect 23842 19836 23848 19848
rect 23532 19808 23848 19836
rect 23532 19796 23538 19808
rect 23842 19796 23848 19808
rect 23900 19836 23906 19848
rect 24581 19839 24639 19845
rect 24581 19836 24593 19839
rect 23900 19808 24593 19836
rect 23900 19796 23906 19808
rect 24581 19805 24593 19808
rect 24627 19805 24639 19839
rect 26786 19836 26792 19848
rect 26747 19808 26792 19836
rect 24581 19799 24639 19805
rect 26786 19796 26792 19808
rect 26844 19796 26850 19848
rect 26896 19845 26924 19876
rect 27338 19864 27344 19876
rect 27396 19904 27402 19916
rect 27586 19904 27614 19944
rect 29730 19932 29736 19944
rect 29788 19932 29794 19984
rect 33778 19972 33784 19984
rect 31726 19944 33784 19972
rect 27396 19876 27614 19904
rect 28077 19907 28135 19913
rect 27396 19864 27402 19876
rect 28077 19873 28089 19907
rect 28123 19904 28135 19907
rect 29181 19907 29239 19913
rect 29181 19904 29193 19907
rect 28123 19876 29193 19904
rect 28123 19873 28135 19876
rect 28077 19867 28135 19873
rect 29181 19873 29193 19876
rect 29227 19873 29239 19907
rect 31726 19904 31754 19944
rect 33778 19932 33784 19944
rect 33836 19932 33842 19984
rect 29181 19867 29239 19873
rect 31588 19876 31754 19904
rect 32493 19907 32551 19913
rect 26881 19839 26939 19845
rect 26881 19805 26893 19839
rect 26927 19805 26939 19839
rect 26881 19799 26939 19805
rect 26973 19839 27031 19845
rect 26973 19805 26985 19839
rect 27019 19805 27031 19839
rect 26973 19799 27031 19805
rect 27157 19839 27215 19845
rect 27157 19805 27169 19839
rect 27203 19836 27215 19839
rect 27890 19836 27896 19848
rect 27203 19808 27896 19836
rect 27203 19805 27215 19808
rect 27157 19799 27215 19805
rect 18322 19768 18328 19780
rect 16163 19740 17816 19768
rect 18283 19740 18328 19768
rect 16163 19737 16175 19740
rect 16117 19731 16175 19737
rect 18322 19728 18328 19740
rect 18380 19728 18386 19780
rect 18785 19771 18843 19777
rect 18785 19737 18797 19771
rect 18831 19768 18843 19771
rect 19674 19771 19732 19777
rect 19674 19768 19686 19771
rect 18831 19740 19686 19768
rect 18831 19737 18843 19740
rect 18785 19731 18843 19737
rect 19674 19737 19686 19740
rect 19720 19737 19732 19771
rect 20070 19768 20076 19780
rect 19674 19731 19732 19737
rect 19812 19740 20076 19768
rect 1946 19660 1952 19712
rect 2004 19700 2010 19712
rect 2133 19703 2191 19709
rect 2133 19700 2145 19703
rect 2004 19672 2145 19700
rect 2004 19660 2010 19672
rect 2133 19669 2145 19672
rect 2179 19669 2191 19703
rect 16666 19700 16672 19712
rect 16627 19672 16672 19700
rect 2133 19663 2191 19669
rect 16666 19660 16672 19672
rect 16724 19660 16730 19712
rect 18417 19703 18475 19709
rect 18417 19669 18429 19703
rect 18463 19700 18475 19703
rect 18598 19700 18604 19712
rect 18463 19672 18604 19700
rect 18463 19669 18475 19672
rect 18417 19663 18475 19669
rect 18598 19660 18604 19672
rect 18656 19660 18662 19712
rect 19334 19660 19340 19712
rect 19392 19700 19398 19712
rect 19812 19700 19840 19740
rect 20070 19728 20076 19740
rect 20128 19768 20134 19780
rect 22640 19771 22698 19777
rect 20128 19740 22094 19768
rect 20128 19728 20134 19740
rect 19392 19672 19840 19700
rect 22066 19700 22094 19740
rect 22640 19737 22652 19771
rect 22686 19768 22698 19771
rect 22922 19768 22928 19780
rect 22686 19740 22928 19768
rect 22686 19737 22698 19740
rect 22640 19731 22698 19737
rect 22922 19728 22928 19740
rect 22980 19728 22986 19780
rect 24848 19771 24906 19777
rect 24848 19737 24860 19771
rect 24894 19737 24906 19771
rect 24848 19731 24906 19737
rect 23014 19700 23020 19712
rect 22066 19672 23020 19700
rect 19392 19660 19398 19672
rect 23014 19660 23020 19672
rect 23072 19660 23078 19712
rect 23750 19700 23756 19712
rect 23711 19672 23756 19700
rect 23750 19660 23756 19672
rect 23808 19660 23814 19712
rect 24762 19660 24768 19712
rect 24820 19700 24826 19712
rect 24872 19700 24900 19731
rect 25590 19728 25596 19780
rect 25648 19768 25654 19780
rect 26988 19768 27016 19799
rect 27890 19796 27896 19808
rect 27948 19796 27954 19848
rect 28169 19839 28227 19845
rect 28169 19805 28181 19839
rect 28215 19836 28227 19839
rect 29270 19836 29276 19848
rect 28215 19808 29276 19836
rect 28215 19805 28227 19808
rect 28169 19799 28227 19805
rect 29270 19796 29276 19808
rect 29328 19796 29334 19848
rect 29733 19839 29791 19845
rect 29733 19805 29745 19839
rect 29779 19836 29791 19839
rect 29822 19836 29828 19848
rect 29779 19808 29828 19836
rect 29779 19805 29791 19808
rect 29733 19799 29791 19805
rect 29822 19796 29828 19808
rect 29880 19796 29886 19848
rect 28353 19771 28411 19777
rect 28353 19768 28365 19771
rect 25648 19740 26648 19768
rect 26988 19740 28365 19768
rect 25648 19728 25654 19740
rect 25958 19700 25964 19712
rect 24820 19672 24900 19700
rect 25919 19672 25964 19700
rect 24820 19660 24826 19672
rect 25958 19660 25964 19672
rect 26016 19660 26022 19712
rect 26620 19700 26648 19740
rect 28353 19737 28365 19740
rect 28399 19737 28411 19771
rect 28810 19768 28816 19780
rect 28771 19740 28816 19768
rect 28353 19731 28411 19737
rect 28810 19728 28816 19740
rect 28868 19728 28874 19780
rect 28902 19728 28908 19780
rect 28960 19768 28966 19780
rect 28997 19771 29055 19777
rect 28997 19768 29009 19771
rect 28960 19740 29009 19768
rect 28960 19728 28966 19740
rect 28997 19737 29009 19740
rect 29043 19737 29055 19771
rect 28997 19731 29055 19737
rect 30000 19771 30058 19777
rect 30000 19737 30012 19771
rect 30046 19768 30058 19771
rect 30834 19768 30840 19780
rect 30046 19740 30840 19768
rect 30046 19737 30058 19740
rect 30000 19731 30058 19737
rect 30834 19728 30840 19740
rect 30892 19728 30898 19780
rect 31588 19777 31616 19876
rect 32493 19873 32505 19907
rect 32539 19904 32551 19907
rect 33410 19904 33416 19916
rect 32539 19876 33416 19904
rect 32539 19873 32551 19876
rect 32493 19867 32551 19873
rect 33410 19864 33416 19876
rect 33468 19864 33474 19916
rect 31754 19796 31760 19848
rect 31812 19836 31818 19848
rect 34330 19836 34336 19848
rect 31812 19808 32352 19836
rect 34291 19808 34336 19836
rect 31812 19796 31818 19808
rect 31573 19771 31631 19777
rect 31573 19737 31585 19771
rect 31619 19737 31631 19771
rect 32214 19768 32220 19780
rect 31573 19731 31631 19737
rect 31680 19740 32220 19768
rect 27706 19700 27712 19712
rect 26620 19672 27712 19700
rect 27706 19660 27712 19672
rect 27764 19660 27770 19712
rect 27798 19660 27804 19712
rect 27856 19700 27862 19712
rect 29086 19700 29092 19712
rect 27856 19672 29092 19700
rect 27856 19660 27862 19672
rect 29086 19660 29092 19672
rect 29144 19700 29150 19712
rect 30190 19700 30196 19712
rect 29144 19672 30196 19700
rect 29144 19660 29150 19672
rect 30190 19660 30196 19672
rect 30248 19700 30254 19712
rect 31113 19703 31171 19709
rect 31113 19700 31125 19703
rect 30248 19672 31125 19700
rect 30248 19660 30254 19672
rect 31113 19669 31125 19672
rect 31159 19669 31171 19703
rect 31113 19663 31171 19669
rect 31386 19660 31392 19712
rect 31444 19700 31450 19712
rect 31680 19700 31708 19740
rect 31444 19672 31708 19700
rect 31772 19709 31800 19740
rect 32214 19728 32220 19740
rect 32272 19728 32278 19780
rect 31772 19703 31831 19709
rect 31772 19672 31785 19703
rect 31444 19660 31450 19672
rect 31773 19669 31785 19672
rect 31819 19669 31831 19703
rect 31773 19663 31831 19669
rect 31941 19703 31999 19709
rect 31941 19669 31953 19703
rect 31987 19700 31999 19703
rect 32324 19700 32352 19808
rect 34330 19796 34336 19808
rect 34388 19796 34394 19848
rect 32677 19771 32735 19777
rect 32677 19737 32689 19771
rect 32723 19768 32735 19771
rect 32766 19768 32772 19780
rect 32723 19740 32772 19768
rect 32723 19737 32735 19740
rect 32677 19731 32735 19737
rect 32766 19728 32772 19740
rect 32824 19728 32830 19780
rect 32950 19728 32956 19780
rect 33008 19768 33014 19780
rect 33318 19768 33324 19780
rect 33008 19740 33324 19768
rect 33008 19728 33014 19740
rect 33318 19728 33324 19740
rect 33376 19728 33382 19780
rect 33042 19700 33048 19712
rect 31987 19672 33048 19700
rect 31987 19669 31999 19672
rect 31941 19663 31999 19669
rect 33042 19660 33048 19672
rect 33100 19660 33106 19712
rect 1104 19610 35027 19632
rect 1104 19558 9390 19610
rect 9442 19558 9454 19610
rect 9506 19558 9518 19610
rect 9570 19558 9582 19610
rect 9634 19558 9646 19610
rect 9698 19558 17831 19610
rect 17883 19558 17895 19610
rect 17947 19558 17959 19610
rect 18011 19558 18023 19610
rect 18075 19558 18087 19610
rect 18139 19558 26272 19610
rect 26324 19558 26336 19610
rect 26388 19558 26400 19610
rect 26452 19558 26464 19610
rect 26516 19558 26528 19610
rect 26580 19558 34713 19610
rect 34765 19558 34777 19610
rect 34829 19558 34841 19610
rect 34893 19558 34905 19610
rect 34957 19558 34969 19610
rect 35021 19558 35027 19610
rect 1104 19536 35027 19558
rect 15562 19496 15568 19508
rect 15304 19468 15568 19496
rect 1946 19428 1952 19440
rect 1907 19400 1952 19428
rect 1946 19388 1952 19400
rect 2004 19388 2010 19440
rect 15304 19369 15332 19468
rect 15562 19456 15568 19468
rect 15620 19456 15626 19508
rect 16022 19456 16028 19508
rect 16080 19496 16086 19508
rect 16301 19499 16359 19505
rect 16301 19496 16313 19499
rect 16080 19468 16313 19496
rect 16080 19456 16086 19468
rect 16301 19465 16313 19468
rect 16347 19465 16359 19499
rect 18598 19496 18604 19508
rect 18559 19468 18604 19496
rect 16301 19459 16359 19465
rect 18598 19456 18604 19468
rect 18656 19456 18662 19508
rect 19889 19499 19947 19505
rect 19889 19465 19901 19499
rect 19935 19496 19947 19499
rect 20438 19496 20444 19508
rect 19935 19468 20444 19496
rect 19935 19465 19947 19468
rect 19889 19459 19947 19465
rect 20438 19456 20444 19468
rect 20496 19456 20502 19508
rect 21450 19456 21456 19508
rect 21508 19496 21514 19508
rect 22462 19496 22468 19508
rect 21508 19468 22324 19496
rect 22423 19468 22468 19496
rect 21508 19456 21514 19468
rect 15381 19431 15439 19437
rect 15381 19397 15393 19431
rect 15427 19428 15439 19431
rect 16206 19428 16212 19440
rect 15427 19400 16212 19428
rect 15427 19397 15439 19400
rect 15381 19391 15439 19397
rect 16206 19388 16212 19400
rect 16264 19388 16270 19440
rect 22296 19428 22324 19468
rect 22462 19456 22468 19468
rect 22520 19456 22526 19508
rect 22922 19496 22928 19508
rect 22883 19468 22928 19496
rect 22922 19456 22928 19468
rect 22980 19456 22986 19508
rect 23658 19496 23664 19508
rect 23032 19468 23664 19496
rect 23032 19428 23060 19468
rect 23658 19456 23664 19468
rect 23716 19496 23722 19508
rect 24486 19496 24492 19508
rect 23716 19468 24492 19496
rect 23716 19456 23722 19468
rect 24486 19456 24492 19468
rect 24544 19456 24550 19508
rect 25958 19496 25964 19508
rect 24964 19468 25964 19496
rect 24964 19440 24992 19468
rect 25958 19456 25964 19468
rect 26016 19456 26022 19508
rect 26326 19456 26332 19508
rect 26384 19496 26390 19508
rect 27709 19499 27767 19505
rect 27709 19496 27721 19499
rect 26384 19468 27721 19496
rect 26384 19456 26390 19468
rect 27709 19465 27721 19468
rect 27755 19465 27767 19499
rect 27709 19459 27767 19465
rect 29089 19499 29147 19505
rect 29089 19465 29101 19499
rect 29135 19496 29147 19499
rect 30098 19496 30104 19508
rect 29135 19468 30104 19496
rect 29135 19465 29147 19468
rect 29089 19459 29147 19465
rect 30098 19456 30104 19468
rect 30156 19456 30162 19508
rect 31386 19456 31392 19508
rect 31444 19496 31450 19508
rect 31444 19468 32720 19496
rect 31444 19456 31450 19468
rect 19812 19400 21036 19428
rect 22296 19400 23060 19428
rect 15289 19363 15347 19369
rect 15289 19329 15301 19363
rect 15335 19329 15347 19363
rect 15289 19323 15347 19329
rect 15473 19363 15531 19369
rect 15473 19329 15485 19363
rect 15519 19329 15531 19363
rect 15473 19323 15531 19329
rect 1762 19292 1768 19304
rect 1723 19264 1768 19292
rect 1762 19252 1768 19264
rect 1820 19252 1826 19304
rect 2222 19292 2228 19304
rect 2183 19264 2228 19292
rect 2222 19252 2228 19264
rect 2280 19252 2286 19304
rect 15482 19292 15510 19323
rect 15562 19320 15568 19372
rect 15620 19360 15626 19372
rect 16117 19363 16175 19369
rect 16117 19360 16129 19363
rect 15620 19332 16129 19360
rect 15620 19320 15626 19332
rect 16117 19329 16129 19332
rect 16163 19360 16175 19363
rect 16574 19360 16580 19372
rect 16163 19332 16580 19360
rect 16163 19329 16175 19332
rect 16117 19323 16175 19329
rect 16574 19320 16580 19332
rect 16632 19320 16638 19372
rect 16666 19320 16672 19372
rect 16724 19360 16730 19372
rect 17037 19363 17095 19369
rect 17037 19360 17049 19363
rect 16724 19332 17049 19360
rect 16724 19320 16730 19332
rect 17037 19329 17049 19332
rect 17083 19329 17095 19363
rect 18414 19360 18420 19372
rect 18375 19332 18420 19360
rect 17037 19323 17095 19329
rect 18414 19320 18420 19332
rect 18472 19360 18478 19372
rect 19153 19363 19211 19369
rect 19153 19360 19165 19363
rect 18472 19332 19165 19360
rect 18472 19320 18478 19332
rect 19153 19329 19165 19332
rect 19199 19329 19211 19363
rect 19334 19360 19340 19372
rect 19295 19332 19340 19360
rect 19153 19323 19211 19329
rect 19334 19320 19340 19332
rect 19392 19320 19398 19372
rect 19812 19369 19840 19400
rect 19797 19363 19855 19369
rect 19797 19329 19809 19363
rect 19843 19329 19855 19363
rect 20622 19360 20628 19372
rect 20583 19332 20628 19360
rect 19797 19323 19855 19329
rect 20622 19320 20628 19332
rect 20680 19320 20686 19372
rect 20806 19360 20812 19372
rect 20767 19332 20812 19360
rect 20806 19320 20812 19332
rect 20864 19320 20870 19372
rect 20901 19363 20959 19369
rect 20901 19329 20913 19363
rect 20947 19329 20959 19363
rect 21008 19360 21036 19400
rect 23934 19388 23940 19440
rect 23992 19428 23998 19440
rect 24946 19428 24952 19440
rect 23992 19400 24256 19428
rect 24859 19400 24952 19428
rect 23992 19388 23998 19400
rect 24228 19372 24256 19400
rect 24946 19388 24952 19400
rect 25004 19388 25010 19440
rect 25038 19388 25044 19440
rect 25096 19428 25102 19440
rect 25149 19431 25207 19437
rect 25149 19428 25161 19431
rect 25096 19400 25161 19428
rect 25096 19388 25102 19400
rect 25149 19397 25161 19400
rect 25195 19397 25207 19431
rect 32306 19428 32312 19440
rect 25149 19391 25207 19397
rect 27172 19400 28028 19428
rect 22370 19360 22376 19372
rect 21008 19332 22376 19360
rect 20901 19323 20959 19329
rect 15933 19295 15991 19301
rect 15933 19292 15945 19295
rect 15482 19264 15945 19292
rect 15933 19261 15945 19264
rect 15979 19261 15991 19295
rect 16942 19292 16948 19304
rect 16903 19264 16948 19292
rect 15933 19255 15991 19261
rect 15948 19156 15976 19255
rect 16942 19252 16948 19264
rect 17000 19252 17006 19304
rect 17405 19227 17463 19233
rect 17405 19193 17417 19227
rect 17451 19224 17463 19227
rect 18322 19224 18328 19236
rect 17451 19196 18328 19224
rect 17451 19193 17463 19196
rect 17405 19187 17463 19193
rect 18322 19184 18328 19196
rect 18380 19184 18386 19236
rect 18690 19184 18696 19236
rect 18748 19224 18754 19236
rect 19153 19227 19211 19233
rect 19153 19224 19165 19227
rect 18748 19196 19165 19224
rect 18748 19184 18754 19196
rect 19153 19193 19165 19196
rect 19199 19193 19211 19227
rect 20916 19224 20944 19323
rect 22370 19320 22376 19332
rect 22428 19320 22434 19372
rect 23106 19360 23112 19372
rect 23067 19332 23112 19360
rect 23106 19320 23112 19332
rect 23164 19320 23170 19372
rect 23290 19320 23296 19372
rect 23348 19360 23354 19372
rect 24029 19363 24087 19369
rect 24029 19360 24041 19363
rect 23348 19332 24041 19360
rect 23348 19320 23354 19332
rect 24029 19329 24041 19332
rect 24075 19329 24087 19363
rect 24210 19360 24216 19372
rect 24171 19332 24216 19360
rect 24029 19323 24087 19329
rect 24210 19320 24216 19332
rect 24268 19320 24274 19372
rect 24854 19320 24860 19372
rect 24912 19360 24918 19372
rect 26050 19360 26056 19372
rect 24912 19332 26056 19360
rect 24912 19320 24918 19332
rect 26050 19320 26056 19332
rect 26108 19320 26114 19372
rect 26142 19320 26148 19372
rect 26200 19360 26206 19372
rect 26421 19363 26479 19369
rect 26200 19332 26245 19360
rect 26200 19320 26206 19332
rect 26421 19329 26433 19363
rect 26467 19360 26479 19363
rect 26786 19360 26792 19372
rect 26467 19332 26792 19360
rect 26467 19329 26479 19332
rect 26421 19323 26479 19329
rect 26786 19320 26792 19332
rect 26844 19360 26850 19372
rect 27172 19369 27200 19400
rect 27157 19363 27215 19369
rect 27157 19360 27169 19363
rect 26844 19332 27169 19360
rect 26844 19320 26850 19332
rect 27157 19329 27169 19332
rect 27203 19329 27215 19363
rect 27338 19360 27344 19372
rect 27299 19332 27344 19360
rect 27157 19323 27215 19329
rect 27338 19320 27344 19332
rect 27396 19320 27402 19372
rect 27433 19363 27491 19369
rect 27433 19329 27445 19363
rect 27479 19329 27491 19363
rect 27549 19363 27607 19369
rect 27549 19360 27561 19363
rect 27433 19323 27491 19329
rect 27540 19329 27561 19360
rect 27595 19329 27607 19363
rect 27798 19360 27804 19372
rect 27540 19323 27607 19329
rect 27724 19332 27804 19360
rect 21818 19252 21824 19304
rect 21876 19292 21882 19304
rect 22005 19295 22063 19301
rect 22005 19292 22017 19295
rect 21876 19264 22017 19292
rect 21876 19252 21882 19264
rect 22005 19261 22017 19264
rect 22051 19292 22063 19295
rect 23385 19295 23443 19301
rect 23385 19292 23397 19295
rect 22051 19264 23397 19292
rect 22051 19261 22063 19264
rect 22005 19255 22063 19261
rect 23385 19261 23397 19264
rect 23431 19292 23443 19295
rect 23750 19292 23756 19304
rect 23431 19264 23756 19292
rect 23431 19261 23443 19264
rect 23385 19255 23443 19261
rect 23750 19252 23756 19264
rect 23808 19292 23814 19304
rect 23845 19295 23903 19301
rect 23845 19292 23857 19295
rect 23808 19264 23857 19292
rect 23808 19252 23814 19264
rect 23845 19261 23857 19264
rect 23891 19261 23903 19295
rect 23845 19255 23903 19261
rect 25866 19252 25872 19304
rect 25924 19292 25930 19304
rect 26329 19295 26387 19301
rect 26329 19292 26341 19295
rect 25924 19264 26341 19292
rect 25924 19252 25930 19264
rect 26329 19261 26341 19264
rect 26375 19261 26387 19295
rect 26329 19255 26387 19261
rect 21266 19224 21272 19236
rect 20916 19196 21272 19224
rect 19153 19187 19211 19193
rect 21266 19184 21272 19196
rect 21324 19184 21330 19236
rect 22373 19227 22431 19233
rect 22373 19193 22385 19227
rect 22419 19224 22431 19227
rect 23014 19224 23020 19236
rect 22419 19196 23020 19224
rect 22419 19193 22431 19196
rect 22373 19187 22431 19193
rect 23014 19184 23020 19196
rect 23072 19184 23078 19236
rect 25774 19224 25780 19236
rect 25148 19196 25780 19224
rect 25148 19168 25176 19196
rect 25774 19184 25780 19196
rect 25832 19184 25838 19236
rect 18414 19156 18420 19168
rect 15948 19128 18420 19156
rect 18414 19116 18420 19128
rect 18472 19116 18478 19168
rect 20625 19159 20683 19165
rect 20625 19125 20637 19159
rect 20671 19156 20683 19159
rect 20714 19156 20720 19168
rect 20671 19128 20720 19156
rect 20671 19125 20683 19128
rect 20625 19119 20683 19125
rect 20714 19116 20720 19128
rect 20772 19116 20778 19168
rect 22646 19116 22652 19168
rect 22704 19156 22710 19168
rect 23290 19156 23296 19168
rect 22704 19128 23296 19156
rect 22704 19116 22710 19128
rect 23290 19116 23296 19128
rect 23348 19116 23354 19168
rect 25130 19156 25136 19168
rect 25043 19128 25136 19156
rect 25130 19116 25136 19128
rect 25188 19116 25194 19168
rect 25314 19156 25320 19168
rect 25275 19128 25320 19156
rect 25314 19116 25320 19128
rect 25372 19116 25378 19168
rect 25869 19159 25927 19165
rect 25869 19125 25881 19159
rect 25915 19156 25927 19159
rect 26142 19156 26148 19168
rect 25915 19128 26148 19156
rect 25915 19125 25927 19128
rect 25869 19119 25927 19125
rect 26142 19116 26148 19128
rect 26200 19116 26206 19168
rect 26344 19156 26372 19255
rect 27246 19252 27252 19304
rect 27304 19292 27310 19304
rect 27448 19292 27476 19323
rect 27540 19306 27592 19323
rect 27304 19264 27476 19292
rect 27304 19252 27310 19264
rect 26970 19184 26976 19236
rect 27028 19224 27034 19236
rect 27564 19224 27592 19306
rect 27724 19304 27752 19332
rect 27798 19320 27804 19332
rect 27856 19320 27862 19372
rect 27706 19252 27712 19304
rect 27764 19252 27770 19304
rect 28000 19292 28028 19400
rect 30392 19400 32312 19428
rect 28445 19363 28503 19369
rect 28445 19329 28457 19363
rect 28491 19360 28503 19363
rect 29270 19360 29276 19372
rect 28491 19332 29276 19360
rect 28491 19329 28503 19332
rect 28445 19323 28503 19329
rect 29270 19320 29276 19332
rect 29328 19320 29334 19372
rect 29362 19320 29368 19372
rect 29420 19360 29426 19372
rect 29549 19363 29607 19369
rect 29549 19360 29561 19363
rect 29420 19332 29561 19360
rect 29420 19320 29426 19332
rect 29549 19329 29561 19332
rect 29595 19329 29607 19363
rect 29549 19323 29607 19329
rect 28718 19292 28724 19304
rect 28000 19264 28724 19292
rect 28718 19252 28724 19264
rect 28776 19292 28782 19304
rect 28813 19295 28871 19301
rect 28813 19292 28825 19295
rect 28776 19264 28825 19292
rect 28776 19252 28782 19264
rect 28813 19261 28825 19264
rect 28859 19261 28871 19295
rect 28813 19255 28871 19261
rect 28905 19295 28963 19301
rect 28905 19261 28917 19295
rect 28951 19261 28963 19295
rect 28905 19255 28963 19261
rect 27028 19196 27592 19224
rect 27028 19184 27034 19196
rect 28350 19184 28356 19236
rect 28408 19224 28414 19236
rect 28920 19224 28948 19255
rect 29822 19252 29828 19304
rect 29880 19292 29886 19304
rect 30392 19301 30420 19400
rect 31772 19372 31800 19400
rect 32306 19388 32312 19400
rect 32364 19388 32370 19440
rect 32692 19437 32720 19468
rect 32677 19431 32735 19437
rect 32677 19397 32689 19431
rect 32723 19397 32735 19431
rect 32677 19391 32735 19397
rect 30644 19363 30702 19369
rect 30644 19329 30656 19363
rect 30690 19360 30702 19363
rect 31018 19360 31024 19372
rect 30690 19332 31024 19360
rect 30690 19329 30702 19332
rect 30644 19323 30702 19329
rect 31018 19320 31024 19332
rect 31076 19320 31082 19372
rect 31754 19320 31760 19372
rect 31812 19320 31818 19372
rect 32122 19320 32128 19372
rect 32180 19360 32186 19372
rect 32493 19363 32551 19369
rect 32493 19360 32505 19363
rect 32180 19332 32505 19360
rect 32180 19320 32186 19332
rect 32493 19329 32505 19332
rect 32539 19329 32551 19363
rect 32493 19323 32551 19329
rect 30377 19295 30435 19301
rect 30377 19292 30389 19295
rect 29880 19264 30389 19292
rect 29880 19252 29886 19264
rect 30377 19261 30389 19264
rect 30423 19261 30435 19295
rect 31938 19292 31944 19304
rect 30377 19255 30435 19261
rect 31772 19264 31944 19292
rect 31772 19233 31800 19264
rect 31938 19252 31944 19264
rect 31996 19292 32002 19304
rect 32306 19292 32312 19304
rect 31996 19264 32312 19292
rect 31996 19252 32002 19264
rect 32306 19252 32312 19264
rect 32364 19252 32370 19304
rect 34330 19292 34336 19304
rect 34291 19264 34336 19292
rect 34330 19252 34336 19264
rect 34388 19252 34394 19304
rect 28408 19196 28948 19224
rect 31757 19227 31815 19233
rect 28408 19184 28414 19196
rect 31757 19193 31769 19227
rect 31803 19193 31815 19227
rect 31757 19187 31815 19193
rect 27338 19156 27344 19168
rect 26344 19128 27344 19156
rect 27338 19116 27344 19128
rect 27396 19116 27402 19168
rect 29730 19156 29736 19168
rect 29691 19128 29736 19156
rect 29730 19116 29736 19128
rect 29788 19116 29794 19168
rect 30742 19116 30748 19168
rect 30800 19156 30806 19168
rect 31018 19156 31024 19168
rect 30800 19128 31024 19156
rect 30800 19116 30806 19128
rect 31018 19116 31024 19128
rect 31076 19116 31082 19168
rect 31110 19116 31116 19168
rect 31168 19156 31174 19168
rect 31938 19156 31944 19168
rect 31168 19128 31944 19156
rect 31168 19116 31174 19128
rect 31938 19116 31944 19128
rect 31996 19116 32002 19168
rect 1104 19066 34868 19088
rect 1104 19014 5170 19066
rect 5222 19014 5234 19066
rect 5286 19014 5298 19066
rect 5350 19014 5362 19066
rect 5414 19014 5426 19066
rect 5478 19014 13611 19066
rect 13663 19014 13675 19066
rect 13727 19014 13739 19066
rect 13791 19014 13803 19066
rect 13855 19014 13867 19066
rect 13919 19014 22052 19066
rect 22104 19014 22116 19066
rect 22168 19014 22180 19066
rect 22232 19014 22244 19066
rect 22296 19014 22308 19066
rect 22360 19014 30493 19066
rect 30545 19014 30557 19066
rect 30609 19014 30621 19066
rect 30673 19014 30685 19066
rect 30737 19014 30749 19066
rect 30801 19014 34868 19066
rect 1104 18992 34868 19014
rect 1762 18912 1768 18964
rect 1820 18952 1826 18964
rect 2041 18955 2099 18961
rect 2041 18952 2053 18955
rect 1820 18924 2053 18952
rect 1820 18912 1826 18924
rect 2041 18921 2053 18924
rect 2087 18921 2099 18955
rect 16942 18952 16948 18964
rect 16903 18924 16948 18952
rect 2041 18915 2099 18921
rect 16942 18912 16948 18924
rect 17000 18912 17006 18964
rect 17681 18955 17739 18961
rect 17681 18921 17693 18955
rect 17727 18952 17739 18955
rect 17727 18924 18736 18952
rect 17727 18921 17739 18924
rect 17681 18915 17739 18921
rect 16574 18844 16580 18896
rect 16632 18844 16638 18896
rect 2038 18776 2044 18828
rect 2096 18816 2102 18828
rect 2222 18816 2228 18828
rect 2096 18788 2228 18816
rect 2096 18776 2102 18788
rect 2222 18776 2228 18788
rect 2280 18776 2286 18828
rect 16592 18816 16620 18844
rect 16669 18819 16727 18825
rect 16669 18816 16681 18819
rect 16592 18788 16681 18816
rect 16669 18785 16681 18788
rect 16715 18785 16727 18819
rect 16669 18779 16727 18785
rect 1762 18708 1768 18760
rect 1820 18748 1826 18760
rect 2685 18751 2743 18757
rect 2685 18748 2697 18751
rect 1820 18720 2697 18748
rect 1820 18708 1826 18720
rect 2685 18717 2697 18720
rect 2731 18717 2743 18751
rect 2685 18711 2743 18717
rect 16577 18751 16635 18757
rect 16577 18717 16589 18751
rect 16623 18748 16635 18751
rect 16758 18748 16764 18760
rect 16623 18720 16764 18748
rect 16623 18717 16635 18720
rect 16577 18711 16635 18717
rect 16758 18708 16764 18720
rect 16816 18708 16822 18760
rect 17402 18708 17408 18760
rect 17460 18748 17466 18760
rect 17589 18751 17647 18757
rect 17589 18748 17601 18751
rect 17460 18720 17601 18748
rect 17460 18708 17466 18720
rect 17589 18717 17601 18720
rect 17635 18717 17647 18751
rect 17589 18711 17647 18717
rect 17773 18751 17831 18757
rect 17773 18717 17785 18751
rect 17819 18717 17831 18751
rect 17773 18711 17831 18717
rect 17788 18680 17816 18711
rect 18414 18708 18420 18760
rect 18472 18757 18478 18760
rect 18472 18751 18521 18757
rect 18472 18717 18475 18751
rect 18509 18717 18521 18751
rect 18598 18748 18604 18760
rect 18559 18720 18604 18748
rect 18472 18711 18521 18717
rect 18472 18708 18478 18711
rect 18598 18708 18604 18720
rect 18656 18708 18662 18760
rect 18708 18757 18736 18924
rect 19978 18912 19984 18964
rect 20036 18952 20042 18964
rect 20036 18924 20760 18952
rect 20036 18912 20042 18924
rect 20732 18884 20760 18924
rect 20806 18912 20812 18964
rect 20864 18952 20870 18964
rect 21085 18955 21143 18961
rect 21085 18952 21097 18955
rect 20864 18924 21097 18952
rect 20864 18912 20870 18924
rect 21085 18921 21097 18924
rect 21131 18952 21143 18955
rect 21358 18952 21364 18964
rect 21131 18924 21364 18952
rect 21131 18921 21143 18924
rect 21085 18915 21143 18921
rect 21358 18912 21364 18924
rect 21416 18952 21422 18964
rect 21729 18955 21787 18961
rect 21729 18952 21741 18955
rect 21416 18924 21741 18952
rect 21416 18912 21422 18924
rect 21729 18921 21741 18924
rect 21775 18921 21787 18955
rect 22554 18952 22560 18964
rect 22515 18924 22560 18952
rect 21729 18915 21787 18921
rect 22554 18912 22560 18924
rect 22612 18912 22618 18964
rect 22646 18912 22652 18964
rect 22704 18952 22710 18964
rect 22741 18955 22799 18961
rect 22741 18952 22753 18955
rect 22704 18924 22753 18952
rect 22704 18912 22710 18924
rect 22741 18921 22753 18924
rect 22787 18921 22799 18955
rect 25406 18952 25412 18964
rect 22741 18915 22799 18921
rect 23584 18924 25412 18952
rect 23584 18896 23612 18924
rect 25406 18912 25412 18924
rect 25464 18912 25470 18964
rect 28442 18912 28448 18964
rect 28500 18952 28506 18964
rect 29089 18955 29147 18961
rect 29089 18952 29101 18955
rect 28500 18924 29101 18952
rect 28500 18912 28506 18924
rect 29089 18921 29101 18924
rect 29135 18921 29147 18955
rect 29089 18915 29147 18921
rect 29454 18912 29460 18964
rect 29512 18952 29518 18964
rect 29733 18955 29791 18961
rect 29733 18952 29745 18955
rect 29512 18924 29745 18952
rect 29512 18912 29518 18924
rect 29733 18921 29745 18924
rect 29779 18921 29791 18955
rect 29733 18915 29791 18921
rect 30834 18912 30840 18964
rect 30892 18952 30898 18964
rect 32953 18955 33011 18961
rect 32953 18952 32965 18955
rect 30892 18924 32965 18952
rect 30892 18912 30898 18924
rect 32953 18921 32965 18924
rect 32999 18921 33011 18955
rect 33686 18952 33692 18964
rect 33647 18924 33692 18952
rect 32953 18915 33011 18921
rect 33686 18912 33692 18924
rect 33744 18912 33750 18964
rect 21174 18884 21180 18896
rect 20732 18856 21180 18884
rect 21174 18844 21180 18856
rect 21232 18884 21238 18896
rect 23566 18884 23572 18896
rect 21232 18856 23572 18884
rect 21232 18844 21238 18856
rect 23566 18844 23572 18856
rect 23624 18844 23630 18896
rect 23750 18884 23756 18896
rect 23711 18856 23756 18884
rect 23750 18844 23756 18856
rect 23808 18844 23814 18896
rect 24670 18844 24676 18896
rect 24728 18884 24734 18896
rect 24857 18887 24915 18893
rect 24857 18884 24869 18887
rect 24728 18856 24869 18884
rect 24728 18844 24734 18856
rect 24857 18853 24869 18856
rect 24903 18853 24915 18887
rect 24857 18847 24915 18853
rect 27246 18844 27252 18896
rect 27304 18844 27310 18896
rect 28718 18884 28724 18896
rect 28092 18856 28724 18884
rect 19426 18776 19432 18828
rect 19484 18816 19490 18828
rect 19705 18819 19763 18825
rect 19705 18816 19717 18819
rect 19484 18788 19717 18816
rect 19484 18776 19490 18788
rect 19705 18785 19717 18788
rect 19751 18785 19763 18819
rect 24946 18816 24952 18828
rect 19705 18779 19763 18785
rect 23768 18788 24952 18816
rect 18693 18751 18751 18757
rect 18693 18717 18705 18751
rect 18739 18717 18751 18751
rect 18874 18748 18880 18760
rect 18835 18720 18880 18748
rect 18693 18711 18751 18717
rect 18874 18708 18880 18720
rect 18932 18708 18938 18760
rect 20346 18708 20352 18760
rect 20404 18748 20410 18760
rect 23768 18757 23796 18788
rect 24946 18776 24952 18788
rect 25004 18776 25010 18828
rect 25777 18819 25835 18825
rect 25777 18785 25789 18819
rect 25823 18816 25835 18819
rect 26973 18819 27031 18825
rect 25823 18788 26740 18816
rect 25823 18785 25835 18788
rect 25777 18779 25835 18785
rect 23753 18751 23811 18757
rect 20404 18720 23704 18748
rect 20404 18708 20410 18720
rect 18616 18680 18644 18708
rect 17788 18652 18644 18680
rect 19972 18683 20030 18689
rect 19972 18649 19984 18683
rect 20018 18680 20030 18683
rect 20254 18680 20260 18692
rect 20018 18652 20260 18680
rect 20018 18649 20030 18652
rect 19972 18643 20030 18649
rect 20254 18640 20260 18652
rect 20312 18640 20318 18692
rect 21082 18640 21088 18692
rect 21140 18680 21146 18692
rect 21450 18680 21456 18692
rect 21140 18652 21456 18680
rect 21140 18640 21146 18652
rect 21450 18640 21456 18652
rect 21508 18680 21514 18692
rect 21545 18683 21603 18689
rect 21545 18680 21557 18683
rect 21508 18652 21557 18680
rect 21508 18640 21514 18652
rect 21545 18649 21557 18652
rect 21591 18649 21603 18683
rect 22370 18680 22376 18692
rect 22331 18652 22376 18680
rect 21545 18643 21603 18649
rect 22370 18640 22376 18652
rect 22428 18640 22434 18692
rect 23676 18680 23704 18720
rect 23753 18717 23765 18751
rect 23799 18717 23811 18751
rect 24029 18751 24087 18757
rect 24029 18748 24041 18751
rect 23753 18711 23811 18717
rect 23860 18720 24041 18748
rect 23860 18680 23888 18720
rect 24029 18717 24041 18720
rect 24075 18717 24087 18751
rect 25130 18748 25136 18760
rect 24029 18711 24087 18717
rect 24320 18720 25136 18748
rect 23676 18652 23888 18680
rect 18233 18615 18291 18621
rect 18233 18581 18245 18615
rect 18279 18612 18291 18615
rect 18506 18612 18512 18624
rect 18279 18584 18512 18612
rect 18279 18581 18291 18584
rect 18233 18575 18291 18581
rect 18506 18572 18512 18584
rect 18564 18572 18570 18624
rect 21266 18572 21272 18624
rect 21324 18612 21330 18624
rect 21634 18612 21640 18624
rect 21324 18584 21640 18612
rect 21324 18572 21330 18584
rect 21634 18572 21640 18584
rect 21692 18612 21698 18624
rect 21745 18615 21803 18621
rect 21745 18612 21757 18615
rect 21692 18584 21757 18612
rect 21692 18572 21698 18584
rect 21745 18581 21757 18584
rect 21791 18581 21803 18615
rect 21745 18575 21803 18581
rect 21913 18615 21971 18621
rect 21913 18581 21925 18615
rect 21959 18612 21971 18615
rect 22462 18612 22468 18624
rect 21959 18584 22468 18612
rect 21959 18581 21971 18584
rect 21913 18575 21971 18581
rect 22462 18572 22468 18584
rect 22520 18612 22526 18624
rect 22573 18615 22631 18621
rect 22573 18612 22585 18615
rect 22520 18584 22585 18612
rect 22520 18572 22526 18584
rect 22573 18581 22585 18584
rect 22619 18581 22631 18615
rect 23860 18612 23888 18652
rect 23937 18683 23995 18689
rect 23937 18649 23949 18683
rect 23983 18680 23995 18683
rect 24320 18680 24348 18720
rect 25130 18708 25136 18720
rect 25188 18708 25194 18760
rect 25961 18751 26019 18757
rect 25961 18717 25973 18751
rect 26007 18717 26019 18751
rect 26142 18748 26148 18760
rect 26103 18720 26148 18748
rect 25961 18711 26019 18717
rect 23983 18652 24348 18680
rect 23983 18649 23995 18652
rect 23937 18643 23995 18649
rect 24578 18640 24584 18692
rect 24636 18680 24642 18692
rect 24673 18683 24731 18689
rect 24673 18680 24685 18683
rect 24636 18652 24685 18680
rect 24636 18640 24642 18652
rect 24673 18649 24685 18652
rect 24719 18649 24731 18683
rect 25976 18680 26004 18711
rect 26142 18708 26148 18720
rect 26200 18708 26206 18760
rect 26237 18751 26295 18757
rect 26237 18717 26249 18751
rect 26283 18748 26295 18751
rect 26602 18748 26608 18760
rect 26283 18720 26608 18748
rect 26283 18717 26295 18720
rect 26237 18711 26295 18717
rect 26602 18708 26608 18720
rect 26660 18708 26666 18760
rect 26712 18757 26740 18788
rect 26973 18785 26985 18819
rect 27019 18816 27031 18819
rect 27264 18816 27292 18844
rect 27706 18816 27712 18828
rect 27019 18788 27712 18816
rect 27019 18785 27031 18788
rect 26973 18779 27031 18785
rect 27706 18776 27712 18788
rect 27764 18776 27770 18828
rect 26697 18751 26755 18757
rect 26697 18717 26709 18751
rect 26743 18717 26755 18751
rect 26697 18711 26755 18717
rect 26881 18751 26939 18757
rect 26881 18717 26893 18751
rect 26927 18717 26939 18751
rect 26881 18711 26939 18717
rect 27065 18751 27123 18757
rect 27065 18717 27077 18751
rect 27111 18748 27123 18751
rect 27154 18748 27160 18760
rect 27111 18720 27160 18748
rect 27111 18717 27123 18720
rect 27065 18711 27123 18717
rect 26326 18680 26332 18692
rect 25976 18652 26332 18680
rect 24673 18643 24731 18649
rect 26326 18640 26332 18652
rect 26384 18640 26390 18692
rect 26896 18680 26924 18711
rect 27154 18708 27160 18720
rect 27212 18708 27218 18760
rect 27249 18751 27307 18757
rect 27249 18717 27261 18751
rect 27295 18748 27307 18751
rect 27614 18748 27620 18760
rect 27295 18720 27620 18748
rect 27295 18717 27307 18720
rect 27249 18711 27307 18717
rect 27614 18708 27620 18720
rect 27672 18708 27678 18760
rect 28092 18757 28120 18856
rect 28718 18844 28724 18856
rect 28776 18884 28782 18896
rect 30101 18887 30159 18893
rect 30101 18884 30113 18887
rect 28776 18856 30113 18884
rect 28776 18844 28782 18856
rect 30101 18853 30113 18856
rect 30147 18853 30159 18887
rect 30101 18847 30159 18853
rect 32398 18844 32404 18896
rect 32456 18884 32462 18896
rect 32493 18887 32551 18893
rect 32493 18884 32505 18887
rect 32456 18856 32505 18884
rect 32456 18844 32462 18856
rect 32493 18853 32505 18856
rect 32539 18853 32551 18887
rect 32493 18847 32551 18853
rect 28169 18819 28227 18825
rect 28169 18785 28181 18819
rect 28215 18816 28227 18819
rect 28350 18816 28356 18828
rect 28215 18788 28356 18816
rect 28215 18785 28227 18788
rect 28169 18779 28227 18785
rect 28350 18776 28356 18788
rect 28408 18776 28414 18828
rect 28445 18819 28503 18825
rect 28445 18785 28457 18819
rect 28491 18816 28503 18819
rect 28810 18816 28816 18828
rect 28491 18788 28816 18816
rect 28491 18785 28503 18788
rect 28445 18779 28503 18785
rect 28810 18776 28816 18788
rect 28868 18816 28874 18828
rect 29086 18816 29092 18828
rect 28868 18788 29092 18816
rect 28868 18776 28874 18788
rect 29086 18776 29092 18788
rect 29144 18776 29150 18828
rect 29181 18819 29239 18825
rect 29181 18785 29193 18819
rect 29227 18785 29239 18819
rect 29181 18779 29239 18785
rect 28077 18751 28135 18757
rect 28077 18717 28089 18751
rect 28123 18717 28135 18751
rect 28077 18711 28135 18717
rect 28258 18708 28264 18760
rect 28316 18748 28322 18760
rect 28905 18751 28963 18757
rect 28905 18748 28917 18751
rect 28316 18720 28917 18748
rect 28316 18708 28322 18720
rect 28905 18717 28917 18720
rect 28951 18717 28963 18751
rect 28905 18711 28963 18717
rect 28994 18708 29000 18760
rect 29052 18748 29058 18760
rect 29052 18720 29097 18748
rect 29052 18708 29058 18720
rect 26970 18680 26976 18692
rect 26896 18652 26976 18680
rect 26970 18640 26976 18652
rect 27028 18640 27034 18692
rect 28534 18640 28540 18692
rect 28592 18680 28598 18692
rect 29196 18680 29224 18779
rect 29638 18776 29644 18828
rect 29696 18816 29702 18828
rect 30190 18816 30196 18828
rect 29696 18788 30196 18816
rect 29696 18776 29702 18788
rect 30190 18776 30196 18788
rect 30248 18776 30254 18828
rect 32674 18776 32680 18828
rect 32732 18816 32738 18828
rect 33781 18819 33839 18825
rect 33781 18816 33793 18819
rect 32732 18788 33793 18816
rect 32732 18776 32738 18788
rect 33781 18785 33793 18788
rect 33827 18785 33839 18819
rect 33781 18779 33839 18785
rect 29917 18751 29975 18757
rect 29917 18748 29929 18751
rect 28592 18652 29224 18680
rect 29288 18720 29929 18748
rect 28592 18640 28598 18652
rect 24946 18612 24952 18624
rect 23860 18584 24952 18612
rect 22573 18575 22631 18581
rect 24946 18572 24952 18584
rect 25004 18572 25010 18624
rect 27338 18572 27344 18624
rect 27396 18612 27402 18624
rect 27433 18615 27491 18621
rect 27433 18612 27445 18615
rect 27396 18584 27445 18612
rect 27396 18572 27402 18584
rect 27433 18581 27445 18584
rect 27479 18581 27491 18615
rect 27433 18575 27491 18581
rect 28350 18572 28356 18624
rect 28408 18612 28414 18624
rect 29288 18612 29316 18720
rect 29917 18717 29929 18720
rect 29963 18717 29975 18751
rect 29917 18711 29975 18717
rect 31113 18751 31171 18757
rect 31113 18717 31125 18751
rect 31159 18748 31171 18751
rect 31662 18748 31668 18760
rect 31159 18720 31668 18748
rect 31159 18717 31171 18720
rect 31113 18711 31171 18717
rect 31662 18708 31668 18720
rect 31720 18708 31726 18760
rect 31754 18708 31760 18760
rect 31812 18748 31818 18760
rect 33137 18751 33195 18757
rect 33137 18748 33149 18751
rect 31812 18720 33149 18748
rect 31812 18708 31818 18720
rect 33137 18717 33149 18720
rect 33183 18717 33195 18751
rect 33137 18711 33195 18717
rect 33226 18708 33232 18760
rect 33284 18748 33290 18760
rect 33689 18751 33747 18757
rect 33284 18720 33329 18748
rect 33284 18708 33290 18720
rect 33689 18717 33701 18751
rect 33735 18717 33747 18751
rect 33689 18711 33747 18717
rect 30834 18640 30840 18692
rect 30892 18680 30898 18692
rect 31358 18683 31416 18689
rect 31358 18680 31370 18683
rect 30892 18652 31370 18680
rect 30892 18640 30898 18652
rect 31358 18649 31370 18652
rect 31404 18649 31416 18683
rect 32953 18683 33011 18689
rect 32953 18680 32965 18683
rect 31358 18643 31416 18649
rect 31496 18652 32965 18680
rect 28408 18584 29316 18612
rect 28408 18572 28414 18584
rect 30282 18572 30288 18624
rect 30340 18612 30346 18624
rect 31496 18612 31524 18652
rect 32953 18649 32965 18652
rect 32999 18649 33011 18683
rect 32953 18643 33011 18649
rect 33042 18640 33048 18692
rect 33100 18680 33106 18692
rect 33704 18680 33732 18711
rect 33100 18652 33732 18680
rect 33965 18683 34023 18689
rect 33100 18640 33106 18652
rect 33965 18649 33977 18683
rect 34011 18649 34023 18683
rect 33965 18643 34023 18649
rect 30340 18584 31524 18612
rect 30340 18572 30346 18584
rect 33686 18572 33692 18624
rect 33744 18612 33750 18624
rect 33980 18612 34008 18643
rect 33744 18584 34008 18612
rect 33744 18572 33750 18584
rect 1104 18522 35027 18544
rect 1104 18470 9390 18522
rect 9442 18470 9454 18522
rect 9506 18470 9518 18522
rect 9570 18470 9582 18522
rect 9634 18470 9646 18522
rect 9698 18470 17831 18522
rect 17883 18470 17895 18522
rect 17947 18470 17959 18522
rect 18011 18470 18023 18522
rect 18075 18470 18087 18522
rect 18139 18470 26272 18522
rect 26324 18470 26336 18522
rect 26388 18470 26400 18522
rect 26452 18470 26464 18522
rect 26516 18470 26528 18522
rect 26580 18470 34713 18522
rect 34765 18470 34777 18522
rect 34829 18470 34841 18522
rect 34893 18470 34905 18522
rect 34957 18470 34969 18522
rect 35021 18470 35027 18522
rect 1104 18448 35027 18470
rect 17402 18408 17408 18420
rect 17363 18380 17408 18408
rect 17402 18368 17408 18380
rect 17460 18368 17466 18420
rect 18414 18368 18420 18420
rect 18472 18408 18478 18420
rect 19794 18408 19800 18420
rect 18472 18380 19800 18408
rect 18472 18368 18478 18380
rect 19794 18368 19800 18380
rect 19852 18368 19858 18420
rect 20254 18408 20260 18420
rect 20215 18380 20260 18408
rect 20254 18368 20260 18380
rect 20312 18368 20318 18420
rect 21358 18408 21364 18420
rect 20732 18380 21364 18408
rect 19426 18340 19432 18352
rect 18432 18312 19432 18340
rect 1762 18272 1768 18284
rect 1723 18244 1768 18272
rect 1762 18232 1768 18244
rect 1820 18232 1826 18284
rect 17034 18272 17040 18284
rect 16995 18244 17040 18272
rect 17034 18232 17040 18244
rect 17092 18232 17098 18284
rect 18432 18281 18460 18312
rect 19426 18300 19432 18312
rect 19484 18300 19490 18352
rect 18417 18275 18475 18281
rect 18417 18241 18429 18275
rect 18463 18241 18475 18275
rect 18417 18235 18475 18241
rect 18506 18232 18512 18284
rect 18564 18272 18570 18284
rect 20732 18281 20760 18380
rect 21358 18368 21364 18380
rect 21416 18368 21422 18420
rect 24946 18368 24952 18420
rect 25004 18408 25010 18420
rect 26602 18408 26608 18420
rect 25004 18380 26608 18408
rect 25004 18368 25010 18380
rect 26602 18368 26608 18380
rect 26660 18408 26666 18420
rect 27982 18408 27988 18420
rect 26660 18380 27752 18408
rect 27943 18380 27988 18408
rect 26660 18368 26666 18380
rect 21174 18340 21180 18352
rect 21135 18312 21180 18340
rect 21174 18300 21180 18312
rect 21232 18300 21238 18352
rect 27246 18300 27252 18352
rect 27304 18340 27310 18352
rect 27617 18343 27675 18349
rect 27617 18340 27629 18343
rect 27304 18312 27629 18340
rect 27304 18300 27310 18312
rect 27617 18309 27629 18312
rect 27663 18309 27675 18343
rect 27724 18340 27752 18380
rect 27982 18368 27988 18380
rect 28040 18368 28046 18420
rect 31294 18368 31300 18420
rect 31352 18408 31358 18420
rect 31352 18380 31754 18408
rect 31352 18368 31358 18380
rect 28994 18340 29000 18352
rect 27724 18312 29000 18340
rect 27617 18303 27675 18309
rect 28994 18300 29000 18312
rect 29052 18300 29058 18352
rect 30926 18340 30932 18352
rect 30300 18312 30932 18340
rect 18673 18275 18731 18281
rect 18673 18272 18685 18275
rect 18564 18244 18685 18272
rect 18564 18232 18570 18244
rect 18673 18241 18685 18244
rect 18719 18241 18731 18275
rect 18673 18235 18731 18241
rect 20441 18275 20499 18281
rect 20441 18241 20453 18275
rect 20487 18241 20499 18275
rect 20441 18235 20499 18241
rect 20717 18275 20775 18281
rect 20717 18241 20729 18275
rect 20763 18241 20775 18275
rect 20717 18235 20775 18241
rect 21453 18278 21511 18281
rect 21453 18275 21588 18278
rect 21453 18241 21465 18275
rect 21499 18272 21588 18275
rect 21634 18272 21640 18284
rect 21499 18250 21640 18272
rect 21499 18241 21511 18250
rect 21560 18244 21640 18250
rect 21453 18235 21511 18241
rect 1946 18204 1952 18216
rect 1907 18176 1952 18204
rect 1946 18164 1952 18176
rect 2004 18164 2010 18216
rect 2774 18204 2780 18216
rect 2735 18176 2780 18204
rect 2774 18164 2780 18176
rect 2832 18164 2838 18216
rect 17126 18204 17132 18216
rect 17087 18176 17132 18204
rect 17126 18164 17132 18176
rect 17184 18164 17190 18216
rect 20456 18136 20484 18235
rect 21634 18232 21640 18244
rect 21692 18232 21698 18284
rect 22272 18275 22330 18281
rect 22272 18241 22284 18275
rect 22318 18272 22330 18275
rect 22830 18272 22836 18284
rect 22318 18244 22836 18272
rect 22318 18241 22330 18244
rect 22272 18235 22330 18241
rect 22830 18232 22836 18244
rect 22888 18232 22894 18284
rect 23842 18272 23848 18284
rect 23803 18244 23848 18272
rect 23842 18232 23848 18244
rect 23900 18232 23906 18284
rect 23934 18232 23940 18284
rect 23992 18272 23998 18284
rect 24101 18275 24159 18281
rect 24101 18272 24113 18275
rect 23992 18244 24113 18272
rect 23992 18232 23998 18244
rect 24101 18241 24113 18244
rect 24147 18241 24159 18275
rect 24101 18235 24159 18241
rect 24578 18232 24584 18284
rect 24636 18272 24642 18284
rect 25314 18272 25320 18284
rect 24636 18244 25320 18272
rect 24636 18232 24642 18244
rect 25314 18232 25320 18244
rect 25372 18272 25378 18284
rect 25869 18275 25927 18281
rect 25869 18272 25881 18275
rect 25372 18244 25881 18272
rect 25372 18232 25378 18244
rect 25869 18241 25881 18244
rect 25915 18241 25927 18275
rect 27338 18272 27344 18284
rect 27299 18244 27344 18272
rect 25869 18235 25927 18241
rect 27338 18232 27344 18244
rect 27396 18232 27402 18284
rect 27489 18275 27547 18281
rect 27489 18241 27501 18275
rect 27535 18272 27547 18275
rect 27706 18272 27712 18284
rect 27535 18241 27568 18272
rect 27667 18244 27712 18272
rect 27489 18235 27568 18241
rect 20625 18207 20683 18213
rect 20625 18173 20637 18207
rect 20671 18204 20683 18207
rect 20806 18204 20812 18216
rect 20671 18176 20812 18204
rect 20671 18173 20683 18176
rect 20625 18167 20683 18173
rect 20806 18164 20812 18176
rect 20864 18204 20870 18216
rect 21266 18204 21272 18216
rect 20864 18176 21272 18204
rect 20864 18164 20870 18176
rect 21266 18164 21272 18176
rect 21324 18164 21330 18216
rect 21542 18164 21548 18216
rect 21600 18204 21606 18216
rect 21910 18204 21916 18216
rect 21600 18176 21916 18204
rect 21600 18164 21606 18176
rect 21910 18164 21916 18176
rect 21968 18204 21974 18216
rect 22005 18207 22063 18213
rect 22005 18204 22017 18207
rect 21968 18176 22017 18204
rect 21968 18164 21974 18176
rect 22005 18173 22017 18176
rect 22051 18173 22063 18207
rect 25685 18207 25743 18213
rect 25685 18204 25697 18207
rect 22005 18167 22063 18173
rect 25240 18176 25697 18204
rect 21177 18139 21235 18145
rect 21177 18136 21189 18139
rect 20456 18108 21189 18136
rect 21177 18105 21189 18108
rect 21223 18105 21235 18139
rect 21177 18099 21235 18105
rect 25130 18096 25136 18148
rect 25188 18136 25194 18148
rect 25240 18145 25268 18176
rect 25685 18173 25697 18176
rect 25731 18173 25743 18207
rect 27540 18204 27568 18235
rect 27706 18232 27712 18244
rect 27764 18232 27770 18284
rect 27847 18275 27905 18281
rect 27847 18241 27859 18275
rect 27893 18272 27905 18275
rect 28074 18272 28080 18284
rect 27893 18244 28080 18272
rect 27893 18241 27905 18244
rect 27847 18235 27905 18241
rect 28074 18232 28080 18244
rect 28132 18232 28138 18284
rect 28350 18232 28356 18284
rect 28408 18272 28414 18284
rect 28701 18275 28759 18281
rect 28701 18272 28713 18275
rect 28408 18244 28713 18272
rect 28408 18232 28414 18244
rect 28701 18241 28713 18244
rect 28747 18241 28759 18275
rect 28701 18235 28759 18241
rect 30190 18232 30196 18284
rect 30248 18272 30254 18284
rect 30300 18281 30328 18312
rect 30926 18300 30932 18312
rect 30984 18300 30990 18352
rect 31110 18300 31116 18352
rect 31168 18340 31174 18352
rect 31726 18340 31754 18380
rect 32398 18368 32404 18420
rect 32456 18408 32462 18420
rect 32456 18380 32720 18408
rect 32456 18368 32462 18380
rect 32309 18343 32367 18349
rect 32309 18340 32321 18343
rect 31168 18312 31616 18340
rect 31726 18312 32321 18340
rect 31168 18300 31174 18312
rect 30285 18275 30343 18281
rect 30285 18272 30297 18275
rect 30248 18244 30297 18272
rect 30248 18232 30254 18244
rect 30285 18241 30297 18244
rect 30331 18241 30343 18275
rect 30285 18235 30343 18241
rect 30377 18275 30435 18281
rect 30377 18241 30389 18275
rect 30423 18272 30435 18275
rect 30423 18244 31064 18272
rect 30423 18241 30435 18244
rect 30377 18235 30435 18241
rect 27614 18204 27620 18216
rect 27527 18176 27620 18204
rect 25685 18167 25743 18173
rect 27614 18164 27620 18176
rect 27672 18204 27678 18216
rect 28258 18204 28264 18216
rect 27672 18176 28264 18204
rect 27672 18164 27678 18176
rect 28258 18164 28264 18176
rect 28316 18164 28322 18216
rect 28442 18204 28448 18216
rect 28403 18176 28448 18204
rect 28442 18164 28448 18176
rect 28500 18164 28506 18216
rect 30561 18207 30619 18213
rect 30561 18173 30573 18207
rect 30607 18204 30619 18207
rect 30926 18204 30932 18216
rect 30607 18176 30932 18204
rect 30607 18173 30619 18176
rect 30561 18167 30619 18173
rect 30926 18164 30932 18176
rect 30984 18164 30990 18216
rect 31036 18204 31064 18244
rect 31294 18232 31300 18284
rect 31352 18272 31358 18284
rect 31481 18275 31539 18281
rect 31481 18272 31493 18275
rect 31352 18244 31493 18272
rect 31352 18232 31358 18244
rect 31481 18241 31493 18244
rect 31527 18241 31539 18275
rect 31588 18272 31616 18312
rect 32309 18309 32321 18312
rect 32355 18309 32367 18343
rect 32490 18340 32496 18352
rect 32451 18312 32496 18340
rect 32309 18303 32367 18309
rect 32490 18300 32496 18312
rect 32548 18300 32554 18352
rect 31665 18275 31723 18281
rect 31665 18272 31677 18275
rect 31588 18244 31677 18272
rect 31481 18235 31539 18241
rect 31665 18241 31677 18244
rect 31711 18241 31723 18275
rect 31665 18235 31723 18241
rect 31757 18275 31815 18281
rect 31757 18241 31769 18275
rect 31803 18272 31815 18275
rect 31938 18272 31944 18284
rect 31803 18244 31944 18272
rect 31803 18241 31815 18244
rect 31757 18235 31815 18241
rect 31938 18232 31944 18244
rect 31996 18232 32002 18284
rect 32585 18275 32643 18281
rect 32585 18241 32597 18275
rect 32631 18272 32643 18275
rect 32692 18272 32720 18380
rect 32950 18368 32956 18420
rect 33008 18408 33014 18420
rect 33045 18411 33103 18417
rect 33045 18408 33057 18411
rect 33008 18380 33057 18408
rect 33008 18368 33014 18380
rect 33045 18377 33057 18380
rect 33091 18377 33103 18411
rect 33045 18371 33103 18377
rect 33321 18343 33379 18349
rect 33321 18309 33333 18343
rect 33367 18340 33379 18343
rect 33686 18340 33692 18352
rect 33367 18312 33692 18340
rect 33367 18309 33379 18312
rect 33321 18303 33379 18309
rect 33686 18300 33692 18312
rect 33744 18300 33750 18352
rect 32631 18244 32720 18272
rect 32631 18241 32643 18244
rect 32585 18235 32643 18241
rect 32858 18232 32864 18284
rect 32916 18272 32922 18284
rect 33045 18275 33103 18281
rect 33045 18272 33057 18275
rect 32916 18244 33057 18272
rect 32916 18232 32922 18244
rect 33045 18241 33057 18244
rect 33091 18272 33103 18275
rect 33091 18244 33364 18272
rect 33091 18241 33103 18244
rect 33045 18235 33103 18241
rect 31846 18204 31852 18216
rect 31036 18176 31852 18204
rect 31846 18164 31852 18176
rect 31904 18164 31910 18216
rect 33226 18204 33232 18216
rect 31956 18176 33232 18204
rect 25225 18139 25283 18145
rect 25225 18136 25237 18139
rect 25188 18108 25237 18136
rect 25188 18096 25194 18108
rect 25225 18105 25237 18108
rect 25271 18105 25283 18139
rect 25225 18099 25283 18105
rect 30469 18139 30527 18145
rect 30469 18105 30481 18139
rect 30515 18136 30527 18139
rect 31956 18136 31984 18176
rect 33226 18164 33232 18176
rect 33284 18164 33290 18216
rect 33336 18204 33364 18244
rect 33594 18232 33600 18284
rect 33652 18272 33658 18284
rect 33781 18275 33839 18281
rect 33781 18272 33793 18275
rect 33652 18244 33793 18272
rect 33652 18232 33658 18244
rect 33781 18241 33793 18244
rect 33827 18241 33839 18275
rect 33781 18235 33839 18241
rect 33873 18207 33931 18213
rect 33873 18204 33885 18207
rect 33336 18176 33885 18204
rect 33873 18173 33885 18176
rect 33919 18173 33931 18207
rect 33873 18167 33931 18173
rect 34057 18207 34115 18213
rect 34057 18173 34069 18207
rect 34103 18173 34115 18207
rect 34057 18167 34115 18173
rect 30515 18108 31984 18136
rect 32309 18139 32367 18145
rect 30515 18105 30527 18108
rect 30469 18099 30527 18105
rect 32309 18105 32321 18139
rect 32355 18136 32367 18139
rect 33137 18139 33195 18145
rect 33137 18136 33149 18139
rect 32355 18108 33149 18136
rect 32355 18105 32367 18108
rect 32309 18099 32367 18105
rect 33137 18105 33149 18108
rect 33183 18105 33195 18139
rect 34072 18136 34100 18167
rect 33137 18099 33195 18105
rect 33244 18108 34100 18136
rect 22370 18028 22376 18080
rect 22428 18068 22434 18080
rect 23385 18071 23443 18077
rect 23385 18068 23397 18071
rect 22428 18040 23397 18068
rect 22428 18028 22434 18040
rect 23385 18037 23397 18040
rect 23431 18037 23443 18071
rect 26050 18068 26056 18080
rect 26011 18040 26056 18068
rect 23385 18031 23443 18037
rect 26050 18028 26056 18040
rect 26108 18028 26114 18080
rect 28258 18028 28264 18080
rect 28316 18068 28322 18080
rect 29825 18071 29883 18077
rect 29825 18068 29837 18071
rect 28316 18040 29837 18068
rect 28316 18028 28322 18040
rect 29825 18037 29837 18040
rect 29871 18037 29883 18071
rect 31478 18068 31484 18080
rect 31439 18040 31484 18068
rect 29825 18031 29883 18037
rect 31478 18028 31484 18040
rect 31536 18028 31542 18080
rect 31846 18028 31852 18080
rect 31904 18068 31910 18080
rect 33244 18068 33272 18108
rect 31904 18040 33272 18068
rect 31904 18028 31910 18040
rect 33962 18028 33968 18080
rect 34020 18068 34026 18080
rect 34020 18040 34065 18068
rect 34020 18028 34026 18040
rect 1104 17978 34868 18000
rect 1104 17926 5170 17978
rect 5222 17926 5234 17978
rect 5286 17926 5298 17978
rect 5350 17926 5362 17978
rect 5414 17926 5426 17978
rect 5478 17926 13611 17978
rect 13663 17926 13675 17978
rect 13727 17926 13739 17978
rect 13791 17926 13803 17978
rect 13855 17926 13867 17978
rect 13919 17926 22052 17978
rect 22104 17926 22116 17978
rect 22168 17926 22180 17978
rect 22232 17926 22244 17978
rect 22296 17926 22308 17978
rect 22360 17926 30493 17978
rect 30545 17926 30557 17978
rect 30609 17926 30621 17978
rect 30673 17926 30685 17978
rect 30737 17926 30749 17978
rect 30801 17926 34868 17978
rect 1104 17904 34868 17926
rect 1946 17824 1952 17876
rect 2004 17864 2010 17876
rect 2133 17867 2191 17873
rect 2133 17864 2145 17867
rect 2004 17836 2145 17864
rect 2004 17824 2010 17836
rect 2133 17833 2145 17836
rect 2179 17833 2191 17867
rect 20806 17864 20812 17876
rect 20767 17836 20812 17864
rect 2133 17827 2191 17833
rect 20806 17824 20812 17836
rect 20864 17824 20870 17876
rect 23845 17867 23903 17873
rect 23845 17833 23857 17867
rect 23891 17864 23903 17867
rect 26050 17864 26056 17876
rect 23891 17836 26056 17864
rect 23891 17833 23903 17836
rect 23845 17827 23903 17833
rect 26050 17824 26056 17836
rect 26108 17824 26114 17876
rect 28350 17864 28356 17876
rect 28311 17836 28356 17864
rect 28350 17824 28356 17836
rect 28408 17824 28414 17876
rect 28442 17824 28448 17876
rect 28500 17864 28506 17876
rect 29822 17864 29828 17876
rect 28500 17836 29828 17864
rect 28500 17824 28506 17836
rect 29822 17824 29828 17836
rect 29880 17824 29886 17876
rect 31202 17824 31208 17876
rect 31260 17864 31266 17876
rect 31665 17867 31723 17873
rect 31665 17864 31677 17867
rect 31260 17836 31677 17864
rect 31260 17824 31266 17836
rect 31665 17833 31677 17836
rect 31711 17833 31723 17867
rect 31665 17827 31723 17833
rect 29454 17796 29460 17808
rect 28736 17768 29460 17796
rect 19426 17728 19432 17740
rect 19387 17700 19432 17728
rect 19426 17688 19432 17700
rect 19484 17688 19490 17740
rect 2041 17663 2099 17669
rect 2041 17629 2053 17663
rect 2087 17660 2099 17663
rect 2130 17660 2136 17672
rect 2087 17632 2136 17660
rect 2087 17629 2099 17632
rect 2041 17623 2099 17629
rect 2130 17620 2136 17632
rect 2188 17620 2194 17672
rect 19444 17660 19472 17688
rect 21542 17660 21548 17672
rect 19444 17632 21548 17660
rect 21542 17620 21548 17632
rect 21600 17620 21606 17672
rect 23658 17660 23664 17672
rect 23619 17632 23664 17660
rect 23658 17620 23664 17632
rect 23716 17620 23722 17672
rect 23937 17663 23995 17669
rect 23937 17629 23949 17663
rect 23983 17629 23995 17663
rect 23937 17623 23995 17629
rect 24581 17663 24639 17669
rect 24581 17629 24593 17663
rect 24627 17660 24639 17663
rect 26421 17663 26479 17669
rect 26421 17660 26433 17663
rect 24627 17632 26433 17660
rect 24627 17629 24639 17632
rect 24581 17623 24639 17629
rect 26421 17629 26433 17632
rect 26467 17660 26479 17663
rect 27154 17660 27160 17672
rect 26467 17632 27160 17660
rect 26467 17629 26479 17632
rect 26421 17623 26479 17629
rect 19334 17552 19340 17604
rect 19392 17592 19398 17604
rect 19674 17595 19732 17601
rect 19674 17592 19686 17595
rect 19392 17564 19686 17592
rect 19392 17552 19398 17564
rect 19674 17561 19686 17564
rect 19720 17561 19732 17595
rect 19674 17555 19732 17561
rect 21634 17552 21640 17604
rect 21692 17592 21698 17604
rect 21790 17595 21848 17601
rect 21790 17592 21802 17595
rect 21692 17564 21802 17592
rect 21692 17552 21698 17564
rect 21790 17561 21802 17564
rect 21836 17561 21848 17595
rect 21790 17555 21848 17561
rect 22554 17484 22560 17536
rect 22612 17524 22618 17536
rect 22925 17527 22983 17533
rect 22925 17524 22937 17527
rect 22612 17496 22937 17524
rect 22612 17484 22618 17496
rect 22925 17493 22937 17496
rect 22971 17493 22983 17527
rect 23474 17524 23480 17536
rect 23435 17496 23480 17524
rect 22925 17487 22983 17493
rect 23474 17484 23480 17496
rect 23532 17484 23538 17536
rect 23952 17524 23980 17623
rect 27154 17620 27160 17632
rect 27212 17660 27218 17672
rect 28442 17660 28448 17672
rect 27212 17632 28448 17660
rect 27212 17620 27218 17632
rect 28442 17620 28448 17632
rect 28500 17620 28506 17672
rect 28736 17669 28764 17768
rect 29454 17756 29460 17768
rect 29512 17796 29518 17808
rect 29730 17796 29736 17808
rect 29512 17768 29736 17796
rect 29512 17756 29518 17768
rect 29730 17756 29736 17768
rect 29788 17756 29794 17808
rect 29840 17737 29868 17824
rect 30926 17756 30932 17808
rect 30984 17796 30990 17808
rect 31846 17796 31852 17808
rect 30984 17768 31852 17796
rect 30984 17756 30990 17768
rect 31846 17756 31852 17768
rect 31904 17756 31910 17808
rect 29825 17731 29883 17737
rect 29825 17697 29837 17731
rect 29871 17697 29883 17731
rect 29825 17691 29883 17697
rect 31018 17688 31024 17740
rect 31076 17728 31082 17740
rect 32677 17731 32735 17737
rect 32677 17728 32689 17731
rect 31076 17700 32689 17728
rect 31076 17688 31082 17700
rect 32677 17697 32689 17700
rect 32723 17697 32735 17731
rect 34330 17728 34336 17740
rect 34291 17700 34336 17728
rect 32677 17691 32735 17697
rect 34330 17688 34336 17700
rect 34388 17688 34394 17740
rect 28629 17663 28687 17669
rect 28629 17629 28641 17663
rect 28675 17629 28687 17663
rect 28629 17623 28687 17629
rect 28721 17663 28779 17669
rect 28721 17629 28733 17663
rect 28767 17629 28779 17663
rect 28721 17623 28779 17629
rect 28813 17663 28871 17669
rect 28813 17629 28825 17663
rect 28859 17660 28871 17663
rect 28902 17660 28908 17672
rect 28859 17632 28908 17660
rect 28859 17629 28871 17632
rect 28813 17623 28871 17629
rect 24848 17595 24906 17601
rect 24848 17561 24860 17595
rect 24894 17592 24906 17595
rect 25314 17592 25320 17604
rect 24894 17564 25320 17592
rect 24894 17561 24906 17564
rect 24848 17555 24906 17561
rect 25314 17552 25320 17564
rect 25372 17552 25378 17604
rect 26694 17601 26700 17604
rect 26688 17555 26700 17601
rect 26752 17592 26758 17604
rect 26752 17564 26788 17592
rect 26694 17552 26700 17555
rect 26752 17552 26758 17564
rect 28258 17552 28264 17604
rect 28316 17592 28322 17604
rect 28644 17592 28672 17623
rect 28902 17620 28908 17632
rect 28960 17620 28966 17672
rect 28997 17663 29055 17669
rect 28997 17629 29009 17663
rect 29043 17629 29055 17663
rect 28997 17623 29055 17629
rect 28316 17564 28672 17592
rect 28316 17552 28322 17564
rect 24946 17524 24952 17536
rect 23952 17496 24952 17524
rect 24946 17484 24952 17496
rect 25004 17484 25010 17536
rect 25682 17484 25688 17536
rect 25740 17524 25746 17536
rect 25961 17527 26019 17533
rect 25961 17524 25973 17527
rect 25740 17496 25973 17524
rect 25740 17484 25746 17496
rect 25961 17493 25973 17496
rect 26007 17493 26019 17527
rect 25961 17487 26019 17493
rect 26142 17484 26148 17536
rect 26200 17524 26206 17536
rect 27801 17527 27859 17533
rect 27801 17524 27813 17527
rect 26200 17496 27813 17524
rect 26200 17484 26206 17496
rect 27801 17493 27813 17496
rect 27847 17493 27859 17527
rect 27801 17487 27859 17493
rect 27890 17484 27896 17536
rect 27948 17524 27954 17536
rect 29012 17524 29040 17623
rect 31202 17620 31208 17672
rect 31260 17660 31266 17672
rect 31665 17663 31723 17669
rect 31665 17660 31677 17663
rect 31260 17632 31677 17660
rect 31260 17620 31266 17632
rect 31665 17629 31677 17632
rect 31711 17629 31723 17663
rect 31665 17623 31723 17629
rect 31846 17620 31852 17672
rect 31904 17660 31910 17672
rect 31941 17663 31999 17669
rect 31941 17660 31953 17663
rect 31904 17632 31953 17660
rect 31904 17620 31910 17632
rect 31941 17629 31953 17632
rect 31987 17660 31999 17663
rect 32214 17660 32220 17672
rect 31987 17632 32220 17660
rect 31987 17629 31999 17632
rect 31941 17623 31999 17629
rect 32214 17620 32220 17632
rect 32272 17620 32278 17672
rect 32493 17663 32551 17669
rect 32493 17629 32505 17663
rect 32539 17629 32551 17663
rect 32493 17623 32551 17629
rect 29730 17552 29736 17604
rect 29788 17592 29794 17604
rect 30070 17595 30128 17601
rect 30070 17592 30082 17595
rect 29788 17564 30082 17592
rect 29788 17552 29794 17564
rect 30070 17561 30082 17564
rect 30116 17561 30128 17595
rect 32508 17592 32536 17623
rect 33226 17592 33232 17604
rect 32508 17564 33232 17592
rect 30070 17555 30128 17561
rect 33226 17552 33232 17564
rect 33284 17552 33290 17604
rect 27948 17496 29040 17524
rect 27948 17484 27954 17496
rect 30650 17484 30656 17536
rect 30708 17524 30714 17536
rect 31205 17527 31263 17533
rect 31205 17524 31217 17527
rect 30708 17496 31217 17524
rect 30708 17484 30714 17496
rect 31205 17493 31217 17496
rect 31251 17493 31263 17527
rect 31205 17487 31263 17493
rect 31849 17527 31907 17533
rect 31849 17493 31861 17527
rect 31895 17524 31907 17527
rect 32214 17524 32220 17536
rect 31895 17496 32220 17524
rect 31895 17493 31907 17496
rect 31849 17487 31907 17493
rect 32214 17484 32220 17496
rect 32272 17524 32278 17536
rect 32950 17524 32956 17536
rect 32272 17496 32956 17524
rect 32272 17484 32278 17496
rect 32950 17484 32956 17496
rect 33008 17484 33014 17536
rect 1104 17434 35027 17456
rect 1104 17382 9390 17434
rect 9442 17382 9454 17434
rect 9506 17382 9518 17434
rect 9570 17382 9582 17434
rect 9634 17382 9646 17434
rect 9698 17382 17831 17434
rect 17883 17382 17895 17434
rect 17947 17382 17959 17434
rect 18011 17382 18023 17434
rect 18075 17382 18087 17434
rect 18139 17382 26272 17434
rect 26324 17382 26336 17434
rect 26388 17382 26400 17434
rect 26452 17382 26464 17434
rect 26516 17382 26528 17434
rect 26580 17382 34713 17434
rect 34765 17382 34777 17434
rect 34829 17382 34841 17434
rect 34893 17382 34905 17434
rect 34957 17382 34969 17434
rect 35021 17382 35027 17434
rect 1104 17360 35027 17382
rect 19334 17320 19340 17332
rect 19295 17292 19340 17320
rect 19334 17280 19340 17292
rect 19392 17280 19398 17332
rect 19426 17280 19432 17332
rect 19484 17280 19490 17332
rect 21450 17320 21456 17332
rect 21411 17292 21456 17320
rect 21450 17280 21456 17292
rect 21508 17280 21514 17332
rect 25682 17320 25688 17332
rect 24872 17292 25688 17320
rect 19058 17212 19064 17264
rect 19116 17252 19122 17264
rect 19444 17252 19472 17280
rect 20806 17252 20812 17264
rect 19116 17224 19380 17252
rect 19444 17224 20116 17252
rect 19116 17212 19122 17224
rect 19245 17187 19303 17193
rect 19245 17153 19257 17187
rect 19291 17153 19303 17187
rect 19352 17184 19380 17224
rect 19426 17184 19432 17196
rect 19352 17156 19432 17184
rect 19245 17147 19303 17153
rect 1762 17116 1768 17128
rect 1723 17088 1768 17116
rect 1762 17076 1768 17088
rect 1820 17076 1826 17128
rect 1949 17119 2007 17125
rect 1949 17085 1961 17119
rect 1995 17116 2007 17119
rect 2590 17116 2596 17128
rect 1995 17088 2596 17116
rect 1995 17085 2007 17088
rect 1949 17079 2007 17085
rect 2590 17076 2596 17088
rect 2648 17076 2654 17128
rect 2774 17116 2780 17128
rect 2735 17088 2780 17116
rect 2774 17076 2780 17088
rect 2832 17076 2838 17128
rect 19260 17116 19288 17147
rect 19426 17144 19432 17156
rect 19484 17184 19490 17196
rect 20088 17193 20116 17224
rect 20272 17224 20812 17252
rect 20073 17187 20131 17193
rect 19484 17156 19577 17184
rect 19484 17144 19490 17156
rect 20073 17153 20085 17187
rect 20119 17153 20131 17187
rect 20272 17184 20300 17224
rect 20806 17212 20812 17224
rect 20864 17212 20870 17264
rect 21542 17212 21548 17264
rect 21600 17252 21606 17264
rect 23100 17255 23158 17261
rect 21600 17224 22876 17252
rect 21600 17212 21606 17224
rect 20073 17147 20131 17153
rect 20180 17156 20300 17184
rect 20340 17187 20398 17193
rect 20180 17116 20208 17156
rect 20340 17153 20352 17187
rect 20386 17184 20398 17187
rect 20622 17184 20628 17196
rect 20386 17156 20628 17184
rect 20386 17153 20398 17156
rect 20340 17147 20398 17153
rect 20622 17144 20628 17156
rect 20680 17144 20686 17196
rect 22094 17144 22100 17196
rect 22152 17184 22158 17196
rect 22189 17187 22247 17193
rect 22189 17184 22201 17187
rect 22152 17156 22201 17184
rect 22152 17144 22158 17156
rect 22189 17153 22201 17156
rect 22235 17184 22247 17187
rect 22462 17184 22468 17196
rect 22235 17156 22468 17184
rect 22235 17153 22247 17156
rect 22189 17147 22247 17153
rect 22462 17144 22468 17156
rect 22520 17144 22526 17196
rect 22848 17193 22876 17224
rect 23100 17221 23112 17255
rect 23146 17252 23158 17255
rect 23474 17252 23480 17264
rect 23146 17224 23480 17252
rect 23146 17221 23158 17224
rect 23100 17215 23158 17221
rect 23474 17212 23480 17224
rect 23532 17212 23538 17264
rect 24872 17261 24900 17292
rect 25682 17280 25688 17292
rect 25740 17280 25746 17332
rect 26878 17280 26884 17332
rect 26936 17320 26942 17332
rect 29822 17320 29828 17332
rect 26936 17292 29828 17320
rect 26936 17280 26942 17292
rect 29822 17280 29828 17292
rect 29880 17280 29886 17332
rect 30282 17320 30288 17332
rect 30243 17292 30288 17320
rect 30282 17280 30288 17292
rect 30340 17280 30346 17332
rect 30374 17280 30380 17332
rect 30432 17320 30438 17332
rect 30432 17292 32720 17320
rect 30432 17280 30438 17292
rect 24857 17255 24915 17261
rect 24857 17221 24869 17255
rect 24903 17221 24915 17255
rect 25038 17252 25044 17264
rect 25096 17261 25102 17264
rect 25096 17255 25131 17261
rect 24983 17224 25044 17252
rect 24857 17215 24915 17221
rect 25038 17212 25044 17224
rect 25119 17252 25131 17255
rect 25590 17252 25596 17264
rect 25119 17224 25596 17252
rect 25119 17221 25131 17224
rect 25096 17215 25131 17221
rect 25096 17212 25102 17215
rect 25590 17212 25596 17224
rect 25648 17252 25654 17264
rect 26050 17252 26056 17264
rect 25648 17224 26056 17252
rect 25648 17212 25654 17224
rect 26050 17212 26056 17224
rect 26108 17212 26114 17264
rect 26145 17255 26203 17261
rect 26145 17221 26157 17255
rect 26191 17252 26203 17255
rect 27402 17255 27460 17261
rect 27402 17252 27414 17255
rect 26191 17224 27414 17252
rect 26191 17221 26203 17224
rect 26145 17215 26203 17221
rect 27402 17221 27414 17224
rect 27448 17221 27460 17255
rect 27402 17215 27460 17221
rect 28442 17212 28448 17264
rect 28500 17252 28506 17264
rect 30650 17252 30656 17264
rect 28500 17224 30656 17252
rect 28500 17212 28506 17224
rect 30650 17212 30656 17224
rect 30708 17218 30714 17264
rect 31665 17255 31723 17261
rect 31665 17221 31677 17255
rect 31711 17252 31723 17255
rect 32214 17252 32220 17264
rect 31711 17224 32220 17252
rect 31711 17221 31723 17224
rect 30708 17215 30798 17218
rect 31665 17215 31723 17221
rect 30708 17212 30813 17215
rect 32214 17212 32220 17224
rect 32272 17212 32278 17264
rect 32692 17261 32720 17292
rect 32677 17255 32735 17261
rect 32677 17221 32689 17255
rect 32723 17221 32735 17255
rect 32677 17215 32735 17221
rect 30668 17209 30813 17212
rect 22833 17187 22891 17193
rect 22833 17153 22845 17187
rect 22879 17153 22891 17187
rect 22833 17147 22891 17153
rect 26329 17187 26387 17193
rect 26329 17153 26341 17187
rect 26375 17184 26387 17187
rect 26786 17184 26792 17196
rect 26375 17156 26792 17184
rect 26375 17153 26387 17156
rect 26329 17147 26387 17153
rect 26786 17144 26792 17156
rect 26844 17144 26850 17196
rect 27154 17184 27160 17196
rect 27115 17156 27160 17184
rect 27154 17144 27160 17156
rect 27212 17144 27218 17196
rect 29178 17184 29184 17196
rect 29139 17156 29184 17184
rect 29178 17144 29184 17156
rect 29236 17144 29242 17196
rect 29638 17144 29644 17196
rect 29696 17184 29702 17196
rect 30009 17187 30067 17193
rect 30009 17184 30021 17187
rect 29696 17156 30021 17184
rect 29696 17144 29702 17156
rect 30009 17153 30021 17156
rect 30055 17153 30067 17187
rect 30466 17184 30472 17196
rect 30009 17147 30067 17153
rect 30116 17156 30472 17184
rect 19260 17088 20208 17116
rect 22005 17119 22063 17125
rect 22005 17085 22017 17119
rect 22051 17116 22063 17119
rect 22554 17116 22560 17128
rect 22051 17088 22560 17116
rect 22051 17085 22063 17088
rect 22005 17079 22063 17085
rect 22554 17076 22560 17088
rect 22612 17076 22618 17128
rect 25866 17076 25872 17128
rect 25924 17116 25930 17128
rect 26050 17116 26056 17128
rect 25924 17088 26056 17116
rect 25924 17076 25930 17088
rect 26050 17076 26056 17088
rect 26108 17076 26114 17128
rect 26605 17119 26663 17125
rect 26605 17085 26617 17119
rect 26651 17085 26663 17119
rect 26605 17079 26663 17085
rect 25498 17048 25504 17060
rect 25056 17020 25504 17048
rect 21818 16940 21824 16992
rect 21876 16980 21882 16992
rect 22370 16980 22376 16992
rect 21876 16952 22376 16980
rect 21876 16940 21882 16952
rect 22370 16940 22376 16952
rect 22428 16940 22434 16992
rect 24213 16983 24271 16989
rect 24213 16949 24225 16983
rect 24259 16980 24271 16983
rect 24946 16980 24952 16992
rect 24259 16952 24952 16980
rect 24259 16949 24271 16952
rect 24213 16943 24271 16949
rect 24946 16940 24952 16952
rect 25004 16980 25010 16992
rect 25056 16989 25084 17020
rect 25498 17008 25504 17020
rect 25556 17008 25562 17060
rect 25041 16983 25099 16989
rect 25041 16980 25053 16983
rect 25004 16952 25053 16980
rect 25004 16940 25010 16952
rect 25041 16949 25053 16952
rect 25087 16949 25099 16983
rect 25222 16980 25228 16992
rect 25183 16952 25228 16980
rect 25041 16943 25099 16949
rect 25222 16940 25228 16952
rect 25280 16940 25286 16992
rect 26510 16980 26516 16992
rect 26471 16952 26516 16980
rect 26510 16940 26516 16952
rect 26568 16940 26574 16992
rect 26620 16980 26648 17079
rect 28810 17076 28816 17128
rect 28868 17116 28874 17128
rect 29089 17119 29147 17125
rect 29089 17116 29101 17119
rect 28868 17088 29101 17116
rect 28868 17076 28874 17088
rect 29089 17085 29101 17088
rect 29135 17085 29147 17119
rect 29089 17079 29147 17085
rect 29362 17076 29368 17128
rect 29420 17116 29426 17128
rect 30116 17125 30144 17156
rect 30466 17144 30472 17156
rect 30524 17144 30530 17196
rect 30668 17190 30767 17209
rect 30755 17175 30767 17190
rect 30801 17175 30813 17209
rect 30755 17169 30813 17175
rect 30926 17144 30932 17196
rect 30984 17144 30990 17196
rect 31481 17187 31539 17193
rect 31481 17184 31493 17187
rect 31404 17156 31493 17184
rect 30101 17119 30159 17125
rect 30101 17116 30113 17119
rect 29420 17088 30113 17116
rect 29420 17076 29426 17088
rect 30101 17085 30113 17088
rect 30147 17085 30159 17119
rect 30285 17119 30343 17125
rect 30285 17116 30297 17119
rect 30101 17079 30159 17085
rect 30208 17088 30297 17116
rect 29549 17051 29607 17057
rect 29549 17017 29561 17051
rect 29595 17048 29607 17051
rect 30006 17048 30012 17060
rect 29595 17020 30012 17048
rect 29595 17017 29607 17020
rect 29549 17011 29607 17017
rect 30006 17008 30012 17020
rect 30064 17008 30070 17060
rect 30208 17048 30236 17088
rect 30285 17085 30297 17088
rect 30331 17116 30343 17119
rect 30944 17116 30972 17144
rect 31021 17119 31079 17125
rect 31021 17116 31033 17119
rect 30331 17088 31033 17116
rect 30331 17085 30343 17088
rect 30285 17079 30343 17085
rect 31021 17085 31033 17088
rect 31067 17085 31079 17119
rect 31021 17079 31079 17085
rect 30116 17020 30236 17048
rect 27798 16980 27804 16992
rect 26620 16952 27804 16980
rect 27798 16940 27804 16952
rect 27856 16980 27862 16992
rect 28537 16983 28595 16989
rect 28537 16980 28549 16983
rect 27856 16952 28549 16980
rect 27856 16940 27862 16952
rect 28537 16949 28549 16952
rect 28583 16949 28595 16983
rect 28537 16943 28595 16949
rect 29362 16940 29368 16992
rect 29420 16980 29426 16992
rect 30116 16980 30144 17020
rect 30374 17008 30380 17060
rect 30432 17048 30438 17060
rect 30929 17051 30987 17057
rect 30929 17048 30941 17051
rect 30432 17020 30941 17048
rect 30432 17008 30438 17020
rect 30929 17017 30941 17020
rect 30975 17017 30987 17051
rect 30929 17011 30987 17017
rect 29420 16952 30144 16980
rect 29420 16940 29426 16952
rect 30466 16940 30472 16992
rect 30524 16980 30530 16992
rect 30837 16983 30895 16989
rect 30837 16980 30849 16983
rect 30524 16952 30849 16980
rect 30524 16940 30530 16952
rect 30837 16949 30849 16952
rect 30883 16949 30895 16983
rect 31404 16980 31432 17156
rect 31481 17153 31493 17156
rect 31527 17153 31539 17187
rect 31481 17147 31539 17153
rect 31757 17187 31815 17193
rect 31757 17153 31769 17187
rect 31803 17184 31815 17187
rect 31846 17184 31852 17196
rect 31803 17156 31852 17184
rect 31803 17153 31815 17156
rect 31757 17147 31815 17153
rect 31846 17144 31852 17156
rect 31904 17144 31910 17196
rect 32490 17116 32496 17128
rect 32451 17088 32496 17116
rect 32490 17076 32496 17088
rect 32548 17076 32554 17128
rect 34330 17116 34336 17128
rect 34291 17088 34336 17116
rect 34330 17076 34336 17088
rect 34388 17076 34394 17128
rect 31481 17051 31539 17057
rect 31481 17017 31493 17051
rect 31527 17048 31539 17051
rect 32674 17048 32680 17060
rect 31527 17020 32680 17048
rect 31527 17017 31539 17020
rect 31481 17011 31539 17017
rect 32674 17008 32680 17020
rect 32732 17008 32738 17060
rect 33778 16980 33784 16992
rect 31404 16952 33784 16980
rect 30837 16943 30895 16949
rect 33778 16940 33784 16952
rect 33836 16940 33842 16992
rect 1104 16890 34868 16912
rect 1104 16838 5170 16890
rect 5222 16838 5234 16890
rect 5286 16838 5298 16890
rect 5350 16838 5362 16890
rect 5414 16838 5426 16890
rect 5478 16838 13611 16890
rect 13663 16838 13675 16890
rect 13727 16838 13739 16890
rect 13791 16838 13803 16890
rect 13855 16838 13867 16890
rect 13919 16838 22052 16890
rect 22104 16838 22116 16890
rect 22168 16838 22180 16890
rect 22232 16838 22244 16890
rect 22296 16838 22308 16890
rect 22360 16838 30493 16890
rect 30545 16838 30557 16890
rect 30609 16838 30621 16890
rect 30673 16838 30685 16890
rect 30737 16838 30749 16890
rect 30801 16838 34868 16890
rect 1104 16816 34868 16838
rect 1762 16736 1768 16788
rect 1820 16776 1826 16788
rect 2041 16779 2099 16785
rect 2041 16776 2053 16779
rect 1820 16748 2053 16776
rect 1820 16736 1826 16748
rect 2041 16745 2053 16748
rect 2087 16745 2099 16779
rect 2590 16776 2596 16788
rect 2551 16748 2596 16776
rect 2041 16739 2099 16745
rect 2590 16736 2596 16748
rect 2648 16736 2654 16788
rect 20622 16776 20628 16788
rect 20583 16748 20628 16776
rect 20622 16736 20628 16748
rect 20680 16736 20686 16788
rect 21634 16776 21640 16788
rect 21595 16748 21640 16776
rect 21634 16736 21640 16748
rect 21692 16736 21698 16788
rect 22370 16776 22376 16788
rect 22331 16748 22376 16776
rect 22370 16736 22376 16748
rect 22428 16736 22434 16788
rect 24302 16776 24308 16788
rect 22480 16748 24308 16776
rect 20714 16708 20720 16720
rect 20675 16680 20720 16708
rect 20714 16668 20720 16680
rect 20772 16668 20778 16720
rect 22480 16708 22508 16748
rect 24302 16736 24308 16748
rect 24360 16736 24366 16788
rect 24762 16776 24768 16788
rect 24723 16748 24768 16776
rect 24762 16736 24768 16748
rect 24820 16736 24826 16788
rect 27525 16779 27583 16785
rect 27525 16745 27537 16779
rect 27571 16776 27583 16779
rect 27706 16776 27712 16788
rect 27571 16748 27712 16776
rect 27571 16745 27583 16748
rect 27525 16739 27583 16745
rect 27706 16736 27712 16748
rect 27764 16776 27770 16788
rect 28442 16776 28448 16788
rect 27764 16748 28448 16776
rect 27764 16736 27770 16748
rect 28442 16736 28448 16748
rect 28500 16736 28506 16788
rect 28810 16776 28816 16788
rect 28771 16748 28816 16776
rect 28810 16736 28816 16748
rect 28868 16736 28874 16788
rect 29730 16776 29736 16788
rect 29691 16748 29736 16776
rect 29730 16736 29736 16748
rect 29788 16736 29794 16788
rect 29822 16736 29828 16788
rect 29880 16776 29886 16788
rect 29880 16748 30328 16776
rect 29880 16736 29886 16748
rect 22646 16708 22652 16720
rect 20916 16680 22508 16708
rect 22572 16680 22652 16708
rect 19426 16600 19432 16652
rect 19484 16640 19490 16652
rect 20916 16649 20944 16680
rect 20901 16643 20959 16649
rect 20901 16640 20913 16643
rect 19484 16612 20913 16640
rect 19484 16600 19490 16612
rect 20901 16609 20913 16612
rect 20947 16609 20959 16643
rect 22370 16640 22376 16652
rect 20901 16603 20959 16609
rect 21652 16612 22376 16640
rect 2498 16572 2504 16584
rect 2459 16544 2504 16572
rect 2498 16532 2504 16544
rect 2556 16532 2562 16584
rect 21652 16581 21680 16612
rect 22370 16600 22376 16612
rect 22428 16600 22434 16652
rect 22572 16649 22600 16680
rect 22646 16668 22652 16680
rect 22704 16708 22710 16720
rect 22704 16680 23520 16708
rect 22704 16668 22710 16680
rect 22557 16643 22615 16649
rect 22557 16609 22569 16643
rect 22603 16609 22615 16643
rect 23382 16640 23388 16652
rect 22557 16603 22615 16609
rect 23032 16612 23388 16640
rect 20625 16575 20683 16581
rect 20625 16541 20637 16575
rect 20671 16572 20683 16575
rect 21637 16575 21695 16581
rect 20671 16544 21588 16572
rect 20671 16541 20683 16544
rect 20625 16535 20683 16541
rect 21560 16504 21588 16544
rect 21637 16541 21649 16575
rect 21683 16541 21695 16575
rect 21818 16572 21824 16584
rect 21779 16544 21824 16572
rect 21637 16535 21695 16541
rect 21818 16532 21824 16544
rect 21876 16532 21882 16584
rect 22281 16575 22339 16581
rect 22281 16541 22293 16575
rect 22327 16572 22339 16575
rect 22462 16572 22468 16584
rect 22327 16544 22468 16572
rect 22327 16541 22339 16544
rect 22281 16535 22339 16541
rect 22462 16532 22468 16544
rect 22520 16532 22526 16584
rect 23032 16581 23060 16612
rect 23382 16600 23388 16612
rect 23440 16600 23446 16652
rect 23492 16640 23520 16680
rect 23750 16668 23756 16720
rect 23808 16708 23814 16720
rect 24673 16711 24731 16717
rect 24673 16708 24685 16711
rect 23808 16680 24685 16708
rect 23808 16668 23814 16680
rect 24673 16677 24685 16680
rect 24719 16677 24731 16711
rect 27154 16708 27160 16720
rect 24673 16671 24731 16677
rect 24780 16680 27160 16708
rect 24029 16643 24087 16649
rect 24029 16640 24041 16643
rect 23492 16612 24041 16640
rect 24029 16609 24041 16612
rect 24075 16640 24087 16643
rect 24394 16640 24400 16652
rect 24075 16612 24400 16640
rect 24075 16609 24087 16612
rect 24029 16603 24087 16609
rect 24394 16600 24400 16612
rect 24452 16640 24458 16652
rect 24780 16640 24808 16680
rect 27154 16668 27160 16680
rect 27212 16708 27218 16720
rect 29362 16708 29368 16720
rect 27212 16680 29368 16708
rect 27212 16668 27218 16680
rect 29362 16668 29368 16680
rect 29420 16668 29426 16720
rect 24452 16612 24808 16640
rect 24452 16600 24458 16612
rect 25222 16600 25228 16652
rect 25280 16640 25286 16652
rect 25280 16612 26372 16640
rect 25280 16600 25286 16612
rect 23017 16575 23075 16581
rect 23017 16541 23029 16575
rect 23063 16541 23075 16575
rect 23017 16535 23075 16541
rect 23753 16575 23811 16581
rect 23753 16541 23765 16575
rect 23799 16541 23811 16575
rect 23753 16535 23811 16541
rect 23845 16575 23903 16581
rect 23845 16541 23857 16575
rect 23891 16572 23903 16575
rect 24578 16572 24584 16584
rect 23891 16544 24584 16572
rect 23891 16541 23903 16544
rect 23845 16535 23903 16541
rect 21910 16504 21916 16516
rect 21560 16476 21916 16504
rect 21910 16464 21916 16476
rect 21968 16504 21974 16516
rect 22186 16504 22192 16516
rect 21968 16476 22192 16504
rect 21968 16464 21974 16476
rect 22186 16464 22192 16476
rect 22244 16464 22250 16516
rect 23109 16507 23167 16513
rect 23109 16504 23121 16507
rect 22480 16476 23121 16504
rect 21726 16396 21732 16448
rect 21784 16436 21790 16448
rect 22480 16436 22508 16476
rect 23109 16473 23121 16476
rect 23155 16473 23167 16507
rect 23768 16504 23796 16535
rect 24578 16532 24584 16544
rect 24636 16532 24642 16584
rect 24762 16572 24768 16584
rect 24688 16544 24768 16572
rect 24688 16504 24716 16544
rect 24762 16532 24768 16544
rect 24820 16572 24826 16584
rect 25130 16572 25136 16584
rect 24820 16544 25136 16572
rect 24820 16532 24826 16544
rect 25130 16532 25136 16544
rect 25188 16532 25194 16584
rect 25498 16572 25504 16584
rect 25459 16544 25504 16572
rect 25498 16532 25504 16544
rect 25556 16532 25562 16584
rect 25590 16532 25596 16584
rect 25648 16572 25654 16584
rect 26142 16572 26148 16584
rect 25648 16544 25693 16572
rect 26103 16544 26148 16572
rect 25648 16532 25654 16544
rect 26142 16532 26148 16544
rect 26200 16532 26206 16584
rect 26344 16581 26372 16612
rect 28166 16600 28172 16652
rect 28224 16640 28230 16652
rect 28353 16643 28411 16649
rect 28353 16640 28365 16643
rect 28224 16612 28365 16640
rect 28224 16600 28230 16612
rect 28353 16609 28365 16612
rect 28399 16640 28411 16643
rect 30300 16640 30328 16748
rect 30466 16668 30472 16720
rect 30524 16708 30530 16720
rect 31665 16711 31723 16717
rect 31665 16708 31677 16711
rect 30524 16680 31677 16708
rect 30524 16668 30530 16680
rect 31665 16677 31677 16680
rect 31711 16677 31723 16711
rect 31665 16671 31723 16677
rect 32493 16643 32551 16649
rect 28399 16612 28948 16640
rect 28399 16609 28411 16612
rect 28353 16603 28411 16609
rect 26329 16575 26387 16581
rect 26329 16541 26341 16575
rect 26375 16541 26387 16575
rect 26329 16535 26387 16541
rect 27341 16575 27399 16581
rect 27341 16541 27353 16575
rect 27387 16572 27399 16575
rect 27798 16572 27804 16584
rect 27387 16544 27804 16572
rect 27387 16541 27399 16544
rect 27341 16535 27399 16541
rect 27798 16532 27804 16544
rect 27856 16532 27862 16584
rect 28442 16572 28448 16584
rect 28403 16544 28448 16572
rect 28442 16532 28448 16544
rect 28500 16532 28506 16584
rect 28920 16572 28948 16612
rect 29840 16612 30144 16640
rect 30300 16612 30972 16640
rect 29840 16572 29868 16612
rect 30006 16572 30012 16584
rect 28920 16544 29868 16572
rect 29967 16544 30012 16572
rect 30006 16532 30012 16544
rect 30064 16532 30070 16584
rect 30116 16572 30144 16612
rect 30944 16581 30972 16612
rect 32493 16609 32505 16643
rect 32539 16640 32551 16643
rect 32858 16640 32864 16652
rect 32539 16612 32864 16640
rect 32539 16609 32551 16612
rect 32493 16603 32551 16609
rect 32858 16600 32864 16612
rect 32916 16600 32922 16652
rect 30745 16575 30803 16581
rect 30745 16572 30757 16575
rect 30116 16544 30757 16572
rect 30745 16541 30757 16544
rect 30791 16541 30803 16575
rect 30745 16535 30803 16541
rect 30929 16575 30987 16581
rect 30929 16541 30941 16575
rect 30975 16541 30987 16575
rect 30929 16535 30987 16541
rect 31202 16532 31208 16584
rect 31260 16572 31266 16584
rect 31573 16575 31631 16581
rect 31573 16572 31585 16575
rect 31260 16544 31585 16572
rect 31260 16532 31266 16544
rect 31573 16541 31585 16544
rect 31619 16541 31631 16575
rect 31754 16572 31760 16584
rect 31715 16544 31760 16572
rect 31573 16535 31631 16541
rect 31754 16532 31760 16544
rect 31812 16532 31818 16584
rect 23768 16476 24716 16504
rect 24857 16507 24915 16513
rect 23109 16467 23167 16473
rect 24857 16473 24869 16507
rect 24903 16504 24915 16507
rect 24946 16504 24952 16516
rect 24903 16476 24952 16504
rect 24903 16473 24915 16476
rect 24857 16467 24915 16473
rect 21784 16408 22508 16436
rect 22557 16439 22615 16445
rect 21784 16396 21790 16408
rect 22557 16405 22569 16439
rect 22603 16436 22615 16439
rect 23014 16436 23020 16448
rect 22603 16408 23020 16436
rect 22603 16405 22615 16408
rect 22557 16399 22615 16405
rect 23014 16396 23020 16408
rect 23072 16396 23078 16448
rect 23842 16396 23848 16448
rect 23900 16436 23906 16448
rect 24029 16439 24087 16445
rect 24029 16436 24041 16439
rect 23900 16408 24041 16436
rect 23900 16396 23906 16408
rect 24029 16405 24041 16408
rect 24075 16405 24087 16439
rect 24029 16399 24087 16405
rect 24302 16396 24308 16448
rect 24360 16436 24366 16448
rect 24670 16436 24676 16448
rect 24360 16408 24676 16436
rect 24360 16396 24366 16408
rect 24670 16396 24676 16408
rect 24728 16436 24734 16448
rect 24872 16436 24900 16467
rect 24946 16464 24952 16476
rect 25004 16464 25010 16516
rect 25317 16507 25375 16513
rect 25317 16473 25329 16507
rect 25363 16504 25375 16507
rect 25682 16504 25688 16516
rect 25363 16476 25688 16504
rect 25363 16473 25375 16476
rect 25317 16467 25375 16473
rect 25682 16464 25688 16476
rect 25740 16464 25746 16516
rect 29086 16464 29092 16516
rect 29144 16504 29150 16516
rect 29546 16504 29552 16516
rect 29144 16476 29552 16504
rect 29144 16464 29150 16476
rect 29546 16464 29552 16476
rect 29604 16464 29610 16516
rect 29733 16507 29791 16513
rect 29733 16473 29745 16507
rect 29779 16504 29791 16507
rect 30374 16504 30380 16516
rect 29779 16476 30380 16504
rect 29779 16473 29791 16476
rect 29733 16467 29791 16473
rect 30374 16464 30380 16476
rect 30432 16464 30438 16516
rect 30466 16464 30472 16516
rect 30524 16504 30530 16516
rect 32214 16504 32220 16516
rect 30524 16476 32220 16504
rect 30524 16464 30530 16476
rect 32214 16464 32220 16476
rect 32272 16464 32278 16516
rect 32674 16504 32680 16516
rect 32635 16476 32680 16504
rect 32674 16464 32680 16476
rect 32732 16464 32738 16516
rect 34333 16507 34391 16513
rect 34333 16473 34345 16507
rect 34379 16504 34391 16507
rect 35158 16504 35164 16516
rect 34379 16476 35164 16504
rect 34379 16473 34391 16476
rect 34333 16467 34391 16473
rect 35158 16464 35164 16476
rect 35216 16464 35222 16516
rect 25406 16436 25412 16448
rect 25464 16445 25470 16448
rect 24728 16408 24900 16436
rect 25373 16408 25412 16436
rect 24728 16396 24734 16408
rect 25406 16396 25412 16408
rect 25464 16399 25473 16445
rect 26510 16436 26516 16448
rect 26423 16408 26516 16436
rect 25464 16396 25470 16399
rect 26510 16396 26516 16408
rect 26568 16436 26574 16448
rect 26878 16436 26884 16448
rect 26568 16408 26884 16436
rect 26568 16396 26574 16408
rect 26878 16396 26884 16408
rect 26936 16396 26942 16448
rect 27801 16439 27859 16445
rect 27801 16405 27813 16439
rect 27847 16436 27859 16439
rect 28534 16436 28540 16448
rect 27847 16408 28540 16436
rect 27847 16405 27859 16408
rect 27801 16399 27859 16405
rect 28534 16396 28540 16408
rect 28592 16396 28598 16448
rect 29454 16396 29460 16448
rect 29512 16436 29518 16448
rect 29917 16439 29975 16445
rect 29917 16436 29929 16439
rect 29512 16408 29929 16436
rect 29512 16396 29518 16408
rect 29917 16405 29929 16408
rect 29963 16405 29975 16439
rect 29917 16399 29975 16405
rect 30006 16396 30012 16448
rect 30064 16436 30070 16448
rect 30837 16439 30895 16445
rect 30837 16436 30849 16439
rect 30064 16408 30849 16436
rect 30064 16396 30070 16408
rect 30837 16405 30849 16408
rect 30883 16405 30895 16439
rect 30837 16399 30895 16405
rect 1104 16346 35027 16368
rect 1104 16294 9390 16346
rect 9442 16294 9454 16346
rect 9506 16294 9518 16346
rect 9570 16294 9582 16346
rect 9634 16294 9646 16346
rect 9698 16294 17831 16346
rect 17883 16294 17895 16346
rect 17947 16294 17959 16346
rect 18011 16294 18023 16346
rect 18075 16294 18087 16346
rect 18139 16294 26272 16346
rect 26324 16294 26336 16346
rect 26388 16294 26400 16346
rect 26452 16294 26464 16346
rect 26516 16294 26528 16346
rect 26580 16294 34713 16346
rect 34765 16294 34777 16346
rect 34829 16294 34841 16346
rect 34893 16294 34905 16346
rect 34957 16294 34969 16346
rect 35021 16294 35027 16346
rect 1104 16272 35027 16294
rect 22370 16232 22376 16244
rect 22331 16204 22376 16232
rect 22370 16192 22376 16204
rect 22428 16192 22434 16244
rect 22738 16192 22744 16244
rect 22796 16232 22802 16244
rect 23017 16235 23075 16241
rect 23017 16232 23029 16235
rect 22796 16204 23029 16232
rect 22796 16192 22802 16204
rect 23017 16201 23029 16204
rect 23063 16201 23075 16235
rect 24026 16232 24032 16244
rect 23017 16195 23075 16201
rect 23124 16204 24032 16232
rect 23124 16164 23152 16204
rect 24026 16192 24032 16204
rect 24084 16192 24090 16244
rect 24486 16232 24492 16244
rect 24447 16204 24492 16232
rect 24486 16192 24492 16204
rect 24544 16192 24550 16244
rect 25314 16232 25320 16244
rect 25275 16204 25320 16232
rect 25314 16192 25320 16204
rect 25372 16192 25378 16244
rect 28902 16192 28908 16244
rect 28960 16232 28966 16244
rect 29917 16235 29975 16241
rect 29917 16232 29929 16235
rect 28960 16204 29929 16232
rect 28960 16192 28966 16204
rect 29917 16201 29929 16204
rect 29963 16201 29975 16235
rect 29917 16195 29975 16201
rect 30653 16235 30711 16241
rect 30653 16201 30665 16235
rect 30699 16232 30711 16235
rect 30742 16232 30748 16244
rect 30699 16204 30748 16232
rect 30699 16201 30711 16204
rect 30653 16195 30711 16201
rect 30742 16192 30748 16204
rect 30800 16192 30806 16244
rect 31478 16232 31484 16244
rect 31439 16204 31484 16232
rect 31478 16192 31484 16204
rect 31536 16192 31542 16244
rect 32398 16232 32404 16244
rect 32359 16204 32404 16232
rect 32398 16192 32404 16204
rect 32456 16192 32462 16244
rect 33045 16235 33103 16241
rect 33045 16201 33057 16235
rect 33091 16232 33103 16235
rect 33502 16232 33508 16244
rect 33091 16204 33508 16232
rect 33091 16201 33103 16204
rect 33045 16195 33103 16201
rect 33502 16192 33508 16204
rect 33560 16192 33566 16244
rect 33781 16235 33839 16241
rect 33781 16201 33793 16235
rect 33827 16232 33839 16235
rect 34514 16232 34520 16244
rect 33827 16204 34520 16232
rect 33827 16201 33839 16204
rect 33781 16195 33839 16201
rect 34514 16192 34520 16204
rect 34572 16192 34578 16244
rect 22940 16136 23152 16164
rect 22094 16096 22100 16108
rect 22055 16068 22100 16096
rect 22094 16056 22100 16068
rect 22152 16056 22158 16108
rect 22940 16105 22968 16136
rect 23566 16124 23572 16176
rect 23624 16164 23630 16176
rect 23661 16167 23719 16173
rect 23661 16164 23673 16167
rect 23624 16136 23673 16164
rect 23624 16124 23630 16136
rect 23661 16133 23673 16136
rect 23707 16133 23719 16167
rect 23661 16127 23719 16133
rect 23845 16167 23903 16173
rect 23845 16133 23857 16167
rect 23891 16164 23903 16167
rect 25498 16164 25504 16176
rect 23891 16136 25504 16164
rect 23891 16133 23903 16136
rect 23845 16127 23903 16133
rect 25498 16124 25504 16136
rect 25556 16124 25562 16176
rect 28258 16164 28264 16176
rect 27448 16136 28264 16164
rect 22925 16099 22983 16105
rect 22925 16065 22937 16099
rect 22971 16065 22983 16099
rect 22925 16059 22983 16065
rect 23109 16099 23167 16105
rect 23109 16065 23121 16099
rect 23155 16065 23167 16099
rect 23109 16059 23167 16065
rect 23937 16099 23995 16105
rect 23937 16065 23949 16099
rect 23983 16096 23995 16099
rect 24026 16096 24032 16108
rect 23983 16068 24032 16096
rect 23983 16065 23995 16068
rect 23937 16059 23995 16065
rect 22186 16028 22192 16040
rect 22147 16000 22192 16028
rect 22186 15988 22192 16000
rect 22244 15988 22250 16040
rect 22373 16031 22431 16037
rect 22373 15997 22385 16031
rect 22419 16028 22431 16031
rect 22646 16028 22652 16040
rect 22419 16000 22652 16028
rect 22419 15997 22431 16000
rect 22373 15991 22431 15997
rect 22646 15988 22652 16000
rect 22704 15988 22710 16040
rect 20530 15920 20536 15972
rect 20588 15960 20594 15972
rect 23124 15960 23152 16059
rect 24026 16056 24032 16068
rect 24084 16056 24090 16108
rect 24397 16099 24455 16105
rect 24397 16065 24409 16099
rect 24443 16065 24455 16099
rect 24397 16059 24455 16065
rect 23658 15960 23664 15972
rect 20588 15932 23152 15960
rect 23619 15932 23664 15960
rect 20588 15920 20594 15932
rect 23658 15920 23664 15932
rect 23716 15920 23722 15972
rect 1578 15852 1584 15904
rect 1636 15892 1642 15904
rect 2041 15895 2099 15901
rect 2041 15892 2053 15895
rect 1636 15864 2053 15892
rect 1636 15852 1642 15864
rect 2041 15861 2053 15864
rect 2087 15861 2099 15895
rect 2041 15855 2099 15861
rect 22094 15852 22100 15904
rect 22152 15892 22158 15904
rect 22554 15892 22560 15904
rect 22152 15864 22560 15892
rect 22152 15852 22158 15864
rect 22554 15852 22560 15864
rect 22612 15892 22618 15904
rect 24412 15892 24440 16059
rect 25222 16056 25228 16108
rect 25280 16096 25286 16108
rect 25317 16099 25375 16105
rect 25317 16096 25329 16099
rect 25280 16068 25329 16096
rect 25280 16056 25286 16068
rect 25317 16065 25329 16068
rect 25363 16065 25375 16099
rect 25317 16059 25375 16065
rect 25332 15960 25360 16059
rect 25406 16056 25412 16108
rect 25464 16096 25470 16108
rect 26053 16099 26111 16105
rect 25464 16068 25509 16096
rect 25464 16056 25470 16068
rect 26053 16065 26065 16099
rect 26099 16096 26111 16099
rect 26142 16096 26148 16108
rect 26099 16068 26148 16096
rect 26099 16065 26111 16068
rect 26053 16059 26111 16065
rect 26142 16056 26148 16068
rect 26200 16056 26206 16108
rect 27448 16105 27476 16136
rect 28258 16124 28264 16136
rect 28316 16164 28322 16176
rect 28810 16164 28816 16176
rect 28316 16136 28816 16164
rect 28316 16124 28322 16136
rect 28810 16124 28816 16136
rect 28868 16124 28874 16176
rect 29270 16164 29276 16176
rect 29231 16136 29276 16164
rect 29270 16124 29276 16136
rect 29328 16124 29334 16176
rect 29454 16124 29460 16176
rect 29512 16164 29518 16176
rect 29512 16136 30052 16164
rect 29512 16124 29518 16136
rect 27433 16099 27491 16105
rect 27433 16065 27445 16099
rect 27479 16065 27491 16099
rect 27433 16059 27491 16065
rect 27525 16099 27583 16105
rect 27525 16065 27537 16099
rect 27571 16096 27583 16099
rect 28166 16096 28172 16108
rect 27571 16068 28172 16096
rect 27571 16065 27583 16068
rect 27525 16059 27583 16065
rect 28166 16056 28172 16068
rect 28224 16056 28230 16108
rect 28350 16096 28356 16108
rect 28311 16068 28356 16096
rect 28350 16056 28356 16068
rect 28408 16056 28414 16108
rect 28718 16056 28724 16108
rect 28776 16096 28782 16108
rect 28776 16094 28994 16096
rect 29086 16094 29092 16108
rect 28776 16068 29092 16094
rect 28776 16056 28782 16068
rect 28966 16066 29092 16068
rect 29086 16056 29092 16066
rect 29144 16056 29150 16108
rect 29181 16099 29239 16105
rect 29181 16065 29193 16099
rect 29227 16096 29239 16099
rect 29227 16068 29316 16096
rect 29227 16065 29239 16068
rect 29181 16059 29239 16065
rect 25590 16028 25596 16040
rect 25503 16000 25596 16028
rect 25590 15988 25596 16000
rect 25648 16028 25654 16040
rect 26329 16031 26387 16037
rect 25648 16000 26280 16028
rect 25648 15988 25654 16000
rect 26145 15963 26203 15969
rect 26145 15960 26157 15963
rect 25332 15932 26157 15960
rect 26145 15929 26157 15932
rect 26191 15929 26203 15963
rect 26252 15960 26280 16000
rect 26329 15997 26341 16031
rect 26375 16028 26387 16031
rect 27154 16028 27160 16040
rect 26375 16000 27160 16028
rect 26375 15997 26387 16000
rect 26329 15991 26387 15997
rect 27154 15988 27160 16000
rect 27212 15988 27218 16040
rect 28445 16031 28503 16037
rect 28445 15997 28457 16031
rect 28491 16028 28503 16031
rect 28626 16028 28632 16040
rect 28491 16000 28632 16028
rect 28491 15997 28503 16000
rect 28445 15991 28503 15997
rect 28626 15988 28632 16000
rect 28684 15988 28690 16040
rect 29288 16028 29316 16068
rect 29362 16056 29368 16108
rect 29420 16096 29426 16108
rect 29822 16096 29828 16108
rect 29420 16068 29465 16096
rect 29783 16068 29828 16096
rect 29420 16056 29426 16068
rect 29822 16056 29828 16068
rect 29880 16056 29886 16108
rect 30024 16105 30052 16136
rect 30190 16124 30196 16176
rect 30248 16164 30254 16176
rect 30248 16136 31432 16164
rect 30248 16124 30254 16136
rect 30009 16099 30067 16105
rect 30009 16065 30021 16099
rect 30055 16065 30067 16099
rect 30466 16096 30472 16108
rect 30427 16068 30472 16096
rect 30009 16059 30067 16065
rect 30466 16056 30472 16068
rect 30524 16056 30530 16108
rect 30650 16096 30656 16108
rect 30611 16068 30656 16096
rect 30650 16056 30656 16068
rect 30708 16056 30714 16108
rect 31404 16105 31432 16136
rect 31938 16124 31944 16176
rect 31996 16164 32002 16176
rect 31996 16136 33916 16164
rect 31996 16124 32002 16136
rect 31389 16099 31447 16105
rect 31389 16065 31401 16099
rect 31435 16065 31447 16099
rect 31389 16059 31447 16065
rect 32309 16099 32367 16105
rect 32309 16065 32321 16099
rect 32355 16065 32367 16099
rect 32950 16096 32956 16108
rect 32911 16068 32956 16096
rect 32309 16059 32367 16065
rect 29546 16028 29552 16040
rect 28736 16000 28994 16028
rect 29288 16000 29552 16028
rect 28736 15969 28764 16000
rect 28721 15963 28779 15969
rect 26252 15932 28580 15960
rect 26145 15923 26203 15929
rect 22612 15864 24440 15892
rect 22612 15852 22618 15864
rect 24946 15852 24952 15904
rect 25004 15892 25010 15904
rect 25590 15892 25596 15904
rect 25004 15864 25596 15892
rect 25004 15852 25010 15864
rect 25590 15852 25596 15864
rect 25648 15852 25654 15904
rect 26237 15895 26295 15901
rect 26237 15861 26249 15895
rect 26283 15892 26295 15895
rect 26602 15892 26608 15904
rect 26283 15864 26608 15892
rect 26283 15861 26295 15864
rect 26237 15855 26295 15861
rect 26602 15852 26608 15864
rect 26660 15852 26666 15904
rect 27709 15895 27767 15901
rect 27709 15861 27721 15895
rect 27755 15892 27767 15895
rect 28442 15892 28448 15904
rect 27755 15864 28448 15892
rect 27755 15861 27767 15864
rect 27709 15855 27767 15861
rect 28442 15852 28448 15864
rect 28500 15852 28506 15904
rect 28552 15892 28580 15932
rect 28721 15929 28733 15963
rect 28767 15929 28779 15963
rect 28966 15960 28994 16000
rect 29546 15988 29552 16000
rect 29604 15988 29610 16040
rect 31110 15988 31116 16040
rect 31168 16028 31174 16040
rect 32324 16028 32352 16059
rect 32950 16056 32956 16068
rect 33008 16056 33014 16108
rect 33318 16056 33324 16108
rect 33376 16096 33382 16108
rect 33888 16105 33916 16136
rect 33689 16099 33747 16105
rect 33689 16096 33701 16099
rect 33376 16068 33701 16096
rect 33376 16056 33382 16068
rect 33689 16065 33701 16068
rect 33735 16065 33747 16099
rect 33689 16059 33747 16065
rect 33873 16099 33931 16105
rect 33873 16065 33885 16099
rect 33919 16065 33931 16099
rect 33873 16059 33931 16065
rect 31168 16000 32352 16028
rect 31168 15988 31174 16000
rect 29086 15960 29092 15972
rect 28966 15932 29092 15960
rect 28721 15923 28779 15929
rect 29086 15920 29092 15932
rect 29144 15920 29150 15972
rect 31202 15920 31208 15972
rect 31260 15960 31266 15972
rect 32674 15960 32680 15972
rect 31260 15932 32680 15960
rect 31260 15920 31266 15932
rect 32674 15920 32680 15932
rect 32732 15920 32738 15972
rect 28994 15892 29000 15904
rect 28552 15864 29000 15892
rect 28994 15852 29000 15864
rect 29052 15852 29058 15904
rect 1104 15802 34868 15824
rect 1104 15750 5170 15802
rect 5222 15750 5234 15802
rect 5286 15750 5298 15802
rect 5350 15750 5362 15802
rect 5414 15750 5426 15802
rect 5478 15750 13611 15802
rect 13663 15750 13675 15802
rect 13727 15750 13739 15802
rect 13791 15750 13803 15802
rect 13855 15750 13867 15802
rect 13919 15750 22052 15802
rect 22104 15750 22116 15802
rect 22168 15750 22180 15802
rect 22232 15750 22244 15802
rect 22296 15750 22308 15802
rect 22360 15750 30493 15802
rect 30545 15750 30557 15802
rect 30609 15750 30621 15802
rect 30673 15750 30685 15802
rect 30737 15750 30749 15802
rect 30801 15750 34868 15802
rect 1104 15728 34868 15750
rect 22830 15648 22836 15700
rect 22888 15688 22894 15700
rect 23017 15691 23075 15697
rect 23017 15688 23029 15691
rect 22888 15660 23029 15688
rect 22888 15648 22894 15660
rect 23017 15657 23029 15660
rect 23063 15657 23075 15691
rect 23017 15651 23075 15657
rect 23845 15691 23903 15697
rect 23845 15657 23857 15691
rect 23891 15688 23903 15691
rect 23934 15688 23940 15700
rect 23891 15660 23940 15688
rect 23891 15657 23903 15660
rect 23845 15651 23903 15657
rect 23934 15648 23940 15660
rect 23992 15648 23998 15700
rect 24118 15648 24124 15700
rect 24176 15688 24182 15700
rect 25133 15691 25191 15697
rect 25133 15688 25145 15691
rect 24176 15660 25145 15688
rect 24176 15648 24182 15660
rect 25133 15657 25145 15660
rect 25179 15657 25191 15691
rect 25133 15651 25191 15657
rect 26605 15691 26663 15697
rect 26605 15657 26617 15691
rect 26651 15688 26663 15691
rect 26786 15688 26792 15700
rect 26651 15660 26792 15688
rect 26651 15657 26663 15660
rect 26605 15651 26663 15657
rect 26786 15648 26792 15660
rect 26844 15648 26850 15700
rect 26970 15648 26976 15700
rect 27028 15688 27034 15700
rect 27433 15691 27491 15697
rect 27433 15688 27445 15691
rect 27028 15660 27445 15688
rect 27028 15648 27034 15660
rect 27433 15657 27445 15660
rect 27479 15657 27491 15691
rect 27433 15651 27491 15657
rect 28261 15691 28319 15697
rect 28261 15657 28273 15691
rect 28307 15688 28319 15691
rect 29178 15688 29184 15700
rect 28307 15660 29184 15688
rect 28307 15657 28319 15660
rect 28261 15651 28319 15657
rect 29178 15648 29184 15660
rect 29236 15648 29242 15700
rect 30653 15691 30711 15697
rect 30653 15657 30665 15691
rect 30699 15688 30711 15691
rect 30834 15688 30840 15700
rect 30699 15660 30840 15688
rect 30699 15657 30711 15660
rect 30653 15651 30711 15657
rect 30834 15648 30840 15660
rect 30892 15648 30898 15700
rect 31389 15691 31447 15697
rect 31389 15657 31401 15691
rect 31435 15688 31447 15691
rect 31570 15688 31576 15700
rect 31435 15660 31576 15688
rect 31435 15657 31447 15660
rect 31389 15651 31447 15657
rect 31570 15648 31576 15660
rect 31628 15648 31634 15700
rect 32030 15688 32036 15700
rect 31991 15660 32036 15688
rect 32030 15648 32036 15660
rect 32088 15648 32094 15700
rect 32585 15691 32643 15697
rect 32585 15657 32597 15691
rect 32631 15688 32643 15691
rect 33134 15688 33140 15700
rect 32631 15660 33140 15688
rect 32631 15657 32643 15660
rect 32585 15651 32643 15657
rect 33134 15648 33140 15660
rect 33192 15648 33198 15700
rect 33873 15691 33931 15697
rect 33873 15657 33885 15691
rect 33919 15688 33931 15691
rect 34054 15688 34060 15700
rect 33919 15660 34060 15688
rect 33919 15657 33931 15660
rect 33873 15651 33931 15657
rect 34054 15648 34060 15660
rect 34112 15648 34118 15700
rect 23106 15580 23112 15632
rect 23164 15620 23170 15632
rect 25777 15623 25835 15629
rect 25777 15620 25789 15623
rect 23164 15592 25789 15620
rect 23164 15580 23170 15592
rect 25777 15589 25789 15592
rect 25823 15589 25835 15623
rect 25777 15583 25835 15589
rect 26418 15580 26424 15632
rect 26476 15620 26482 15632
rect 31294 15620 31300 15632
rect 26476 15592 31300 15620
rect 26476 15580 26482 15592
rect 31294 15580 31300 15592
rect 31352 15580 31358 15632
rect 31846 15580 31852 15632
rect 31904 15620 31910 15632
rect 32674 15620 32680 15632
rect 31904 15592 32680 15620
rect 31904 15580 31910 15592
rect 32674 15580 32680 15592
rect 32732 15580 32738 15632
rect 1578 15552 1584 15564
rect 1539 15524 1584 15552
rect 1578 15512 1584 15524
rect 1636 15512 1642 15564
rect 2774 15552 2780 15564
rect 2735 15524 2780 15552
rect 2774 15512 2780 15524
rect 2832 15512 2838 15564
rect 24210 15512 24216 15564
rect 24268 15552 24274 15564
rect 24268 15524 25452 15552
rect 24268 15512 24274 15524
rect 23014 15484 23020 15496
rect 22975 15456 23020 15484
rect 23014 15444 23020 15456
rect 23072 15444 23078 15496
rect 23201 15487 23259 15493
rect 23201 15453 23213 15487
rect 23247 15484 23259 15487
rect 23290 15484 23296 15496
rect 23247 15456 23296 15484
rect 23247 15453 23259 15456
rect 23201 15447 23259 15453
rect 23290 15444 23296 15456
rect 23348 15444 23354 15496
rect 23842 15484 23848 15496
rect 23803 15456 23848 15484
rect 23842 15444 23848 15456
rect 23900 15444 23906 15496
rect 24026 15444 24032 15496
rect 24084 15484 24090 15496
rect 25038 15484 25044 15496
rect 24084 15456 25044 15484
rect 24084 15444 24090 15456
rect 25038 15444 25044 15456
rect 25096 15444 25102 15496
rect 25133 15487 25191 15493
rect 25133 15453 25145 15487
rect 25179 15484 25191 15487
rect 25317 15487 25375 15493
rect 25179 15456 25268 15484
rect 25179 15453 25191 15456
rect 25133 15447 25191 15453
rect 1762 15416 1768 15428
rect 1723 15388 1768 15416
rect 1762 15376 1768 15388
rect 1820 15376 1826 15428
rect 25240 15348 25268 15456
rect 25317 15453 25329 15487
rect 25363 15453 25375 15487
rect 25424 15484 25452 15524
rect 25682 15512 25688 15564
rect 25740 15552 25746 15564
rect 32306 15552 32312 15564
rect 25740 15524 27384 15552
rect 25740 15512 25746 15524
rect 25777 15487 25835 15493
rect 25777 15484 25789 15487
rect 25424 15456 25789 15484
rect 25317 15447 25375 15453
rect 25777 15453 25789 15456
rect 25823 15453 25835 15487
rect 25777 15447 25835 15453
rect 25332 15416 25360 15447
rect 25866 15444 25872 15496
rect 25924 15484 25930 15496
rect 25961 15487 26019 15493
rect 25961 15484 25973 15487
rect 25924 15456 25973 15484
rect 25924 15444 25930 15456
rect 25961 15453 25973 15456
rect 26007 15484 26019 15487
rect 26878 15484 26884 15496
rect 26007 15456 26740 15484
rect 26839 15456 26884 15484
rect 26007 15453 26019 15456
rect 25961 15447 26019 15453
rect 25590 15416 25596 15428
rect 25332 15388 25596 15416
rect 25590 15376 25596 15388
rect 25648 15376 25654 15428
rect 26418 15376 26424 15428
rect 26476 15416 26482 15428
rect 26605 15419 26663 15425
rect 26605 15416 26617 15419
rect 26476 15388 26617 15416
rect 26476 15376 26482 15388
rect 26605 15385 26617 15388
rect 26651 15385 26663 15419
rect 26605 15379 26663 15385
rect 25406 15348 25412 15360
rect 25240 15320 25412 15348
rect 25406 15308 25412 15320
rect 25464 15348 25470 15360
rect 26510 15348 26516 15360
rect 25464 15320 26516 15348
rect 25464 15308 25470 15320
rect 26510 15308 26516 15320
rect 26568 15308 26574 15360
rect 26712 15348 26740 15456
rect 26878 15444 26884 15456
rect 26936 15444 26942 15496
rect 27356 15493 27384 15524
rect 27908 15524 30052 15552
rect 27341 15487 27399 15493
rect 27341 15453 27353 15487
rect 27387 15453 27399 15487
rect 27341 15447 27399 15453
rect 26789 15419 26847 15425
rect 26789 15385 26801 15419
rect 26835 15416 26847 15419
rect 27798 15416 27804 15428
rect 26835 15388 27804 15416
rect 26835 15385 26847 15388
rect 26789 15379 26847 15385
rect 27798 15376 27804 15388
rect 27856 15376 27862 15428
rect 27908 15348 27936 15524
rect 28442 15484 28448 15496
rect 28403 15456 28448 15484
rect 28442 15444 28448 15456
rect 28500 15444 28506 15496
rect 28626 15444 28632 15496
rect 28684 15484 28690 15496
rect 28721 15487 28779 15493
rect 28721 15484 28733 15487
rect 28684 15456 28733 15484
rect 28684 15444 28690 15456
rect 28721 15453 28733 15456
rect 28767 15453 28779 15487
rect 28721 15447 28779 15453
rect 29733 15487 29791 15493
rect 29733 15453 29745 15487
rect 29779 15453 29791 15487
rect 29733 15447 29791 15453
rect 28460 15416 28488 15444
rect 29748 15416 29776 15447
rect 29822 15444 29828 15496
rect 29880 15484 29886 15496
rect 29917 15487 29975 15493
rect 29917 15484 29929 15487
rect 29880 15456 29929 15484
rect 29880 15444 29886 15456
rect 29917 15453 29929 15456
rect 29963 15453 29975 15487
rect 29917 15447 29975 15453
rect 28460 15388 29776 15416
rect 30024 15416 30052 15524
rect 31312 15524 32312 15552
rect 30374 15444 30380 15496
rect 30432 15484 30438 15496
rect 30653 15487 30711 15493
rect 30653 15484 30665 15487
rect 30432 15456 30665 15484
rect 30432 15444 30438 15456
rect 30653 15453 30665 15456
rect 30699 15453 30711 15487
rect 30834 15484 30840 15496
rect 30795 15456 30840 15484
rect 30653 15447 30711 15453
rect 30834 15444 30840 15456
rect 30892 15444 30898 15496
rect 31312 15493 31340 15524
rect 32306 15512 32312 15524
rect 32364 15512 32370 15564
rect 33962 15552 33968 15564
rect 32600 15524 33968 15552
rect 31297 15487 31355 15493
rect 31297 15453 31309 15487
rect 31343 15453 31355 15487
rect 31297 15447 31355 15453
rect 31662 15444 31668 15496
rect 31720 15484 31726 15496
rect 32600 15493 32628 15524
rect 33962 15512 33968 15524
rect 34020 15512 34026 15564
rect 31941 15487 31999 15493
rect 31941 15484 31953 15487
rect 31720 15456 31953 15484
rect 31720 15444 31726 15456
rect 31941 15453 31953 15456
rect 31987 15453 31999 15487
rect 31941 15447 31999 15453
rect 32585 15487 32643 15493
rect 32585 15453 32597 15487
rect 32631 15453 32643 15487
rect 32585 15447 32643 15453
rect 32674 15444 32680 15496
rect 32732 15484 32738 15496
rect 32769 15487 32827 15493
rect 32769 15484 32781 15487
rect 32732 15456 32781 15484
rect 32732 15444 32738 15456
rect 32769 15453 32781 15456
rect 32815 15453 32827 15487
rect 33778 15484 33784 15496
rect 33739 15456 33784 15484
rect 32769 15447 32827 15453
rect 33778 15444 33784 15456
rect 33836 15444 33842 15496
rect 34238 15416 34244 15428
rect 30024 15388 34244 15416
rect 34238 15376 34244 15388
rect 34296 15376 34302 15428
rect 26712 15320 27936 15348
rect 28350 15308 28356 15360
rect 28408 15348 28414 15360
rect 28629 15351 28687 15357
rect 28629 15348 28641 15351
rect 28408 15320 28641 15348
rect 28408 15308 28414 15320
rect 28629 15317 28641 15320
rect 28675 15348 28687 15351
rect 29825 15351 29883 15357
rect 29825 15348 29837 15351
rect 28675 15320 29837 15348
rect 28675 15317 28687 15320
rect 28629 15311 28687 15317
rect 29825 15317 29837 15320
rect 29871 15317 29883 15351
rect 29825 15311 29883 15317
rect 1104 15258 35027 15280
rect 1104 15206 9390 15258
rect 9442 15206 9454 15258
rect 9506 15206 9518 15258
rect 9570 15206 9582 15258
rect 9634 15206 9646 15258
rect 9698 15206 17831 15258
rect 17883 15206 17895 15258
rect 17947 15206 17959 15258
rect 18011 15206 18023 15258
rect 18075 15206 18087 15258
rect 18139 15206 26272 15258
rect 26324 15206 26336 15258
rect 26388 15206 26400 15258
rect 26452 15206 26464 15258
rect 26516 15206 26528 15258
rect 26580 15206 34713 15258
rect 34765 15206 34777 15258
rect 34829 15206 34841 15258
rect 34893 15206 34905 15258
rect 34957 15206 34969 15258
rect 35021 15206 35027 15258
rect 1104 15184 35027 15206
rect 1762 15104 1768 15156
rect 1820 15144 1826 15156
rect 2225 15147 2283 15153
rect 2225 15144 2237 15147
rect 1820 15116 2237 15144
rect 1820 15104 1826 15116
rect 2225 15113 2237 15116
rect 2271 15113 2283 15147
rect 24854 15144 24860 15156
rect 24815 15116 24860 15144
rect 2225 15107 2283 15113
rect 24854 15104 24860 15116
rect 24912 15104 24918 15156
rect 25590 15144 25596 15156
rect 25551 15116 25596 15144
rect 25590 15104 25596 15116
rect 25648 15104 25654 15156
rect 26145 15147 26203 15153
rect 26145 15113 26157 15147
rect 26191 15144 26203 15147
rect 27062 15144 27068 15156
rect 26191 15116 27068 15144
rect 26191 15113 26203 15116
rect 26145 15107 26203 15113
rect 27062 15104 27068 15116
rect 27120 15104 27126 15156
rect 27246 15144 27252 15156
rect 27207 15116 27252 15144
rect 27246 15104 27252 15116
rect 27304 15104 27310 15156
rect 28074 15144 28080 15156
rect 28035 15116 28080 15144
rect 28074 15104 28080 15116
rect 28132 15104 28138 15156
rect 29362 15144 29368 15156
rect 29323 15116 29368 15144
rect 29362 15104 29368 15116
rect 29420 15104 29426 15156
rect 30009 15147 30067 15153
rect 30009 15113 30021 15147
rect 30055 15144 30067 15147
rect 30282 15144 30288 15156
rect 30055 15116 30288 15144
rect 30055 15113 30067 15116
rect 30009 15107 30067 15113
rect 30282 15104 30288 15116
rect 30340 15104 30346 15156
rect 32401 15147 32459 15153
rect 32401 15113 32413 15147
rect 32447 15144 32459 15147
rect 32766 15144 32772 15156
rect 32447 15116 32772 15144
rect 32447 15113 32459 15116
rect 32401 15107 32459 15113
rect 32766 15104 32772 15116
rect 32824 15104 32830 15156
rect 33042 15144 33048 15156
rect 33003 15116 33048 15144
rect 33042 15104 33048 15116
rect 33100 15104 33106 15156
rect 28721 15079 28779 15085
rect 28721 15045 28733 15079
rect 28767 15076 28779 15079
rect 29822 15076 29828 15088
rect 28767 15048 29828 15076
rect 28767 15045 28779 15048
rect 28721 15039 28779 15045
rect 29822 15036 29828 15048
rect 29880 15036 29886 15088
rect 30098 15036 30104 15088
rect 30156 15076 30162 15088
rect 31297 15079 31355 15085
rect 31297 15076 31309 15079
rect 30156 15048 31309 15076
rect 30156 15036 30162 15048
rect 31297 15045 31309 15048
rect 31343 15045 31355 15079
rect 31297 15039 31355 15045
rect 2133 15011 2191 15017
rect 2133 14977 2145 15011
rect 2179 14977 2191 15011
rect 2133 14971 2191 14977
rect 2777 15011 2835 15017
rect 2777 14977 2789 15011
rect 2823 15008 2835 15011
rect 2866 15008 2872 15020
rect 2823 14980 2872 15008
rect 2823 14977 2835 14980
rect 2777 14971 2835 14977
rect 2148 14940 2176 14971
rect 2866 14968 2872 14980
rect 2924 14968 2930 15020
rect 22002 15008 22008 15020
rect 6886 14980 22008 15008
rect 6886 14940 6914 14980
rect 22002 14968 22008 14980
rect 22060 14968 22066 15020
rect 24762 15008 24768 15020
rect 24723 14980 24768 15008
rect 24762 14968 24768 14980
rect 24820 14968 24826 15020
rect 25406 15008 25412 15020
rect 25367 14980 25412 15008
rect 25406 14968 25412 14980
rect 25464 14968 25470 15020
rect 25590 15008 25596 15020
rect 25551 14980 25596 15008
rect 25590 14968 25596 14980
rect 25648 14968 25654 15020
rect 25774 14968 25780 15020
rect 25832 15008 25838 15020
rect 26053 15011 26111 15017
rect 26053 15008 26065 15011
rect 25832 14980 26065 15008
rect 25832 14968 25838 14980
rect 26053 14977 26065 14980
rect 26099 14977 26111 15011
rect 26053 14971 26111 14977
rect 26142 14968 26148 15020
rect 26200 15008 26206 15020
rect 27157 15011 27215 15017
rect 27157 15008 27169 15011
rect 26200 14980 27169 15008
rect 26200 14968 26206 14980
rect 27157 14977 27169 14980
rect 27203 14977 27215 15011
rect 27157 14971 27215 14977
rect 27798 14968 27804 15020
rect 27856 15008 27862 15020
rect 27985 15011 28043 15017
rect 27985 15008 27997 15011
rect 27856 14980 27997 15008
rect 27856 14968 27862 14980
rect 27985 14977 27997 14980
rect 28031 14977 28043 15011
rect 27985 14971 28043 14977
rect 28166 14968 28172 15020
rect 28224 15008 28230 15020
rect 28629 15011 28687 15017
rect 28629 15008 28641 15011
rect 28224 14980 28641 15008
rect 28224 14968 28230 14980
rect 28629 14977 28641 14980
rect 28675 14977 28687 15011
rect 28810 15008 28816 15020
rect 28771 14980 28816 15008
rect 28629 14971 28687 14977
rect 28810 14968 28816 14980
rect 28868 14968 28874 15020
rect 29273 15011 29331 15017
rect 29273 14977 29285 15011
rect 29319 14977 29331 15011
rect 29273 14971 29331 14977
rect 29917 15011 29975 15017
rect 29917 14977 29929 15011
rect 29963 15008 29975 15011
rect 30926 15008 30932 15020
rect 29963 14980 30932 15008
rect 29963 14977 29975 14980
rect 29917 14971 29975 14977
rect 2148 14912 6914 14940
rect 15286 14900 15292 14952
rect 15344 14940 15350 14952
rect 28994 14940 29000 14952
rect 15344 14912 29000 14940
rect 15344 14900 15350 14912
rect 28994 14900 29000 14912
rect 29052 14940 29058 14952
rect 29288 14940 29316 14971
rect 30926 14968 30932 14980
rect 30984 14968 30990 15020
rect 31205 15011 31263 15017
rect 31205 14977 31217 15011
rect 31251 15008 31263 15011
rect 31662 15008 31668 15020
rect 31251 14980 31668 15008
rect 31251 14977 31263 14980
rect 31205 14971 31263 14977
rect 31662 14968 31668 14980
rect 31720 14968 31726 15020
rect 32309 15011 32367 15017
rect 32309 14977 32321 15011
rect 32355 15008 32367 15011
rect 32766 15008 32772 15020
rect 32355 14980 32772 15008
rect 32355 14977 32367 14980
rect 32309 14971 32367 14977
rect 32766 14968 32772 14980
rect 32824 14968 32830 15020
rect 32953 15011 33011 15017
rect 32953 14977 32965 15011
rect 32999 15008 33011 15011
rect 33594 15008 33600 15020
rect 32999 14980 33600 15008
rect 32999 14977 33011 14980
rect 32953 14971 33011 14977
rect 33594 14968 33600 14980
rect 33652 14968 33658 15020
rect 33778 15008 33784 15020
rect 33739 14980 33784 15008
rect 33778 14968 33784 14980
rect 33836 14968 33842 15020
rect 29052 14912 29316 14940
rect 30745 14943 30803 14949
rect 29052 14900 29058 14912
rect 30745 14909 30757 14943
rect 30791 14940 30803 14943
rect 32122 14940 32128 14952
rect 30791 14912 32128 14940
rect 30791 14909 30803 14912
rect 30745 14903 30803 14909
rect 32122 14900 32128 14912
rect 32180 14900 32186 14952
rect 1762 14764 1768 14816
rect 1820 14804 1826 14816
rect 2869 14807 2927 14813
rect 2869 14804 2881 14807
rect 1820 14776 2881 14804
rect 1820 14764 1826 14776
rect 2869 14773 2881 14776
rect 2915 14773 2927 14807
rect 2869 14767 2927 14773
rect 1104 14714 34868 14736
rect 1104 14662 5170 14714
rect 5222 14662 5234 14714
rect 5286 14662 5298 14714
rect 5350 14662 5362 14714
rect 5414 14662 5426 14714
rect 5478 14662 13611 14714
rect 13663 14662 13675 14714
rect 13727 14662 13739 14714
rect 13791 14662 13803 14714
rect 13855 14662 13867 14714
rect 13919 14662 22052 14714
rect 22104 14662 22116 14714
rect 22168 14662 22180 14714
rect 22232 14662 22244 14714
rect 22296 14662 22308 14714
rect 22360 14662 30493 14714
rect 30545 14662 30557 14714
rect 30609 14662 30621 14714
rect 30673 14662 30685 14714
rect 30737 14662 30749 14714
rect 30801 14662 34868 14714
rect 1104 14640 34868 14662
rect 26605 14603 26663 14609
rect 26605 14569 26617 14603
rect 26651 14600 26663 14603
rect 26694 14600 26700 14612
rect 26651 14572 26700 14600
rect 26651 14569 26663 14572
rect 26605 14563 26663 14569
rect 26694 14560 26700 14572
rect 26752 14560 26758 14612
rect 31018 14600 31024 14612
rect 30979 14572 31024 14600
rect 31018 14560 31024 14572
rect 31076 14560 31082 14612
rect 31757 14603 31815 14609
rect 31757 14569 31769 14603
rect 31803 14600 31815 14603
rect 32490 14600 32496 14612
rect 31803 14572 32496 14600
rect 31803 14569 31815 14572
rect 31757 14563 31815 14569
rect 32490 14560 32496 14572
rect 32548 14560 32554 14612
rect 26053 14535 26111 14541
rect 26053 14501 26065 14535
rect 26099 14532 26111 14535
rect 27430 14532 27436 14544
rect 26099 14504 27436 14532
rect 26099 14501 26111 14504
rect 26053 14495 26111 14501
rect 27430 14492 27436 14504
rect 27488 14492 27494 14544
rect 1762 14464 1768 14476
rect 1723 14436 1768 14464
rect 1762 14424 1768 14436
rect 1820 14424 1826 14476
rect 2774 14464 2780 14476
rect 2735 14436 2780 14464
rect 2774 14424 2780 14436
rect 2832 14424 2838 14476
rect 30469 14467 30527 14473
rect 30469 14433 30481 14467
rect 30515 14464 30527 14467
rect 32493 14467 32551 14473
rect 32493 14464 32505 14467
rect 30515 14436 32505 14464
rect 30515 14433 30527 14436
rect 30469 14427 30527 14433
rect 32493 14433 32505 14436
rect 32539 14433 32551 14467
rect 32493 14427 32551 14433
rect 1578 14396 1584 14408
rect 1539 14368 1584 14396
rect 1578 14356 1584 14368
rect 1636 14356 1642 14408
rect 25133 14399 25191 14405
rect 25133 14365 25145 14399
rect 25179 14396 25191 14399
rect 25498 14396 25504 14408
rect 25179 14368 25504 14396
rect 25179 14365 25191 14368
rect 25133 14359 25191 14365
rect 25498 14356 25504 14368
rect 25556 14356 25562 14408
rect 25958 14396 25964 14408
rect 25919 14368 25964 14396
rect 25958 14356 25964 14368
rect 26016 14356 26022 14408
rect 26602 14396 26608 14408
rect 26563 14368 26608 14396
rect 26602 14356 26608 14368
rect 26660 14356 26666 14408
rect 26789 14399 26847 14405
rect 26789 14365 26801 14399
rect 26835 14396 26847 14399
rect 26878 14396 26884 14408
rect 26835 14368 26884 14396
rect 26835 14365 26847 14368
rect 26789 14359 26847 14365
rect 26878 14356 26884 14368
rect 26936 14356 26942 14408
rect 30929 14399 30987 14405
rect 30929 14365 30941 14399
rect 30975 14396 30987 14399
rect 34330 14396 34336 14408
rect 30975 14368 31754 14396
rect 34291 14368 34336 14396
rect 30975 14365 30987 14368
rect 30929 14359 30987 14365
rect 25225 14331 25283 14337
rect 25225 14297 25237 14331
rect 25271 14328 25283 14331
rect 26050 14328 26056 14340
rect 25271 14300 26056 14328
rect 25271 14297 25283 14300
rect 25225 14291 25283 14297
rect 26050 14288 26056 14300
rect 26108 14288 26114 14340
rect 31726 14260 31754 14368
rect 34330 14356 34336 14368
rect 34388 14356 34394 14408
rect 32674 14328 32680 14340
rect 32635 14300 32680 14328
rect 32674 14288 32680 14300
rect 32732 14288 32738 14340
rect 33502 14260 33508 14272
rect 31726 14232 33508 14260
rect 33502 14220 33508 14232
rect 33560 14220 33566 14272
rect 1104 14170 35027 14192
rect 1104 14118 9390 14170
rect 9442 14118 9454 14170
rect 9506 14118 9518 14170
rect 9570 14118 9582 14170
rect 9634 14118 9646 14170
rect 9698 14118 17831 14170
rect 17883 14118 17895 14170
rect 17947 14118 17959 14170
rect 18011 14118 18023 14170
rect 18075 14118 18087 14170
rect 18139 14118 26272 14170
rect 26324 14118 26336 14170
rect 26388 14118 26400 14170
rect 26452 14118 26464 14170
rect 26516 14118 26528 14170
rect 26580 14118 34713 14170
rect 34765 14118 34777 14170
rect 34829 14118 34841 14170
rect 34893 14118 34905 14170
rect 34957 14118 34969 14170
rect 35021 14118 35027 14170
rect 1104 14096 35027 14118
rect 30377 14059 30435 14065
rect 30377 14025 30389 14059
rect 30423 14056 30435 14059
rect 30834 14056 30840 14068
rect 30423 14028 30840 14056
rect 30423 14025 30435 14028
rect 30377 14019 30435 14025
rect 30834 14016 30840 14028
rect 30892 14016 30898 14068
rect 31386 14016 31392 14068
rect 31444 14056 31450 14068
rect 31665 14059 31723 14065
rect 31665 14056 31677 14059
rect 31444 14028 31677 14056
rect 31444 14016 31450 14028
rect 31665 14025 31677 14028
rect 31711 14025 31723 14059
rect 31665 14019 31723 14025
rect 31021 13991 31079 13997
rect 31021 13957 31033 13991
rect 31067 13988 31079 13991
rect 32677 13991 32735 13997
rect 32677 13988 32689 13991
rect 31067 13960 32689 13988
rect 31067 13957 31079 13960
rect 31021 13951 31079 13957
rect 32677 13957 32689 13960
rect 32723 13957 32735 13991
rect 32677 13951 32735 13957
rect 30282 13920 30288 13932
rect 30243 13892 30288 13920
rect 30282 13880 30288 13892
rect 30340 13880 30346 13932
rect 30926 13920 30932 13932
rect 30887 13892 30932 13920
rect 30926 13880 30932 13892
rect 30984 13880 30990 13932
rect 31570 13920 31576 13932
rect 31531 13892 31576 13920
rect 31570 13880 31576 13892
rect 31628 13880 31634 13932
rect 1762 13852 1768 13864
rect 1723 13824 1768 13852
rect 1762 13812 1768 13824
rect 1820 13812 1826 13864
rect 1946 13852 1952 13864
rect 1907 13824 1952 13852
rect 1946 13812 1952 13824
rect 2004 13812 2010 13864
rect 2774 13852 2780 13864
rect 2735 13824 2780 13852
rect 2774 13812 2780 13824
rect 2832 13812 2838 13864
rect 32490 13852 32496 13864
rect 32451 13824 32496 13852
rect 32490 13812 32496 13824
rect 32548 13812 32554 13864
rect 34330 13852 34336 13864
rect 34291 13824 34336 13852
rect 34330 13812 34336 13824
rect 34388 13812 34394 13864
rect 1104 13626 34868 13648
rect 1104 13574 5170 13626
rect 5222 13574 5234 13626
rect 5286 13574 5298 13626
rect 5350 13574 5362 13626
rect 5414 13574 5426 13626
rect 5478 13574 13611 13626
rect 13663 13574 13675 13626
rect 13727 13574 13739 13626
rect 13791 13574 13803 13626
rect 13855 13574 13867 13626
rect 13919 13574 22052 13626
rect 22104 13574 22116 13626
rect 22168 13574 22180 13626
rect 22232 13574 22244 13626
rect 22296 13574 22308 13626
rect 22360 13574 30493 13626
rect 30545 13574 30557 13626
rect 30609 13574 30621 13626
rect 30673 13574 30685 13626
rect 30737 13574 30749 13626
rect 30801 13574 34868 13626
rect 1104 13552 34868 13574
rect 1762 13472 1768 13524
rect 1820 13512 1826 13524
rect 2685 13515 2743 13521
rect 2685 13512 2697 13515
rect 1820 13484 2697 13512
rect 1820 13472 1826 13484
rect 2685 13481 2697 13484
rect 2731 13481 2743 13515
rect 31202 13512 31208 13524
rect 31163 13484 31208 13512
rect 2685 13475 2743 13481
rect 31202 13472 31208 13484
rect 31260 13472 31266 13524
rect 31846 13512 31852 13524
rect 31807 13484 31852 13512
rect 31846 13472 31852 13484
rect 31904 13472 31910 13524
rect 32582 13512 32588 13524
rect 32543 13484 32588 13512
rect 32582 13472 32588 13484
rect 32640 13472 32646 13524
rect 33594 13512 33600 13524
rect 33555 13484 33600 13512
rect 33594 13472 33600 13484
rect 33652 13472 33658 13524
rect 1578 13404 1584 13456
rect 1636 13444 1642 13456
rect 2041 13447 2099 13453
rect 2041 13444 2053 13447
rect 1636 13416 2053 13444
rect 1636 13404 1642 13416
rect 2041 13413 2053 13416
rect 2087 13413 2099 13447
rect 2041 13407 2099 13413
rect 30374 13268 30380 13320
rect 30432 13308 30438 13320
rect 31113 13311 31171 13317
rect 31113 13308 31125 13311
rect 30432 13280 31125 13308
rect 30432 13268 30438 13280
rect 31113 13277 31125 13280
rect 31159 13277 31171 13311
rect 31113 13271 31171 13277
rect 31754 13268 31760 13320
rect 31812 13308 31818 13320
rect 33778 13308 33784 13320
rect 31812 13280 31857 13308
rect 33739 13280 33784 13308
rect 31812 13268 31818 13280
rect 33778 13268 33784 13280
rect 33836 13268 33842 13320
rect 1104 13082 35027 13104
rect 1104 13030 9390 13082
rect 9442 13030 9454 13082
rect 9506 13030 9518 13082
rect 9570 13030 9582 13082
rect 9634 13030 9646 13082
rect 9698 13030 17831 13082
rect 17883 13030 17895 13082
rect 17947 13030 17959 13082
rect 18011 13030 18023 13082
rect 18075 13030 18087 13082
rect 18139 13030 26272 13082
rect 26324 13030 26336 13082
rect 26388 13030 26400 13082
rect 26452 13030 26464 13082
rect 26516 13030 26528 13082
rect 26580 13030 34713 13082
rect 34765 13030 34777 13082
rect 34829 13030 34841 13082
rect 34893 13030 34905 13082
rect 34957 13030 34969 13082
rect 35021 13030 35027 13082
rect 1104 13008 35027 13030
rect 1946 12928 1952 12980
rect 2004 12968 2010 12980
rect 2133 12971 2191 12977
rect 2133 12968 2145 12971
rect 2004 12940 2145 12968
rect 2004 12928 2010 12940
rect 2133 12937 2145 12940
rect 2179 12937 2191 12971
rect 2133 12931 2191 12937
rect 34330 12900 34336 12912
rect 34291 12872 34336 12900
rect 34330 12860 34336 12872
rect 34388 12860 34394 12912
rect 2041 12835 2099 12841
rect 2041 12801 2053 12835
rect 2087 12832 2099 12835
rect 2222 12832 2228 12844
rect 2087 12804 2228 12832
rect 2087 12801 2099 12804
rect 2041 12795 2099 12801
rect 2222 12792 2228 12804
rect 2280 12832 2286 12844
rect 2682 12832 2688 12844
rect 2280 12804 2688 12832
rect 2280 12792 2286 12804
rect 2682 12792 2688 12804
rect 2740 12832 2746 12844
rect 30926 12832 30932 12844
rect 2740 12804 30932 12832
rect 2740 12792 2746 12804
rect 30926 12792 30932 12804
rect 30984 12832 30990 12844
rect 31478 12832 31484 12844
rect 30984 12804 31484 12832
rect 30984 12792 30990 12804
rect 31478 12792 31484 12804
rect 31536 12792 31542 12844
rect 31389 12767 31447 12773
rect 31389 12733 31401 12767
rect 31435 12764 31447 12767
rect 32493 12767 32551 12773
rect 32493 12764 32505 12767
rect 31435 12736 32505 12764
rect 31435 12733 31447 12736
rect 31389 12727 31447 12733
rect 32493 12733 32505 12736
rect 32539 12733 32551 12767
rect 32493 12727 32551 12733
rect 32677 12767 32735 12773
rect 32677 12733 32689 12767
rect 32723 12764 32735 12767
rect 33134 12764 33140 12776
rect 32723 12736 33140 12764
rect 32723 12733 32735 12736
rect 32677 12727 32735 12733
rect 33134 12724 33140 12736
rect 33192 12724 33198 12776
rect 1104 12538 34868 12560
rect 1104 12486 5170 12538
rect 5222 12486 5234 12538
rect 5286 12486 5298 12538
rect 5350 12486 5362 12538
rect 5414 12486 5426 12538
rect 5478 12486 13611 12538
rect 13663 12486 13675 12538
rect 13727 12486 13739 12538
rect 13791 12486 13803 12538
rect 13855 12486 13867 12538
rect 13919 12486 22052 12538
rect 22104 12486 22116 12538
rect 22168 12486 22180 12538
rect 22232 12486 22244 12538
rect 22296 12486 22308 12538
rect 22360 12486 30493 12538
rect 30545 12486 30557 12538
rect 30609 12486 30621 12538
rect 30673 12486 30685 12538
rect 30737 12486 30749 12538
rect 30801 12486 34868 12538
rect 1104 12464 34868 12486
rect 32033 12427 32091 12433
rect 32033 12393 32045 12427
rect 32079 12424 32091 12427
rect 32490 12424 32496 12436
rect 32079 12396 32496 12424
rect 32079 12393 32091 12396
rect 32033 12387 32091 12393
rect 32490 12384 32496 12396
rect 32548 12384 32554 12436
rect 32493 12291 32551 12297
rect 32493 12257 32505 12291
rect 32539 12288 32551 12291
rect 33318 12288 33324 12300
rect 32539 12260 33324 12288
rect 32539 12257 32551 12260
rect 32493 12251 32551 12257
rect 33318 12248 33324 12260
rect 33376 12248 33382 12300
rect 34330 12288 34336 12300
rect 34291 12260 34336 12288
rect 34330 12248 34336 12260
rect 34388 12248 34394 12300
rect 2041 12223 2099 12229
rect 2041 12189 2053 12223
rect 2087 12220 2099 12223
rect 2130 12220 2136 12232
rect 2087 12192 2136 12220
rect 2087 12189 2099 12192
rect 2041 12183 2099 12189
rect 2130 12180 2136 12192
rect 2188 12220 2194 12232
rect 14366 12220 14372 12232
rect 2188 12192 14372 12220
rect 2188 12180 2194 12192
rect 14366 12180 14372 12192
rect 14424 12180 14430 12232
rect 31205 12223 31263 12229
rect 31205 12189 31217 12223
rect 31251 12220 31263 12223
rect 31570 12220 31576 12232
rect 31251 12192 31576 12220
rect 31251 12189 31263 12192
rect 31205 12183 31263 12189
rect 31570 12180 31576 12192
rect 31628 12180 31634 12232
rect 31297 12155 31355 12161
rect 31297 12121 31309 12155
rect 31343 12152 31355 12155
rect 32677 12155 32735 12161
rect 32677 12152 32689 12155
rect 31343 12124 32689 12152
rect 31343 12121 31355 12124
rect 31297 12115 31355 12121
rect 32677 12121 32689 12124
rect 32723 12121 32735 12155
rect 32677 12115 32735 12121
rect 1946 12044 1952 12096
rect 2004 12084 2010 12096
rect 2133 12087 2191 12093
rect 2133 12084 2145 12087
rect 2004 12056 2145 12084
rect 2004 12044 2010 12056
rect 2133 12053 2145 12056
rect 2179 12053 2191 12087
rect 2133 12047 2191 12053
rect 1104 11994 35027 12016
rect 1104 11942 9390 11994
rect 9442 11942 9454 11994
rect 9506 11942 9518 11994
rect 9570 11942 9582 11994
rect 9634 11942 9646 11994
rect 9698 11942 17831 11994
rect 17883 11942 17895 11994
rect 17947 11942 17959 11994
rect 18011 11942 18023 11994
rect 18075 11942 18087 11994
rect 18139 11942 26272 11994
rect 26324 11942 26336 11994
rect 26388 11942 26400 11994
rect 26452 11942 26464 11994
rect 26516 11942 26528 11994
rect 26580 11942 34713 11994
rect 34765 11942 34777 11994
rect 34829 11942 34841 11994
rect 34893 11942 34905 11994
rect 34957 11942 34969 11994
rect 35021 11942 35027 11994
rect 1104 11920 35027 11942
rect 1946 11812 1952 11824
rect 1907 11784 1952 11812
rect 1946 11772 1952 11784
rect 2004 11772 2010 11824
rect 32677 11747 32735 11753
rect 32677 11713 32689 11747
rect 32723 11744 32735 11747
rect 32858 11744 32864 11756
rect 32723 11716 32864 11744
rect 32723 11713 32735 11716
rect 32677 11707 32735 11713
rect 32858 11704 32864 11716
rect 32916 11704 32922 11756
rect 33226 11704 33232 11756
rect 33284 11744 33290 11756
rect 33321 11747 33379 11753
rect 33321 11744 33333 11747
rect 33284 11716 33333 11744
rect 33284 11704 33290 11716
rect 33321 11713 33333 11716
rect 33367 11713 33379 11747
rect 33962 11744 33968 11756
rect 33923 11716 33968 11744
rect 33321 11707 33379 11713
rect 33962 11704 33968 11716
rect 34020 11704 34026 11756
rect 1765 11679 1823 11685
rect 1765 11645 1777 11679
rect 1811 11676 1823 11679
rect 2038 11676 2044 11688
rect 1811 11648 2044 11676
rect 1811 11645 1823 11648
rect 1765 11639 1823 11645
rect 2038 11636 2044 11648
rect 2096 11636 2102 11688
rect 2774 11676 2780 11688
rect 2735 11648 2780 11676
rect 2774 11636 2780 11648
rect 2832 11636 2838 11688
rect 1104 11450 34868 11472
rect 1104 11398 5170 11450
rect 5222 11398 5234 11450
rect 5286 11398 5298 11450
rect 5350 11398 5362 11450
rect 5414 11398 5426 11450
rect 5478 11398 13611 11450
rect 13663 11398 13675 11450
rect 13727 11398 13739 11450
rect 13791 11398 13803 11450
rect 13855 11398 13867 11450
rect 13919 11398 22052 11450
rect 22104 11398 22116 11450
rect 22168 11398 22180 11450
rect 22232 11398 22244 11450
rect 22296 11398 22308 11450
rect 22360 11398 30493 11450
rect 30545 11398 30557 11450
rect 30609 11398 30621 11450
rect 30673 11398 30685 11450
rect 30737 11398 30749 11450
rect 30801 11398 34868 11450
rect 1104 11376 34868 11398
rect 2038 11336 2044 11348
rect 1999 11308 2044 11336
rect 2038 11296 2044 11308
rect 2096 11296 2102 11348
rect 33134 11296 33140 11348
rect 33192 11336 33198 11348
rect 33229 11339 33287 11345
rect 33229 11336 33241 11339
rect 33192 11308 33241 11336
rect 33192 11296 33198 11308
rect 33229 11305 33241 11308
rect 33275 11305 33287 11339
rect 33229 11299 33287 11305
rect 33410 11296 33416 11348
rect 33468 11336 33474 11348
rect 33965 11339 34023 11345
rect 33965 11336 33977 11339
rect 33468 11308 33977 11336
rect 33468 11296 33474 11308
rect 33965 11305 33977 11308
rect 34011 11305 34023 11339
rect 33965 11299 34023 11305
rect 1762 11092 1768 11144
rect 1820 11132 1826 11144
rect 2685 11135 2743 11141
rect 2685 11132 2697 11135
rect 1820 11104 2697 11132
rect 1820 11092 1826 11104
rect 2685 11101 2697 11104
rect 2731 11101 2743 11135
rect 2685 11095 2743 11101
rect 33137 11135 33195 11141
rect 33137 11101 33149 11135
rect 33183 11132 33195 11135
rect 33502 11132 33508 11144
rect 33183 11104 33508 11132
rect 33183 11101 33195 11104
rect 33137 11095 33195 11101
rect 33502 11092 33508 11104
rect 33560 11092 33566 11144
rect 1104 10906 35027 10928
rect 1104 10854 9390 10906
rect 9442 10854 9454 10906
rect 9506 10854 9518 10906
rect 9570 10854 9582 10906
rect 9634 10854 9646 10906
rect 9698 10854 17831 10906
rect 17883 10854 17895 10906
rect 17947 10854 17959 10906
rect 18011 10854 18023 10906
rect 18075 10854 18087 10906
rect 18139 10854 26272 10906
rect 26324 10854 26336 10906
rect 26388 10854 26400 10906
rect 26452 10854 26464 10906
rect 26516 10854 26528 10906
rect 26580 10854 34713 10906
rect 34765 10854 34777 10906
rect 34829 10854 34841 10906
rect 34893 10854 34905 10906
rect 34957 10854 34969 10906
rect 35021 10854 35027 10906
rect 1104 10832 35027 10854
rect 32674 10752 32680 10804
rect 32732 10792 32738 10804
rect 33873 10795 33931 10801
rect 33873 10792 33885 10795
rect 32732 10764 33885 10792
rect 32732 10752 32738 10764
rect 33873 10761 33885 10764
rect 33919 10761 33931 10795
rect 33873 10755 33931 10761
rect 1762 10656 1768 10668
rect 1723 10628 1768 10656
rect 1762 10616 1768 10628
rect 1820 10616 1826 10668
rect 33318 10656 33324 10668
rect 33279 10628 33324 10656
rect 33318 10616 33324 10628
rect 33376 10616 33382 10668
rect 33781 10659 33839 10665
rect 33781 10625 33793 10659
rect 33827 10625 33839 10659
rect 33781 10619 33839 10625
rect 1949 10591 2007 10597
rect 1949 10557 1961 10591
rect 1995 10588 2007 10591
rect 2038 10588 2044 10600
rect 1995 10560 2044 10588
rect 1995 10557 2007 10560
rect 1949 10551 2007 10557
rect 2038 10548 2044 10560
rect 2096 10548 2102 10600
rect 2774 10588 2780 10600
rect 2735 10560 2780 10588
rect 2774 10548 2780 10560
rect 2832 10548 2838 10600
rect 31478 10548 31484 10600
rect 31536 10588 31542 10600
rect 33796 10588 33824 10619
rect 31536 10560 33824 10588
rect 31536 10548 31542 10560
rect 1104 10362 34868 10384
rect 1104 10310 5170 10362
rect 5222 10310 5234 10362
rect 5286 10310 5298 10362
rect 5350 10310 5362 10362
rect 5414 10310 5426 10362
rect 5478 10310 13611 10362
rect 13663 10310 13675 10362
rect 13727 10310 13739 10362
rect 13791 10310 13803 10362
rect 13855 10310 13867 10362
rect 13919 10310 22052 10362
rect 22104 10310 22116 10362
rect 22168 10310 22180 10362
rect 22232 10310 22244 10362
rect 22296 10310 22308 10362
rect 22360 10310 30493 10362
rect 30545 10310 30557 10362
rect 30609 10310 30621 10362
rect 30673 10310 30685 10362
rect 30737 10310 30749 10362
rect 30801 10310 34868 10362
rect 1104 10288 34868 10310
rect 2038 10248 2044 10260
rect 1999 10220 2044 10248
rect 2038 10208 2044 10220
rect 2096 10208 2102 10260
rect 34238 10248 34244 10260
rect 34199 10220 34244 10248
rect 34238 10208 34244 10220
rect 34296 10208 34302 10260
rect 1949 10047 2007 10053
rect 1949 10013 1961 10047
rect 1995 10044 2007 10047
rect 4706 10044 4712 10056
rect 1995 10016 4712 10044
rect 1995 10013 2007 10016
rect 1949 10007 2007 10013
rect 4706 10004 4712 10016
rect 4764 10004 4770 10056
rect 34054 10044 34060 10056
rect 34015 10016 34060 10044
rect 34054 10004 34060 10016
rect 34112 10004 34118 10056
rect 1104 9818 35027 9840
rect 1104 9766 9390 9818
rect 9442 9766 9454 9818
rect 9506 9766 9518 9818
rect 9570 9766 9582 9818
rect 9634 9766 9646 9818
rect 9698 9766 17831 9818
rect 17883 9766 17895 9818
rect 17947 9766 17959 9818
rect 18011 9766 18023 9818
rect 18075 9766 18087 9818
rect 18139 9766 26272 9818
rect 26324 9766 26336 9818
rect 26388 9766 26400 9818
rect 26452 9766 26464 9818
rect 26516 9766 26528 9818
rect 26580 9766 34713 9818
rect 34765 9766 34777 9818
rect 34829 9766 34841 9818
rect 34893 9766 34905 9818
rect 34957 9766 34969 9818
rect 35021 9766 35027 9818
rect 1104 9744 35027 9766
rect 2501 9571 2559 9577
rect 2501 9537 2513 9571
rect 2547 9568 2559 9571
rect 2866 9568 2872 9580
rect 2547 9540 2872 9568
rect 2547 9537 2559 9540
rect 2501 9531 2559 9537
rect 2866 9528 2872 9540
rect 2924 9568 2930 9580
rect 9122 9568 9128 9580
rect 2924 9540 9128 9568
rect 2924 9528 2930 9540
rect 9122 9528 9128 9540
rect 9180 9528 9186 9580
rect 1578 9324 1584 9376
rect 1636 9364 1642 9376
rect 2041 9367 2099 9373
rect 2041 9364 2053 9367
rect 1636 9336 2053 9364
rect 1636 9324 1642 9336
rect 2041 9333 2053 9336
rect 2087 9333 2099 9367
rect 2590 9364 2596 9376
rect 2551 9336 2596 9364
rect 2041 9327 2099 9333
rect 2590 9324 2596 9336
rect 2648 9324 2654 9376
rect 1104 9274 34868 9296
rect 1104 9222 5170 9274
rect 5222 9222 5234 9274
rect 5286 9222 5298 9274
rect 5350 9222 5362 9274
rect 5414 9222 5426 9274
rect 5478 9222 13611 9274
rect 13663 9222 13675 9274
rect 13727 9222 13739 9274
rect 13791 9222 13803 9274
rect 13855 9222 13867 9274
rect 13919 9222 22052 9274
rect 22104 9222 22116 9274
rect 22168 9222 22180 9274
rect 22232 9222 22244 9274
rect 22296 9222 22308 9274
rect 22360 9222 30493 9274
rect 30545 9222 30557 9274
rect 30609 9222 30621 9274
rect 30673 9222 30685 9274
rect 30737 9222 30749 9274
rect 30801 9222 34868 9274
rect 1104 9200 34868 9222
rect 1578 9024 1584 9036
rect 1539 8996 1584 9024
rect 1578 8984 1584 8996
rect 1636 8984 1642 9036
rect 1765 9027 1823 9033
rect 1765 8993 1777 9027
rect 1811 9024 1823 9027
rect 2590 9024 2596 9036
rect 1811 8996 2596 9024
rect 1811 8993 1823 8996
rect 1765 8987 1823 8993
rect 2590 8984 2596 8996
rect 2648 8984 2654 9036
rect 2774 9024 2780 9036
rect 2735 8996 2780 9024
rect 2774 8984 2780 8996
rect 2832 8984 2838 9036
rect 32490 8916 32496 8968
rect 32548 8956 32554 8968
rect 33965 8959 34023 8965
rect 33965 8956 33977 8959
rect 32548 8928 33977 8956
rect 32548 8916 32554 8928
rect 33965 8925 33977 8928
rect 34011 8925 34023 8959
rect 33965 8919 34023 8925
rect 1104 8730 35027 8752
rect 1104 8678 9390 8730
rect 9442 8678 9454 8730
rect 9506 8678 9518 8730
rect 9570 8678 9582 8730
rect 9634 8678 9646 8730
rect 9698 8678 17831 8730
rect 17883 8678 17895 8730
rect 17947 8678 17959 8730
rect 18011 8678 18023 8730
rect 18075 8678 18087 8730
rect 18139 8678 26272 8730
rect 26324 8678 26336 8730
rect 26388 8678 26400 8730
rect 26452 8678 26464 8730
rect 26516 8678 26528 8730
rect 26580 8678 34713 8730
rect 34765 8678 34777 8730
rect 34829 8678 34841 8730
rect 34893 8678 34905 8730
rect 34957 8678 34969 8730
rect 35021 8678 35027 8730
rect 1104 8656 35027 8678
rect 34330 8548 34336 8560
rect 34291 8520 34336 8548
rect 34330 8508 34336 8520
rect 34388 8508 34394 8560
rect 32490 8480 32496 8492
rect 32451 8452 32496 8480
rect 32490 8440 32496 8452
rect 32548 8440 32554 8492
rect 1762 8412 1768 8424
rect 1723 8384 1768 8412
rect 1762 8372 1768 8384
rect 1820 8372 1826 8424
rect 1949 8415 2007 8421
rect 1949 8381 1961 8415
rect 1995 8412 2007 8415
rect 2590 8412 2596 8424
rect 1995 8384 2596 8412
rect 1995 8381 2007 8384
rect 1949 8375 2007 8381
rect 2590 8372 2596 8384
rect 2648 8372 2654 8424
rect 2774 8412 2780 8424
rect 2735 8384 2780 8412
rect 2774 8372 2780 8384
rect 2832 8372 2838 8424
rect 32677 8415 32735 8421
rect 32677 8381 32689 8415
rect 32723 8412 32735 8415
rect 33870 8412 33876 8424
rect 32723 8384 33876 8412
rect 32723 8381 32735 8384
rect 32677 8375 32735 8381
rect 33870 8372 33876 8384
rect 33928 8372 33934 8424
rect 1104 8186 34868 8208
rect 1104 8134 5170 8186
rect 5222 8134 5234 8186
rect 5286 8134 5298 8186
rect 5350 8134 5362 8186
rect 5414 8134 5426 8186
rect 5478 8134 13611 8186
rect 13663 8134 13675 8186
rect 13727 8134 13739 8186
rect 13791 8134 13803 8186
rect 13855 8134 13867 8186
rect 13919 8134 22052 8186
rect 22104 8134 22116 8186
rect 22168 8134 22180 8186
rect 22232 8134 22244 8186
rect 22296 8134 22308 8186
rect 22360 8134 30493 8186
rect 30545 8134 30557 8186
rect 30609 8134 30621 8186
rect 30673 8134 30685 8186
rect 30737 8134 30749 8186
rect 30801 8134 34868 8186
rect 1104 8112 34868 8134
rect 1762 8032 1768 8084
rect 1820 8072 1826 8084
rect 2041 8075 2099 8081
rect 2041 8072 2053 8075
rect 1820 8044 2053 8072
rect 1820 8032 1826 8044
rect 2041 8041 2053 8044
rect 2087 8041 2099 8075
rect 2590 8072 2596 8084
rect 2551 8044 2596 8072
rect 2041 8035 2099 8041
rect 2590 8032 2596 8044
rect 2648 8032 2654 8084
rect 31662 8032 31668 8084
rect 31720 8072 31726 8084
rect 33134 8072 33140 8084
rect 31720 8044 33140 8072
rect 31720 8032 31726 8044
rect 33134 8032 33140 8044
rect 33192 8032 33198 8084
rect 33870 8072 33876 8084
rect 33831 8044 33876 8072
rect 33870 8032 33876 8044
rect 33928 8032 33934 8084
rect 7190 7936 7196 7948
rect 2516 7908 7196 7936
rect 2516 7877 2544 7908
rect 7190 7896 7196 7908
rect 7248 7936 7254 7948
rect 7374 7936 7380 7948
rect 7248 7908 7380 7936
rect 7248 7896 7254 7908
rect 7374 7896 7380 7908
rect 7432 7896 7438 7948
rect 2501 7871 2559 7877
rect 2501 7837 2513 7871
rect 2547 7837 2559 7871
rect 2501 7831 2559 7837
rect 3329 7871 3387 7877
rect 3329 7837 3341 7871
rect 3375 7837 3387 7871
rect 33318 7868 33324 7880
rect 33279 7840 33324 7868
rect 3329 7831 3387 7837
rect 1762 7760 1768 7812
rect 1820 7800 1826 7812
rect 3344 7800 3372 7831
rect 33318 7828 33324 7840
rect 33376 7828 33382 7880
rect 33778 7868 33784 7880
rect 33739 7840 33784 7868
rect 33778 7828 33784 7840
rect 33836 7828 33842 7880
rect 1820 7772 3372 7800
rect 1820 7760 1826 7772
rect 1104 7642 35027 7664
rect 1104 7590 9390 7642
rect 9442 7590 9454 7642
rect 9506 7590 9518 7642
rect 9570 7590 9582 7642
rect 9634 7590 9646 7642
rect 9698 7590 17831 7642
rect 17883 7590 17895 7642
rect 17947 7590 17959 7642
rect 18011 7590 18023 7642
rect 18075 7590 18087 7642
rect 18139 7590 26272 7642
rect 26324 7590 26336 7642
rect 26388 7590 26400 7642
rect 26452 7590 26464 7642
rect 26516 7590 26528 7642
rect 26580 7590 34713 7642
rect 34765 7590 34777 7642
rect 34829 7590 34841 7642
rect 34893 7590 34905 7642
rect 34957 7590 34969 7642
rect 35021 7590 35027 7642
rect 1104 7568 35027 7590
rect 1762 7392 1768 7404
rect 1723 7364 1768 7392
rect 1762 7352 1768 7364
rect 1820 7352 1826 7404
rect 33137 7395 33195 7401
rect 33137 7361 33149 7395
rect 33183 7392 33195 7395
rect 33502 7392 33508 7404
rect 33183 7364 33508 7392
rect 33183 7361 33195 7364
rect 33137 7355 33195 7361
rect 33502 7352 33508 7364
rect 33560 7352 33566 7404
rect 1946 7324 1952 7336
rect 1907 7296 1952 7324
rect 1946 7284 1952 7296
rect 2004 7284 2010 7336
rect 2774 7324 2780 7336
rect 2735 7296 2780 7324
rect 2774 7284 2780 7296
rect 2832 7284 2838 7336
rect 4246 7188 4252 7200
rect 4207 7160 4252 7188
rect 4246 7148 4252 7160
rect 4304 7148 4310 7200
rect 33226 7188 33232 7200
rect 33187 7160 33232 7188
rect 33226 7148 33232 7160
rect 33284 7148 33290 7200
rect 33962 7188 33968 7200
rect 33923 7160 33968 7188
rect 33962 7148 33968 7160
rect 34020 7148 34026 7200
rect 1104 7098 34868 7120
rect 1104 7046 5170 7098
rect 5222 7046 5234 7098
rect 5286 7046 5298 7098
rect 5350 7046 5362 7098
rect 5414 7046 5426 7098
rect 5478 7046 13611 7098
rect 13663 7046 13675 7098
rect 13727 7046 13739 7098
rect 13791 7046 13803 7098
rect 13855 7046 13867 7098
rect 13919 7046 22052 7098
rect 22104 7046 22116 7098
rect 22168 7046 22180 7098
rect 22232 7046 22244 7098
rect 22296 7046 22308 7098
rect 22360 7046 30493 7098
rect 30545 7046 30557 7098
rect 30609 7046 30621 7098
rect 30673 7046 30685 7098
rect 30737 7046 30749 7098
rect 30801 7046 34868 7098
rect 1104 7024 34868 7046
rect 1946 6944 1952 6996
rect 2004 6984 2010 6996
rect 2133 6987 2191 6993
rect 2133 6984 2145 6987
rect 2004 6956 2145 6984
rect 2004 6944 2010 6956
rect 2133 6953 2145 6956
rect 2179 6953 2191 6987
rect 2133 6947 2191 6953
rect 32677 6851 32735 6857
rect 32677 6817 32689 6851
rect 32723 6848 32735 6851
rect 33226 6848 33232 6860
rect 32723 6820 33232 6848
rect 32723 6817 32735 6820
rect 32677 6811 32735 6817
rect 33226 6808 33232 6820
rect 33284 6808 33290 6860
rect 34330 6848 34336 6860
rect 34291 6820 34336 6848
rect 34330 6808 34336 6820
rect 34388 6808 34394 6860
rect 2041 6783 2099 6789
rect 2041 6749 2053 6783
rect 2087 6780 2099 6783
rect 2314 6780 2320 6792
rect 2087 6752 2320 6780
rect 2087 6749 2099 6752
rect 2041 6743 2099 6749
rect 2314 6740 2320 6752
rect 2372 6740 2378 6792
rect 2682 6780 2688 6792
rect 2643 6752 2688 6780
rect 2682 6740 2688 6752
rect 2740 6740 2746 6792
rect 4157 6783 4215 6789
rect 4157 6749 4169 6783
rect 4203 6749 4215 6783
rect 4157 6743 4215 6749
rect 1762 6672 1768 6724
rect 1820 6712 1826 6724
rect 4172 6712 4200 6743
rect 4338 6740 4344 6792
rect 4396 6780 4402 6792
rect 4617 6783 4675 6789
rect 4617 6780 4629 6783
rect 4396 6752 4629 6780
rect 4396 6740 4402 6752
rect 4617 6749 4629 6752
rect 4663 6749 4675 6783
rect 4617 6743 4675 6749
rect 4890 6740 4896 6792
rect 4948 6780 4954 6792
rect 5445 6783 5503 6789
rect 5445 6780 5457 6783
rect 4948 6752 5457 6780
rect 4948 6740 4954 6752
rect 5445 6749 5457 6752
rect 5491 6749 5503 6783
rect 5445 6743 5503 6749
rect 9122 6740 9128 6792
rect 9180 6780 9186 6792
rect 9309 6783 9367 6789
rect 9309 6780 9321 6783
rect 9180 6752 9321 6780
rect 9180 6740 9186 6752
rect 9309 6749 9321 6752
rect 9355 6780 9367 6783
rect 19978 6780 19984 6792
rect 9355 6752 19984 6780
rect 9355 6749 9367 6752
rect 9309 6743 9367 6749
rect 19978 6740 19984 6752
rect 20036 6740 20042 6792
rect 31849 6783 31907 6789
rect 31849 6749 31861 6783
rect 31895 6780 31907 6783
rect 31938 6780 31944 6792
rect 31895 6752 31944 6780
rect 31895 6749 31907 6752
rect 31849 6743 31907 6749
rect 31938 6740 31944 6752
rect 31996 6740 32002 6792
rect 32493 6783 32551 6789
rect 32493 6749 32505 6783
rect 32539 6749 32551 6783
rect 32493 6743 32551 6749
rect 1820 6684 4200 6712
rect 1820 6672 1826 6684
rect 7190 6672 7196 6724
rect 7248 6712 7254 6724
rect 9953 6715 10011 6721
rect 9953 6712 9965 6715
rect 7248 6684 9965 6712
rect 7248 6672 7254 6684
rect 9953 6681 9965 6684
rect 9999 6712 10011 6715
rect 30282 6712 30288 6724
rect 9999 6684 30288 6712
rect 9999 6681 10011 6684
rect 9953 6675 10011 6681
rect 30282 6672 30288 6684
rect 30340 6672 30346 6724
rect 32508 6712 32536 6743
rect 33962 6712 33968 6724
rect 32508 6684 33968 6712
rect 33962 6672 33968 6684
rect 34020 6672 34026 6724
rect 1946 6604 1952 6656
rect 2004 6644 2010 6656
rect 2777 6647 2835 6653
rect 2777 6644 2789 6647
rect 2004 6616 2789 6644
rect 2004 6604 2010 6616
rect 2777 6613 2789 6616
rect 2823 6613 2835 6647
rect 2777 6607 2835 6613
rect 2958 6604 2964 6656
rect 3016 6644 3022 6656
rect 4709 6647 4767 6653
rect 4709 6644 4721 6647
rect 3016 6616 4721 6644
rect 3016 6604 3022 6616
rect 4709 6613 4721 6616
rect 4755 6613 4767 6647
rect 4709 6607 4767 6613
rect 31941 6647 31999 6653
rect 31941 6613 31953 6647
rect 31987 6644 31999 6647
rect 32674 6644 32680 6656
rect 31987 6616 32680 6644
rect 31987 6613 31999 6616
rect 31941 6607 31999 6613
rect 32674 6604 32680 6616
rect 32732 6604 32738 6656
rect 1104 6554 35027 6576
rect 1104 6502 9390 6554
rect 9442 6502 9454 6554
rect 9506 6502 9518 6554
rect 9570 6502 9582 6554
rect 9634 6502 9646 6554
rect 9698 6502 17831 6554
rect 17883 6502 17895 6554
rect 17947 6502 17959 6554
rect 18011 6502 18023 6554
rect 18075 6502 18087 6554
rect 18139 6502 26272 6554
rect 26324 6502 26336 6554
rect 26388 6502 26400 6554
rect 26452 6502 26464 6554
rect 26516 6502 26528 6554
rect 26580 6502 34713 6554
rect 34765 6502 34777 6554
rect 34829 6502 34841 6554
rect 34893 6502 34905 6554
rect 34957 6502 34969 6554
rect 35021 6502 35027 6554
rect 1104 6480 35027 6502
rect 1946 6372 1952 6384
rect 1907 6344 1952 6372
rect 1946 6332 1952 6344
rect 2004 6332 2010 6384
rect 31665 6375 31723 6381
rect 31665 6341 31677 6375
rect 31711 6372 31723 6375
rect 32677 6375 32735 6381
rect 32677 6372 32689 6375
rect 31711 6344 32689 6372
rect 31711 6341 31723 6344
rect 31665 6335 31723 6341
rect 32677 6341 32689 6344
rect 32723 6341 32735 6375
rect 32677 6335 32735 6341
rect 1762 6304 1768 6316
rect 1723 6276 1768 6304
rect 1762 6264 1768 6276
rect 1820 6264 1826 6316
rect 3878 6264 3884 6316
rect 3936 6304 3942 6316
rect 4709 6307 4767 6313
rect 4709 6304 4721 6307
rect 3936 6276 4721 6304
rect 3936 6264 3942 6276
rect 4709 6273 4721 6276
rect 4755 6304 4767 6307
rect 10502 6304 10508 6316
rect 4755 6276 10508 6304
rect 4755 6273 4767 6276
rect 4709 6267 4767 6273
rect 10502 6264 10508 6276
rect 10560 6264 10566 6316
rect 31478 6264 31484 6316
rect 31536 6304 31542 6316
rect 31573 6307 31631 6313
rect 31573 6304 31585 6307
rect 31536 6276 31585 6304
rect 31536 6264 31542 6276
rect 31573 6273 31585 6276
rect 31619 6273 31631 6307
rect 31573 6267 31631 6273
rect 2866 6236 2872 6248
rect 2827 6208 2872 6236
rect 2866 6196 2872 6208
rect 2924 6196 2930 6248
rect 32493 6239 32551 6245
rect 32493 6205 32505 6239
rect 32539 6236 32551 6239
rect 33318 6236 33324 6248
rect 32539 6208 33324 6236
rect 32539 6205 32551 6208
rect 32493 6199 32551 6205
rect 33318 6196 33324 6208
rect 33376 6196 33382 6248
rect 34330 6236 34336 6248
rect 34291 6208 34336 6236
rect 34330 6196 34336 6208
rect 34388 6196 34394 6248
rect 3050 6128 3056 6180
rect 3108 6168 3114 6180
rect 5537 6171 5595 6177
rect 5537 6168 5549 6171
rect 3108 6140 5549 6168
rect 3108 6128 3114 6140
rect 5537 6137 5549 6140
rect 5583 6137 5595 6171
rect 5537 6131 5595 6137
rect 1578 6060 1584 6112
rect 1636 6100 1642 6112
rect 4249 6103 4307 6109
rect 4249 6100 4261 6103
rect 1636 6072 4261 6100
rect 1636 6060 1642 6072
rect 4249 6069 4261 6072
rect 4295 6069 4307 6103
rect 4798 6100 4804 6112
rect 4759 6072 4804 6100
rect 4249 6063 4307 6069
rect 4798 6060 4804 6072
rect 4856 6060 4862 6112
rect 1104 6010 34868 6032
rect 1104 5958 5170 6010
rect 5222 5958 5234 6010
rect 5286 5958 5298 6010
rect 5350 5958 5362 6010
rect 5414 5958 5426 6010
rect 5478 5958 13611 6010
rect 13663 5958 13675 6010
rect 13727 5958 13739 6010
rect 13791 5958 13803 6010
rect 13855 5958 13867 6010
rect 13919 5958 22052 6010
rect 22104 5958 22116 6010
rect 22168 5958 22180 6010
rect 22232 5958 22244 6010
rect 22296 5958 22308 6010
rect 22360 5958 30493 6010
rect 30545 5958 30557 6010
rect 30609 5958 30621 6010
rect 30673 5958 30685 6010
rect 30737 5958 30749 6010
rect 30801 5958 34868 6010
rect 1104 5936 34868 5958
rect 2314 5788 2320 5840
rect 2372 5828 2378 5840
rect 2372 5800 6592 5828
rect 2372 5788 2378 5800
rect 1578 5760 1584 5772
rect 1539 5732 1584 5760
rect 1578 5720 1584 5732
rect 1636 5720 1642 5772
rect 1765 5763 1823 5769
rect 1765 5729 1777 5763
rect 1811 5760 1823 5763
rect 4065 5763 4123 5769
rect 4065 5760 4077 5763
rect 1811 5732 4077 5760
rect 1811 5729 1823 5732
rect 1765 5723 1823 5729
rect 4065 5729 4077 5732
rect 4111 5729 4123 5763
rect 6454 5760 6460 5772
rect 4065 5723 4123 5729
rect 4632 5732 6460 5760
rect 4632 5704 4660 5732
rect 6454 5720 6460 5732
rect 6512 5720 6518 5772
rect 6564 5704 6592 5800
rect 28810 5720 28816 5772
rect 28868 5760 28874 5772
rect 32493 5763 32551 5769
rect 32493 5760 32505 5763
rect 28868 5732 32505 5760
rect 28868 5720 28874 5732
rect 32493 5729 32505 5732
rect 32539 5729 32551 5763
rect 32493 5723 32551 5729
rect 3973 5695 4031 5701
rect 3973 5661 3985 5695
rect 4019 5692 4031 5695
rect 4338 5692 4344 5704
rect 4019 5664 4344 5692
rect 4019 5661 4031 5664
rect 3973 5655 4031 5661
rect 4338 5652 4344 5664
rect 4396 5652 4402 5704
rect 4614 5692 4620 5704
rect 4575 5664 4620 5692
rect 4614 5652 4620 5664
rect 4672 5652 4678 5704
rect 5074 5652 5080 5704
rect 5132 5692 5138 5704
rect 5261 5695 5319 5701
rect 5261 5692 5273 5695
rect 5132 5664 5273 5692
rect 5132 5652 5138 5664
rect 5261 5661 5273 5664
rect 5307 5692 5319 5695
rect 5626 5692 5632 5704
rect 5307 5664 5632 5692
rect 5307 5661 5319 5664
rect 5261 5655 5319 5661
rect 5626 5652 5632 5664
rect 5684 5652 5690 5704
rect 6086 5692 6092 5704
rect 6047 5664 6092 5692
rect 6086 5652 6092 5664
rect 6144 5652 6150 5704
rect 6546 5692 6552 5704
rect 6459 5664 6552 5692
rect 6546 5652 6552 5664
rect 6604 5652 6610 5704
rect 7374 5692 7380 5704
rect 7335 5664 7380 5692
rect 7374 5652 7380 5664
rect 7432 5652 7438 5704
rect 30745 5695 30803 5701
rect 30745 5661 30757 5695
rect 30791 5692 30803 5695
rect 31294 5692 31300 5704
rect 30791 5664 31300 5692
rect 30791 5661 30803 5664
rect 30745 5655 30803 5661
rect 31294 5652 31300 5664
rect 31352 5652 31358 5704
rect 31389 5695 31447 5701
rect 31389 5661 31401 5695
rect 31435 5692 31447 5695
rect 31846 5692 31852 5704
rect 31435 5664 31852 5692
rect 31435 5661 31447 5664
rect 31389 5655 31447 5661
rect 31846 5652 31852 5664
rect 31904 5652 31910 5704
rect 32030 5692 32036 5704
rect 31991 5664 32036 5692
rect 32030 5652 32036 5664
rect 32088 5652 32094 5704
rect 3418 5624 3424 5636
rect 3379 5596 3424 5624
rect 3418 5584 3424 5596
rect 3476 5584 3482 5636
rect 4154 5584 4160 5636
rect 4212 5624 4218 5636
rect 5353 5627 5411 5633
rect 5353 5624 5365 5627
rect 4212 5596 5365 5624
rect 4212 5584 4218 5596
rect 5353 5593 5365 5596
rect 5399 5593 5411 5627
rect 5353 5587 5411 5593
rect 32122 5584 32128 5636
rect 32180 5624 32186 5636
rect 32677 5627 32735 5633
rect 32677 5624 32689 5627
rect 32180 5596 32689 5624
rect 32180 5584 32186 5596
rect 32677 5593 32689 5596
rect 32723 5593 32735 5627
rect 32677 5587 32735 5593
rect 34333 5627 34391 5633
rect 34333 5593 34345 5627
rect 34379 5624 34391 5627
rect 34606 5624 34612 5636
rect 34379 5596 34612 5624
rect 34379 5593 34391 5596
rect 34333 5587 34391 5593
rect 34606 5584 34612 5596
rect 34664 5584 34670 5636
rect 4706 5556 4712 5568
rect 4667 5528 4712 5556
rect 4706 5516 4712 5528
rect 4764 5516 4770 5568
rect 6641 5559 6699 5565
rect 6641 5525 6653 5559
rect 6687 5556 6699 5559
rect 6730 5556 6736 5568
rect 6687 5528 6736 5556
rect 6687 5525 6699 5528
rect 6641 5519 6699 5525
rect 6730 5516 6736 5528
rect 6788 5516 6794 5568
rect 1104 5466 35027 5488
rect 1104 5414 9390 5466
rect 9442 5414 9454 5466
rect 9506 5414 9518 5466
rect 9570 5414 9582 5466
rect 9634 5414 9646 5466
rect 9698 5414 17831 5466
rect 17883 5414 17895 5466
rect 17947 5414 17959 5466
rect 18011 5414 18023 5466
rect 18075 5414 18087 5466
rect 18139 5414 26272 5466
rect 26324 5414 26336 5466
rect 26388 5414 26400 5466
rect 26452 5414 26464 5466
rect 26516 5414 26528 5466
rect 26580 5414 34713 5466
rect 34765 5414 34777 5466
rect 34829 5414 34841 5466
rect 34893 5414 34905 5466
rect 34957 5414 34969 5466
rect 35021 5414 35027 5466
rect 1104 5392 35027 5414
rect 4706 5352 4712 5364
rect 1964 5324 4712 5352
rect 1964 5293 1992 5324
rect 4706 5312 4712 5324
rect 4764 5312 4770 5364
rect 1949 5287 2007 5293
rect 1949 5253 1961 5287
rect 1995 5253 2007 5287
rect 1949 5247 2007 5253
rect 4249 5287 4307 5293
rect 4249 5253 4261 5287
rect 4295 5284 4307 5287
rect 7285 5287 7343 5293
rect 7285 5284 7297 5287
rect 4295 5256 7297 5284
rect 4295 5253 4307 5256
rect 4249 5247 4307 5253
rect 7285 5253 7297 5256
rect 7331 5253 7343 5287
rect 7285 5247 7343 5253
rect 32677 5287 32735 5293
rect 32677 5253 32689 5287
rect 32723 5284 32735 5287
rect 34054 5284 34060 5296
rect 32723 5256 34060 5284
rect 32723 5253 32735 5256
rect 32677 5247 32735 5253
rect 34054 5244 34060 5256
rect 34112 5244 34118 5296
rect 6454 5176 6460 5228
rect 6512 5216 6518 5228
rect 6549 5219 6607 5225
rect 6549 5216 6561 5219
rect 6512 5188 6561 5216
rect 6512 5176 6518 5188
rect 6549 5185 6561 5188
rect 6595 5216 6607 5219
rect 7190 5216 7196 5228
rect 6595 5188 6914 5216
rect 7151 5188 7196 5216
rect 6595 5185 6607 5188
rect 6549 5179 6607 5185
rect 1762 5148 1768 5160
rect 1723 5120 1768 5148
rect 1762 5108 1768 5120
rect 1820 5108 1826 5160
rect 2774 5148 2780 5160
rect 2735 5120 2780 5148
rect 2774 5108 2780 5120
rect 2832 5108 2838 5160
rect 4065 5151 4123 5157
rect 4065 5117 4077 5151
rect 4111 5148 4123 5151
rect 4890 5148 4896 5160
rect 4111 5120 4896 5148
rect 4111 5117 4123 5120
rect 4065 5111 4123 5117
rect 4890 5108 4896 5120
rect 4948 5108 4954 5160
rect 4985 5151 5043 5157
rect 4985 5117 4997 5151
rect 5031 5117 5043 5151
rect 6886 5148 6914 5188
rect 7190 5176 7196 5188
rect 7248 5176 7254 5228
rect 28074 5176 28080 5228
rect 28132 5216 28138 5228
rect 29917 5219 29975 5225
rect 29917 5216 29929 5219
rect 28132 5188 29929 5216
rect 28132 5176 28138 5188
rect 29917 5185 29929 5188
rect 29963 5185 29975 5219
rect 29917 5179 29975 5185
rect 32030 5176 32036 5228
rect 32088 5216 32094 5228
rect 32493 5219 32551 5225
rect 32493 5216 32505 5219
rect 32088 5188 32505 5216
rect 32088 5176 32094 5188
rect 32493 5185 32505 5188
rect 32539 5185 32551 5219
rect 32493 5179 32551 5185
rect 13170 5148 13176 5160
rect 6886 5120 13176 5148
rect 4985 5111 5043 5117
rect 4430 5040 4436 5092
rect 4488 5080 4494 5092
rect 5000 5080 5028 5111
rect 13170 5108 13176 5120
rect 13228 5108 13234 5160
rect 33042 5148 33048 5160
rect 33003 5120 33048 5148
rect 33042 5108 33048 5120
rect 33100 5108 33106 5160
rect 4488 5052 5028 5080
rect 4488 5040 4494 5052
rect 1854 4972 1860 5024
rect 1912 5012 1918 5024
rect 6641 5015 6699 5021
rect 6641 5012 6653 5015
rect 1912 4984 6653 5012
rect 1912 4972 1918 4984
rect 6641 4981 6653 4984
rect 6687 4981 6699 5015
rect 6641 4975 6699 4981
rect 30009 5015 30067 5021
rect 30009 4981 30021 5015
rect 30055 5012 30067 5015
rect 31018 5012 31024 5024
rect 30055 4984 31024 5012
rect 30055 4981 30067 4984
rect 30009 4975 30067 4981
rect 31018 4972 31024 4984
rect 31076 4972 31082 5024
rect 31202 5012 31208 5024
rect 31163 4984 31208 5012
rect 31202 4972 31208 4984
rect 31260 4972 31266 5024
rect 1104 4922 34868 4944
rect 1104 4870 5170 4922
rect 5222 4870 5234 4922
rect 5286 4870 5298 4922
rect 5350 4870 5362 4922
rect 5414 4870 5426 4922
rect 5478 4870 13611 4922
rect 13663 4870 13675 4922
rect 13727 4870 13739 4922
rect 13791 4870 13803 4922
rect 13855 4870 13867 4922
rect 13919 4870 22052 4922
rect 22104 4870 22116 4922
rect 22168 4870 22180 4922
rect 22232 4870 22244 4922
rect 22296 4870 22308 4922
rect 22360 4870 30493 4922
rect 30545 4870 30557 4922
rect 30609 4870 30621 4922
rect 30673 4870 30685 4922
rect 30737 4870 30749 4922
rect 30801 4870 34868 4922
rect 1104 4848 34868 4870
rect 6086 4740 6092 4752
rect 1596 4712 6092 4740
rect 1596 4681 1624 4712
rect 6086 4700 6092 4712
rect 6144 4700 6150 4752
rect 1581 4675 1639 4681
rect 1581 4641 1593 4675
rect 1627 4641 1639 4675
rect 1581 4635 1639 4641
rect 1765 4675 1823 4681
rect 1765 4641 1777 4675
rect 1811 4672 1823 4675
rect 1854 4672 1860 4684
rect 1811 4644 1860 4672
rect 1811 4641 1823 4644
rect 1765 4635 1823 4641
rect 1854 4632 1860 4644
rect 1912 4632 1918 4684
rect 2774 4672 2780 4684
rect 2735 4644 2780 4672
rect 2774 4632 2780 4644
rect 2832 4632 2838 4684
rect 4157 4675 4215 4681
rect 4157 4641 4169 4675
rect 4203 4672 4215 4675
rect 4798 4672 4804 4684
rect 4203 4644 4804 4672
rect 4203 4641 4215 4644
rect 4157 4635 4215 4641
rect 4798 4632 4804 4644
rect 4856 4632 4862 4684
rect 4890 4632 4896 4684
rect 4948 4672 4954 4684
rect 4948 4644 4993 4672
rect 4948 4632 4954 4644
rect 5074 4632 5080 4684
rect 5132 4672 5138 4684
rect 8018 4672 8024 4684
rect 5132 4644 8024 4672
rect 5132 4632 5138 4644
rect 3973 4607 4031 4613
rect 3973 4573 3985 4607
rect 4019 4573 4031 4607
rect 6454 4604 6460 4616
rect 6415 4576 6460 4604
rect 3973 4567 4031 4573
rect 3988 4536 4016 4567
rect 6454 4564 6460 4576
rect 6512 4564 6518 4616
rect 6932 4613 6960 4644
rect 8018 4632 8024 4644
rect 8076 4632 8082 4684
rect 31846 4632 31852 4684
rect 31904 4672 31910 4684
rect 32493 4675 32551 4681
rect 32493 4672 32505 4675
rect 31904 4644 32505 4672
rect 31904 4632 31910 4644
rect 32493 4641 32505 4644
rect 32539 4641 32551 4675
rect 32674 4672 32680 4684
rect 32635 4644 32680 4672
rect 32493 4635 32551 4641
rect 32674 4632 32680 4644
rect 32732 4632 32738 4684
rect 6917 4607 6975 4613
rect 6917 4573 6929 4607
rect 6963 4604 6975 4607
rect 6963 4576 6997 4604
rect 6963 4573 6975 4576
rect 6917 4567 6975 4573
rect 7190 4564 7196 4616
rect 7248 4604 7254 4616
rect 7561 4607 7619 4613
rect 7561 4604 7573 4607
rect 7248 4576 7573 4604
rect 7248 4564 7254 4576
rect 7561 4573 7573 4576
rect 7607 4573 7619 4607
rect 8386 4604 8392 4616
rect 8347 4576 8392 4604
rect 7561 4567 7619 4573
rect 8386 4564 8392 4576
rect 8444 4564 8450 4616
rect 19978 4604 19984 4616
rect 19891 4576 19984 4604
rect 19978 4564 19984 4576
rect 20036 4604 20042 4616
rect 28074 4604 28080 4616
rect 20036 4576 28080 4604
rect 20036 4564 20042 4576
rect 28074 4564 28080 4576
rect 28132 4564 28138 4616
rect 29181 4607 29239 4613
rect 29181 4573 29193 4607
rect 29227 4604 29239 4607
rect 30193 4607 30251 4613
rect 30193 4604 30205 4607
rect 29227 4576 30205 4604
rect 29227 4573 29239 4576
rect 29181 4567 29239 4573
rect 30193 4573 30205 4576
rect 30239 4573 30251 4607
rect 30193 4567 30251 4573
rect 5534 4536 5540 4548
rect 3988 4508 5540 4536
rect 5534 4496 5540 4508
rect 5592 4496 5598 4548
rect 5810 4496 5816 4548
rect 5868 4536 5874 4548
rect 7653 4539 7711 4545
rect 7653 4536 7665 4539
rect 5868 4508 7665 4536
rect 5868 4496 5874 4508
rect 7653 4505 7665 4508
rect 7699 4505 7711 4539
rect 7653 4499 7711 4505
rect 30377 4539 30435 4545
rect 30377 4505 30389 4539
rect 30423 4536 30435 4539
rect 30834 4536 30840 4548
rect 30423 4508 30840 4536
rect 30423 4505 30435 4508
rect 30377 4499 30435 4505
rect 30834 4496 30840 4508
rect 30892 4496 30898 4548
rect 32033 4539 32091 4545
rect 32033 4505 32045 4539
rect 32079 4505 32091 4539
rect 34330 4536 34336 4548
rect 34291 4508 34336 4536
rect 32033 4499 32091 4505
rect 6914 4428 6920 4480
rect 6972 4468 6978 4480
rect 7009 4471 7067 4477
rect 7009 4468 7021 4471
rect 6972 4440 7021 4468
rect 6972 4428 6978 4440
rect 7009 4437 7021 4440
rect 7055 4437 7067 4471
rect 7009 4431 7067 4437
rect 19794 4428 19800 4480
rect 19852 4468 19858 4480
rect 20073 4471 20131 4477
rect 20073 4468 20085 4471
rect 19852 4440 20085 4468
rect 19852 4428 19858 4440
rect 20073 4437 20085 4440
rect 20119 4437 20131 4471
rect 32048 4468 32076 4499
rect 34330 4496 34336 4508
rect 34388 4496 34394 4548
rect 34514 4468 34520 4480
rect 32048 4440 34520 4468
rect 20073 4431 20131 4437
rect 34514 4428 34520 4440
rect 34572 4428 34578 4480
rect 1104 4378 35027 4400
rect 1104 4326 9390 4378
rect 9442 4326 9454 4378
rect 9506 4326 9518 4378
rect 9570 4326 9582 4378
rect 9634 4326 9646 4378
rect 9698 4326 17831 4378
rect 17883 4326 17895 4378
rect 17947 4326 17959 4378
rect 18011 4326 18023 4378
rect 18075 4326 18087 4378
rect 18139 4326 26272 4378
rect 26324 4326 26336 4378
rect 26388 4326 26400 4378
rect 26452 4326 26464 4378
rect 26516 4326 26528 4378
rect 26580 4326 34713 4378
rect 34765 4326 34777 4378
rect 34829 4326 34841 4378
rect 34893 4326 34905 4378
rect 34957 4326 34969 4378
rect 35021 4326 35027 4378
rect 1104 4304 35027 4326
rect 19794 4196 19800 4208
rect 6472 4168 6776 4196
rect 19755 4168 19800 4196
rect 1762 4088 1768 4140
rect 1820 4128 1826 4140
rect 2041 4131 2099 4137
rect 2041 4128 2053 4131
rect 1820 4100 2053 4128
rect 1820 4088 1826 4100
rect 2041 4097 2053 4100
rect 2087 4097 2099 4131
rect 2041 4091 2099 4097
rect 3970 4088 3976 4140
rect 4028 4128 4034 4140
rect 4028 4100 4292 4128
rect 4028 4088 4034 4100
rect 2593 4063 2651 4069
rect 2593 4029 2605 4063
rect 2639 4029 2651 4063
rect 2593 4023 2651 4029
rect 2777 4063 2835 4069
rect 2777 4029 2789 4063
rect 2823 4060 2835 4063
rect 4154 4060 4160 4072
rect 2823 4032 4160 4060
rect 2823 4029 2835 4032
rect 2777 4023 2835 4029
rect 2608 3992 2636 4023
rect 4154 4020 4160 4032
rect 4212 4020 4218 4072
rect 4264 4069 4292 4100
rect 4338 4088 4344 4140
rect 4396 4128 4402 4140
rect 4985 4131 5043 4137
rect 4985 4128 4997 4131
rect 4396 4100 4997 4128
rect 4396 4088 4402 4100
rect 4985 4097 4997 4100
rect 5031 4097 5043 4131
rect 5626 4128 5632 4140
rect 5587 4100 5632 4128
rect 4985 4091 5043 4097
rect 5626 4088 5632 4100
rect 5684 4128 5690 4140
rect 6472 4128 6500 4168
rect 5684 4100 6500 4128
rect 5684 4088 5690 4100
rect 6546 4088 6552 4140
rect 6604 4128 6610 4140
rect 6748 4128 6776 4168
rect 19794 4156 19800 4168
rect 19852 4156 19858 4208
rect 6604 4100 6649 4128
rect 6748 4100 7972 4128
rect 6604 4088 6610 4100
rect 4249 4063 4307 4069
rect 4249 4029 4261 4063
rect 4295 4029 4307 4063
rect 4249 4023 4307 4029
rect 5534 4020 5540 4072
rect 5592 4060 5598 4072
rect 7377 4063 7435 4069
rect 7377 4060 7389 4063
rect 5592 4032 7389 4060
rect 5592 4020 5598 4032
rect 7377 4029 7389 4032
rect 7423 4029 7435 4063
rect 7944 4060 7972 4100
rect 8018 4088 8024 4140
rect 8076 4128 8082 4140
rect 9122 4128 9128 4140
rect 8076 4100 8121 4128
rect 9083 4100 9128 4128
rect 8076 4088 8082 4100
rect 9122 4088 9128 4100
rect 9180 4088 9186 4140
rect 28810 4128 28816 4140
rect 28771 4100 28816 4128
rect 28810 4088 28816 4100
rect 28868 4088 28874 4140
rect 31294 4088 31300 4140
rect 31352 4128 31358 4140
rect 32493 4131 32551 4137
rect 32493 4128 32505 4131
rect 31352 4100 32505 4128
rect 31352 4088 31358 4100
rect 32493 4097 32505 4100
rect 32539 4097 32551 4131
rect 32493 4091 32551 4097
rect 9140 4060 9168 4088
rect 13078 4060 13084 4072
rect 7944 4032 9168 4060
rect 13039 4032 13084 4060
rect 7377 4023 7435 4029
rect 13078 4020 13084 4032
rect 13136 4020 13142 4072
rect 13262 4060 13268 4072
rect 13223 4032 13268 4060
rect 13262 4020 13268 4032
rect 13320 4020 13326 4072
rect 13446 4020 13452 4072
rect 13504 4060 13510 4072
rect 13541 4063 13599 4069
rect 13541 4060 13553 4063
rect 13504 4032 13553 4060
rect 13504 4020 13510 4032
rect 13541 4029 13553 4032
rect 13587 4029 13599 4063
rect 13541 4023 13599 4029
rect 19613 4063 19671 4069
rect 19613 4029 19625 4063
rect 19659 4060 19671 4063
rect 20254 4060 20260 4072
rect 19659 4032 20260 4060
rect 19659 4029 19671 4032
rect 19613 4023 19671 4029
rect 20254 4020 20260 4032
rect 20312 4020 20318 4072
rect 20622 4060 20628 4072
rect 20583 4032 20628 4060
rect 20622 4020 20628 4032
rect 20680 4020 20686 4072
rect 27890 4020 27896 4072
rect 27948 4060 27954 4072
rect 29917 4063 29975 4069
rect 29917 4060 29929 4063
rect 27948 4032 29929 4060
rect 27948 4020 27954 4032
rect 29917 4029 29929 4032
rect 29963 4029 29975 4063
rect 30098 4060 30104 4072
rect 30059 4032 30104 4060
rect 29917 4023 29975 4029
rect 30098 4020 30104 4032
rect 30156 4020 30162 4072
rect 31757 4063 31815 4069
rect 31757 4029 31769 4063
rect 31803 4060 31815 4063
rect 31846 4060 31852 4072
rect 31803 4032 31852 4060
rect 31803 4029 31815 4032
rect 31757 4023 31815 4029
rect 31846 4020 31852 4032
rect 31904 4020 31910 4072
rect 32674 4060 32680 4072
rect 32635 4032 32680 4060
rect 32674 4020 32680 4032
rect 32732 4020 32738 4072
rect 34333 4063 34391 4069
rect 34333 4029 34345 4063
rect 34379 4060 34391 4063
rect 35434 4060 35440 4072
rect 34379 4032 35440 4060
rect 34379 4029 34391 4032
rect 34333 4023 34391 4029
rect 35434 4020 35440 4032
rect 35492 4020 35498 4072
rect 6454 3992 6460 4004
rect 2608 3964 6460 3992
rect 6454 3952 6460 3964
rect 6512 3952 6518 4004
rect 6546 3952 6552 4004
rect 6604 3992 6610 4004
rect 15654 3992 15660 4004
rect 6604 3964 15660 3992
rect 6604 3952 6610 3964
rect 15654 3952 15660 3964
rect 15712 3952 15718 4004
rect 27706 3952 27712 4004
rect 27764 3992 27770 4004
rect 33134 3992 33140 4004
rect 27764 3964 33140 3992
rect 27764 3952 27770 3964
rect 33134 3952 33140 3964
rect 33192 3952 33198 4004
rect 4338 3884 4344 3936
rect 4396 3924 4402 3936
rect 5077 3927 5135 3933
rect 5077 3924 5089 3927
rect 4396 3896 5089 3924
rect 4396 3884 4402 3896
rect 5077 3893 5089 3896
rect 5123 3893 5135 3927
rect 5718 3924 5724 3936
rect 5679 3896 5724 3924
rect 5077 3887 5135 3893
rect 5718 3884 5724 3896
rect 5776 3884 5782 3936
rect 6086 3884 6092 3936
rect 6144 3924 6150 3936
rect 6641 3927 6699 3933
rect 6641 3924 6653 3927
rect 6144 3896 6653 3924
rect 6144 3884 6150 3896
rect 6641 3893 6653 3896
rect 6687 3893 6699 3927
rect 6641 3887 6699 3893
rect 7190 3884 7196 3936
rect 7248 3924 7254 3936
rect 8113 3927 8171 3933
rect 8113 3924 8125 3927
rect 7248 3896 8125 3924
rect 7248 3884 7254 3896
rect 8113 3893 8125 3896
rect 8159 3893 8171 3927
rect 9214 3924 9220 3936
rect 9175 3896 9220 3924
rect 8113 3887 8171 3893
rect 9214 3884 9220 3896
rect 9272 3884 9278 3936
rect 15562 3884 15568 3936
rect 15620 3924 15626 3936
rect 15749 3927 15807 3933
rect 15749 3924 15761 3927
rect 15620 3896 15761 3924
rect 15620 3884 15626 3896
rect 15749 3893 15761 3896
rect 15795 3893 15807 3927
rect 15749 3887 15807 3893
rect 16850 3884 16856 3936
rect 16908 3924 16914 3936
rect 17037 3927 17095 3933
rect 17037 3924 17049 3927
rect 16908 3896 17049 3924
rect 16908 3884 16914 3896
rect 17037 3893 17049 3896
rect 17083 3893 17095 3927
rect 17037 3887 17095 3893
rect 20070 3884 20076 3936
rect 20128 3924 20134 3936
rect 27614 3924 27620 3936
rect 20128 3896 27620 3924
rect 20128 3884 20134 3896
rect 27614 3884 27620 3896
rect 27672 3884 27678 3936
rect 29457 3927 29515 3933
rect 29457 3893 29469 3927
rect 29503 3924 29515 3927
rect 31662 3924 31668 3936
rect 29503 3896 31668 3924
rect 29503 3893 29515 3896
rect 29457 3887 29515 3893
rect 31662 3884 31668 3896
rect 31720 3884 31726 3936
rect 1104 3834 34868 3856
rect 1104 3782 5170 3834
rect 5222 3782 5234 3834
rect 5286 3782 5298 3834
rect 5350 3782 5362 3834
rect 5414 3782 5426 3834
rect 5478 3782 13611 3834
rect 13663 3782 13675 3834
rect 13727 3782 13739 3834
rect 13791 3782 13803 3834
rect 13855 3782 13867 3834
rect 13919 3782 22052 3834
rect 22104 3782 22116 3834
rect 22168 3782 22180 3834
rect 22232 3782 22244 3834
rect 22296 3782 22308 3834
rect 22360 3782 30493 3834
rect 30545 3782 30557 3834
rect 30609 3782 30621 3834
rect 30673 3782 30685 3834
rect 30737 3782 30749 3834
rect 30801 3782 34868 3834
rect 1104 3760 34868 3782
rect 13078 3720 13084 3732
rect 13039 3692 13084 3720
rect 13078 3680 13084 3692
rect 13136 3680 13142 3732
rect 20070 3720 20076 3732
rect 13188 3692 20076 3720
rect 8386 3652 8392 3664
rect 1596 3624 8392 3652
rect 1596 3593 1624 3624
rect 8386 3612 8392 3624
rect 8444 3612 8450 3664
rect 10502 3612 10508 3664
rect 10560 3652 10566 3664
rect 13188 3652 13216 3692
rect 20070 3680 20076 3692
rect 20128 3680 20134 3732
rect 20254 3720 20260 3732
rect 20215 3692 20260 3720
rect 20254 3680 20260 3692
rect 20312 3680 20318 3732
rect 23750 3680 23756 3732
rect 23808 3720 23814 3732
rect 27706 3720 27712 3732
rect 23808 3692 27712 3720
rect 23808 3680 23814 3692
rect 27706 3680 27712 3692
rect 27764 3680 27770 3732
rect 27890 3720 27896 3732
rect 27851 3692 27896 3720
rect 27890 3680 27896 3692
rect 27948 3680 27954 3732
rect 28445 3723 28503 3729
rect 28445 3689 28457 3723
rect 28491 3720 28503 3723
rect 30098 3720 30104 3732
rect 28491 3692 30104 3720
rect 28491 3689 28503 3692
rect 28445 3683 28503 3689
rect 30098 3680 30104 3692
rect 30156 3680 30162 3732
rect 31938 3720 31944 3732
rect 30208 3692 31944 3720
rect 10560 3624 13216 3652
rect 10560 3612 10566 3624
rect 14366 3612 14372 3664
rect 14424 3652 14430 3664
rect 14424 3624 26234 3652
rect 14424 3612 14430 3624
rect 1581 3587 1639 3593
rect 1581 3553 1593 3587
rect 1627 3553 1639 3587
rect 2774 3584 2780 3596
rect 2735 3556 2780 3584
rect 1581 3547 1639 3553
rect 2774 3544 2780 3556
rect 2832 3544 2838 3596
rect 6086 3584 6092 3596
rect 6047 3556 6092 3584
rect 6086 3544 6092 3556
rect 6144 3544 6150 3596
rect 6454 3584 6460 3596
rect 6415 3556 6460 3584
rect 6454 3544 6460 3556
rect 6512 3544 6518 3596
rect 15562 3584 15568 3596
rect 15523 3556 15568 3584
rect 15562 3544 15568 3556
rect 15620 3544 15626 3596
rect 16114 3584 16120 3596
rect 16075 3556 16120 3584
rect 16114 3544 16120 3556
rect 16172 3544 16178 3596
rect 21266 3584 21272 3596
rect 21227 3556 21272 3584
rect 21266 3544 21272 3556
rect 21324 3544 21330 3596
rect 4154 3516 4160 3528
rect 4115 3488 4160 3516
rect 4154 3476 4160 3488
rect 4212 3476 4218 3528
rect 4798 3516 4804 3528
rect 4759 3488 4804 3516
rect 4798 3476 4804 3488
rect 4856 3476 4862 3528
rect 5445 3519 5503 3525
rect 5445 3485 5457 3519
rect 5491 3516 5503 3519
rect 5905 3519 5963 3525
rect 5905 3516 5917 3519
rect 5491 3488 5917 3516
rect 5491 3485 5503 3488
rect 5445 3479 5503 3485
rect 5905 3485 5917 3488
rect 5951 3485 5963 3519
rect 5905 3479 5963 3485
rect 8389 3519 8447 3525
rect 8389 3485 8401 3519
rect 8435 3485 8447 3519
rect 9306 3516 9312 3528
rect 9267 3488 9312 3516
rect 8389 3479 8447 3485
rect 1765 3451 1823 3457
rect 1765 3417 1777 3451
rect 1811 3448 1823 3451
rect 2958 3448 2964 3460
rect 1811 3420 2964 3448
rect 1811 3417 1823 3420
rect 1765 3411 1823 3417
rect 2958 3408 2964 3420
rect 3016 3408 3022 3460
rect 7006 3408 7012 3460
rect 7064 3448 7070 3460
rect 8404 3448 8432 3479
rect 9306 3476 9312 3488
rect 9364 3476 9370 3528
rect 10042 3516 10048 3528
rect 10003 3488 10048 3516
rect 10042 3476 10048 3488
rect 10100 3476 10106 3528
rect 10502 3516 10508 3528
rect 10463 3488 10508 3516
rect 10502 3476 10508 3488
rect 10560 3476 10566 3528
rect 13725 3519 13783 3525
rect 13725 3485 13737 3519
rect 13771 3516 13783 3519
rect 14274 3516 14280 3528
rect 13771 3488 14280 3516
rect 13771 3485 13783 3488
rect 13725 3479 13783 3485
rect 14274 3476 14280 3488
rect 14332 3476 14338 3528
rect 14366 3476 14372 3528
rect 14424 3516 14430 3528
rect 14424 3488 14469 3516
rect 14424 3476 14430 3488
rect 19426 3476 19432 3528
rect 19484 3516 19490 3528
rect 19613 3519 19671 3525
rect 19613 3516 19625 3519
rect 19484 3488 19625 3516
rect 19484 3476 19490 3488
rect 19613 3485 19625 3488
rect 19659 3485 19671 3519
rect 20714 3516 20720 3528
rect 20675 3488 20720 3516
rect 19613 3479 19671 3485
rect 20714 3476 20720 3488
rect 20772 3476 20778 3528
rect 23750 3476 23756 3528
rect 23808 3516 23814 3528
rect 23845 3519 23903 3525
rect 23845 3516 23857 3519
rect 23808 3488 23857 3516
rect 23808 3476 23814 3488
rect 23845 3485 23857 3488
rect 23891 3485 23903 3519
rect 24762 3516 24768 3528
rect 24723 3488 24768 3516
rect 23845 3479 23903 3485
rect 24762 3476 24768 3488
rect 24820 3476 24826 3528
rect 26206 3516 26234 3624
rect 30208 3584 30236 3692
rect 31938 3680 31944 3692
rect 31996 3680 32002 3732
rect 34054 3720 34060 3732
rect 34015 3692 34060 3720
rect 34054 3680 34060 3692
rect 34112 3680 34118 3732
rect 31754 3652 31760 3664
rect 29012 3556 30236 3584
rect 30300 3624 31760 3652
rect 28353 3519 28411 3525
rect 28353 3516 28365 3519
rect 26206 3488 28365 3516
rect 28353 3485 28365 3488
rect 28399 3485 28411 3519
rect 28353 3479 28411 3485
rect 7064 3420 8432 3448
rect 7064 3408 7070 3420
rect 9122 3408 9128 3460
rect 9180 3448 9186 3460
rect 15746 3448 15752 3460
rect 9180 3420 14596 3448
rect 15707 3420 15752 3448
rect 9180 3408 9186 3420
rect 9766 3340 9772 3392
rect 9824 3380 9830 3392
rect 10597 3383 10655 3389
rect 10597 3380 10609 3383
rect 9824 3352 10609 3380
rect 9824 3340 9830 3352
rect 10597 3349 10609 3352
rect 10643 3349 10655 3383
rect 14458 3380 14464 3392
rect 14419 3352 14464 3380
rect 10597 3343 10655 3349
rect 14458 3340 14464 3352
rect 14516 3340 14522 3392
rect 14568 3380 14596 3420
rect 15746 3408 15752 3420
rect 15804 3408 15810 3460
rect 20901 3451 20959 3457
rect 20901 3417 20913 3451
rect 20947 3448 20959 3451
rect 22094 3448 22100 3460
rect 20947 3420 22100 3448
rect 20947 3417 20959 3420
rect 20901 3411 20959 3417
rect 22094 3408 22100 3420
rect 22152 3408 22158 3460
rect 27706 3448 27712 3460
rect 22664 3420 27712 3448
rect 22664 3380 22692 3420
rect 27706 3408 27712 3420
rect 27764 3408 27770 3460
rect 28368 3448 28396 3479
rect 28442 3476 28448 3528
rect 28500 3516 28506 3528
rect 29012 3525 29040 3556
rect 28997 3519 29055 3525
rect 28997 3516 29009 3519
rect 28500 3488 29009 3516
rect 28500 3476 28506 3488
rect 28997 3485 29009 3488
rect 29043 3485 29055 3519
rect 28997 3479 29055 3485
rect 29638 3476 29644 3528
rect 29696 3516 29702 3528
rect 29917 3519 29975 3525
rect 29917 3516 29929 3519
rect 29696 3488 29929 3516
rect 29696 3476 29702 3488
rect 29917 3485 29929 3488
rect 29963 3485 29975 3519
rect 29917 3479 29975 3485
rect 30300 3448 30328 3624
rect 31754 3612 31760 3624
rect 31812 3612 31818 3664
rect 33134 3612 33140 3664
rect 33192 3652 33198 3664
rect 33192 3624 34008 3652
rect 33192 3612 33198 3624
rect 31021 3587 31079 3593
rect 31021 3553 31033 3587
rect 31067 3584 31079 3587
rect 31202 3584 31208 3596
rect 31067 3556 31208 3584
rect 31067 3553 31079 3556
rect 31021 3547 31079 3553
rect 31202 3544 31208 3556
rect 31260 3544 31266 3596
rect 31294 3544 31300 3596
rect 31352 3584 31358 3596
rect 33778 3584 33784 3596
rect 31352 3556 33784 3584
rect 31352 3544 31358 3556
rect 33778 3544 33784 3556
rect 33836 3544 33842 3596
rect 30374 3476 30380 3528
rect 30432 3516 30438 3528
rect 30561 3519 30619 3525
rect 30561 3516 30573 3519
rect 30432 3488 30573 3516
rect 30432 3476 30438 3488
rect 30561 3485 30573 3488
rect 30607 3485 30619 3519
rect 33502 3516 33508 3528
rect 33463 3488 33508 3516
rect 30561 3479 30619 3485
rect 33502 3476 33508 3488
rect 33560 3476 33566 3528
rect 33980 3525 34008 3624
rect 33965 3519 34023 3525
rect 33965 3485 33977 3519
rect 34011 3485 34023 3519
rect 33965 3479 34023 3485
rect 28368 3420 30328 3448
rect 31018 3408 31024 3460
rect 31076 3448 31082 3460
rect 31205 3451 31263 3457
rect 31205 3448 31217 3451
rect 31076 3420 31217 3448
rect 31076 3408 31082 3420
rect 31205 3417 31217 3420
rect 31251 3417 31263 3451
rect 31205 3411 31263 3417
rect 32861 3451 32919 3457
rect 32861 3417 32873 3451
rect 32907 3448 32919 3451
rect 35894 3448 35900 3460
rect 32907 3420 35900 3448
rect 32907 3417 32919 3420
rect 32861 3411 32919 3417
rect 35894 3408 35900 3420
rect 35952 3408 35958 3460
rect 14568 3352 22692 3380
rect 23937 3383 23995 3389
rect 23937 3349 23949 3383
rect 23983 3380 23995 3383
rect 24026 3380 24032 3392
rect 23983 3352 24032 3380
rect 23983 3349 23995 3352
rect 23937 3343 23995 3349
rect 24026 3340 24032 3352
rect 24084 3340 24090 3392
rect 29089 3383 29147 3389
rect 29089 3349 29101 3383
rect 29135 3380 29147 3383
rect 32490 3380 32496 3392
rect 29135 3352 32496 3380
rect 29135 3349 29147 3352
rect 29089 3343 29147 3349
rect 32490 3340 32496 3352
rect 32548 3340 32554 3392
rect 1104 3290 35027 3312
rect 1104 3238 9390 3290
rect 9442 3238 9454 3290
rect 9506 3238 9518 3290
rect 9570 3238 9582 3290
rect 9634 3238 9646 3290
rect 9698 3238 17831 3290
rect 17883 3238 17895 3290
rect 17947 3238 17959 3290
rect 18011 3238 18023 3290
rect 18075 3238 18087 3290
rect 18139 3238 26272 3290
rect 26324 3238 26336 3290
rect 26388 3238 26400 3290
rect 26452 3238 26464 3290
rect 26516 3238 26528 3290
rect 26580 3238 34713 3290
rect 34765 3238 34777 3290
rect 34829 3238 34841 3290
rect 34893 3238 34905 3290
rect 34957 3238 34969 3290
rect 35021 3238 35027 3290
rect 1104 3216 35027 3238
rect 6914 3176 6920 3188
rect 2056 3148 6920 3176
rect 2056 3117 2084 3148
rect 6914 3136 6920 3148
rect 6972 3136 6978 3188
rect 8018 3136 8024 3188
rect 8076 3176 8082 3188
rect 13262 3176 13268 3188
rect 8076 3148 9904 3176
rect 13223 3148 13268 3176
rect 8076 3136 8082 3148
rect 2041 3111 2099 3117
rect 2041 3077 2053 3111
rect 2087 3077 2099 3111
rect 4338 3108 4344 3120
rect 4299 3080 4344 3108
rect 2041 3071 2099 3077
rect 4338 3068 4344 3080
rect 4396 3068 4402 3120
rect 7190 3108 7196 3120
rect 7151 3080 7196 3108
rect 7190 3068 7196 3080
rect 7248 3068 7254 3120
rect 9493 3111 9551 3117
rect 9493 3077 9505 3111
rect 9539 3108 9551 3111
rect 9766 3108 9772 3120
rect 9539 3080 9772 3108
rect 9539 3077 9551 3080
rect 9493 3071 9551 3077
rect 9766 3068 9772 3080
rect 9824 3068 9830 3120
rect 9876 3108 9904 3148
rect 13262 3136 13268 3148
rect 13320 3136 13326 3188
rect 19334 3176 19340 3188
rect 13372 3148 19340 3176
rect 13372 3108 13400 3148
rect 19334 3136 19340 3148
rect 19392 3136 19398 3188
rect 22094 3176 22100 3188
rect 22055 3148 22100 3176
rect 22094 3136 22100 3148
rect 22152 3136 22158 3188
rect 24762 3176 24768 3188
rect 23860 3148 24768 3176
rect 14458 3108 14464 3120
rect 9876 3080 13400 3108
rect 14419 3080 14464 3108
rect 14458 3068 14464 3080
rect 14516 3068 14522 3120
rect 23750 3108 23756 3120
rect 16546 3080 23756 3108
rect 7006 3040 7012 3052
rect 6967 3012 7012 3040
rect 7006 3000 7012 3012
rect 7064 3000 7070 3052
rect 13170 3040 13176 3052
rect 13131 3012 13176 3040
rect 13170 3000 13176 3012
rect 13228 3000 13234 3052
rect 14274 3040 14280 3052
rect 14235 3012 14280 3040
rect 14274 3000 14280 3012
rect 14332 3000 14338 3052
rect 1857 2975 1915 2981
rect 1857 2941 1869 2975
rect 1903 2972 1915 2975
rect 3050 2972 3056 2984
rect 1903 2944 3056 2972
rect 1903 2941 1915 2944
rect 1857 2935 1915 2941
rect 3050 2932 3056 2944
rect 3108 2932 3114 2984
rect 3234 2972 3240 2984
rect 3195 2944 3240 2972
rect 3234 2932 3240 2944
rect 3292 2932 3298 2984
rect 4157 2975 4215 2981
rect 4157 2941 4169 2975
rect 4203 2972 4215 2975
rect 4798 2972 4804 2984
rect 4203 2944 4804 2972
rect 4203 2941 4215 2944
rect 4157 2935 4215 2941
rect 4798 2932 4804 2944
rect 4856 2932 4862 2984
rect 5074 2972 5080 2984
rect 5035 2944 5080 2972
rect 5074 2932 5080 2944
rect 5132 2932 5138 2984
rect 8386 2972 8392 2984
rect 8347 2944 8392 2972
rect 8386 2932 8392 2944
rect 8444 2932 8450 2984
rect 9309 2975 9367 2981
rect 9309 2941 9321 2975
rect 9355 2972 9367 2975
rect 10042 2972 10048 2984
rect 9355 2944 10048 2972
rect 9355 2941 9367 2944
rect 9309 2935 9367 2941
rect 10042 2932 10048 2944
rect 10100 2932 10106 2984
rect 10318 2972 10324 2984
rect 10279 2944 10324 2972
rect 10318 2932 10324 2944
rect 10376 2932 10382 2984
rect 3878 2864 3884 2916
rect 3936 2904 3942 2916
rect 4890 2904 4896 2916
rect 3936 2876 4896 2904
rect 3936 2864 3942 2876
rect 4890 2864 4896 2876
rect 4948 2864 4954 2916
rect 13188 2904 13216 3000
rect 14826 2972 14832 2984
rect 14787 2944 14832 2972
rect 14826 2932 14832 2944
rect 14884 2932 14890 2984
rect 16546 2904 16574 3080
rect 23750 3068 23756 3080
rect 23808 3068 23814 3120
rect 16850 3040 16856 3052
rect 16811 3012 16856 3040
rect 16850 3000 16856 3012
rect 16908 3000 16914 3052
rect 19426 3040 19432 3052
rect 19387 3012 19432 3040
rect 19426 3000 19432 3012
rect 19484 3000 19490 3052
rect 21910 3000 21916 3052
rect 21968 3040 21974 3052
rect 23860 3049 23888 3148
rect 24762 3136 24768 3148
rect 24820 3136 24826 3188
rect 27801 3179 27859 3185
rect 27801 3145 27813 3179
rect 27847 3176 27859 3179
rect 32674 3176 32680 3188
rect 27847 3148 32680 3176
rect 27847 3145 27859 3148
rect 27801 3139 27859 3145
rect 32674 3136 32680 3148
rect 32732 3136 32738 3188
rect 24026 3108 24032 3120
rect 23987 3080 24032 3108
rect 24026 3068 24032 3080
rect 24084 3068 24090 3120
rect 27614 3068 27620 3120
rect 27672 3108 27678 3120
rect 28534 3108 28540 3120
rect 27672 3080 28540 3108
rect 27672 3068 27678 3080
rect 27724 3049 27752 3080
rect 28534 3068 28540 3080
rect 28592 3068 28598 3120
rect 29089 3111 29147 3117
rect 29089 3077 29101 3111
rect 29135 3108 29147 3111
rect 29825 3111 29883 3117
rect 29825 3108 29837 3111
rect 29135 3080 29837 3108
rect 29135 3077 29147 3080
rect 29089 3071 29147 3077
rect 29825 3077 29837 3080
rect 29871 3077 29883 3111
rect 29825 3071 29883 3077
rect 29914 3068 29920 3120
rect 29972 3108 29978 3120
rect 31294 3108 31300 3120
rect 29972 3080 31300 3108
rect 29972 3068 29978 3080
rect 31294 3068 31300 3080
rect 31352 3068 31358 3120
rect 32490 3108 32496 3120
rect 32451 3080 32496 3108
rect 32490 3068 32496 3080
rect 32548 3068 32554 3120
rect 22005 3043 22063 3049
rect 22005 3040 22017 3043
rect 21968 3012 22017 3040
rect 21968 3000 21974 3012
rect 22005 3009 22017 3012
rect 22051 3009 22063 3043
rect 22005 3003 22063 3009
rect 23845 3043 23903 3049
rect 23845 3009 23857 3043
rect 23891 3009 23903 3043
rect 23845 3003 23903 3009
rect 27709 3043 27767 3049
rect 27709 3009 27721 3043
rect 27755 3009 27767 3043
rect 27709 3003 27767 3009
rect 28353 3043 28411 3049
rect 28353 3009 28365 3043
rect 28399 3040 28411 3043
rect 28442 3040 28448 3052
rect 28399 3012 28448 3040
rect 28399 3009 28411 3012
rect 28353 3003 28411 3009
rect 17034 2972 17040 2984
rect 16995 2944 17040 2972
rect 17034 2932 17040 2944
rect 17092 2932 17098 2984
rect 17402 2972 17408 2984
rect 17363 2944 17408 2972
rect 17402 2932 17408 2944
rect 17460 2932 17466 2984
rect 19610 2972 19616 2984
rect 19571 2944 19616 2972
rect 19610 2932 19616 2944
rect 19668 2932 19674 2984
rect 19978 2972 19984 2984
rect 19939 2944 19984 2972
rect 19978 2932 19984 2944
rect 20036 2932 20042 2984
rect 13188 2876 16574 2904
rect 22020 2904 22048 3003
rect 24486 2972 24492 2984
rect 24447 2944 24492 2972
rect 24486 2932 24492 2944
rect 24544 2932 24550 2984
rect 28368 2904 28396 3003
rect 28442 3000 28448 3012
rect 28500 3000 28506 3052
rect 28997 3043 29055 3049
rect 28997 3009 29009 3043
rect 29043 3009 29055 3043
rect 29638 3040 29644 3052
rect 29599 3012 29644 3040
rect 28997 3003 29055 3009
rect 29012 2972 29040 3003
rect 29638 3000 29644 3012
rect 29696 3000 29702 3052
rect 29086 2972 29092 2984
rect 28999 2944 29092 2972
rect 29086 2932 29092 2944
rect 29144 2972 29150 2984
rect 29914 2972 29920 2984
rect 29144 2944 29920 2972
rect 29144 2932 29150 2944
rect 29914 2932 29920 2944
rect 29972 2932 29978 2984
rect 30282 2972 30288 2984
rect 30243 2944 30288 2972
rect 30282 2932 30288 2944
rect 30340 2932 30346 2984
rect 32309 2975 32367 2981
rect 32309 2941 32321 2975
rect 32355 2972 32367 2975
rect 33502 2972 33508 2984
rect 32355 2944 33508 2972
rect 32355 2941 32367 2944
rect 32309 2935 32367 2941
rect 33502 2932 33508 2944
rect 33560 2932 33566 2984
rect 33689 2975 33747 2981
rect 33689 2941 33701 2975
rect 33735 2941 33747 2975
rect 33689 2935 33747 2941
rect 22020 2876 28396 2904
rect 28534 2864 28540 2916
rect 28592 2904 28598 2916
rect 28592 2876 30328 2904
rect 28592 2864 28598 2876
rect 658 2796 664 2848
rect 716 2836 722 2848
rect 6822 2836 6828 2848
rect 716 2808 6828 2836
rect 716 2796 722 2808
rect 6822 2796 6828 2808
rect 6880 2796 6886 2848
rect 28445 2839 28503 2845
rect 28445 2805 28457 2839
rect 28491 2836 28503 2839
rect 30190 2836 30196 2848
rect 28491 2808 30196 2836
rect 28491 2805 28503 2808
rect 28445 2799 28503 2805
rect 30190 2796 30196 2808
rect 30248 2796 30254 2848
rect 30300 2836 30328 2876
rect 32214 2864 32220 2916
rect 32272 2904 32278 2916
rect 33704 2904 33732 2935
rect 32272 2876 33732 2904
rect 32272 2864 32278 2876
rect 32766 2836 32772 2848
rect 30300 2808 32772 2836
rect 32766 2796 32772 2808
rect 32824 2796 32830 2848
rect 1104 2746 34868 2768
rect 1104 2694 5170 2746
rect 5222 2694 5234 2746
rect 5286 2694 5298 2746
rect 5350 2694 5362 2746
rect 5414 2694 5426 2746
rect 5478 2694 13611 2746
rect 13663 2694 13675 2746
rect 13727 2694 13739 2746
rect 13791 2694 13803 2746
rect 13855 2694 13867 2746
rect 13919 2694 22052 2746
rect 22104 2694 22116 2746
rect 22168 2694 22180 2746
rect 22232 2694 22244 2746
rect 22296 2694 22308 2746
rect 22360 2694 30493 2746
rect 30545 2694 30557 2746
rect 30609 2694 30621 2746
rect 30673 2694 30685 2746
rect 30737 2694 30749 2746
rect 30801 2694 34868 2746
rect 1104 2672 34868 2694
rect 15746 2632 15752 2644
rect 15707 2604 15752 2632
rect 15746 2592 15752 2604
rect 15804 2592 15810 2644
rect 17034 2632 17040 2644
rect 16995 2604 17040 2632
rect 17034 2592 17040 2604
rect 17092 2592 17098 2644
rect 18141 2635 18199 2641
rect 18141 2601 18153 2635
rect 18187 2632 18199 2635
rect 19058 2632 19064 2644
rect 18187 2604 19064 2632
rect 18187 2601 18199 2604
rect 18141 2595 18199 2601
rect 19058 2592 19064 2604
rect 19116 2592 19122 2644
rect 19521 2635 19579 2641
rect 19521 2601 19533 2635
rect 19567 2632 19579 2635
rect 19610 2632 19616 2644
rect 19567 2604 19616 2632
rect 19567 2601 19579 2604
rect 19521 2595 19579 2601
rect 19610 2592 19616 2604
rect 19668 2592 19674 2644
rect 20714 2592 20720 2644
rect 20772 2632 20778 2644
rect 20993 2635 21051 2641
rect 20993 2632 21005 2635
rect 20772 2604 21005 2632
rect 20772 2592 20778 2604
rect 20993 2601 21005 2604
rect 21039 2601 21051 2635
rect 20993 2595 21051 2601
rect 27801 2635 27859 2641
rect 27801 2601 27813 2635
rect 27847 2632 27859 2635
rect 30834 2632 30840 2644
rect 27847 2604 30840 2632
rect 27847 2601 27859 2604
rect 27801 2595 27859 2601
rect 30834 2592 30840 2604
rect 30892 2592 30898 2644
rect 4246 2564 4252 2576
rect 1596 2536 4252 2564
rect 1596 2505 1624 2536
rect 4246 2524 4252 2536
rect 4304 2524 4310 2576
rect 7374 2564 7380 2576
rect 6564 2536 7380 2564
rect 1581 2499 1639 2505
rect 1581 2465 1593 2499
rect 1627 2465 1639 2499
rect 2590 2496 2596 2508
rect 2551 2468 2596 2496
rect 1581 2459 1639 2465
rect 2590 2456 2596 2468
rect 2648 2456 2654 2508
rect 4154 2496 4160 2508
rect 4115 2468 4160 2496
rect 4154 2456 4160 2468
rect 4212 2456 4218 2508
rect 4522 2456 4528 2508
rect 4580 2496 4586 2508
rect 6564 2505 6592 2536
rect 7374 2524 7380 2536
rect 7432 2524 7438 2576
rect 28445 2567 28503 2573
rect 28445 2533 28457 2567
rect 28491 2564 28503 2567
rect 32122 2564 32128 2576
rect 28491 2536 32128 2564
rect 28491 2533 28503 2536
rect 28445 2527 28503 2533
rect 32122 2524 32128 2536
rect 32180 2524 32186 2576
rect 4617 2499 4675 2505
rect 4617 2496 4629 2499
rect 4580 2468 4629 2496
rect 4580 2456 4586 2468
rect 4617 2465 4629 2468
rect 4663 2465 4675 2499
rect 4617 2459 4675 2465
rect 6549 2499 6607 2505
rect 6549 2465 6561 2499
rect 6595 2465 6607 2499
rect 6730 2496 6736 2508
rect 6691 2468 6736 2496
rect 6549 2459 6607 2465
rect 6730 2456 6736 2468
rect 6788 2456 6794 2508
rect 6822 2456 6828 2508
rect 6880 2496 6886 2508
rect 7009 2499 7067 2505
rect 7009 2496 7021 2499
rect 6880 2468 7021 2496
rect 6880 2456 6886 2468
rect 7009 2465 7021 2468
rect 7055 2465 7067 2499
rect 7009 2459 7067 2465
rect 9125 2499 9183 2505
rect 9125 2465 9137 2499
rect 9171 2496 9183 2499
rect 9306 2496 9312 2508
rect 9171 2468 9312 2496
rect 9171 2465 9183 2468
rect 9125 2459 9183 2465
rect 9306 2456 9312 2468
rect 9364 2456 9370 2508
rect 9766 2496 9772 2508
rect 9727 2468 9772 2496
rect 9766 2456 9772 2468
rect 9824 2456 9830 2508
rect 29086 2496 29092 2508
rect 26206 2468 29092 2496
rect 15654 2428 15660 2440
rect 15615 2400 15660 2428
rect 15654 2388 15660 2400
rect 15712 2428 15718 2440
rect 16945 2431 17003 2437
rect 16945 2428 16957 2431
rect 15712 2400 16957 2428
rect 15712 2388 15718 2400
rect 16945 2397 16957 2400
rect 16991 2397 17003 2431
rect 16945 2391 17003 2397
rect 18230 2388 18236 2440
rect 18288 2428 18294 2440
rect 18325 2431 18383 2437
rect 18325 2428 18337 2431
rect 18288 2400 18337 2428
rect 18288 2388 18294 2400
rect 18325 2397 18337 2400
rect 18371 2397 18383 2431
rect 18325 2391 18383 2397
rect 19334 2388 19340 2440
rect 19392 2428 19398 2440
rect 19429 2431 19487 2437
rect 19429 2428 19441 2431
rect 19392 2400 19441 2428
rect 19392 2388 19398 2400
rect 19429 2397 19441 2400
rect 19475 2428 19487 2431
rect 26206 2428 26234 2468
rect 29086 2456 29092 2468
rect 29144 2456 29150 2508
rect 29917 2499 29975 2505
rect 29917 2465 29929 2499
rect 29963 2496 29975 2499
rect 30374 2496 30380 2508
rect 29963 2468 30380 2496
rect 29963 2465 29975 2468
rect 29917 2459 29975 2465
rect 30374 2456 30380 2468
rect 30432 2456 30438 2508
rect 30926 2496 30932 2508
rect 30887 2468 30932 2496
rect 30926 2456 30932 2468
rect 30984 2456 30990 2508
rect 31662 2456 31668 2508
rect 31720 2496 31726 2508
rect 32309 2499 32367 2505
rect 32309 2496 32321 2499
rect 31720 2468 32321 2496
rect 31720 2456 31726 2468
rect 32309 2465 32321 2468
rect 32355 2465 32367 2499
rect 32858 2496 32864 2508
rect 32819 2468 32864 2496
rect 32309 2459 32367 2465
rect 32858 2456 32864 2468
rect 32916 2456 32922 2508
rect 27706 2428 27712 2440
rect 19475 2400 26234 2428
rect 27619 2400 27712 2428
rect 19475 2397 19487 2400
rect 19429 2391 19487 2397
rect 27706 2388 27712 2400
rect 27764 2388 27770 2440
rect 28353 2431 28411 2437
rect 28353 2397 28365 2431
rect 28399 2428 28411 2431
rect 28534 2428 28540 2440
rect 28399 2400 28540 2428
rect 28399 2397 28411 2400
rect 28353 2391 28411 2397
rect 28534 2388 28540 2400
rect 28592 2388 28598 2440
rect 28994 2428 29000 2440
rect 28955 2400 29000 2428
rect 28994 2388 29000 2400
rect 29052 2388 29058 2440
rect 1765 2363 1823 2369
rect 1765 2329 1777 2363
rect 1811 2329 1823 2363
rect 1765 2323 1823 2329
rect 4341 2363 4399 2369
rect 4341 2329 4353 2363
rect 4387 2360 4399 2363
rect 5718 2360 5724 2372
rect 4387 2332 5724 2360
rect 4387 2329 4399 2332
rect 4341 2323 4399 2329
rect 1780 2292 1808 2323
rect 5718 2320 5724 2332
rect 5776 2320 5782 2372
rect 9306 2360 9312 2372
rect 9267 2332 9312 2360
rect 9306 2320 9312 2332
rect 9364 2320 9370 2372
rect 5810 2292 5816 2304
rect 1780 2264 5816 2292
rect 5810 2252 5816 2264
rect 5868 2252 5874 2304
rect 27724 2292 27752 2388
rect 29089 2363 29147 2369
rect 29089 2329 29101 2363
rect 29135 2360 29147 2363
rect 30101 2363 30159 2369
rect 30101 2360 30113 2363
rect 29135 2332 30113 2360
rect 29135 2329 29147 2332
rect 29089 2323 29147 2329
rect 30101 2329 30113 2332
rect 30147 2329 30159 2363
rect 30101 2323 30159 2329
rect 30190 2320 30196 2372
rect 30248 2360 30254 2372
rect 32493 2363 32551 2369
rect 32493 2360 32505 2363
rect 30248 2332 32505 2360
rect 30248 2320 30254 2332
rect 32493 2329 32505 2332
rect 32539 2329 32551 2363
rect 32493 2323 32551 2329
rect 33410 2292 33416 2304
rect 27724 2264 33416 2292
rect 33410 2252 33416 2264
rect 33468 2252 33474 2304
rect 1104 2202 35027 2224
rect 1104 2150 9390 2202
rect 9442 2150 9454 2202
rect 9506 2150 9518 2202
rect 9570 2150 9582 2202
rect 9634 2150 9646 2202
rect 9698 2150 17831 2202
rect 17883 2150 17895 2202
rect 17947 2150 17959 2202
rect 18011 2150 18023 2202
rect 18075 2150 18087 2202
rect 18139 2150 26272 2202
rect 26324 2150 26336 2202
rect 26388 2150 26400 2202
rect 26452 2150 26464 2202
rect 26516 2150 26528 2202
rect 26580 2150 34713 2202
rect 34765 2150 34777 2202
rect 34829 2150 34841 2202
rect 34893 2150 34905 2202
rect 34957 2150 34969 2202
rect 35021 2150 35027 2202
rect 1104 2128 35027 2150
rect 34514 1096 34520 1148
rect 34572 1136 34578 1148
rect 34790 1136 34796 1148
rect 34572 1108 34796 1136
rect 34572 1096 34578 1108
rect 34790 1096 34796 1108
rect 34848 1096 34854 1148
<< via1 >>
rect 20352 39992 20404 40044
rect 32496 39992 32548 40044
rect 23940 39788 23992 39840
rect 32588 39788 32640 39840
rect 5170 39686 5222 39738
rect 5234 39686 5286 39738
rect 5298 39686 5350 39738
rect 5362 39686 5414 39738
rect 5426 39686 5478 39738
rect 13611 39686 13663 39738
rect 13675 39686 13727 39738
rect 13739 39686 13791 39738
rect 13803 39686 13855 39738
rect 13867 39686 13919 39738
rect 22052 39686 22104 39738
rect 22116 39686 22168 39738
rect 22180 39686 22232 39738
rect 22244 39686 22296 39738
rect 22308 39686 22360 39738
rect 30493 39686 30545 39738
rect 30557 39686 30609 39738
rect 30621 39686 30673 39738
rect 30685 39686 30737 39738
rect 30749 39686 30801 39738
rect 18972 39584 19024 39636
rect 23940 39627 23992 39636
rect 23940 39593 23949 39627
rect 23949 39593 23983 39627
rect 23983 39593 23992 39627
rect 23940 39584 23992 39593
rect 25228 39584 25280 39636
rect 29460 39516 29512 39568
rect 32404 39584 32456 39636
rect 31300 39516 31352 39568
rect 7104 39491 7156 39500
rect 3884 39380 3936 39432
rect 4160 39380 4212 39432
rect 1308 39312 1360 39364
rect 3240 39244 3292 39296
rect 7104 39457 7113 39491
rect 7113 39457 7147 39491
rect 7147 39457 7156 39491
rect 7104 39448 7156 39457
rect 14832 39491 14884 39500
rect 14832 39457 14841 39491
rect 14841 39457 14875 39491
rect 14875 39457 14884 39491
rect 14832 39448 14884 39457
rect 9312 39423 9364 39432
rect 9312 39389 9321 39423
rect 9321 39389 9355 39423
rect 9355 39389 9364 39423
rect 9312 39380 9364 39389
rect 13728 39423 13780 39432
rect 13728 39389 13737 39423
rect 13737 39389 13771 39423
rect 13771 39389 13780 39423
rect 13728 39380 13780 39389
rect 14004 39380 14056 39432
rect 16856 39423 16908 39432
rect 16856 39389 16865 39423
rect 16865 39389 16899 39423
rect 16899 39389 16908 39423
rect 16856 39380 16908 39389
rect 6736 39355 6788 39364
rect 6736 39321 6745 39355
rect 6745 39321 6779 39355
rect 6779 39321 6788 39355
rect 6736 39312 6788 39321
rect 14464 39355 14516 39364
rect 14464 39321 14473 39355
rect 14473 39321 14507 39355
rect 14507 39321 14516 39355
rect 14464 39312 14516 39321
rect 17316 39380 17368 39432
rect 18696 39380 18748 39432
rect 19156 39380 19208 39432
rect 20260 39423 20312 39432
rect 20260 39389 20269 39423
rect 20269 39389 20303 39423
rect 20303 39389 20312 39423
rect 20260 39380 20312 39389
rect 21456 39380 21508 39432
rect 22100 39380 22152 39432
rect 23388 39423 23440 39432
rect 23388 39389 23397 39423
rect 23397 39389 23431 39423
rect 23431 39389 23440 39423
rect 23388 39380 23440 39389
rect 23848 39423 23900 39432
rect 23848 39389 23857 39423
rect 23857 39389 23891 39423
rect 23891 39389 23900 39423
rect 23848 39380 23900 39389
rect 26056 39423 26108 39432
rect 24400 39312 24452 39364
rect 26056 39389 26065 39423
rect 26065 39389 26099 39423
rect 26099 39389 26108 39423
rect 26056 39380 26108 39389
rect 7288 39244 7340 39296
rect 13452 39244 13504 39296
rect 16580 39244 16632 39296
rect 17040 39244 17092 39296
rect 18328 39244 18380 39296
rect 22192 39244 22244 39296
rect 24584 39244 24636 39296
rect 28448 39380 28500 39432
rect 28264 39312 28316 39364
rect 28632 39380 28684 39432
rect 29828 39380 29880 39432
rect 30564 39423 30616 39432
rect 30564 39389 30573 39423
rect 30573 39389 30607 39423
rect 30607 39389 30616 39423
rect 30564 39380 30616 39389
rect 30196 39312 30248 39364
rect 28540 39244 28592 39296
rect 29644 39244 29696 39296
rect 30380 39287 30432 39296
rect 30380 39253 30389 39287
rect 30389 39253 30423 39287
rect 30423 39253 30432 39287
rect 30380 39244 30432 39253
rect 32496 39423 32548 39432
rect 32496 39389 32505 39423
rect 32505 39389 32539 39423
rect 32539 39389 32548 39423
rect 32496 39380 32548 39389
rect 34336 39355 34388 39364
rect 34336 39321 34345 39355
rect 34345 39321 34379 39355
rect 34379 39321 34388 39355
rect 34336 39312 34388 39321
rect 30932 39244 30984 39296
rect 9390 39142 9442 39194
rect 9454 39142 9506 39194
rect 9518 39142 9570 39194
rect 9582 39142 9634 39194
rect 9646 39142 9698 39194
rect 17831 39142 17883 39194
rect 17895 39142 17947 39194
rect 17959 39142 18011 39194
rect 18023 39142 18075 39194
rect 18087 39142 18139 39194
rect 26272 39142 26324 39194
rect 26336 39142 26388 39194
rect 26400 39142 26452 39194
rect 26464 39142 26516 39194
rect 26528 39142 26580 39194
rect 34713 39142 34765 39194
rect 34777 39142 34829 39194
rect 34841 39142 34893 39194
rect 34905 39142 34957 39194
rect 34969 39142 35021 39194
rect 3516 39040 3568 39092
rect 5080 38972 5132 39024
rect 4160 38947 4212 38956
rect 4160 38913 4169 38947
rect 4169 38913 4203 38947
rect 4203 38913 4212 38947
rect 4160 38904 4212 38913
rect 23388 39040 23440 39092
rect 17040 39015 17092 39024
rect 17040 38981 17049 39015
rect 17049 38981 17083 39015
rect 17083 38981 17092 39015
rect 17040 38972 17092 38981
rect 22192 39015 22244 39024
rect 22192 38981 22201 39015
rect 22201 38981 22235 39015
rect 22235 38981 22244 39015
rect 22192 38972 22244 38981
rect 24584 39015 24636 39024
rect 24584 38981 24593 39015
rect 24593 38981 24627 39015
rect 24627 38981 24636 39015
rect 24584 38972 24636 38981
rect 26976 38972 27028 39024
rect 28264 38972 28316 39024
rect 29644 39015 29696 39024
rect 29644 38981 29653 39015
rect 29653 38981 29687 39015
rect 29687 38981 29696 39015
rect 29644 38972 29696 38981
rect 14004 38947 14056 38956
rect 2780 38879 2832 38888
rect 2780 38845 2789 38879
rect 2789 38845 2823 38879
rect 2823 38845 2832 38879
rect 2780 38836 2832 38845
rect 5540 38836 5592 38888
rect 5816 38879 5868 38888
rect 5816 38845 5825 38879
rect 5825 38845 5859 38879
rect 5859 38845 5868 38879
rect 5816 38836 5868 38845
rect 3976 38768 4028 38820
rect 14004 38913 14013 38947
rect 14013 38913 14047 38947
rect 14047 38913 14056 38947
rect 14004 38904 14056 38913
rect 19156 38947 19208 38956
rect 19156 38913 19165 38947
rect 19165 38913 19199 38947
rect 19199 38913 19208 38947
rect 19156 38904 19208 38913
rect 24400 38947 24452 38956
rect 24400 38913 24409 38947
rect 24409 38913 24443 38947
rect 24443 38913 24452 38947
rect 24400 38904 24452 38913
rect 29460 38947 29512 38956
rect 29460 38913 29469 38947
rect 29469 38913 29503 38947
rect 29503 38913 29512 38947
rect 29460 38904 29512 38913
rect 32588 39015 32640 39024
rect 32588 38981 32597 39015
rect 32597 38981 32631 39015
rect 32631 38981 32640 39015
rect 32588 38972 32640 38981
rect 8576 38879 8628 38888
rect 8576 38845 8585 38879
rect 8585 38845 8619 38879
rect 8619 38845 8628 38879
rect 8576 38836 8628 38845
rect 9036 38879 9088 38888
rect 9036 38845 9045 38879
rect 9045 38845 9079 38879
rect 9079 38845 9088 38879
rect 9036 38836 9088 38845
rect 3884 38700 3936 38752
rect 14372 38768 14424 38820
rect 15200 38836 15252 38888
rect 16120 38879 16172 38888
rect 16120 38845 16129 38879
rect 16129 38845 16163 38879
rect 16163 38845 16172 38879
rect 16120 38836 16172 38845
rect 17684 38836 17736 38888
rect 18236 38879 18288 38888
rect 18236 38845 18245 38879
rect 18245 38845 18279 38879
rect 18279 38845 18288 38879
rect 18236 38836 18288 38845
rect 19340 38879 19392 38888
rect 19340 38845 19349 38879
rect 19349 38845 19383 38879
rect 19383 38845 19392 38879
rect 19340 38836 19392 38845
rect 19984 38879 20036 38888
rect 19984 38845 19993 38879
rect 19993 38845 20027 38879
rect 20027 38845 20036 38879
rect 19984 38836 20036 38845
rect 22376 38836 22428 38888
rect 22560 38879 22612 38888
rect 22560 38845 22569 38879
rect 22569 38845 22603 38879
rect 22603 38845 22612 38879
rect 22560 38836 22612 38845
rect 25136 38879 25188 38888
rect 25136 38845 25145 38879
rect 25145 38845 25179 38879
rect 25179 38845 25188 38879
rect 25136 38836 25188 38845
rect 27344 38879 27396 38888
rect 15660 38768 15712 38820
rect 20536 38768 20588 38820
rect 27344 38845 27353 38879
rect 27353 38845 27387 38879
rect 27387 38845 27396 38879
rect 27344 38836 27396 38845
rect 8116 38700 8168 38752
rect 16672 38700 16724 38752
rect 23848 38700 23900 38752
rect 26976 38700 27028 38752
rect 27068 38700 27120 38752
rect 28356 38768 28408 38820
rect 30564 38836 30616 38888
rect 31852 38836 31904 38888
rect 32864 38879 32916 38888
rect 32864 38845 32873 38879
rect 32873 38845 32907 38879
rect 32907 38845 32916 38879
rect 32864 38836 32916 38845
rect 28448 38700 28500 38752
rect 32772 38700 32824 38752
rect 5170 38598 5222 38650
rect 5234 38598 5286 38650
rect 5298 38598 5350 38650
rect 5362 38598 5414 38650
rect 5426 38598 5478 38650
rect 13611 38598 13663 38650
rect 13675 38598 13727 38650
rect 13739 38598 13791 38650
rect 13803 38598 13855 38650
rect 13867 38598 13919 38650
rect 22052 38598 22104 38650
rect 22116 38598 22168 38650
rect 22180 38598 22232 38650
rect 22244 38598 22296 38650
rect 22308 38598 22360 38650
rect 30493 38598 30545 38650
rect 30557 38598 30609 38650
rect 30621 38598 30673 38650
rect 30685 38598 30737 38650
rect 30749 38598 30801 38650
rect 6736 38496 6788 38548
rect 8576 38496 8628 38548
rect 14464 38496 14516 38548
rect 15200 38539 15252 38548
rect 15200 38505 15209 38539
rect 15209 38505 15243 38539
rect 15243 38505 15252 38539
rect 15200 38496 15252 38505
rect 19340 38496 19392 38548
rect 22376 38496 22428 38548
rect 29368 38496 29420 38548
rect 16028 38428 16080 38480
rect 25044 38428 25096 38480
rect 25780 38428 25832 38480
rect 7748 38403 7800 38412
rect 664 38224 716 38276
rect 4160 38292 4212 38344
rect 4896 38292 4948 38344
rect 4436 38224 4488 38276
rect 7748 38369 7757 38403
rect 7757 38369 7791 38403
rect 7791 38369 7800 38403
rect 7748 38360 7800 38369
rect 16580 38403 16632 38412
rect 16580 38369 16589 38403
rect 16589 38369 16623 38403
rect 16623 38369 16632 38403
rect 16580 38360 16632 38369
rect 17408 38403 17460 38412
rect 17408 38369 17417 38403
rect 17417 38369 17451 38403
rect 17451 38369 17460 38403
rect 17408 38360 17460 38369
rect 20260 38360 20312 38412
rect 20628 38360 20680 38412
rect 26056 38360 26108 38412
rect 26424 38428 26476 38480
rect 9128 38335 9180 38344
rect 9128 38301 9137 38335
rect 9137 38301 9171 38335
rect 9171 38301 9180 38335
rect 9128 38292 9180 38301
rect 14280 38335 14332 38344
rect 14280 38301 14289 38335
rect 14289 38301 14323 38335
rect 14323 38301 14332 38335
rect 14280 38292 14332 38301
rect 14372 38292 14424 38344
rect 4068 38199 4120 38208
rect 4068 38165 4077 38199
rect 4077 38165 4111 38199
rect 4111 38165 4120 38199
rect 4068 38156 4120 38165
rect 7196 38224 7248 38276
rect 18604 38292 18656 38344
rect 24860 38292 24912 38344
rect 16856 38224 16908 38276
rect 20168 38267 20220 38276
rect 20168 38233 20177 38267
rect 20177 38233 20211 38267
rect 20211 38233 20220 38267
rect 20168 38224 20220 38233
rect 25136 38267 25188 38276
rect 25136 38233 25145 38267
rect 25145 38233 25179 38267
rect 25179 38233 25188 38267
rect 25136 38224 25188 38233
rect 7472 38156 7524 38208
rect 18236 38156 18288 38208
rect 24308 38156 24360 38208
rect 24492 38156 24544 38208
rect 27436 38335 27488 38344
rect 27436 38301 27445 38335
rect 27445 38301 27479 38335
rect 27479 38301 27488 38335
rect 27436 38292 27488 38301
rect 27620 38292 27672 38344
rect 28080 38199 28132 38208
rect 28080 38165 28089 38199
rect 28089 38165 28123 38199
rect 28123 38165 28132 38199
rect 28080 38156 28132 38165
rect 28356 38156 28408 38208
rect 29368 38360 29420 38412
rect 34152 38403 34204 38412
rect 34152 38369 34161 38403
rect 34161 38369 34195 38403
rect 34195 38369 34204 38403
rect 34152 38360 34204 38369
rect 32220 38292 32272 38344
rect 30288 38224 30340 38276
rect 31208 38156 31260 38208
rect 9390 38054 9442 38106
rect 9454 38054 9506 38106
rect 9518 38054 9570 38106
rect 9582 38054 9634 38106
rect 9646 38054 9698 38106
rect 17831 38054 17883 38106
rect 17895 38054 17947 38106
rect 17959 38054 18011 38106
rect 18023 38054 18075 38106
rect 18087 38054 18139 38106
rect 26272 38054 26324 38106
rect 26336 38054 26388 38106
rect 26400 38054 26452 38106
rect 26464 38054 26516 38106
rect 26528 38054 26580 38106
rect 34713 38054 34765 38106
rect 34777 38054 34829 38106
rect 34841 38054 34893 38106
rect 34905 38054 34957 38106
rect 34969 38054 35021 38106
rect 5540 37995 5592 38004
rect 5540 37961 5549 37995
rect 5549 37961 5583 37995
rect 5583 37961 5592 37995
rect 5540 37952 5592 37961
rect 7196 37995 7248 38004
rect 7196 37961 7205 37995
rect 7205 37961 7239 37995
rect 7239 37961 7248 37995
rect 7196 37952 7248 37961
rect 9128 37952 9180 38004
rect 18696 37952 18748 38004
rect 20168 37995 20220 38004
rect 20168 37961 20177 37995
rect 20177 37961 20211 37995
rect 20211 37961 20220 37995
rect 20168 37952 20220 37961
rect 3240 37927 3292 37936
rect 3240 37893 3249 37927
rect 3249 37893 3283 37927
rect 3283 37893 3292 37927
rect 3240 37884 3292 37893
rect 4896 37884 4948 37936
rect 8116 37927 8168 37936
rect 1676 37859 1728 37868
rect 1676 37825 1685 37859
rect 1685 37825 1719 37859
rect 1719 37825 1728 37859
rect 1676 37816 1728 37825
rect 2964 37816 3016 37868
rect 4804 37816 4856 37868
rect 6368 37816 6420 37868
rect 8116 37893 8125 37927
rect 8125 37893 8159 37927
rect 8159 37893 8168 37927
rect 8116 37884 8168 37893
rect 8392 37884 8444 37936
rect 3056 37791 3108 37800
rect 3056 37757 3065 37791
rect 3065 37757 3099 37791
rect 3099 37757 3108 37791
rect 3056 37748 3108 37757
rect 3424 37748 3476 37800
rect 9312 37748 9364 37800
rect 18604 37884 18656 37936
rect 23480 37952 23532 38004
rect 24492 37995 24544 38004
rect 24492 37961 24501 37995
rect 24501 37961 24535 37995
rect 24535 37961 24544 37995
rect 24492 37952 24544 37961
rect 22192 37884 22244 37936
rect 30288 37952 30340 38004
rect 25136 37927 25188 37936
rect 25136 37893 25145 37927
rect 25145 37893 25179 37927
rect 25179 37893 25188 37927
rect 25136 37884 25188 37893
rect 25320 37884 25372 37936
rect 30012 37884 30064 37936
rect 30104 37884 30156 37936
rect 34336 37927 34388 37936
rect 34336 37893 34345 37927
rect 34345 37893 34379 37927
rect 34379 37893 34388 37927
rect 34336 37884 34388 37893
rect 15660 37859 15712 37868
rect 15660 37825 15669 37859
rect 15669 37825 15703 37859
rect 15703 37825 15712 37859
rect 15660 37816 15712 37825
rect 16396 37816 16448 37868
rect 17132 37859 17184 37868
rect 17132 37825 17141 37859
rect 17141 37825 17175 37859
rect 17175 37825 17184 37859
rect 17132 37816 17184 37825
rect 17684 37816 17736 37868
rect 18972 37859 19024 37868
rect 18972 37825 18981 37859
rect 18981 37825 19015 37859
rect 19015 37825 19024 37859
rect 18972 37816 19024 37825
rect 20444 37816 20496 37868
rect 18696 37748 18748 37800
rect 23480 37816 23532 37868
rect 24400 37859 24452 37868
rect 24400 37825 24409 37859
rect 24409 37825 24443 37859
rect 24443 37825 24452 37859
rect 24400 37816 24452 37825
rect 25044 37859 25096 37868
rect 25044 37825 25053 37859
rect 25053 37825 25087 37859
rect 25087 37825 25096 37859
rect 25044 37816 25096 37825
rect 25320 37748 25372 37800
rect 27160 37859 27212 37868
rect 27160 37825 27169 37859
rect 27169 37825 27203 37859
rect 27203 37825 27212 37859
rect 27160 37816 27212 37825
rect 27436 37816 27488 37868
rect 31576 37859 31628 37868
rect 31576 37825 31585 37859
rect 31585 37825 31619 37859
rect 31619 37825 31628 37859
rect 31576 37816 31628 37825
rect 27528 37748 27580 37800
rect 27620 37748 27672 37800
rect 29000 37791 29052 37800
rect 29000 37757 29009 37791
rect 29009 37757 29043 37791
rect 29043 37757 29052 37791
rect 29000 37748 29052 37757
rect 29644 37748 29696 37800
rect 30932 37748 30984 37800
rect 31392 37791 31444 37800
rect 31392 37757 31401 37791
rect 31401 37757 31435 37791
rect 31435 37757 31444 37791
rect 31392 37748 31444 37757
rect 32496 37791 32548 37800
rect 16580 37680 16632 37732
rect 22192 37680 22244 37732
rect 5724 37612 5776 37664
rect 16028 37612 16080 37664
rect 16120 37655 16172 37664
rect 16120 37621 16129 37655
rect 16129 37621 16163 37655
rect 16163 37621 16172 37655
rect 16120 37612 16172 37621
rect 21180 37612 21232 37664
rect 21456 37655 21508 37664
rect 21456 37621 21465 37655
rect 21465 37621 21499 37655
rect 21499 37621 21508 37655
rect 21456 37612 21508 37621
rect 23756 37612 23808 37664
rect 24124 37612 24176 37664
rect 24308 37680 24360 37732
rect 25780 37612 25832 37664
rect 25964 37655 26016 37664
rect 25964 37621 25973 37655
rect 25973 37621 26007 37655
rect 26007 37621 26016 37655
rect 25964 37612 26016 37621
rect 27344 37680 27396 37732
rect 32496 37757 32505 37791
rect 32505 37757 32539 37791
rect 32539 37757 32548 37791
rect 32496 37748 32548 37757
rect 32588 37680 32640 37732
rect 5170 37510 5222 37562
rect 5234 37510 5286 37562
rect 5298 37510 5350 37562
rect 5362 37510 5414 37562
rect 5426 37510 5478 37562
rect 13611 37510 13663 37562
rect 13675 37510 13727 37562
rect 13739 37510 13791 37562
rect 13803 37510 13855 37562
rect 13867 37510 13919 37562
rect 22052 37510 22104 37562
rect 22116 37510 22168 37562
rect 22180 37510 22232 37562
rect 22244 37510 22296 37562
rect 22308 37510 22360 37562
rect 30493 37510 30545 37562
rect 30557 37510 30609 37562
rect 30621 37510 30673 37562
rect 30685 37510 30737 37562
rect 30749 37510 30801 37562
rect 3056 37408 3108 37460
rect 6368 37408 6420 37460
rect 3976 37340 4028 37392
rect 14280 37408 14332 37460
rect 15292 37408 15344 37460
rect 19248 37340 19300 37392
rect 2044 37315 2096 37324
rect 2044 37281 2053 37315
rect 2053 37281 2087 37315
rect 2087 37281 2096 37315
rect 2044 37272 2096 37281
rect 3332 37272 3384 37324
rect 2964 37204 3016 37256
rect 3976 37247 4028 37256
rect 3976 37213 3985 37247
rect 3985 37213 4019 37247
rect 4019 37213 4028 37247
rect 3976 37204 4028 37213
rect 5540 37204 5592 37256
rect 4068 37136 4120 37188
rect 4620 37136 4672 37188
rect 6736 37204 6788 37256
rect 19156 37272 19208 37324
rect 20352 37408 20404 37460
rect 21364 37451 21416 37460
rect 21364 37417 21373 37451
rect 21373 37417 21407 37451
rect 21407 37417 21416 37451
rect 21364 37408 21416 37417
rect 19432 37340 19484 37392
rect 24400 37408 24452 37460
rect 24860 37408 24912 37460
rect 25688 37408 25740 37460
rect 25780 37408 25832 37460
rect 30104 37408 30156 37460
rect 34060 37408 34112 37460
rect 7380 37247 7432 37256
rect 7380 37213 7389 37247
rect 7389 37213 7423 37247
rect 7423 37213 7432 37247
rect 7380 37204 7432 37213
rect 7472 37247 7524 37256
rect 7472 37213 7481 37247
rect 7481 37213 7515 37247
rect 7515 37213 7524 37247
rect 17408 37247 17460 37256
rect 7472 37204 7524 37213
rect 17408 37213 17417 37247
rect 17417 37213 17451 37247
rect 17451 37213 17460 37247
rect 17408 37204 17460 37213
rect 18604 37204 18656 37256
rect 18880 37247 18932 37256
rect 18880 37213 18889 37247
rect 18889 37213 18923 37247
rect 18923 37213 18932 37247
rect 18880 37204 18932 37213
rect 20444 37204 20496 37256
rect 21456 37272 21508 37324
rect 32496 37340 32548 37392
rect 21916 37204 21968 37256
rect 22468 37204 22520 37256
rect 22744 37204 22796 37256
rect 29920 37272 29972 37324
rect 30748 37272 30800 37324
rect 31484 37272 31536 37324
rect 33048 37315 33100 37324
rect 33048 37281 33057 37315
rect 33057 37281 33091 37315
rect 33091 37281 33100 37315
rect 33048 37272 33100 37281
rect 24032 37247 24084 37256
rect 24032 37213 24041 37247
rect 24041 37213 24075 37247
rect 24075 37213 24084 37247
rect 24032 37204 24084 37213
rect 24676 37247 24728 37256
rect 24676 37213 24685 37247
rect 24685 37213 24719 37247
rect 24719 37213 24728 37247
rect 24676 37204 24728 37213
rect 25320 37247 25372 37256
rect 25320 37213 25329 37247
rect 25329 37213 25363 37247
rect 25363 37213 25372 37247
rect 25320 37204 25372 37213
rect 26056 37204 26108 37256
rect 26976 37204 27028 37256
rect 28172 37247 28224 37256
rect 28172 37213 28181 37247
rect 28181 37213 28215 37247
rect 28215 37213 28224 37247
rect 28172 37204 28224 37213
rect 29184 37247 29236 37256
rect 29184 37213 29193 37247
rect 29193 37213 29227 37247
rect 29227 37213 29236 37247
rect 29184 37204 29236 37213
rect 30104 37247 30156 37256
rect 30104 37213 30113 37247
rect 30113 37213 30147 37247
rect 30147 37213 30156 37247
rect 30104 37204 30156 37213
rect 30288 37204 30340 37256
rect 4160 37068 4212 37120
rect 6828 37068 6880 37120
rect 14280 37068 14332 37120
rect 17500 37111 17552 37120
rect 17500 37077 17509 37111
rect 17509 37077 17543 37111
rect 17543 37077 17552 37111
rect 17500 37068 17552 37077
rect 19064 37068 19116 37120
rect 20720 37111 20772 37120
rect 20720 37077 20729 37111
rect 20729 37077 20763 37111
rect 20763 37077 20772 37111
rect 20720 37068 20772 37077
rect 30012 37136 30064 37188
rect 31576 37204 31628 37256
rect 32496 37247 32548 37256
rect 32496 37213 32505 37247
rect 32505 37213 32539 37247
rect 32539 37213 32548 37247
rect 32496 37204 32548 37213
rect 31116 37136 31168 37188
rect 32680 37179 32732 37188
rect 32680 37145 32689 37179
rect 32689 37145 32723 37179
rect 32723 37145 32732 37179
rect 32680 37136 32732 37145
rect 23572 37068 23624 37120
rect 24768 37111 24820 37120
rect 24768 37077 24777 37111
rect 24777 37077 24811 37111
rect 24811 37077 24820 37111
rect 24768 37068 24820 37077
rect 25412 37111 25464 37120
rect 25412 37077 25421 37111
rect 25421 37077 25455 37111
rect 25455 37077 25464 37111
rect 25412 37068 25464 37077
rect 26976 37068 27028 37120
rect 27160 37111 27212 37120
rect 27160 37077 27169 37111
rect 27169 37077 27203 37111
rect 27203 37077 27212 37111
rect 27160 37068 27212 37077
rect 27988 37111 28040 37120
rect 27988 37077 27997 37111
rect 27997 37077 28031 37111
rect 28031 37077 28040 37111
rect 27988 37068 28040 37077
rect 29368 37068 29420 37120
rect 29736 37068 29788 37120
rect 30564 37068 30616 37120
rect 30932 37068 30984 37120
rect 32036 37111 32088 37120
rect 32036 37077 32045 37111
rect 32045 37077 32079 37111
rect 32079 37077 32088 37111
rect 32036 37068 32088 37077
rect 9390 36966 9442 37018
rect 9454 36966 9506 37018
rect 9518 36966 9570 37018
rect 9582 36966 9634 37018
rect 9646 36966 9698 37018
rect 17831 36966 17883 37018
rect 17895 36966 17947 37018
rect 17959 36966 18011 37018
rect 18023 36966 18075 37018
rect 18087 36966 18139 37018
rect 26272 36966 26324 37018
rect 26336 36966 26388 37018
rect 26400 36966 26452 37018
rect 26464 36966 26516 37018
rect 26528 36966 26580 37018
rect 34713 36966 34765 37018
rect 34777 36966 34829 37018
rect 34841 36966 34893 37018
rect 34905 36966 34957 37018
rect 34969 36966 35021 37018
rect 5540 36864 5592 36916
rect 7288 36907 7340 36916
rect 7288 36873 7297 36907
rect 7297 36873 7331 36907
rect 7331 36873 7340 36907
rect 7288 36864 7340 36873
rect 20720 36864 20772 36916
rect 32680 36864 32732 36916
rect 3976 36728 4028 36780
rect 5540 36771 5592 36780
rect 5540 36737 5549 36771
rect 5549 36737 5583 36771
rect 5583 36737 5592 36771
rect 5540 36728 5592 36737
rect 5724 36728 5776 36780
rect 6552 36771 6604 36780
rect 6552 36737 6561 36771
rect 6561 36737 6595 36771
rect 6595 36737 6604 36771
rect 6552 36728 6604 36737
rect 7380 36728 7432 36780
rect 17316 36728 17368 36780
rect 17592 36771 17644 36780
rect 17592 36737 17601 36771
rect 17601 36737 17635 36771
rect 17635 36737 17644 36771
rect 17592 36728 17644 36737
rect 18236 36771 18288 36780
rect 18236 36737 18245 36771
rect 18245 36737 18279 36771
rect 18279 36737 18288 36771
rect 18236 36728 18288 36737
rect 18696 36771 18748 36780
rect 18696 36737 18705 36771
rect 18705 36737 18739 36771
rect 18739 36737 18748 36771
rect 18696 36728 18748 36737
rect 19340 36771 19392 36780
rect 19340 36737 19349 36771
rect 19349 36737 19383 36771
rect 19383 36737 19392 36771
rect 19340 36728 19392 36737
rect 20536 36728 20588 36780
rect 2780 36703 2832 36712
rect 2780 36669 2789 36703
rect 2789 36669 2823 36703
rect 2823 36669 2832 36703
rect 2780 36660 2832 36669
rect 4436 36703 4488 36712
rect 4436 36669 4445 36703
rect 4445 36669 4479 36703
rect 4479 36669 4488 36703
rect 4436 36660 4488 36669
rect 4988 36660 5040 36712
rect 5080 36660 5132 36712
rect 20444 36660 20496 36712
rect 20628 36703 20680 36712
rect 20628 36669 20637 36703
rect 20637 36669 20671 36703
rect 20671 36669 20680 36703
rect 20628 36660 20680 36669
rect 27620 36796 27672 36848
rect 22376 36771 22428 36780
rect 22376 36737 22385 36771
rect 22385 36737 22419 36771
rect 22419 36737 22428 36771
rect 22376 36728 22428 36737
rect 22928 36728 22980 36780
rect 24492 36771 24544 36780
rect 24492 36737 24501 36771
rect 24501 36737 24535 36771
rect 24535 36737 24544 36771
rect 24492 36728 24544 36737
rect 25136 36771 25188 36780
rect 25136 36737 25145 36771
rect 25145 36737 25179 36771
rect 25179 36737 25188 36771
rect 25136 36728 25188 36737
rect 25872 36771 25924 36780
rect 25872 36737 25881 36771
rect 25881 36737 25915 36771
rect 25915 36737 25924 36771
rect 25872 36728 25924 36737
rect 26424 36771 26476 36780
rect 26424 36737 26433 36771
rect 26433 36737 26467 36771
rect 26467 36737 26476 36771
rect 26424 36728 26476 36737
rect 26516 36728 26568 36780
rect 28540 36728 28592 36780
rect 30012 36796 30064 36848
rect 30564 36796 30616 36848
rect 29092 36771 29144 36780
rect 29092 36737 29101 36771
rect 29101 36737 29135 36771
rect 29135 36737 29144 36771
rect 29092 36728 29144 36737
rect 29460 36728 29512 36780
rect 29552 36728 29604 36780
rect 25320 36660 25372 36712
rect 31208 36839 31260 36848
rect 31208 36805 31217 36839
rect 31217 36805 31251 36839
rect 31251 36805 31260 36839
rect 31208 36796 31260 36805
rect 30840 36703 30892 36712
rect 30840 36669 30849 36703
rect 30849 36669 30883 36703
rect 30883 36669 30892 36703
rect 30840 36660 30892 36669
rect 31944 36660 31996 36712
rect 33508 36703 33560 36712
rect 33508 36669 33517 36703
rect 33517 36669 33551 36703
rect 33551 36669 33560 36703
rect 33508 36660 33560 36669
rect 27896 36592 27948 36644
rect 30932 36592 30984 36644
rect 17684 36524 17736 36576
rect 18972 36524 19024 36576
rect 20536 36524 20588 36576
rect 22560 36524 22612 36576
rect 23388 36524 23440 36576
rect 23664 36567 23716 36576
rect 23664 36533 23673 36567
rect 23673 36533 23707 36567
rect 23707 36533 23716 36567
rect 23664 36524 23716 36533
rect 24308 36567 24360 36576
rect 24308 36533 24317 36567
rect 24317 36533 24351 36567
rect 24351 36533 24360 36567
rect 24308 36524 24360 36533
rect 24860 36524 24912 36576
rect 25688 36567 25740 36576
rect 25688 36533 25697 36567
rect 25697 36533 25731 36567
rect 25731 36533 25740 36567
rect 25688 36524 25740 36533
rect 26148 36524 26200 36576
rect 26516 36524 26568 36576
rect 27160 36567 27212 36576
rect 27160 36533 27169 36567
rect 27169 36533 27203 36567
rect 27203 36533 27212 36567
rect 27160 36524 27212 36533
rect 27252 36524 27304 36576
rect 28448 36567 28500 36576
rect 28448 36533 28457 36567
rect 28457 36533 28491 36567
rect 28491 36533 28500 36567
rect 28448 36524 28500 36533
rect 28540 36524 28592 36576
rect 29276 36524 29328 36576
rect 29920 36524 29972 36576
rect 30288 36524 30340 36576
rect 32956 36524 33008 36576
rect 5170 36422 5222 36474
rect 5234 36422 5286 36474
rect 5298 36422 5350 36474
rect 5362 36422 5414 36474
rect 5426 36422 5478 36474
rect 13611 36422 13663 36474
rect 13675 36422 13727 36474
rect 13739 36422 13791 36474
rect 13803 36422 13855 36474
rect 13867 36422 13919 36474
rect 22052 36422 22104 36474
rect 22116 36422 22168 36474
rect 22180 36422 22232 36474
rect 22244 36422 22296 36474
rect 22308 36422 22360 36474
rect 30493 36422 30545 36474
rect 30557 36422 30609 36474
rect 30621 36422 30673 36474
rect 30685 36422 30737 36474
rect 30749 36422 30801 36474
rect 22744 36320 22796 36372
rect 22928 36363 22980 36372
rect 22928 36329 22937 36363
rect 22937 36329 22971 36363
rect 22971 36329 22980 36363
rect 22928 36320 22980 36329
rect 26056 36363 26108 36372
rect 26056 36329 26065 36363
rect 26065 36329 26099 36363
rect 26099 36329 26108 36363
rect 26056 36320 26108 36329
rect 27068 36320 27120 36372
rect 27528 36320 27580 36372
rect 30196 36363 30248 36372
rect 30196 36329 30205 36363
rect 30205 36329 30239 36363
rect 30239 36329 30248 36363
rect 30196 36320 30248 36329
rect 31024 36363 31076 36372
rect 31024 36329 31033 36363
rect 31033 36329 31067 36363
rect 31067 36329 31076 36363
rect 31024 36320 31076 36329
rect 31760 36320 31812 36372
rect 32220 36320 32272 36372
rect 19340 36252 19392 36304
rect 3240 36227 3292 36236
rect 3240 36193 3249 36227
rect 3249 36193 3283 36227
rect 3283 36193 3292 36227
rect 3240 36184 3292 36193
rect 1768 36116 1820 36168
rect 2044 36116 2096 36168
rect 4804 36184 4856 36236
rect 3976 36159 4028 36168
rect 3976 36125 3985 36159
rect 3985 36125 4019 36159
rect 4019 36125 4028 36159
rect 3976 36116 4028 36125
rect 4804 36091 4856 36100
rect 4804 36057 4813 36091
rect 4813 36057 4847 36091
rect 4847 36057 4856 36091
rect 9128 36116 9180 36168
rect 18420 36159 18472 36168
rect 18420 36125 18429 36159
rect 18429 36125 18463 36159
rect 18463 36125 18472 36159
rect 18420 36116 18472 36125
rect 19800 36159 19852 36168
rect 19800 36125 19809 36159
rect 19809 36125 19843 36159
rect 19843 36125 19852 36159
rect 19800 36116 19852 36125
rect 25228 36252 25280 36304
rect 25320 36252 25372 36304
rect 28724 36252 28776 36304
rect 30288 36252 30340 36304
rect 20628 36159 20680 36168
rect 20628 36125 20637 36159
rect 20637 36125 20671 36159
rect 20671 36125 20680 36159
rect 20628 36116 20680 36125
rect 21272 36159 21324 36168
rect 21272 36125 21281 36159
rect 21281 36125 21315 36159
rect 21315 36125 21324 36159
rect 21272 36116 21324 36125
rect 21916 36159 21968 36168
rect 21916 36125 21925 36159
rect 21925 36125 21959 36159
rect 21959 36125 21968 36159
rect 21916 36116 21968 36125
rect 22652 36159 22704 36168
rect 22652 36125 22661 36159
rect 22661 36125 22695 36159
rect 22695 36125 22704 36159
rect 22652 36116 22704 36125
rect 22744 36159 22796 36168
rect 22744 36125 22753 36159
rect 22753 36125 22787 36159
rect 22787 36125 22796 36159
rect 22744 36116 22796 36125
rect 23296 36116 23348 36168
rect 23572 36159 23624 36168
rect 23572 36125 23581 36159
rect 23581 36125 23615 36159
rect 23615 36125 23624 36159
rect 23572 36116 23624 36125
rect 25780 36159 25832 36168
rect 25780 36125 25789 36159
rect 25789 36125 25823 36159
rect 25823 36125 25832 36159
rect 25780 36116 25832 36125
rect 26608 36184 26660 36236
rect 29184 36227 29236 36236
rect 27344 36159 27396 36168
rect 4804 36048 4856 36057
rect 6552 35980 6604 36032
rect 17408 36048 17460 36100
rect 27344 36125 27353 36159
rect 27353 36125 27387 36159
rect 27387 36125 27396 36159
rect 27344 36116 27396 36125
rect 29184 36193 29193 36227
rect 29193 36193 29227 36227
rect 29227 36193 29236 36227
rect 30840 36252 30892 36304
rect 29184 36184 29236 36193
rect 27804 36116 27856 36168
rect 28264 36116 28316 36168
rect 28908 36159 28960 36168
rect 28908 36125 28917 36159
rect 28917 36125 28951 36159
rect 28951 36125 28960 36159
rect 28908 36116 28960 36125
rect 29920 36159 29972 36168
rect 29920 36125 29929 36159
rect 29929 36125 29963 36159
rect 29963 36125 29972 36159
rect 29920 36116 29972 36125
rect 31116 36184 31168 36236
rect 34336 36227 34388 36236
rect 34336 36193 34345 36227
rect 34345 36193 34379 36227
rect 34379 36193 34388 36227
rect 34336 36184 34388 36193
rect 18236 36023 18288 36032
rect 18236 35989 18245 36023
rect 18245 35989 18279 36023
rect 18279 35989 18288 36023
rect 18236 35980 18288 35989
rect 19892 36023 19944 36032
rect 19892 35989 19901 36023
rect 19901 35989 19935 36023
rect 19935 35989 19944 36023
rect 19892 35980 19944 35989
rect 20168 35980 20220 36032
rect 21088 36023 21140 36032
rect 21088 35989 21097 36023
rect 21097 35989 21131 36023
rect 21131 35989 21140 36023
rect 21088 35980 21140 35989
rect 22468 35980 22520 36032
rect 24676 35980 24728 36032
rect 26884 36023 26936 36032
rect 26884 35989 26893 36023
rect 26893 35989 26927 36023
rect 26927 35989 26936 36023
rect 29092 36048 29144 36100
rect 26884 35980 26936 35989
rect 27436 35980 27488 36032
rect 28724 35980 28776 36032
rect 29368 35980 29420 36032
rect 30196 36048 30248 36100
rect 31576 36116 31628 36168
rect 32036 36048 32088 36100
rect 9390 35878 9442 35930
rect 9454 35878 9506 35930
rect 9518 35878 9570 35930
rect 9582 35878 9634 35930
rect 9646 35878 9698 35930
rect 17831 35878 17883 35930
rect 17895 35878 17947 35930
rect 17959 35878 18011 35930
rect 18023 35878 18075 35930
rect 18087 35878 18139 35930
rect 26272 35878 26324 35930
rect 26336 35878 26388 35930
rect 26400 35878 26452 35930
rect 26464 35878 26516 35930
rect 26528 35878 26580 35930
rect 34713 35878 34765 35930
rect 34777 35878 34829 35930
rect 34841 35878 34893 35930
rect 34905 35878 34957 35930
rect 34969 35878 35021 35930
rect 21272 35776 21324 35828
rect 22376 35776 22428 35828
rect 25136 35776 25188 35828
rect 28172 35776 28224 35828
rect 29184 35776 29236 35828
rect 30012 35776 30064 35828
rect 18236 35708 18288 35760
rect 24308 35708 24360 35760
rect 25780 35708 25832 35760
rect 2504 35640 2556 35692
rect 3976 35640 4028 35692
rect 16580 35640 16632 35692
rect 17684 35640 17736 35692
rect 2044 35615 2096 35624
rect 2044 35581 2053 35615
rect 2053 35581 2087 35615
rect 2087 35581 2096 35615
rect 2044 35572 2096 35581
rect 3884 35615 3936 35624
rect 3884 35581 3893 35615
rect 3893 35581 3927 35615
rect 3927 35581 3936 35615
rect 3884 35572 3936 35581
rect 6552 35572 6604 35624
rect 17592 35479 17644 35488
rect 17592 35445 17601 35479
rect 17601 35445 17635 35479
rect 17635 35445 17644 35479
rect 17592 35436 17644 35445
rect 19248 35436 19300 35488
rect 19524 35479 19576 35488
rect 19524 35445 19533 35479
rect 19533 35445 19567 35479
rect 19567 35445 19576 35479
rect 19524 35436 19576 35445
rect 19984 35479 20036 35488
rect 19984 35445 19993 35479
rect 19993 35445 20027 35479
rect 20027 35445 20036 35479
rect 19984 35436 20036 35445
rect 20720 35640 20772 35692
rect 20996 35683 21048 35692
rect 20996 35649 21005 35683
rect 21005 35649 21039 35683
rect 21039 35649 21048 35683
rect 20996 35640 21048 35649
rect 21272 35640 21324 35692
rect 22744 35640 22796 35692
rect 25228 35683 25280 35692
rect 20628 35572 20680 35624
rect 22928 35572 22980 35624
rect 23388 35615 23440 35624
rect 23388 35581 23397 35615
rect 23397 35581 23431 35615
rect 23431 35581 23440 35615
rect 23388 35572 23440 35581
rect 25228 35649 25237 35683
rect 25237 35649 25271 35683
rect 25271 35649 25280 35683
rect 25228 35640 25280 35649
rect 26608 35640 26660 35692
rect 25136 35572 25188 35624
rect 27068 35640 27120 35692
rect 27896 35708 27948 35760
rect 31944 35708 31996 35760
rect 29920 35683 29972 35692
rect 29920 35649 29929 35683
rect 29929 35649 29963 35683
rect 29963 35649 29972 35683
rect 29920 35640 29972 35649
rect 30196 35640 30248 35692
rect 26792 35572 26844 35624
rect 27344 35572 27396 35624
rect 28080 35572 28132 35624
rect 28540 35572 28592 35624
rect 28816 35572 28868 35624
rect 29184 35572 29236 35624
rect 31024 35572 31076 35624
rect 31668 35640 31720 35692
rect 31760 35640 31812 35692
rect 32956 35640 33008 35692
rect 34060 35751 34112 35760
rect 34060 35717 34069 35751
rect 34069 35717 34103 35751
rect 34103 35717 34112 35751
rect 34060 35708 34112 35717
rect 28632 35504 28684 35556
rect 30840 35504 30892 35556
rect 31852 35572 31904 35624
rect 32864 35572 32916 35624
rect 33508 35572 33560 35624
rect 23112 35436 23164 35488
rect 25504 35436 25556 35488
rect 26056 35436 26108 35488
rect 26516 35436 26568 35488
rect 27528 35479 27580 35488
rect 27528 35445 27537 35479
rect 27537 35445 27571 35479
rect 27571 35445 27580 35479
rect 27528 35436 27580 35445
rect 27620 35436 27672 35488
rect 30932 35436 30984 35488
rect 31760 35479 31812 35488
rect 31760 35445 31769 35479
rect 31769 35445 31803 35479
rect 31803 35445 31812 35479
rect 31760 35436 31812 35445
rect 32772 35479 32824 35488
rect 32772 35445 32781 35479
rect 32781 35445 32815 35479
rect 32815 35445 32824 35479
rect 32772 35436 32824 35445
rect 33140 35436 33192 35488
rect 33692 35436 33744 35488
rect 5170 35334 5222 35386
rect 5234 35334 5286 35386
rect 5298 35334 5350 35386
rect 5362 35334 5414 35386
rect 5426 35334 5478 35386
rect 13611 35334 13663 35386
rect 13675 35334 13727 35386
rect 13739 35334 13791 35386
rect 13803 35334 13855 35386
rect 13867 35334 13919 35386
rect 22052 35334 22104 35386
rect 22116 35334 22168 35386
rect 22180 35334 22232 35386
rect 22244 35334 22296 35386
rect 22308 35334 22360 35386
rect 30493 35334 30545 35386
rect 30557 35334 30609 35386
rect 30621 35334 30673 35386
rect 30685 35334 30737 35386
rect 30749 35334 30801 35386
rect 18420 35232 18472 35284
rect 20628 35232 20680 35284
rect 22376 35232 22428 35284
rect 22928 35275 22980 35284
rect 22928 35241 22937 35275
rect 22937 35241 22971 35275
rect 22971 35241 22980 35275
rect 22928 35232 22980 35241
rect 2780 35139 2832 35148
rect 2780 35105 2789 35139
rect 2789 35105 2823 35139
rect 2823 35105 2832 35139
rect 2780 35096 2832 35105
rect 16672 35096 16724 35148
rect 21364 35164 21416 35216
rect 23296 35232 23348 35284
rect 25872 35232 25924 35284
rect 27160 35232 27212 35284
rect 23112 35164 23164 35216
rect 29000 35164 29052 35216
rect 29368 35164 29420 35216
rect 29644 35164 29696 35216
rect 29828 35164 29880 35216
rect 3976 35071 4028 35080
rect 3976 35037 3985 35071
rect 3985 35037 4019 35071
rect 4019 35037 4028 35071
rect 3976 35028 4028 35037
rect 2136 34960 2188 35012
rect 2504 34960 2556 35012
rect 4712 34960 4764 35012
rect 5540 34960 5592 35012
rect 18328 35071 18380 35080
rect 18328 35037 18337 35071
rect 18337 35037 18371 35071
rect 18371 35037 18380 35071
rect 18328 35028 18380 35037
rect 19524 35071 19576 35080
rect 19524 35037 19533 35071
rect 19533 35037 19567 35071
rect 19567 35037 19576 35071
rect 19524 35028 19576 35037
rect 20996 35028 21048 35080
rect 21456 35096 21508 35148
rect 22192 35071 22244 35080
rect 20260 35003 20312 35012
rect 2872 34892 2924 34944
rect 18328 34892 18380 34944
rect 19800 34935 19852 34944
rect 19800 34901 19809 34935
rect 19809 34901 19843 34935
rect 19843 34901 19852 34935
rect 19800 34892 19852 34901
rect 20260 34969 20269 35003
rect 20269 34969 20303 35003
rect 20303 34969 20312 35003
rect 20260 34960 20312 34969
rect 22192 35037 22201 35071
rect 22201 35037 22235 35071
rect 22235 35037 22244 35071
rect 22192 35028 22244 35037
rect 22744 35096 22796 35148
rect 24584 35139 24636 35148
rect 24584 35105 24593 35139
rect 24593 35105 24627 35139
rect 24627 35105 24636 35139
rect 24584 35096 24636 35105
rect 28632 35096 28684 35148
rect 23296 35028 23348 35080
rect 24860 35071 24912 35080
rect 22376 34960 22428 35012
rect 20444 34935 20496 34944
rect 20444 34901 20453 34935
rect 20453 34901 20487 34935
rect 20487 34901 20496 34935
rect 20444 34892 20496 34901
rect 20628 34935 20680 34944
rect 20628 34901 20637 34935
rect 20637 34901 20671 34935
rect 20671 34901 20680 34935
rect 20628 34892 20680 34901
rect 20812 34935 20864 34944
rect 20812 34901 20821 34935
rect 20821 34901 20855 34935
rect 20855 34901 20864 34935
rect 20812 34892 20864 34901
rect 21640 34935 21692 34944
rect 21640 34901 21649 34935
rect 21649 34901 21683 34935
rect 21683 34901 21692 34935
rect 21640 34892 21692 34901
rect 22192 34892 22244 34944
rect 23572 34960 23624 35012
rect 24860 35037 24894 35071
rect 24894 35037 24912 35071
rect 24860 35028 24912 35037
rect 26516 35071 26568 35080
rect 26516 35037 26525 35071
rect 26525 35037 26559 35071
rect 26559 35037 26568 35071
rect 26516 35028 26568 35037
rect 27160 35028 27212 35080
rect 29828 35071 29880 35080
rect 22744 34892 22796 34944
rect 24860 34892 24912 34944
rect 25872 34892 25924 34944
rect 27712 34960 27764 35012
rect 27988 34960 28040 35012
rect 29828 35037 29837 35071
rect 29837 35037 29871 35071
rect 29871 35037 29880 35071
rect 29828 35028 29880 35037
rect 29920 35071 29972 35080
rect 29920 35037 29929 35071
rect 29929 35037 29963 35071
rect 29963 35037 29972 35071
rect 29920 35028 29972 35037
rect 30104 34960 30156 35012
rect 32128 35028 32180 35080
rect 27620 34892 27672 34944
rect 28264 34892 28316 34944
rect 28816 34892 28868 34944
rect 29368 34892 29420 34944
rect 34612 34960 34664 35012
rect 31668 34892 31720 34944
rect 32036 34935 32088 34944
rect 32036 34901 32045 34935
rect 32045 34901 32079 34935
rect 32079 34901 32088 34935
rect 32036 34892 32088 34901
rect 9390 34790 9442 34842
rect 9454 34790 9506 34842
rect 9518 34790 9570 34842
rect 9582 34790 9634 34842
rect 9646 34790 9698 34842
rect 17831 34790 17883 34842
rect 17895 34790 17947 34842
rect 17959 34790 18011 34842
rect 18023 34790 18075 34842
rect 18087 34790 18139 34842
rect 26272 34790 26324 34842
rect 26336 34790 26388 34842
rect 26400 34790 26452 34842
rect 26464 34790 26516 34842
rect 26528 34790 26580 34842
rect 34713 34790 34765 34842
rect 34777 34790 34829 34842
rect 34841 34790 34893 34842
rect 34905 34790 34957 34842
rect 34969 34790 35021 34842
rect 17132 34688 17184 34740
rect 1768 34595 1820 34604
rect 1768 34561 1777 34595
rect 1777 34561 1811 34595
rect 1811 34561 1820 34595
rect 1768 34552 1820 34561
rect 18236 34620 18288 34672
rect 20260 34688 20312 34740
rect 20628 34731 20680 34740
rect 20628 34697 20637 34731
rect 20637 34697 20671 34731
rect 20671 34697 20680 34731
rect 20628 34688 20680 34697
rect 20720 34688 20772 34740
rect 22652 34688 22704 34740
rect 23296 34688 23348 34740
rect 23940 34688 23992 34740
rect 24584 34688 24636 34740
rect 25412 34688 25464 34740
rect 28540 34731 28592 34740
rect 19340 34620 19392 34672
rect 19984 34620 20036 34672
rect 18696 34552 18748 34604
rect 19248 34595 19300 34604
rect 19248 34561 19257 34595
rect 19257 34561 19291 34595
rect 19291 34561 19300 34595
rect 19248 34552 19300 34561
rect 21272 34595 21324 34604
rect 21272 34561 21281 34595
rect 21281 34561 21315 34595
rect 21315 34561 21324 34595
rect 21272 34552 21324 34561
rect 21456 34552 21508 34604
rect 21732 34552 21784 34604
rect 23664 34620 23716 34672
rect 24216 34620 24268 34672
rect 26976 34620 27028 34672
rect 22560 34552 22612 34604
rect 23388 34552 23440 34604
rect 23940 34552 23992 34604
rect 24400 34552 24452 34604
rect 25780 34552 25832 34604
rect 28540 34697 28549 34731
rect 28549 34697 28583 34731
rect 28583 34697 28592 34731
rect 28540 34688 28592 34697
rect 29276 34688 29328 34740
rect 29828 34688 29880 34740
rect 31208 34688 31260 34740
rect 31300 34688 31352 34740
rect 31760 34688 31812 34740
rect 29920 34620 29972 34672
rect 30104 34620 30156 34672
rect 1952 34527 2004 34536
rect 1952 34493 1961 34527
rect 1961 34493 1995 34527
rect 1995 34493 2004 34527
rect 1952 34484 2004 34493
rect 2780 34527 2832 34536
rect 2780 34493 2789 34527
rect 2789 34493 2823 34527
rect 2823 34493 2832 34527
rect 2780 34484 2832 34493
rect 20996 34484 21048 34536
rect 26424 34484 26476 34536
rect 27160 34527 27212 34536
rect 27160 34493 27169 34527
rect 27169 34493 27203 34527
rect 27203 34493 27212 34527
rect 27160 34484 27212 34493
rect 28816 34552 28868 34604
rect 30012 34552 30064 34604
rect 30564 34620 30616 34672
rect 34336 34663 34388 34672
rect 34336 34629 34345 34663
rect 34345 34629 34379 34663
rect 34379 34629 34388 34663
rect 34336 34620 34388 34629
rect 32496 34595 32548 34604
rect 20536 34416 20588 34468
rect 21824 34416 21876 34468
rect 16120 34348 16172 34400
rect 21272 34348 21324 34400
rect 21548 34348 21600 34400
rect 23756 34416 23808 34468
rect 25044 34416 25096 34468
rect 29368 34484 29420 34536
rect 32496 34561 32505 34595
rect 32505 34561 32539 34595
rect 32539 34561 32548 34595
rect 32496 34552 32548 34561
rect 23020 34348 23072 34400
rect 29828 34348 29880 34400
rect 30104 34348 30156 34400
rect 31576 34348 31628 34400
rect 5170 34246 5222 34298
rect 5234 34246 5286 34298
rect 5298 34246 5350 34298
rect 5362 34246 5414 34298
rect 5426 34246 5478 34298
rect 13611 34246 13663 34298
rect 13675 34246 13727 34298
rect 13739 34246 13791 34298
rect 13803 34246 13855 34298
rect 13867 34246 13919 34298
rect 22052 34246 22104 34298
rect 22116 34246 22168 34298
rect 22180 34246 22232 34298
rect 22244 34246 22296 34298
rect 22308 34246 22360 34298
rect 30493 34246 30545 34298
rect 30557 34246 30609 34298
rect 30621 34246 30673 34298
rect 30685 34246 30737 34298
rect 30749 34246 30801 34298
rect 1952 34144 2004 34196
rect 18696 34187 18748 34196
rect 18696 34153 18705 34187
rect 18705 34153 18739 34187
rect 18739 34153 18748 34187
rect 18696 34144 18748 34153
rect 4436 34008 4488 34060
rect 6552 34008 6604 34060
rect 21548 34144 21600 34196
rect 21824 34144 21876 34196
rect 22008 34144 22060 34196
rect 20812 34076 20864 34128
rect 22376 34144 22428 34196
rect 22652 34076 22704 34128
rect 2504 33983 2556 33992
rect 2504 33949 2513 33983
rect 2513 33949 2547 33983
rect 2547 33949 2556 33983
rect 2504 33940 2556 33949
rect 18328 33940 18380 33992
rect 19800 33940 19852 33992
rect 3056 33915 3108 33924
rect 3056 33881 3065 33915
rect 3065 33881 3099 33915
rect 3099 33881 3108 33915
rect 3056 33872 3108 33881
rect 4896 33872 4948 33924
rect 18420 33804 18472 33856
rect 19800 33804 19852 33856
rect 20076 33804 20128 33856
rect 20352 33983 20404 33992
rect 20352 33949 20361 33983
rect 20361 33949 20395 33983
rect 20395 33949 20404 33983
rect 20352 33940 20404 33949
rect 23020 34008 23072 34060
rect 20996 33940 21048 33992
rect 21088 33872 21140 33924
rect 21272 33872 21324 33924
rect 22008 33872 22060 33924
rect 23112 33915 23164 33924
rect 23112 33881 23121 33915
rect 23121 33881 23155 33915
rect 23155 33881 23164 33915
rect 23112 33872 23164 33881
rect 24216 33940 24268 33992
rect 24584 33983 24636 33992
rect 24584 33949 24593 33983
rect 24593 33949 24627 33983
rect 24627 33949 24636 33983
rect 24584 33940 24636 33949
rect 24676 33940 24728 33992
rect 22928 33804 22980 33856
rect 23572 33872 23624 33924
rect 25044 33872 25096 33924
rect 23848 33847 23900 33856
rect 23848 33813 23857 33847
rect 23857 33813 23891 33847
rect 23891 33813 23900 33847
rect 23848 33804 23900 33813
rect 26608 34144 26660 34196
rect 27436 34144 27488 34196
rect 27620 34076 27672 34128
rect 30104 34144 30156 34196
rect 31116 34187 31168 34196
rect 31116 34153 31125 34187
rect 31125 34153 31159 34187
rect 31159 34153 31168 34187
rect 31116 34144 31168 34153
rect 29092 34076 29144 34128
rect 26424 34051 26476 34060
rect 26424 34017 26433 34051
rect 26433 34017 26467 34051
rect 26467 34017 26476 34051
rect 26424 34008 26476 34017
rect 29460 34008 29512 34060
rect 25964 33872 26016 33924
rect 28080 33940 28132 33992
rect 28540 33940 28592 33992
rect 27344 33872 27396 33924
rect 28264 33915 28316 33924
rect 27068 33804 27120 33856
rect 27436 33804 27488 33856
rect 28264 33881 28273 33915
rect 28273 33881 28307 33915
rect 28307 33881 28316 33915
rect 28264 33872 28316 33881
rect 29092 33872 29144 33924
rect 28540 33847 28592 33856
rect 28540 33813 28549 33847
rect 28549 33813 28583 33847
rect 28583 33813 28592 33847
rect 28540 33804 28592 33813
rect 28632 33847 28684 33856
rect 28632 33813 28641 33847
rect 28641 33813 28675 33847
rect 28675 33813 28684 33847
rect 28632 33804 28684 33813
rect 29184 33804 29236 33856
rect 29736 34076 29788 34128
rect 31576 34076 31628 34128
rect 29736 33983 29788 33992
rect 29736 33949 29745 33983
rect 29745 33949 29779 33983
rect 29779 33949 29788 33983
rect 29736 33940 29788 33949
rect 31300 34008 31352 34060
rect 31760 34008 31812 34060
rect 30932 33940 30984 33992
rect 31116 33940 31168 33992
rect 32036 34008 32088 34060
rect 30104 33872 30156 33924
rect 30840 33872 30892 33924
rect 32128 33872 32180 33924
rect 34336 33915 34388 33924
rect 34336 33881 34345 33915
rect 34345 33881 34379 33915
rect 34379 33881 34388 33915
rect 34336 33872 34388 33881
rect 30564 33804 30616 33856
rect 31944 33804 31996 33856
rect 9390 33702 9442 33754
rect 9454 33702 9506 33754
rect 9518 33702 9570 33754
rect 9582 33702 9634 33754
rect 9646 33702 9698 33754
rect 17831 33702 17883 33754
rect 17895 33702 17947 33754
rect 17959 33702 18011 33754
rect 18023 33702 18075 33754
rect 18087 33702 18139 33754
rect 26272 33702 26324 33754
rect 26336 33702 26388 33754
rect 26400 33702 26452 33754
rect 26464 33702 26516 33754
rect 26528 33702 26580 33754
rect 34713 33702 34765 33754
rect 34777 33702 34829 33754
rect 34841 33702 34893 33754
rect 34905 33702 34957 33754
rect 34969 33702 35021 33754
rect 2136 33643 2188 33652
rect 2136 33609 2145 33643
rect 2145 33609 2179 33643
rect 2179 33609 2188 33643
rect 2136 33600 2188 33609
rect 19064 33600 19116 33652
rect 19984 33600 20036 33652
rect 20352 33600 20404 33652
rect 21456 33600 21508 33652
rect 21732 33600 21784 33652
rect 31300 33643 31352 33652
rect 3240 33532 3292 33584
rect 16212 33532 16264 33584
rect 2320 33464 2372 33516
rect 2872 33507 2924 33516
rect 2872 33473 2881 33507
rect 2881 33473 2915 33507
rect 2915 33473 2924 33507
rect 2872 33464 2924 33473
rect 18236 33464 18288 33516
rect 18420 33507 18472 33516
rect 18420 33473 18454 33507
rect 18454 33473 18472 33507
rect 18420 33464 18472 33473
rect 18972 33464 19024 33516
rect 19524 33303 19576 33312
rect 19524 33269 19533 33303
rect 19533 33269 19567 33303
rect 19567 33269 19576 33303
rect 19524 33260 19576 33269
rect 20260 33464 20312 33516
rect 20444 33507 20496 33516
rect 20444 33473 20453 33507
rect 20453 33473 20487 33507
rect 20487 33473 20496 33507
rect 20444 33464 20496 33473
rect 20628 33507 20680 33516
rect 20628 33473 20637 33507
rect 20637 33473 20671 33507
rect 20671 33473 20680 33507
rect 21272 33507 21324 33516
rect 20628 33464 20680 33473
rect 21272 33473 21281 33507
rect 21281 33473 21315 33507
rect 21315 33473 21324 33507
rect 21272 33464 21324 33473
rect 21824 33464 21876 33516
rect 22468 33532 22520 33584
rect 24032 33507 24084 33516
rect 24032 33473 24041 33507
rect 24041 33473 24075 33507
rect 24075 33473 24084 33507
rect 24032 33464 24084 33473
rect 25688 33532 25740 33584
rect 25780 33532 25832 33584
rect 21640 33396 21692 33448
rect 24492 33439 24544 33448
rect 24492 33405 24501 33439
rect 24501 33405 24535 33439
rect 24535 33405 24544 33439
rect 24492 33396 24544 33405
rect 26700 33464 26752 33516
rect 27344 33507 27396 33516
rect 27344 33473 27353 33507
rect 27353 33473 27387 33507
rect 27387 33473 27396 33507
rect 27344 33464 27396 33473
rect 29736 33532 29788 33584
rect 31300 33609 31309 33643
rect 31309 33609 31343 33643
rect 31343 33609 31352 33643
rect 31300 33600 31352 33609
rect 30564 33532 30616 33584
rect 32128 33532 32180 33584
rect 32312 33532 32364 33584
rect 34428 33532 34480 33584
rect 29276 33464 29328 33516
rect 29460 33464 29512 33516
rect 27620 33396 27672 33448
rect 29920 33439 29972 33448
rect 29920 33405 29929 33439
rect 29929 33405 29963 33439
rect 29963 33405 29972 33439
rect 29920 33396 29972 33405
rect 23296 33260 23348 33312
rect 23480 33260 23532 33312
rect 26608 33260 26660 33312
rect 26700 33260 26752 33312
rect 29276 33328 29328 33380
rect 29184 33303 29236 33312
rect 29184 33269 29193 33303
rect 29193 33269 29227 33303
rect 29227 33269 29236 33303
rect 29184 33260 29236 33269
rect 29828 33260 29880 33312
rect 32680 33260 32732 33312
rect 5170 33158 5222 33210
rect 5234 33158 5286 33210
rect 5298 33158 5350 33210
rect 5362 33158 5414 33210
rect 5426 33158 5478 33210
rect 13611 33158 13663 33210
rect 13675 33158 13727 33210
rect 13739 33158 13791 33210
rect 13803 33158 13855 33210
rect 13867 33158 13919 33210
rect 22052 33158 22104 33210
rect 22116 33158 22168 33210
rect 22180 33158 22232 33210
rect 22244 33158 22296 33210
rect 22308 33158 22360 33210
rect 30493 33158 30545 33210
rect 30557 33158 30609 33210
rect 30621 33158 30673 33210
rect 30685 33158 30737 33210
rect 30749 33158 30801 33210
rect 1676 33056 1728 33108
rect 19708 33056 19760 33108
rect 20628 33056 20680 33108
rect 21916 33056 21968 33108
rect 24032 33056 24084 33108
rect 26148 33056 26200 33108
rect 13452 32988 13504 33040
rect 19432 32988 19484 33040
rect 18420 32920 18472 32972
rect 19248 32920 19300 32972
rect 2964 32852 3016 32904
rect 18880 32895 18932 32904
rect 18880 32861 18889 32895
rect 18889 32861 18923 32895
rect 18923 32861 18932 32895
rect 18880 32852 18932 32861
rect 19800 32895 19852 32904
rect 19800 32861 19834 32895
rect 19834 32861 19852 32895
rect 19800 32852 19852 32861
rect 28816 33056 28868 33108
rect 29276 33056 29328 33108
rect 32588 33056 32640 33108
rect 29828 32988 29880 33040
rect 29920 32988 29972 33040
rect 20628 32920 20680 32972
rect 21548 32895 21600 32904
rect 21548 32861 21557 32895
rect 21557 32861 21591 32895
rect 21591 32861 21600 32895
rect 22836 32895 22888 32904
rect 21548 32852 21600 32861
rect 22836 32861 22845 32895
rect 22845 32861 22879 32895
rect 22879 32861 22888 32895
rect 22836 32852 22888 32861
rect 16028 32716 16080 32768
rect 22376 32784 22428 32836
rect 22468 32784 22520 32836
rect 23388 32784 23440 32836
rect 23664 32827 23716 32836
rect 23664 32793 23673 32827
rect 23673 32793 23707 32827
rect 23707 32793 23716 32827
rect 23664 32784 23716 32793
rect 24124 32784 24176 32836
rect 20168 32716 20220 32768
rect 20628 32716 20680 32768
rect 20904 32759 20956 32768
rect 20904 32725 20913 32759
rect 20913 32725 20947 32759
rect 20947 32725 20956 32759
rect 20904 32716 20956 32725
rect 22836 32716 22888 32768
rect 23296 32716 23348 32768
rect 24952 32852 25004 32904
rect 26608 32852 26660 32904
rect 29184 32852 29236 32904
rect 29920 32895 29972 32904
rect 29920 32861 29929 32895
rect 29929 32861 29963 32895
rect 29963 32861 29972 32895
rect 29920 32852 29972 32861
rect 25412 32784 25464 32836
rect 25596 32784 25648 32836
rect 27436 32716 27488 32768
rect 28448 32784 28500 32836
rect 30748 32852 30800 32904
rect 31300 32852 31352 32904
rect 31576 32784 31628 32836
rect 33784 32784 33836 32836
rect 34244 32784 34296 32836
rect 29828 32716 29880 32768
rect 30932 32716 30984 32768
rect 31116 32716 31168 32768
rect 31484 32716 31536 32768
rect 34060 32759 34112 32768
rect 34060 32725 34069 32759
rect 34069 32725 34103 32759
rect 34103 32725 34112 32759
rect 34060 32716 34112 32725
rect 9390 32614 9442 32666
rect 9454 32614 9506 32666
rect 9518 32614 9570 32666
rect 9582 32614 9634 32666
rect 9646 32614 9698 32666
rect 17831 32614 17883 32666
rect 17895 32614 17947 32666
rect 17959 32614 18011 32666
rect 18023 32614 18075 32666
rect 18087 32614 18139 32666
rect 26272 32614 26324 32666
rect 26336 32614 26388 32666
rect 26400 32614 26452 32666
rect 26464 32614 26516 32666
rect 26528 32614 26580 32666
rect 34713 32614 34765 32666
rect 34777 32614 34829 32666
rect 34841 32614 34893 32666
rect 34905 32614 34957 32666
rect 34969 32614 35021 32666
rect 16304 32512 16356 32564
rect 17408 32444 17460 32496
rect 18880 32512 18932 32564
rect 20628 32512 20680 32564
rect 23020 32512 23072 32564
rect 23112 32512 23164 32564
rect 25596 32555 25648 32564
rect 21272 32444 21324 32496
rect 23848 32444 23900 32496
rect 18236 32376 18288 32428
rect 20444 32376 20496 32428
rect 21088 32419 21140 32428
rect 21088 32385 21097 32419
rect 21097 32385 21131 32419
rect 21131 32385 21140 32419
rect 21088 32376 21140 32385
rect 19616 32308 19668 32360
rect 20904 32308 20956 32360
rect 23940 32376 23992 32428
rect 24952 32444 25004 32496
rect 25228 32444 25280 32496
rect 25596 32521 25605 32555
rect 25605 32521 25639 32555
rect 25639 32521 25648 32555
rect 25596 32512 25648 32521
rect 26056 32512 26108 32564
rect 26148 32512 26200 32564
rect 26884 32444 26936 32496
rect 28632 32444 28684 32496
rect 27344 32419 27396 32428
rect 22468 32308 22520 32360
rect 22652 32351 22704 32360
rect 22652 32317 22661 32351
rect 22661 32317 22695 32351
rect 22695 32317 22704 32351
rect 22652 32308 22704 32317
rect 23848 32308 23900 32360
rect 25688 32308 25740 32360
rect 25780 32240 25832 32292
rect 25872 32240 25924 32292
rect 27344 32385 27353 32419
rect 27353 32385 27387 32419
rect 27387 32385 27396 32419
rect 27344 32376 27396 32385
rect 27528 32376 27580 32428
rect 28264 32376 28316 32428
rect 29460 32512 29512 32564
rect 30196 32512 30248 32564
rect 31576 32512 31628 32564
rect 31668 32512 31720 32564
rect 31760 32555 31812 32564
rect 31760 32521 31769 32555
rect 31769 32521 31803 32555
rect 31803 32521 31812 32555
rect 31760 32512 31812 32521
rect 29184 32444 29236 32496
rect 31300 32487 31352 32496
rect 31300 32453 31309 32487
rect 31309 32453 31343 32487
rect 31343 32453 31352 32487
rect 31300 32444 31352 32453
rect 31392 32444 31444 32496
rect 32680 32487 32732 32496
rect 26056 32240 26108 32292
rect 28540 32308 28592 32360
rect 27436 32240 27488 32292
rect 19064 32172 19116 32224
rect 19340 32172 19392 32224
rect 20720 32172 20772 32224
rect 21456 32172 21508 32224
rect 24032 32215 24084 32224
rect 24032 32181 24041 32215
rect 24041 32181 24075 32215
rect 24075 32181 24084 32215
rect 24032 32172 24084 32181
rect 24676 32172 24728 32224
rect 27988 32172 28040 32224
rect 28080 32172 28132 32224
rect 29828 32376 29880 32428
rect 31484 32419 31536 32428
rect 31484 32385 31493 32419
rect 31493 32385 31527 32419
rect 31527 32385 31536 32419
rect 31484 32376 31536 32385
rect 32680 32453 32689 32487
rect 32689 32453 32723 32487
rect 32723 32453 32732 32487
rect 32680 32444 32732 32453
rect 29460 32308 29512 32360
rect 30840 32308 30892 32360
rect 33416 32308 33468 32360
rect 34336 32351 34388 32360
rect 34336 32317 34345 32351
rect 34345 32317 34379 32351
rect 34379 32317 34388 32351
rect 34336 32308 34388 32317
rect 29736 32240 29788 32292
rect 32312 32240 32364 32292
rect 29460 32215 29512 32224
rect 29460 32181 29469 32215
rect 29469 32181 29503 32215
rect 29503 32181 29512 32215
rect 29460 32172 29512 32181
rect 31208 32172 31260 32224
rect 31392 32172 31444 32224
rect 5170 32070 5222 32122
rect 5234 32070 5286 32122
rect 5298 32070 5350 32122
rect 5362 32070 5414 32122
rect 5426 32070 5478 32122
rect 13611 32070 13663 32122
rect 13675 32070 13727 32122
rect 13739 32070 13791 32122
rect 13803 32070 13855 32122
rect 13867 32070 13919 32122
rect 22052 32070 22104 32122
rect 22116 32070 22168 32122
rect 22180 32070 22232 32122
rect 22244 32070 22296 32122
rect 22308 32070 22360 32122
rect 30493 32070 30545 32122
rect 30557 32070 30609 32122
rect 30621 32070 30673 32122
rect 30685 32070 30737 32122
rect 30749 32070 30801 32122
rect 17408 32011 17460 32020
rect 17408 31977 17417 32011
rect 17417 31977 17451 32011
rect 17451 31977 17460 32011
rect 17408 31968 17460 31977
rect 17592 31968 17644 32020
rect 21272 31968 21324 32020
rect 17684 31900 17736 31952
rect 1768 31764 1820 31816
rect 19064 31764 19116 31816
rect 19248 31900 19300 31952
rect 23112 32011 23164 32020
rect 23112 31977 23121 32011
rect 23121 31977 23155 32011
rect 23155 31977 23164 32011
rect 23112 31968 23164 31977
rect 23940 31968 23992 32020
rect 24492 31968 24544 32020
rect 25504 31968 25556 32020
rect 25780 31968 25832 32020
rect 26148 31968 26200 32020
rect 27620 31968 27672 32020
rect 29828 31968 29880 32020
rect 30104 32011 30156 32020
rect 19524 31832 19576 31884
rect 20352 31832 20404 31884
rect 19616 31764 19668 31816
rect 20444 31764 20496 31816
rect 22376 31764 22428 31816
rect 22652 31832 22704 31884
rect 23572 31832 23624 31884
rect 24216 31832 24268 31884
rect 24676 31875 24728 31884
rect 24676 31841 24685 31875
rect 24685 31841 24719 31875
rect 24719 31841 24728 31875
rect 25504 31875 25556 31884
rect 24676 31832 24728 31841
rect 25504 31841 25513 31875
rect 25513 31841 25547 31875
rect 25547 31841 25556 31875
rect 25504 31832 25556 31841
rect 22928 31764 22980 31816
rect 23848 31807 23900 31816
rect 23848 31773 23857 31807
rect 23857 31773 23891 31807
rect 23891 31773 23900 31807
rect 23848 31764 23900 31773
rect 18512 31696 18564 31748
rect 17500 31628 17552 31680
rect 20628 31696 20680 31748
rect 20812 31696 20864 31748
rect 19156 31628 19208 31680
rect 22468 31696 22520 31748
rect 23296 31696 23348 31748
rect 25688 31807 25740 31816
rect 25688 31773 25697 31807
rect 25697 31773 25731 31807
rect 25731 31773 25740 31807
rect 25688 31764 25740 31773
rect 24400 31696 24452 31748
rect 22192 31628 22244 31680
rect 22560 31628 22612 31680
rect 23388 31628 23440 31680
rect 23848 31628 23900 31680
rect 25044 31671 25096 31680
rect 25044 31637 25053 31671
rect 25053 31637 25087 31671
rect 25087 31637 25096 31671
rect 25044 31628 25096 31637
rect 26608 31807 26660 31816
rect 26608 31773 26617 31807
rect 26617 31773 26651 31807
rect 26651 31773 26660 31807
rect 26608 31764 26660 31773
rect 27160 31764 27212 31816
rect 27436 31696 27488 31748
rect 28172 31764 28224 31816
rect 28448 31764 28500 31816
rect 28264 31696 28316 31748
rect 28816 31696 28868 31748
rect 29368 31696 29420 31748
rect 30104 31977 30113 32011
rect 30113 31977 30147 32011
rect 30147 31977 30156 32011
rect 30104 31968 30156 31977
rect 30656 31968 30708 32020
rect 31760 31968 31812 32020
rect 31300 31900 31352 31952
rect 30656 31764 30708 31816
rect 31116 31832 31168 31884
rect 31576 31832 31628 31884
rect 31668 31807 31720 31816
rect 30932 31739 30984 31748
rect 30932 31705 30941 31739
rect 30941 31705 30975 31739
rect 30975 31705 30984 31739
rect 30932 31696 30984 31705
rect 31024 31739 31076 31748
rect 31208 31742 31260 31794
rect 31668 31773 31677 31807
rect 31677 31773 31711 31807
rect 31711 31773 31720 31807
rect 31668 31764 31720 31773
rect 32220 31832 32272 31884
rect 32312 31832 32364 31884
rect 32680 31807 32732 31816
rect 32680 31773 32714 31807
rect 32714 31773 32732 31807
rect 32680 31764 32732 31773
rect 31024 31705 31059 31739
rect 31059 31705 31076 31739
rect 31024 31696 31076 31705
rect 27620 31628 27672 31680
rect 27896 31628 27948 31680
rect 32404 31628 32456 31680
rect 9390 31526 9442 31578
rect 9454 31526 9506 31578
rect 9518 31526 9570 31578
rect 9582 31526 9634 31578
rect 9646 31526 9698 31578
rect 17831 31526 17883 31578
rect 17895 31526 17947 31578
rect 17959 31526 18011 31578
rect 18023 31526 18075 31578
rect 18087 31526 18139 31578
rect 26272 31526 26324 31578
rect 26336 31526 26388 31578
rect 26400 31526 26452 31578
rect 26464 31526 26516 31578
rect 26528 31526 26580 31578
rect 34713 31526 34765 31578
rect 34777 31526 34829 31578
rect 34841 31526 34893 31578
rect 34905 31526 34957 31578
rect 34969 31526 35021 31578
rect 20812 31424 20864 31476
rect 22100 31424 22152 31476
rect 22468 31424 22520 31476
rect 25136 31424 25188 31476
rect 1768 31331 1820 31340
rect 1768 31297 1777 31331
rect 1777 31297 1811 31331
rect 1811 31297 1820 31331
rect 1768 31288 1820 31297
rect 20720 31356 20772 31408
rect 21088 31399 21140 31408
rect 21088 31365 21097 31399
rect 21097 31365 21131 31399
rect 21131 31365 21140 31399
rect 21088 31356 21140 31365
rect 23480 31356 23532 31408
rect 24860 31399 24912 31408
rect 24860 31365 24894 31399
rect 24894 31365 24912 31399
rect 24860 31356 24912 31365
rect 27068 31356 27120 31408
rect 31208 31424 31260 31476
rect 31576 31467 31628 31476
rect 31576 31433 31585 31467
rect 31585 31433 31619 31467
rect 31619 31433 31628 31467
rect 31576 31424 31628 31433
rect 31760 31467 31812 31476
rect 31760 31433 31769 31467
rect 31769 31433 31803 31467
rect 31803 31433 31812 31467
rect 31760 31424 31812 31433
rect 17592 31288 17644 31340
rect 18604 31331 18656 31340
rect 18604 31297 18638 31331
rect 18638 31297 18656 31331
rect 18604 31288 18656 31297
rect 20536 31288 20588 31340
rect 2136 31220 2188 31272
rect 2780 31263 2832 31272
rect 2780 31229 2789 31263
rect 2789 31229 2823 31263
rect 2823 31229 2832 31263
rect 2780 31220 2832 31229
rect 18236 31220 18288 31272
rect 22652 31288 22704 31340
rect 24584 31263 24636 31272
rect 21364 31152 21416 31204
rect 18604 31084 18656 31136
rect 19248 31084 19300 31136
rect 19892 31084 19944 31136
rect 21916 31084 21968 31136
rect 24584 31229 24593 31263
rect 24593 31229 24627 31263
rect 24627 31229 24636 31263
rect 24584 31220 24636 31229
rect 26424 31331 26476 31340
rect 26424 31297 26433 31331
rect 26433 31297 26467 31331
rect 26467 31297 26476 31331
rect 26424 31288 26476 31297
rect 26976 31288 27028 31340
rect 27252 31288 27304 31340
rect 27804 31288 27856 31340
rect 28724 31288 28776 31340
rect 29828 31356 29880 31408
rect 31484 31399 31536 31408
rect 31484 31365 31493 31399
rect 31493 31365 31527 31399
rect 31527 31365 31536 31399
rect 31484 31356 31536 31365
rect 31852 31356 31904 31408
rect 27068 31220 27120 31272
rect 30748 31220 30800 31272
rect 23848 31152 23900 31204
rect 24400 31152 24452 31204
rect 23572 31084 23624 31136
rect 23756 31084 23808 31136
rect 24768 31084 24820 31136
rect 25872 31084 25924 31136
rect 26792 31084 26844 31136
rect 29368 31152 29420 31204
rect 31392 31331 31444 31340
rect 31392 31297 31401 31331
rect 31401 31297 31435 31331
rect 31435 31297 31444 31331
rect 32496 31331 32548 31340
rect 31392 31288 31444 31297
rect 32496 31297 32505 31331
rect 32505 31297 32539 31331
rect 32539 31297 32548 31331
rect 32496 31288 32548 31297
rect 34336 31331 34388 31340
rect 34336 31297 34345 31331
rect 34345 31297 34379 31331
rect 34379 31297 34388 31331
rect 34336 31288 34388 31297
rect 31484 31220 31536 31272
rect 33508 31220 33560 31272
rect 28724 31084 28776 31136
rect 30380 31084 30432 31136
rect 30932 31084 30984 31136
rect 33692 31152 33744 31204
rect 34060 31084 34112 31136
rect 5170 30982 5222 31034
rect 5234 30982 5286 31034
rect 5298 30982 5350 31034
rect 5362 30982 5414 31034
rect 5426 30982 5478 31034
rect 13611 30982 13663 31034
rect 13675 30982 13727 31034
rect 13739 30982 13791 31034
rect 13803 30982 13855 31034
rect 13867 30982 13919 31034
rect 22052 30982 22104 31034
rect 22116 30982 22168 31034
rect 22180 30982 22232 31034
rect 22244 30982 22296 31034
rect 22308 30982 22360 31034
rect 30493 30982 30545 31034
rect 30557 30982 30609 31034
rect 30621 30982 30673 31034
rect 30685 30982 30737 31034
rect 30749 30982 30801 31034
rect 2136 30923 2188 30932
rect 2136 30889 2145 30923
rect 2145 30889 2179 30923
rect 2179 30889 2188 30923
rect 2136 30880 2188 30889
rect 17776 30880 17828 30932
rect 19524 30923 19576 30932
rect 18420 30812 18472 30864
rect 19524 30889 19533 30923
rect 19533 30889 19567 30923
rect 19567 30889 19576 30923
rect 19524 30880 19576 30889
rect 21088 30880 21140 30932
rect 19340 30812 19392 30864
rect 19984 30812 20036 30864
rect 2136 30676 2188 30728
rect 18512 30744 18564 30796
rect 19248 30744 19300 30796
rect 20352 30787 20404 30796
rect 20352 30753 20361 30787
rect 20361 30753 20395 30787
rect 20395 30753 20404 30787
rect 20352 30744 20404 30753
rect 17776 30719 17828 30728
rect 17776 30685 17785 30719
rect 17785 30685 17819 30719
rect 17819 30685 17828 30719
rect 17776 30676 17828 30685
rect 19064 30676 19116 30728
rect 19432 30719 19484 30728
rect 19432 30685 19441 30719
rect 19441 30685 19475 30719
rect 19475 30685 19484 30719
rect 19432 30676 19484 30685
rect 21456 30676 21508 30728
rect 21916 30880 21968 30932
rect 22652 30880 22704 30932
rect 25136 30880 25188 30932
rect 28908 30880 28960 30932
rect 29368 30880 29420 30932
rect 29644 30880 29696 30932
rect 31484 30880 31536 30932
rect 23296 30812 23348 30864
rect 29184 30812 29236 30864
rect 22560 30744 22612 30796
rect 18512 30651 18564 30660
rect 18512 30617 18521 30651
rect 18521 30617 18555 30651
rect 18555 30617 18564 30651
rect 18512 30608 18564 30617
rect 19892 30608 19944 30660
rect 21364 30608 21416 30660
rect 22928 30676 22980 30728
rect 24492 30744 24544 30796
rect 26424 30744 26476 30796
rect 27160 30744 27212 30796
rect 24032 30676 24084 30728
rect 24676 30719 24728 30728
rect 24676 30685 24685 30719
rect 24685 30685 24719 30719
rect 24719 30685 24728 30719
rect 24676 30676 24728 30685
rect 29092 30744 29144 30796
rect 32312 30880 32364 30932
rect 32956 30880 33008 30932
rect 33416 30923 33468 30932
rect 33416 30889 33425 30923
rect 33425 30889 33459 30923
rect 33459 30889 33468 30923
rect 33416 30880 33468 30889
rect 30748 30744 30800 30796
rect 31760 30744 31812 30796
rect 32036 30787 32088 30796
rect 32036 30753 32045 30787
rect 32045 30753 32079 30787
rect 32079 30753 32088 30787
rect 32036 30744 32088 30753
rect 23848 30651 23900 30660
rect 23848 30617 23857 30651
rect 23857 30617 23891 30651
rect 23891 30617 23900 30651
rect 23848 30608 23900 30617
rect 23940 30608 23992 30660
rect 18972 30540 19024 30592
rect 19800 30583 19852 30592
rect 19800 30549 19809 30583
rect 19809 30549 19843 30583
rect 19843 30549 19852 30583
rect 19800 30540 19852 30549
rect 20168 30540 20220 30592
rect 23020 30540 23072 30592
rect 28448 30719 28500 30728
rect 28448 30685 28457 30719
rect 28457 30685 28491 30719
rect 28491 30685 28500 30719
rect 28448 30676 28500 30685
rect 28816 30676 28868 30728
rect 28172 30608 28224 30660
rect 28264 30651 28316 30660
rect 28264 30617 28273 30651
rect 28273 30617 28307 30651
rect 28307 30617 28316 30651
rect 28264 30608 28316 30617
rect 28540 30608 28592 30660
rect 30932 30719 30984 30728
rect 30932 30685 30941 30719
rect 30941 30685 30975 30719
rect 30975 30685 30984 30719
rect 30932 30676 30984 30685
rect 31300 30676 31352 30728
rect 33416 30676 33468 30728
rect 34060 30719 34112 30728
rect 34060 30685 34069 30719
rect 34069 30685 34103 30719
rect 34103 30685 34112 30719
rect 34060 30676 34112 30685
rect 27344 30583 27396 30592
rect 27344 30549 27353 30583
rect 27353 30549 27387 30583
rect 27387 30549 27396 30583
rect 27344 30540 27396 30549
rect 28080 30540 28132 30592
rect 28724 30540 28776 30592
rect 30748 30540 30800 30592
rect 31024 30608 31076 30660
rect 32128 30540 32180 30592
rect 34244 30583 34296 30592
rect 34244 30549 34253 30583
rect 34253 30549 34287 30583
rect 34287 30549 34296 30583
rect 34244 30540 34296 30549
rect 9390 30438 9442 30490
rect 9454 30438 9506 30490
rect 9518 30438 9570 30490
rect 9582 30438 9634 30490
rect 9646 30438 9698 30490
rect 17831 30438 17883 30490
rect 17895 30438 17947 30490
rect 17959 30438 18011 30490
rect 18023 30438 18075 30490
rect 18087 30438 18139 30490
rect 26272 30438 26324 30490
rect 26336 30438 26388 30490
rect 26400 30438 26452 30490
rect 26464 30438 26516 30490
rect 26528 30438 26580 30490
rect 34713 30438 34765 30490
rect 34777 30438 34829 30490
rect 34841 30438 34893 30490
rect 34905 30438 34957 30490
rect 34969 30438 35021 30490
rect 21364 30379 21416 30388
rect 18972 30268 19024 30320
rect 21364 30345 21373 30379
rect 21373 30345 21407 30379
rect 21407 30345 21416 30379
rect 21364 30336 21416 30345
rect 19616 30268 19668 30320
rect 22652 30336 22704 30388
rect 23296 30336 23348 30388
rect 24860 30336 24912 30388
rect 18144 30243 18196 30252
rect 18144 30209 18153 30243
rect 18153 30209 18187 30243
rect 18187 30209 18196 30243
rect 18144 30200 18196 30209
rect 21916 30268 21968 30320
rect 22468 30268 22520 30320
rect 19248 30132 19300 30184
rect 22836 30200 22888 30252
rect 23848 30175 23900 30184
rect 19156 30064 19208 30116
rect 17500 29996 17552 30048
rect 18512 29996 18564 30048
rect 18788 29996 18840 30048
rect 19248 29996 19300 30048
rect 19524 30039 19576 30048
rect 19524 30005 19533 30039
rect 19533 30005 19567 30039
rect 19567 30005 19576 30039
rect 19524 29996 19576 30005
rect 23848 30141 23857 30175
rect 23857 30141 23891 30175
rect 23891 30141 23900 30175
rect 23848 30132 23900 30141
rect 24584 30200 24636 30252
rect 24860 30200 24912 30252
rect 25320 30268 25372 30320
rect 25596 30336 25648 30388
rect 25688 30268 25740 30320
rect 27988 30336 28040 30388
rect 30380 30336 30432 30388
rect 30472 30336 30524 30388
rect 31668 30336 31720 30388
rect 26056 30268 26108 30320
rect 28356 30268 28408 30320
rect 30012 30200 30064 30252
rect 31576 30268 31628 30320
rect 33232 30311 33284 30320
rect 33232 30277 33266 30311
rect 33266 30277 33284 30311
rect 33232 30268 33284 30277
rect 26056 30132 26108 30184
rect 27344 30132 27396 30184
rect 28540 30132 28592 30184
rect 29920 30132 29972 30184
rect 30472 30132 30524 30184
rect 30932 30175 30984 30184
rect 30932 30141 30941 30175
rect 30941 30141 30975 30175
rect 30975 30141 30984 30175
rect 30932 30132 30984 30141
rect 31668 30200 31720 30252
rect 32496 30243 32548 30252
rect 32496 30209 32505 30243
rect 32505 30209 32539 30243
rect 32539 30209 32548 30243
rect 32496 30200 32548 30209
rect 32956 30243 33008 30252
rect 32956 30209 32965 30243
rect 32965 30209 32999 30243
rect 32999 30209 33008 30243
rect 32956 30200 33008 30209
rect 33048 30200 33100 30252
rect 25780 30064 25832 30116
rect 28632 30064 28684 30116
rect 31392 30064 31444 30116
rect 22744 29996 22796 30048
rect 23020 29996 23072 30048
rect 27712 29996 27764 30048
rect 28448 29996 28500 30048
rect 29092 29996 29144 30048
rect 31484 29996 31536 30048
rect 5170 29894 5222 29946
rect 5234 29894 5286 29946
rect 5298 29894 5350 29946
rect 5362 29894 5414 29946
rect 5426 29894 5478 29946
rect 13611 29894 13663 29946
rect 13675 29894 13727 29946
rect 13739 29894 13791 29946
rect 13803 29894 13855 29946
rect 13867 29894 13919 29946
rect 22052 29894 22104 29946
rect 22116 29894 22168 29946
rect 22180 29894 22232 29946
rect 22244 29894 22296 29946
rect 22308 29894 22360 29946
rect 30493 29894 30545 29946
rect 30557 29894 30609 29946
rect 30621 29894 30673 29946
rect 30685 29894 30737 29946
rect 30749 29894 30801 29946
rect 16212 29835 16264 29844
rect 16212 29801 16221 29835
rect 16221 29801 16255 29835
rect 16255 29801 16264 29835
rect 16212 29792 16264 29801
rect 22928 29792 22980 29844
rect 26148 29792 26200 29844
rect 28632 29792 28684 29844
rect 29276 29792 29328 29844
rect 29552 29792 29604 29844
rect 17500 29767 17552 29776
rect 17500 29733 17509 29767
rect 17509 29733 17543 29767
rect 17543 29733 17552 29767
rect 17500 29724 17552 29733
rect 16856 29631 16908 29640
rect 16856 29597 16865 29631
rect 16865 29597 16899 29631
rect 16899 29597 16908 29631
rect 16856 29588 16908 29597
rect 19616 29724 19668 29776
rect 19800 29724 19852 29776
rect 20168 29767 20220 29776
rect 20168 29733 20177 29767
rect 20177 29733 20211 29767
rect 20211 29733 20220 29767
rect 20168 29724 20220 29733
rect 21824 29724 21876 29776
rect 25964 29767 26016 29776
rect 25964 29733 25973 29767
rect 25973 29733 26007 29767
rect 26007 29733 26016 29767
rect 25964 29724 26016 29733
rect 27712 29767 27764 29776
rect 27712 29733 27721 29767
rect 27721 29733 27755 29767
rect 27755 29733 27764 29767
rect 27712 29724 27764 29733
rect 17868 29588 17920 29640
rect 18420 29631 18472 29640
rect 18420 29597 18429 29631
rect 18429 29597 18463 29631
rect 18463 29597 18472 29631
rect 18420 29588 18472 29597
rect 18696 29656 18748 29708
rect 19524 29656 19576 29708
rect 17592 29520 17644 29572
rect 18696 29563 18748 29572
rect 18696 29529 18731 29563
rect 18731 29529 18748 29563
rect 18696 29520 18748 29529
rect 16672 29495 16724 29504
rect 16672 29461 16681 29495
rect 16681 29461 16715 29495
rect 16715 29461 16724 29495
rect 16672 29452 16724 29461
rect 18604 29452 18656 29504
rect 18972 29588 19024 29640
rect 19984 29631 20036 29640
rect 19984 29597 19993 29631
rect 19993 29597 20027 29631
rect 20027 29597 20036 29631
rect 23388 29656 23440 29708
rect 19984 29588 20036 29597
rect 19248 29520 19300 29572
rect 22284 29520 22336 29572
rect 22652 29631 22704 29640
rect 22652 29597 22661 29631
rect 22661 29597 22695 29631
rect 22695 29597 22704 29631
rect 22652 29588 22704 29597
rect 22836 29631 22888 29640
rect 22836 29597 22845 29631
rect 22845 29597 22879 29631
rect 22879 29597 22888 29631
rect 23572 29631 23624 29640
rect 22836 29588 22888 29597
rect 23572 29597 23581 29631
rect 23581 29597 23615 29631
rect 23615 29597 23624 29631
rect 23572 29588 23624 29597
rect 24860 29656 24912 29708
rect 25044 29656 25096 29708
rect 27436 29656 27488 29708
rect 27988 29656 28040 29708
rect 28724 29656 28776 29708
rect 24768 29631 24820 29640
rect 24768 29597 24777 29631
rect 24777 29597 24811 29631
rect 24811 29597 24820 29631
rect 24768 29588 24820 29597
rect 24952 29631 25004 29640
rect 24952 29597 24961 29631
rect 24961 29597 24995 29631
rect 24995 29597 25004 29631
rect 24952 29588 25004 29597
rect 25596 29588 25648 29640
rect 25872 29631 25924 29640
rect 25872 29597 25881 29631
rect 25881 29597 25915 29631
rect 25915 29597 25924 29631
rect 25872 29588 25924 29597
rect 25964 29588 26016 29640
rect 27344 29631 27396 29640
rect 27344 29597 27353 29631
rect 27353 29597 27387 29631
rect 27387 29597 27396 29631
rect 27344 29588 27396 29597
rect 22744 29520 22796 29572
rect 23204 29520 23256 29572
rect 19340 29452 19392 29504
rect 20260 29452 20312 29504
rect 23848 29452 23900 29504
rect 26884 29520 26936 29572
rect 28540 29588 28592 29640
rect 29092 29631 29144 29640
rect 29092 29597 29101 29631
rect 29101 29597 29135 29631
rect 29135 29597 29144 29631
rect 29092 29588 29144 29597
rect 29184 29631 29236 29640
rect 29184 29597 29193 29631
rect 29193 29597 29227 29631
rect 29227 29597 29236 29631
rect 29184 29588 29236 29597
rect 29644 29588 29696 29640
rect 34244 29792 34296 29844
rect 33232 29767 33284 29776
rect 33232 29733 33241 29767
rect 33241 29733 33275 29767
rect 33275 29733 33284 29767
rect 33232 29724 33284 29733
rect 30104 29656 30156 29708
rect 32404 29656 32456 29708
rect 32588 29656 32640 29708
rect 34244 29656 34296 29708
rect 28816 29520 28868 29572
rect 25320 29452 25372 29504
rect 25412 29452 25464 29504
rect 25964 29452 26016 29504
rect 27896 29452 27948 29504
rect 28264 29452 28316 29504
rect 28724 29452 28776 29504
rect 30380 29588 30432 29640
rect 30196 29520 30248 29572
rect 32036 29588 32088 29640
rect 30748 29495 30800 29504
rect 30748 29461 30757 29495
rect 30757 29461 30791 29495
rect 30791 29461 30800 29495
rect 30748 29452 30800 29461
rect 31116 29452 31168 29504
rect 32036 29452 32088 29504
rect 33324 29588 33376 29640
rect 33600 29631 33652 29640
rect 33600 29597 33609 29631
rect 33609 29597 33643 29631
rect 33643 29597 33652 29631
rect 33600 29588 33652 29597
rect 33784 29588 33836 29640
rect 34060 29588 34112 29640
rect 34336 29631 34388 29640
rect 34336 29597 34345 29631
rect 34345 29597 34379 29631
rect 34379 29597 34388 29631
rect 34336 29588 34388 29597
rect 32220 29520 32272 29572
rect 32772 29495 32824 29504
rect 32772 29461 32781 29495
rect 32781 29461 32815 29495
rect 32815 29461 32824 29495
rect 32772 29452 32824 29461
rect 33784 29452 33836 29504
rect 9390 29350 9442 29402
rect 9454 29350 9506 29402
rect 9518 29350 9570 29402
rect 9582 29350 9634 29402
rect 9646 29350 9698 29402
rect 17831 29350 17883 29402
rect 17895 29350 17947 29402
rect 17959 29350 18011 29402
rect 18023 29350 18075 29402
rect 18087 29350 18139 29402
rect 26272 29350 26324 29402
rect 26336 29350 26388 29402
rect 26400 29350 26452 29402
rect 26464 29350 26516 29402
rect 26528 29350 26580 29402
rect 34713 29350 34765 29402
rect 34777 29350 34829 29402
rect 34841 29350 34893 29402
rect 34905 29350 34957 29402
rect 34969 29350 35021 29402
rect 16672 29248 16724 29300
rect 20536 29291 20588 29300
rect 18420 29180 18472 29232
rect 20536 29257 20545 29291
rect 20545 29257 20579 29291
rect 20579 29257 20588 29291
rect 20536 29248 20588 29257
rect 20628 29248 20680 29300
rect 21272 29248 21324 29300
rect 20076 29180 20128 29232
rect 17592 29155 17644 29164
rect 17592 29121 17626 29155
rect 17626 29121 17644 29155
rect 17592 29112 17644 29121
rect 18144 29112 18196 29164
rect 19156 29155 19208 29164
rect 19156 29121 19165 29155
rect 19165 29121 19199 29155
rect 19199 29121 19208 29155
rect 19156 29112 19208 29121
rect 19248 29112 19300 29164
rect 20444 29180 20496 29232
rect 21180 29180 21232 29232
rect 18972 29044 19024 29096
rect 22008 29112 22060 29164
rect 23572 29248 23624 29300
rect 24676 29248 24728 29300
rect 27436 29248 27488 29300
rect 27712 29248 27764 29300
rect 30748 29248 30800 29300
rect 31116 29291 31168 29300
rect 31116 29257 31125 29291
rect 31125 29257 31159 29291
rect 31159 29257 31168 29291
rect 31116 29248 31168 29257
rect 31300 29248 31352 29300
rect 31576 29248 31628 29300
rect 24124 29180 24176 29232
rect 26424 29180 26476 29232
rect 22560 29112 22612 29164
rect 22836 29112 22888 29164
rect 23480 29155 23532 29164
rect 23480 29121 23514 29155
rect 23514 29121 23532 29155
rect 23480 29112 23532 29121
rect 23020 29044 23072 29096
rect 23204 29087 23256 29096
rect 23204 29053 23213 29087
rect 23213 29053 23247 29087
rect 23247 29053 23256 29087
rect 23204 29044 23256 29053
rect 26884 29112 26936 29164
rect 27252 29112 27304 29164
rect 27804 29155 27856 29164
rect 27804 29121 27813 29155
rect 27813 29121 27847 29155
rect 27847 29121 27856 29155
rect 27804 29112 27856 29121
rect 27896 29112 27948 29164
rect 28172 29180 28224 29232
rect 28816 29112 28868 29164
rect 29092 29112 29144 29164
rect 30840 29112 30892 29164
rect 31116 29112 31168 29164
rect 31481 29158 31533 29167
rect 31481 29124 31490 29158
rect 31490 29124 31524 29158
rect 31524 29124 31533 29158
rect 31481 29115 31533 29124
rect 33140 29248 33192 29300
rect 33968 29248 34020 29300
rect 31852 29180 31904 29232
rect 18972 28908 19024 28960
rect 21824 28976 21876 29028
rect 30104 29044 30156 29096
rect 26424 29019 26476 29028
rect 26424 28985 26433 29019
rect 26433 28985 26467 29019
rect 26467 28985 26476 29019
rect 26424 28976 26476 28985
rect 27896 28976 27948 29028
rect 27988 28976 28040 29028
rect 29552 28976 29604 29028
rect 30288 28976 30340 29028
rect 31668 28976 31720 29028
rect 31944 29112 31996 29164
rect 32128 29112 32180 29164
rect 32404 29112 32456 29164
rect 33048 29112 33100 29164
rect 33324 29112 33376 29164
rect 33784 29155 33836 29164
rect 33784 29121 33793 29155
rect 33793 29121 33827 29155
rect 33827 29121 33836 29155
rect 33784 29112 33836 29121
rect 32404 28976 32456 29028
rect 33232 28976 33284 29028
rect 21272 28908 21324 28960
rect 23388 28908 23440 28960
rect 23480 28908 23532 28960
rect 28080 28908 28132 28960
rect 28448 28908 28500 28960
rect 29184 28908 29236 28960
rect 29736 28908 29788 28960
rect 30196 28908 30248 28960
rect 31576 28908 31628 28960
rect 34336 28976 34388 29028
rect 5170 28806 5222 28858
rect 5234 28806 5286 28858
rect 5298 28806 5350 28858
rect 5362 28806 5414 28858
rect 5426 28806 5478 28858
rect 13611 28806 13663 28858
rect 13675 28806 13727 28858
rect 13739 28806 13791 28858
rect 13803 28806 13855 28858
rect 13867 28806 13919 28858
rect 22052 28806 22104 28858
rect 22116 28806 22168 28858
rect 22180 28806 22232 28858
rect 22244 28806 22296 28858
rect 22308 28806 22360 28858
rect 30493 28806 30545 28858
rect 30557 28806 30609 28858
rect 30621 28806 30673 28858
rect 30685 28806 30737 28858
rect 30749 28806 30801 28858
rect 21272 28704 21324 28756
rect 22376 28704 22428 28756
rect 25964 28747 26016 28756
rect 25964 28713 25973 28747
rect 25973 28713 26007 28747
rect 26007 28713 26016 28747
rect 25964 28704 26016 28713
rect 27344 28704 27396 28756
rect 27804 28747 27856 28756
rect 27804 28713 27813 28747
rect 27813 28713 27847 28747
rect 27847 28713 27856 28747
rect 27804 28704 27856 28713
rect 29000 28704 29052 28756
rect 31944 28704 31996 28756
rect 32128 28704 32180 28756
rect 32864 28704 32916 28756
rect 33876 28747 33928 28756
rect 33876 28713 33885 28747
rect 33885 28713 33919 28747
rect 33919 28713 33928 28747
rect 33876 28704 33928 28713
rect 18788 28636 18840 28688
rect 22744 28636 22796 28688
rect 16304 28543 16356 28552
rect 16304 28509 16313 28543
rect 16313 28509 16347 28543
rect 16347 28509 16356 28543
rect 16304 28500 16356 28509
rect 19248 28568 19300 28620
rect 17592 28543 17644 28552
rect 17592 28509 17601 28543
rect 17601 28509 17635 28543
rect 17635 28509 17644 28543
rect 17592 28500 17644 28509
rect 18144 28543 18196 28552
rect 18144 28509 18153 28543
rect 18153 28509 18187 28543
rect 18187 28509 18196 28543
rect 18144 28500 18196 28509
rect 17132 28432 17184 28484
rect 18972 28500 19024 28552
rect 23204 28568 23256 28620
rect 29000 28611 29052 28620
rect 29000 28577 29009 28611
rect 29009 28577 29043 28611
rect 29043 28577 29052 28611
rect 31116 28636 31168 28688
rect 33324 28636 33376 28688
rect 29000 28568 29052 28577
rect 31852 28568 31904 28620
rect 19524 28543 19576 28552
rect 19524 28509 19533 28543
rect 19533 28509 19567 28543
rect 19567 28509 19576 28543
rect 19524 28500 19576 28509
rect 24032 28543 24084 28552
rect 16764 28407 16816 28416
rect 16764 28373 16773 28407
rect 16773 28373 16807 28407
rect 16807 28373 16816 28407
rect 16764 28364 16816 28373
rect 18604 28364 18656 28416
rect 19064 28364 19116 28416
rect 24032 28509 24041 28543
rect 24041 28509 24075 28543
rect 24075 28509 24084 28543
rect 24032 28500 24084 28509
rect 24584 28543 24636 28552
rect 24584 28509 24593 28543
rect 24593 28509 24627 28543
rect 24627 28509 24636 28543
rect 24584 28500 24636 28509
rect 24860 28543 24912 28552
rect 24860 28509 24894 28543
rect 24894 28509 24912 28543
rect 24860 28500 24912 28509
rect 26056 28500 26108 28552
rect 26700 28543 26752 28552
rect 26700 28509 26734 28543
rect 26734 28509 26752 28543
rect 26700 28500 26752 28509
rect 29092 28543 29144 28552
rect 20812 28475 20864 28484
rect 20812 28441 20821 28475
rect 20821 28441 20855 28475
rect 20855 28441 20864 28475
rect 20812 28432 20864 28441
rect 22100 28432 22152 28484
rect 22560 28432 22612 28484
rect 23112 28432 23164 28484
rect 24400 28432 24452 28484
rect 29092 28509 29101 28543
rect 29101 28509 29135 28543
rect 29135 28509 29144 28543
rect 29092 28500 29144 28509
rect 29736 28543 29788 28552
rect 29736 28509 29745 28543
rect 29745 28509 29779 28543
rect 29779 28509 29788 28543
rect 29736 28500 29788 28509
rect 29828 28500 29880 28552
rect 30288 28500 30340 28552
rect 29184 28432 29236 28484
rect 29644 28432 29696 28484
rect 30012 28475 30064 28484
rect 30012 28441 30046 28475
rect 30046 28441 30064 28475
rect 30012 28432 30064 28441
rect 31484 28432 31536 28484
rect 32864 28500 32916 28552
rect 21180 28364 21232 28416
rect 22928 28364 22980 28416
rect 23480 28364 23532 28416
rect 24492 28364 24544 28416
rect 27252 28364 27304 28416
rect 28448 28364 28500 28416
rect 29552 28364 29604 28416
rect 29828 28364 29880 28416
rect 30104 28364 30156 28416
rect 30840 28364 30892 28416
rect 32128 28364 32180 28416
rect 33784 28432 33836 28484
rect 33600 28364 33652 28416
rect 9390 28262 9442 28314
rect 9454 28262 9506 28314
rect 9518 28262 9570 28314
rect 9582 28262 9634 28314
rect 9646 28262 9698 28314
rect 17831 28262 17883 28314
rect 17895 28262 17947 28314
rect 17959 28262 18011 28314
rect 18023 28262 18075 28314
rect 18087 28262 18139 28314
rect 26272 28262 26324 28314
rect 26336 28262 26388 28314
rect 26400 28262 26452 28314
rect 26464 28262 26516 28314
rect 26528 28262 26580 28314
rect 34713 28262 34765 28314
rect 34777 28262 34829 28314
rect 34841 28262 34893 28314
rect 34905 28262 34957 28314
rect 34969 28262 35021 28314
rect 16764 28160 16816 28212
rect 20168 28160 20220 28212
rect 17684 28092 17736 28144
rect 18420 28092 18472 28144
rect 16120 28067 16172 28076
rect 16120 28033 16129 28067
rect 16129 28033 16163 28067
rect 16163 28033 16172 28067
rect 16120 28024 16172 28033
rect 17040 28024 17092 28076
rect 17132 28067 17184 28076
rect 17132 28033 17141 28067
rect 17141 28033 17175 28067
rect 17175 28033 17184 28067
rect 19156 28092 19208 28144
rect 20628 28160 20680 28212
rect 20444 28135 20496 28144
rect 17132 28024 17184 28033
rect 19064 28024 19116 28076
rect 20444 28101 20453 28135
rect 20453 28101 20487 28135
rect 20487 28101 20496 28135
rect 20444 28092 20496 28101
rect 23296 28160 23348 28212
rect 23572 28160 23624 28212
rect 22008 28024 22060 28076
rect 22468 28092 22520 28144
rect 23204 28092 23256 28144
rect 24124 28067 24176 28076
rect 24124 28033 24133 28067
rect 24133 28033 24167 28067
rect 24167 28033 24176 28067
rect 24124 28024 24176 28033
rect 26056 28160 26108 28212
rect 27068 28160 27120 28212
rect 30932 28160 30984 28212
rect 31668 28160 31720 28212
rect 34060 28160 34112 28212
rect 25044 28092 25096 28144
rect 28816 28092 28868 28144
rect 16304 27820 16356 27872
rect 17408 27820 17460 27872
rect 18236 27888 18288 27940
rect 20168 27888 20220 27940
rect 23388 27956 23440 28008
rect 26148 28024 26200 28076
rect 27528 28024 27580 28076
rect 27160 27999 27212 28008
rect 27160 27965 27169 27999
rect 27169 27965 27203 27999
rect 27203 27965 27212 27999
rect 27160 27956 27212 27965
rect 28356 27999 28408 28008
rect 28356 27965 28365 27999
rect 28365 27965 28399 27999
rect 28399 27965 28408 27999
rect 28356 27956 28408 27965
rect 18420 27820 18472 27872
rect 18512 27820 18564 27872
rect 22376 27820 22428 27872
rect 22836 27820 22888 27872
rect 24492 27888 24544 27940
rect 25596 27888 25648 27940
rect 23572 27820 23624 27872
rect 24952 27820 25004 27872
rect 26884 27888 26936 27940
rect 28080 27820 28132 27872
rect 29000 28024 29052 28076
rect 29644 28092 29696 28144
rect 30012 28135 30064 28144
rect 30012 28101 30021 28135
rect 30021 28101 30055 28135
rect 30055 28101 30064 28135
rect 30012 28092 30064 28101
rect 29092 27956 29144 28008
rect 29828 28067 29880 28076
rect 31024 28092 31076 28144
rect 29828 28033 29848 28067
rect 29848 28033 29880 28067
rect 29828 28024 29880 28033
rect 29644 27999 29696 28008
rect 29644 27965 29653 27999
rect 29653 27965 29687 27999
rect 29687 27965 29696 27999
rect 31116 28024 31168 28076
rect 32680 28135 32732 28144
rect 32680 28101 32689 28135
rect 32689 28101 32723 28135
rect 32723 28101 32732 28135
rect 32680 28092 32732 28101
rect 32496 28067 32548 28076
rect 32496 28033 32505 28067
rect 32505 28033 32539 28067
rect 32539 28033 32548 28067
rect 32496 28024 32548 28033
rect 29644 27956 29696 27965
rect 30932 27956 30984 28008
rect 31576 27999 31628 28008
rect 31576 27965 31585 27999
rect 31585 27965 31619 27999
rect 31619 27965 31628 27999
rect 31576 27956 31628 27965
rect 32404 27956 32456 28008
rect 34336 27999 34388 28008
rect 34336 27965 34345 27999
rect 34345 27965 34379 27999
rect 34379 27965 34388 27999
rect 34336 27956 34388 27965
rect 32864 27888 32916 27940
rect 29368 27820 29420 27872
rect 29552 27820 29604 27872
rect 30380 27820 30432 27872
rect 31300 27820 31352 27872
rect 31852 27820 31904 27872
rect 32404 27820 32456 27872
rect 5170 27718 5222 27770
rect 5234 27718 5286 27770
rect 5298 27718 5350 27770
rect 5362 27718 5414 27770
rect 5426 27718 5478 27770
rect 13611 27718 13663 27770
rect 13675 27718 13727 27770
rect 13739 27718 13791 27770
rect 13803 27718 13855 27770
rect 13867 27718 13919 27770
rect 22052 27718 22104 27770
rect 22116 27718 22168 27770
rect 22180 27718 22232 27770
rect 22244 27718 22296 27770
rect 22308 27718 22360 27770
rect 30493 27718 30545 27770
rect 30557 27718 30609 27770
rect 30621 27718 30673 27770
rect 30685 27718 30737 27770
rect 30749 27718 30801 27770
rect 17040 27616 17092 27668
rect 22836 27616 22888 27668
rect 22928 27616 22980 27668
rect 25872 27616 25924 27668
rect 27528 27616 27580 27668
rect 17592 27548 17644 27600
rect 7656 27480 7708 27532
rect 6644 27387 6696 27396
rect 6644 27353 6653 27387
rect 6653 27353 6687 27387
rect 6687 27353 6696 27387
rect 6644 27344 6696 27353
rect 3516 27276 3568 27328
rect 17040 27480 17092 27532
rect 18512 27548 18564 27600
rect 22652 27548 22704 27600
rect 25504 27548 25556 27600
rect 17868 27523 17920 27532
rect 17868 27489 17902 27523
rect 17902 27489 17920 27523
rect 17868 27480 17920 27489
rect 19064 27480 19116 27532
rect 16028 27455 16080 27464
rect 16028 27421 16037 27455
rect 16037 27421 16071 27455
rect 16071 27421 16080 27455
rect 16028 27412 16080 27421
rect 17408 27455 17460 27464
rect 17408 27421 17417 27455
rect 17417 27421 17451 27455
rect 17451 27421 17460 27455
rect 17408 27412 17460 27421
rect 18328 27412 18380 27464
rect 18604 27455 18656 27464
rect 18604 27421 18613 27455
rect 18613 27421 18647 27455
rect 18647 27421 18656 27455
rect 18604 27412 18656 27421
rect 19156 27412 19208 27464
rect 19432 27455 19484 27464
rect 19432 27421 19441 27455
rect 19441 27421 19475 27455
rect 19475 27421 19484 27455
rect 19432 27412 19484 27421
rect 22468 27412 22520 27464
rect 17408 27276 17460 27328
rect 18236 27276 18288 27328
rect 19340 27276 19392 27328
rect 19524 27344 19576 27396
rect 21916 27344 21968 27396
rect 20444 27276 20496 27328
rect 22836 27276 22888 27328
rect 23848 27480 23900 27532
rect 24124 27480 24176 27532
rect 26056 27480 26108 27532
rect 29460 27548 29512 27600
rect 30012 27616 30064 27668
rect 34244 27616 34296 27668
rect 29736 27548 29788 27600
rect 29092 27480 29144 27532
rect 29920 27523 29972 27532
rect 23296 27412 23348 27464
rect 24676 27455 24728 27464
rect 24676 27421 24685 27455
rect 24685 27421 24719 27455
rect 24719 27421 24728 27455
rect 24676 27412 24728 27421
rect 24768 27412 24820 27464
rect 27160 27412 27212 27464
rect 27988 27455 28040 27464
rect 27988 27421 27997 27455
rect 27997 27421 28031 27455
rect 28031 27421 28040 27455
rect 27988 27412 28040 27421
rect 28264 27455 28316 27464
rect 28264 27421 28273 27455
rect 28273 27421 28307 27455
rect 28307 27421 28316 27455
rect 28264 27412 28316 27421
rect 28908 27455 28960 27464
rect 28908 27421 28917 27455
rect 28917 27421 28951 27455
rect 28951 27421 28960 27455
rect 28908 27412 28960 27421
rect 29184 27455 29236 27464
rect 29184 27421 29193 27455
rect 29193 27421 29227 27455
rect 29227 27421 29236 27455
rect 29184 27412 29236 27421
rect 29920 27489 29929 27523
rect 29929 27489 29963 27523
rect 29963 27489 29972 27523
rect 29920 27480 29972 27489
rect 30196 27523 30248 27532
rect 30196 27489 30205 27523
rect 30205 27489 30239 27523
rect 30239 27489 30248 27523
rect 30196 27480 30248 27489
rect 30288 27480 30340 27532
rect 31300 27523 31352 27532
rect 31300 27489 31309 27523
rect 31309 27489 31343 27523
rect 31343 27489 31352 27523
rect 31300 27480 31352 27489
rect 31668 27480 31720 27532
rect 32220 27480 32272 27532
rect 29828 27412 29880 27464
rect 30104 27455 30156 27464
rect 30104 27421 30113 27455
rect 30113 27421 30147 27455
rect 30147 27421 30156 27455
rect 30104 27412 30156 27421
rect 31116 27412 31168 27464
rect 31484 27412 31536 27464
rect 32036 27455 32088 27464
rect 32036 27421 32045 27455
rect 32045 27421 32079 27455
rect 32079 27421 32088 27455
rect 32036 27412 32088 27421
rect 23204 27344 23256 27396
rect 24860 27344 24912 27396
rect 25964 27344 26016 27396
rect 23756 27276 23808 27328
rect 25596 27319 25648 27328
rect 25596 27285 25605 27319
rect 25605 27285 25639 27319
rect 25639 27285 25648 27319
rect 25596 27276 25648 27285
rect 27068 27344 27120 27396
rect 28080 27344 28132 27396
rect 26148 27276 26200 27328
rect 27620 27276 27672 27328
rect 28724 27319 28776 27328
rect 28724 27285 28733 27319
rect 28733 27285 28767 27319
rect 28767 27285 28776 27319
rect 28724 27276 28776 27285
rect 29460 27276 29512 27328
rect 31576 27344 31628 27396
rect 31668 27344 31720 27396
rect 32496 27412 32548 27464
rect 30104 27276 30156 27328
rect 32588 27319 32640 27328
rect 32588 27285 32597 27319
rect 32597 27285 32631 27319
rect 32631 27285 32640 27319
rect 32588 27276 32640 27285
rect 9390 27174 9442 27226
rect 9454 27174 9506 27226
rect 9518 27174 9570 27226
rect 9582 27174 9634 27226
rect 9646 27174 9698 27226
rect 17831 27174 17883 27226
rect 17895 27174 17947 27226
rect 17959 27174 18011 27226
rect 18023 27174 18075 27226
rect 18087 27174 18139 27226
rect 26272 27174 26324 27226
rect 26336 27174 26388 27226
rect 26400 27174 26452 27226
rect 26464 27174 26516 27226
rect 26528 27174 26580 27226
rect 34713 27174 34765 27226
rect 34777 27174 34829 27226
rect 34841 27174 34893 27226
rect 34905 27174 34957 27226
rect 34969 27174 35021 27226
rect 6644 27115 6696 27124
rect 6644 27081 6653 27115
rect 6653 27081 6687 27115
rect 6687 27081 6696 27115
rect 6644 27072 6696 27081
rect 7656 27072 7708 27124
rect 2136 26936 2188 26988
rect 6552 26979 6604 26988
rect 6552 26945 6561 26979
rect 6561 26945 6595 26979
rect 6595 26945 6604 26979
rect 6552 26936 6604 26945
rect 8944 26979 8996 26988
rect 8944 26945 8953 26979
rect 8953 26945 8987 26979
rect 8987 26945 8996 26979
rect 8944 26936 8996 26945
rect 16304 26979 16356 26988
rect 16304 26945 16313 26979
rect 16313 26945 16347 26979
rect 16347 26945 16356 26979
rect 16304 26936 16356 26945
rect 18328 27072 18380 27124
rect 16764 27004 16816 27056
rect 17040 26979 17092 26988
rect 17040 26945 17049 26979
rect 17049 26945 17083 26979
rect 17083 26945 17092 26979
rect 17040 26936 17092 26945
rect 18236 27004 18288 27056
rect 16948 26868 17000 26920
rect 18052 26979 18104 26988
rect 18052 26945 18061 26979
rect 18061 26945 18095 26979
rect 18095 26945 18104 26979
rect 18512 26979 18564 26988
rect 18052 26936 18104 26945
rect 18512 26945 18521 26979
rect 18521 26945 18555 26979
rect 18555 26945 18564 26979
rect 18512 26936 18564 26945
rect 18788 27004 18840 27056
rect 19708 27047 19760 27056
rect 19432 26979 19484 26988
rect 19432 26945 19441 26979
rect 19441 26945 19475 26979
rect 19475 26945 19484 26979
rect 19432 26936 19484 26945
rect 19708 27013 19742 27047
rect 19742 27013 19760 27047
rect 19708 27004 19760 27013
rect 21456 26979 21508 26988
rect 21456 26945 21465 26979
rect 21465 26945 21499 26979
rect 21499 26945 21508 26979
rect 21456 26936 21508 26945
rect 22468 27004 22520 27056
rect 22652 27004 22704 27056
rect 23020 27004 23072 27056
rect 23296 27004 23348 27056
rect 28172 27072 28224 27124
rect 28540 27072 28592 27124
rect 32588 27072 32640 27124
rect 28724 27004 28776 27056
rect 23572 26936 23624 26988
rect 18144 26868 18196 26920
rect 18420 26868 18472 26920
rect 23020 26868 23072 26920
rect 24584 26936 24636 26988
rect 23756 26868 23808 26920
rect 27160 26979 27212 26988
rect 27160 26945 27169 26979
rect 27169 26945 27203 26979
rect 27203 26945 27212 26979
rect 27160 26936 27212 26945
rect 29368 26936 29420 26988
rect 29644 26979 29696 26988
rect 29644 26945 29653 26979
rect 29653 26945 29687 26979
rect 29687 26945 29696 26979
rect 29644 26936 29696 26945
rect 18236 26800 18288 26852
rect 20444 26800 20496 26852
rect 24400 26843 24452 26852
rect 16120 26775 16172 26784
rect 16120 26741 16129 26775
rect 16129 26741 16163 26775
rect 16163 26741 16172 26775
rect 16120 26732 16172 26741
rect 17040 26732 17092 26784
rect 17868 26732 17920 26784
rect 21272 26775 21324 26784
rect 21272 26741 21281 26775
rect 21281 26741 21315 26775
rect 21315 26741 21324 26775
rect 21272 26732 21324 26741
rect 24400 26809 24409 26843
rect 24409 26809 24443 26843
rect 24443 26809 24452 26843
rect 24400 26800 24452 26809
rect 23388 26775 23440 26784
rect 23388 26741 23397 26775
rect 23397 26741 23431 26775
rect 23431 26741 23440 26775
rect 24124 26775 24176 26784
rect 23388 26732 23440 26741
rect 24124 26741 24133 26775
rect 24133 26741 24167 26775
rect 24167 26741 24176 26775
rect 24124 26732 24176 26741
rect 24584 26732 24636 26784
rect 29184 26868 29236 26920
rect 29552 26868 29604 26920
rect 26332 26800 26384 26852
rect 27988 26800 28040 26852
rect 28172 26800 28224 26852
rect 31116 26936 31168 26988
rect 32956 27004 33008 27056
rect 31760 26979 31812 26988
rect 31760 26945 31769 26979
rect 31769 26945 31803 26979
rect 31803 26945 31812 26979
rect 31760 26936 31812 26945
rect 33600 27004 33652 27056
rect 34244 27004 34296 27056
rect 33508 26979 33560 26988
rect 33508 26945 33517 26979
rect 33517 26945 33551 26979
rect 33551 26945 33560 26979
rect 33508 26936 33560 26945
rect 33692 26979 33744 26988
rect 33692 26945 33701 26979
rect 33701 26945 33735 26979
rect 33735 26945 33744 26979
rect 33692 26936 33744 26945
rect 32128 26868 32180 26920
rect 32404 26911 32456 26920
rect 32404 26877 32413 26911
rect 32413 26877 32447 26911
rect 32447 26877 32456 26911
rect 32404 26868 32456 26877
rect 32864 26911 32916 26920
rect 32864 26877 32873 26911
rect 32873 26877 32907 26911
rect 32907 26877 32916 26911
rect 32864 26868 32916 26877
rect 33048 26868 33100 26920
rect 30932 26800 30984 26852
rect 34244 26800 34296 26852
rect 27068 26732 27120 26784
rect 29368 26775 29420 26784
rect 29368 26741 29377 26775
rect 29377 26741 29411 26775
rect 29411 26741 29420 26775
rect 29368 26732 29420 26741
rect 29644 26732 29696 26784
rect 29920 26732 29972 26784
rect 32404 26732 32456 26784
rect 33324 26775 33376 26784
rect 33324 26741 33333 26775
rect 33333 26741 33367 26775
rect 33367 26741 33376 26775
rect 33324 26732 33376 26741
rect 5170 26630 5222 26682
rect 5234 26630 5286 26682
rect 5298 26630 5350 26682
rect 5362 26630 5414 26682
rect 5426 26630 5478 26682
rect 13611 26630 13663 26682
rect 13675 26630 13727 26682
rect 13739 26630 13791 26682
rect 13803 26630 13855 26682
rect 13867 26630 13919 26682
rect 22052 26630 22104 26682
rect 22116 26630 22168 26682
rect 22180 26630 22232 26682
rect 22244 26630 22296 26682
rect 22308 26630 22360 26682
rect 30493 26630 30545 26682
rect 30557 26630 30609 26682
rect 30621 26630 30673 26682
rect 30685 26630 30737 26682
rect 30749 26630 30801 26682
rect 16948 26528 17000 26580
rect 19064 26528 19116 26580
rect 26148 26571 26200 26580
rect 26148 26537 26157 26571
rect 26157 26537 26191 26571
rect 26191 26537 26200 26571
rect 26148 26528 26200 26537
rect 16120 26460 16172 26512
rect 18972 26460 19024 26512
rect 19432 26503 19484 26512
rect 19432 26469 19441 26503
rect 19441 26469 19475 26503
rect 19475 26469 19484 26503
rect 19432 26460 19484 26469
rect 24400 26460 24452 26512
rect 24768 26460 24820 26512
rect 25044 26460 25096 26512
rect 29184 26528 29236 26580
rect 28264 26460 28316 26512
rect 28448 26460 28500 26512
rect 29644 26460 29696 26512
rect 17868 26435 17920 26444
rect 17868 26401 17877 26435
rect 17877 26401 17911 26435
rect 17911 26401 17920 26435
rect 17868 26392 17920 26401
rect 18788 26392 18840 26444
rect 22468 26435 22520 26444
rect 16764 26367 16816 26376
rect 16764 26333 16773 26367
rect 16773 26333 16807 26367
rect 16807 26333 16816 26367
rect 16764 26324 16816 26333
rect 17040 26367 17092 26376
rect 17040 26333 17049 26367
rect 17049 26333 17083 26367
rect 17083 26333 17092 26367
rect 17040 26324 17092 26333
rect 17316 26324 17368 26376
rect 17500 26367 17552 26376
rect 17500 26333 17509 26367
rect 17509 26333 17543 26367
rect 17543 26333 17552 26367
rect 17500 26324 17552 26333
rect 17684 26367 17736 26376
rect 17684 26333 17693 26367
rect 17693 26333 17727 26367
rect 17727 26333 17736 26367
rect 17684 26324 17736 26333
rect 16028 26256 16080 26308
rect 17408 26256 17460 26308
rect 18144 26324 18196 26376
rect 18604 26324 18656 26376
rect 18880 26367 18932 26376
rect 18880 26333 18889 26367
rect 18889 26333 18923 26367
rect 18923 26333 18932 26367
rect 18880 26324 18932 26333
rect 19340 26324 19392 26376
rect 22468 26401 22477 26435
rect 22477 26401 22511 26435
rect 22511 26401 22520 26435
rect 22468 26392 22520 26401
rect 23848 26392 23900 26444
rect 24860 26392 24912 26444
rect 26608 26392 26660 26444
rect 20812 26367 20864 26376
rect 20812 26333 20821 26367
rect 20821 26333 20855 26367
rect 20855 26333 20864 26367
rect 20812 26324 20864 26333
rect 23204 26367 23256 26376
rect 23204 26333 23213 26367
rect 23213 26333 23247 26367
rect 23247 26333 23256 26367
rect 23204 26324 23256 26333
rect 23480 26367 23532 26376
rect 23480 26333 23515 26367
rect 23515 26333 23532 26367
rect 23480 26324 23532 26333
rect 18328 26256 18380 26308
rect 20536 26256 20588 26308
rect 23296 26299 23348 26308
rect 23296 26265 23305 26299
rect 23305 26265 23339 26299
rect 23339 26265 23348 26299
rect 23296 26256 23348 26265
rect 23388 26299 23440 26308
rect 23388 26265 23397 26299
rect 23397 26265 23431 26299
rect 23431 26265 23440 26299
rect 23388 26256 23440 26265
rect 25412 26256 25464 26308
rect 26792 26324 26844 26376
rect 29736 26392 29788 26444
rect 30196 26528 30248 26580
rect 33692 26528 33744 26580
rect 29920 26460 29972 26512
rect 30288 26367 30340 26376
rect 26056 26256 26108 26308
rect 27528 26256 27580 26308
rect 30288 26333 30297 26367
rect 30297 26333 30331 26367
rect 30331 26333 30340 26367
rect 30288 26324 30340 26333
rect 30840 26392 30892 26444
rect 31576 26324 31628 26376
rect 31760 26367 31812 26376
rect 31760 26333 31769 26367
rect 31769 26333 31803 26367
rect 31803 26333 31812 26367
rect 31760 26324 31812 26333
rect 32680 26460 32732 26512
rect 32404 26392 32456 26444
rect 32128 26367 32180 26376
rect 18420 26188 18472 26240
rect 23020 26231 23072 26240
rect 23020 26197 23029 26231
rect 23029 26197 23063 26231
rect 23063 26197 23072 26231
rect 23020 26188 23072 26197
rect 25596 26188 25648 26240
rect 26884 26188 26936 26240
rect 30932 26256 30984 26308
rect 32128 26333 32137 26367
rect 32137 26333 32171 26367
rect 32171 26333 32180 26367
rect 32128 26324 32180 26333
rect 32312 26324 32364 26376
rect 32404 26256 32456 26308
rect 32680 26256 32732 26308
rect 33416 26256 33468 26308
rect 27804 26188 27856 26240
rect 28264 26188 28316 26240
rect 28724 26188 28776 26240
rect 29552 26188 29604 26240
rect 29736 26188 29788 26240
rect 31024 26188 31076 26240
rect 31484 26188 31536 26240
rect 32128 26188 32180 26240
rect 33232 26188 33284 26240
rect 9390 26086 9442 26138
rect 9454 26086 9506 26138
rect 9518 26086 9570 26138
rect 9582 26086 9634 26138
rect 9646 26086 9698 26138
rect 17831 26086 17883 26138
rect 17895 26086 17947 26138
rect 17959 26086 18011 26138
rect 18023 26086 18075 26138
rect 18087 26086 18139 26138
rect 26272 26086 26324 26138
rect 26336 26086 26388 26138
rect 26400 26086 26452 26138
rect 26464 26086 26516 26138
rect 26528 26086 26580 26138
rect 34713 26086 34765 26138
rect 34777 26086 34829 26138
rect 34841 26086 34893 26138
rect 34905 26086 34957 26138
rect 34969 26086 35021 26138
rect 25780 25984 25832 26036
rect 18144 25916 18196 25968
rect 18236 25916 18288 25968
rect 17592 25891 17644 25900
rect 17592 25857 17601 25891
rect 17601 25857 17635 25891
rect 17635 25857 17644 25891
rect 17592 25848 17644 25857
rect 17684 25891 17736 25900
rect 17684 25857 17693 25891
rect 17693 25857 17727 25891
rect 17727 25857 17736 25891
rect 17684 25848 17736 25857
rect 18328 25848 18380 25900
rect 18604 25891 18656 25900
rect 18604 25857 18613 25891
rect 18613 25857 18647 25891
rect 18647 25857 18656 25891
rect 18604 25848 18656 25857
rect 18788 25891 18840 25900
rect 18788 25857 18797 25891
rect 18797 25857 18831 25891
rect 18831 25857 18840 25891
rect 18788 25848 18840 25857
rect 20720 25916 20772 25968
rect 19432 25848 19484 25900
rect 17408 25780 17460 25832
rect 19340 25712 19392 25764
rect 20444 25712 20496 25764
rect 1584 25644 1636 25696
rect 17408 25644 17460 25696
rect 19616 25644 19668 25696
rect 20904 25644 20956 25696
rect 21180 25687 21232 25696
rect 21180 25653 21189 25687
rect 21189 25653 21223 25687
rect 21223 25653 21232 25687
rect 21180 25644 21232 25653
rect 22376 25848 22428 25900
rect 22468 25848 22520 25900
rect 23020 25916 23072 25968
rect 23848 25916 23900 25968
rect 25412 25916 25464 25968
rect 27436 25984 27488 26036
rect 27528 25959 27580 25968
rect 24584 25848 24636 25900
rect 25872 25848 25924 25900
rect 24308 25780 24360 25832
rect 27528 25925 27537 25959
rect 27537 25925 27571 25959
rect 27571 25925 27580 25959
rect 27528 25916 27580 25925
rect 27344 25848 27396 25900
rect 27620 25848 27672 25900
rect 27804 25891 27856 25900
rect 27804 25857 27813 25891
rect 27813 25857 27847 25891
rect 27847 25857 27856 25891
rect 27804 25848 27856 25857
rect 27988 25891 28040 25900
rect 27988 25857 27997 25891
rect 27997 25857 28031 25891
rect 28031 25857 28040 25891
rect 27988 25848 28040 25857
rect 28172 25891 28224 25900
rect 28172 25857 28181 25891
rect 28181 25857 28215 25891
rect 28215 25857 28224 25891
rect 28172 25848 28224 25857
rect 29092 25916 29144 25968
rect 31760 25916 31812 25968
rect 28724 25848 28776 25900
rect 29368 25848 29420 25900
rect 31024 25891 31076 25900
rect 31024 25857 31033 25891
rect 31033 25857 31067 25891
rect 31067 25857 31076 25891
rect 31024 25848 31076 25857
rect 31392 25891 31444 25900
rect 31392 25857 31401 25891
rect 31401 25857 31435 25891
rect 31435 25857 31444 25891
rect 31392 25848 31444 25857
rect 31484 25891 31536 25900
rect 31484 25857 31498 25891
rect 31498 25857 31532 25891
rect 31532 25857 31536 25891
rect 31484 25848 31536 25857
rect 34336 25891 34388 25900
rect 34336 25857 34345 25891
rect 34345 25857 34379 25891
rect 34379 25857 34388 25891
rect 34336 25848 34388 25857
rect 22008 25755 22060 25764
rect 22008 25721 22017 25755
rect 22017 25721 22051 25755
rect 22051 25721 22060 25755
rect 22008 25712 22060 25721
rect 24400 25712 24452 25764
rect 25688 25712 25740 25764
rect 26976 25712 27028 25764
rect 27252 25712 27304 25764
rect 27896 25712 27948 25764
rect 28172 25712 28224 25764
rect 31944 25780 31996 25832
rect 24492 25644 24544 25696
rect 26424 25644 26476 25696
rect 29920 25644 29972 25696
rect 31208 25644 31260 25696
rect 31668 25687 31720 25696
rect 31668 25653 31677 25687
rect 31677 25653 31711 25687
rect 31711 25653 31720 25687
rect 31668 25644 31720 25653
rect 5170 25542 5222 25594
rect 5234 25542 5286 25594
rect 5298 25542 5350 25594
rect 5362 25542 5414 25594
rect 5426 25542 5478 25594
rect 13611 25542 13663 25594
rect 13675 25542 13727 25594
rect 13739 25542 13791 25594
rect 13803 25542 13855 25594
rect 13867 25542 13919 25594
rect 22052 25542 22104 25594
rect 22116 25542 22168 25594
rect 22180 25542 22232 25594
rect 22244 25542 22296 25594
rect 22308 25542 22360 25594
rect 30493 25542 30545 25594
rect 30557 25542 30609 25594
rect 30621 25542 30673 25594
rect 30685 25542 30737 25594
rect 30749 25542 30801 25594
rect 18880 25440 18932 25492
rect 19432 25483 19484 25492
rect 19432 25449 19441 25483
rect 19441 25449 19475 25483
rect 19475 25449 19484 25483
rect 19432 25440 19484 25449
rect 23296 25440 23348 25492
rect 24952 25483 25004 25492
rect 24952 25449 24961 25483
rect 24961 25449 24995 25483
rect 24995 25449 25004 25483
rect 24952 25440 25004 25449
rect 27988 25440 28040 25492
rect 28356 25440 28408 25492
rect 29276 25440 29328 25492
rect 31024 25440 31076 25492
rect 1584 25347 1636 25356
rect 1584 25313 1593 25347
rect 1593 25313 1627 25347
rect 1627 25313 1636 25347
rect 1584 25304 1636 25313
rect 2780 25347 2832 25356
rect 2780 25313 2789 25347
rect 2789 25313 2823 25347
rect 2823 25313 2832 25347
rect 2780 25304 2832 25313
rect 15292 25279 15344 25288
rect 15292 25245 15301 25279
rect 15301 25245 15335 25279
rect 15335 25245 15344 25279
rect 15292 25236 15344 25245
rect 20628 25372 20680 25424
rect 26056 25372 26108 25424
rect 18420 25347 18472 25356
rect 16580 25279 16632 25288
rect 16580 25245 16589 25279
rect 16589 25245 16623 25279
rect 16623 25245 16632 25279
rect 16580 25236 16632 25245
rect 17040 25236 17092 25288
rect 17132 25236 17184 25288
rect 17408 25279 17460 25288
rect 17408 25245 17417 25279
rect 17417 25245 17451 25279
rect 17451 25245 17460 25279
rect 17408 25236 17460 25245
rect 1768 25211 1820 25220
rect 1768 25177 1777 25211
rect 1777 25177 1811 25211
rect 1811 25177 1820 25211
rect 1768 25168 1820 25177
rect 16856 25168 16908 25220
rect 18052 25168 18104 25220
rect 18420 25313 18429 25347
rect 18429 25313 18463 25347
rect 18463 25313 18472 25347
rect 18420 25304 18472 25313
rect 22468 25304 22520 25356
rect 22836 25347 22888 25356
rect 22836 25313 22845 25347
rect 22845 25313 22879 25347
rect 22879 25313 22888 25347
rect 22836 25304 22888 25313
rect 26148 25304 26200 25356
rect 26332 25304 26384 25356
rect 26516 25304 26568 25356
rect 26700 25304 26752 25356
rect 27528 25372 27580 25424
rect 29001 25372 29053 25424
rect 31576 25347 31628 25356
rect 18788 25236 18840 25288
rect 19616 25236 19668 25288
rect 18604 25168 18656 25220
rect 19064 25168 19116 25220
rect 19892 25279 19944 25288
rect 19892 25245 19906 25279
rect 19906 25245 19940 25279
rect 19940 25245 19944 25279
rect 19892 25236 19944 25245
rect 20076 25279 20128 25288
rect 20076 25245 20085 25279
rect 20085 25245 20119 25279
rect 20119 25245 20128 25279
rect 20076 25236 20128 25245
rect 20720 25236 20772 25288
rect 21916 25236 21968 25288
rect 23020 25236 23072 25288
rect 23388 25236 23440 25288
rect 24216 25236 24268 25288
rect 25688 25279 25740 25288
rect 25688 25245 25697 25279
rect 25697 25245 25731 25279
rect 25731 25245 25740 25279
rect 25688 25236 25740 25245
rect 26056 25279 26108 25288
rect 21272 25168 21324 25220
rect 23296 25168 23348 25220
rect 24584 25168 24636 25220
rect 25412 25168 25464 25220
rect 26056 25245 26065 25279
rect 26065 25245 26099 25279
rect 26099 25245 26108 25279
rect 26056 25236 26108 25245
rect 26608 25236 26660 25288
rect 17592 25143 17644 25152
rect 17592 25109 17601 25143
rect 17601 25109 17635 25143
rect 17635 25109 17644 25143
rect 17592 25100 17644 25109
rect 18880 25100 18932 25152
rect 22928 25100 22980 25152
rect 23572 25100 23624 25152
rect 26792 25236 26844 25288
rect 31576 25313 31585 25347
rect 31585 25313 31619 25347
rect 31619 25313 31628 25347
rect 31576 25304 31628 25313
rect 31760 25304 31812 25356
rect 32036 25304 32088 25356
rect 32864 25304 32916 25356
rect 26976 25168 27028 25220
rect 27436 25279 27488 25288
rect 27436 25245 27445 25279
rect 27445 25245 27479 25279
rect 27479 25245 27488 25279
rect 28080 25279 28132 25288
rect 27436 25236 27488 25245
rect 28080 25245 28089 25279
rect 28089 25245 28123 25279
rect 28123 25245 28132 25279
rect 28080 25236 28132 25245
rect 28356 25279 28408 25288
rect 28356 25245 28365 25279
rect 28365 25245 28399 25279
rect 28399 25245 28408 25279
rect 28356 25236 28408 25245
rect 27252 25168 27304 25220
rect 26884 25143 26936 25152
rect 26884 25109 26893 25143
rect 26893 25109 26927 25143
rect 26927 25109 26936 25143
rect 26884 25100 26936 25109
rect 28356 25100 28408 25152
rect 28448 25100 28500 25152
rect 30104 25236 30156 25288
rect 30656 25279 30708 25288
rect 30656 25245 30665 25279
rect 30665 25245 30699 25279
rect 30699 25245 30708 25279
rect 30656 25236 30708 25245
rect 31116 25236 31168 25288
rect 30380 25168 30432 25220
rect 29644 25100 29696 25152
rect 30748 25168 30800 25220
rect 31944 25236 31996 25288
rect 34060 25168 34112 25220
rect 34336 25211 34388 25220
rect 34336 25177 34345 25211
rect 34345 25177 34379 25211
rect 34379 25177 34388 25211
rect 34336 25168 34388 25177
rect 31576 25100 31628 25152
rect 9390 24998 9442 25050
rect 9454 24998 9506 25050
rect 9518 24998 9570 25050
rect 9582 24998 9634 25050
rect 9646 24998 9698 25050
rect 17831 24998 17883 25050
rect 17895 24998 17947 25050
rect 17959 24998 18011 25050
rect 18023 24998 18075 25050
rect 18087 24998 18139 25050
rect 26272 24998 26324 25050
rect 26336 24998 26388 25050
rect 26400 24998 26452 25050
rect 26464 24998 26516 25050
rect 26528 24998 26580 25050
rect 34713 24998 34765 25050
rect 34777 24998 34829 25050
rect 34841 24998 34893 25050
rect 34905 24998 34957 25050
rect 34969 24998 35021 25050
rect 1768 24896 1820 24948
rect 16580 24896 16632 24948
rect 17316 24896 17368 24948
rect 19616 24896 19668 24948
rect 23020 24896 23072 24948
rect 23204 24896 23256 24948
rect 26608 24896 26660 24948
rect 26976 24896 27028 24948
rect 27620 24896 27672 24948
rect 28356 24896 28408 24948
rect 31944 24896 31996 24948
rect 17408 24871 17460 24880
rect 17408 24837 17417 24871
rect 17417 24837 17451 24871
rect 17451 24837 17460 24871
rect 17408 24828 17460 24837
rect 17500 24828 17552 24880
rect 19892 24828 19944 24880
rect 2044 24803 2096 24812
rect 2044 24769 2053 24803
rect 2053 24769 2087 24803
rect 2087 24769 2096 24803
rect 2044 24760 2096 24769
rect 3056 24760 3108 24812
rect 16028 24803 16080 24812
rect 16028 24769 16037 24803
rect 16037 24769 16071 24803
rect 16071 24769 16080 24803
rect 16028 24760 16080 24769
rect 17224 24760 17276 24812
rect 18328 24760 18380 24812
rect 18880 24803 18932 24812
rect 18880 24769 18889 24803
rect 18889 24769 18923 24803
rect 18923 24769 18932 24803
rect 18880 24760 18932 24769
rect 19064 24803 19116 24812
rect 19064 24769 19073 24803
rect 19073 24769 19107 24803
rect 19107 24769 19116 24803
rect 19064 24760 19116 24769
rect 20720 24828 20772 24880
rect 18604 24692 18656 24744
rect 21180 24760 21232 24812
rect 22560 24828 22612 24880
rect 21456 24803 21508 24812
rect 21456 24769 21465 24803
rect 21465 24769 21499 24803
rect 21499 24769 21508 24803
rect 21456 24760 21508 24769
rect 21916 24760 21968 24812
rect 22744 24803 22796 24812
rect 22744 24769 22778 24803
rect 22778 24769 22796 24803
rect 24676 24828 24728 24880
rect 25504 24828 25556 24880
rect 24308 24803 24360 24812
rect 22744 24760 22796 24769
rect 24308 24769 24317 24803
rect 24317 24769 24351 24803
rect 24351 24769 24360 24803
rect 24308 24760 24360 24769
rect 20536 24692 20588 24744
rect 20996 24692 21048 24744
rect 22376 24692 22428 24744
rect 26700 24828 26752 24880
rect 27068 24828 27120 24880
rect 28448 24828 28500 24880
rect 26792 24760 26844 24812
rect 28172 24760 28224 24812
rect 29736 24828 29788 24880
rect 17316 24556 17368 24608
rect 17684 24556 17736 24608
rect 18328 24599 18380 24608
rect 18328 24565 18337 24599
rect 18337 24565 18371 24599
rect 18371 24565 18380 24599
rect 18328 24556 18380 24565
rect 20628 24556 20680 24608
rect 30564 24828 30616 24880
rect 30656 24828 30708 24880
rect 30196 24760 30248 24812
rect 23848 24599 23900 24608
rect 23848 24565 23857 24599
rect 23857 24565 23891 24599
rect 23891 24565 23900 24599
rect 23848 24556 23900 24565
rect 27068 24556 27120 24608
rect 29552 24692 29604 24744
rect 31024 24760 31076 24812
rect 31576 24828 31628 24880
rect 31852 24828 31904 24880
rect 33600 24871 33652 24880
rect 33600 24837 33609 24871
rect 33609 24837 33643 24871
rect 33643 24837 33652 24871
rect 33600 24828 33652 24837
rect 31484 24760 31536 24812
rect 31208 24692 31260 24744
rect 30748 24624 30800 24676
rect 31484 24624 31536 24676
rect 32128 24624 32180 24676
rect 32404 24624 32456 24676
rect 32680 24803 32732 24812
rect 32680 24769 32689 24803
rect 32689 24769 32723 24803
rect 32723 24769 32732 24803
rect 32680 24760 32732 24769
rect 33232 24760 33284 24812
rect 33416 24760 33468 24812
rect 34060 24760 34112 24812
rect 33508 24624 33560 24676
rect 29092 24556 29144 24608
rect 29736 24556 29788 24608
rect 29920 24556 29972 24608
rect 31116 24599 31168 24608
rect 31116 24565 31125 24599
rect 31125 24565 31159 24599
rect 31159 24565 31168 24599
rect 31116 24556 31168 24565
rect 31852 24556 31904 24608
rect 5170 24454 5222 24506
rect 5234 24454 5286 24506
rect 5298 24454 5350 24506
rect 5362 24454 5414 24506
rect 5426 24454 5478 24506
rect 13611 24454 13663 24506
rect 13675 24454 13727 24506
rect 13739 24454 13791 24506
rect 13803 24454 13855 24506
rect 13867 24454 13919 24506
rect 22052 24454 22104 24506
rect 22116 24454 22168 24506
rect 22180 24454 22232 24506
rect 22244 24454 22296 24506
rect 22308 24454 22360 24506
rect 30493 24454 30545 24506
rect 30557 24454 30609 24506
rect 30621 24454 30673 24506
rect 30685 24454 30737 24506
rect 30749 24454 30801 24506
rect 16856 24352 16908 24404
rect 17224 24395 17276 24404
rect 17224 24361 17233 24395
rect 17233 24361 17267 24395
rect 17267 24361 17276 24395
rect 17224 24352 17276 24361
rect 18420 24352 18472 24404
rect 16028 24216 16080 24268
rect 15752 24191 15804 24200
rect 15752 24157 15761 24191
rect 15761 24157 15795 24191
rect 15795 24157 15804 24191
rect 16764 24216 16816 24268
rect 15752 24148 15804 24157
rect 17500 24148 17552 24200
rect 17316 24080 17368 24132
rect 16672 24012 16724 24064
rect 17408 24012 17460 24064
rect 18604 24191 18656 24200
rect 18604 24157 18613 24191
rect 18613 24157 18647 24191
rect 18647 24157 18656 24191
rect 18604 24148 18656 24157
rect 20076 24352 20128 24404
rect 20996 24352 21048 24404
rect 22376 24352 22428 24404
rect 22468 24352 22520 24404
rect 22928 24395 22980 24404
rect 22928 24361 22937 24395
rect 22937 24361 22971 24395
rect 22971 24361 22980 24395
rect 22928 24352 22980 24361
rect 23112 24395 23164 24404
rect 23112 24361 23121 24395
rect 23121 24361 23155 24395
rect 23155 24361 23164 24395
rect 23112 24352 23164 24361
rect 24032 24352 24084 24404
rect 26976 24352 27028 24404
rect 27436 24352 27488 24404
rect 31392 24352 31444 24404
rect 33048 24352 33100 24404
rect 21180 24216 21232 24268
rect 22468 24216 22520 24268
rect 18880 24191 18932 24200
rect 18880 24157 18889 24191
rect 18889 24157 18923 24191
rect 18923 24157 18932 24191
rect 18880 24148 18932 24157
rect 19064 24148 19116 24200
rect 21732 24148 21784 24200
rect 22284 24148 22336 24200
rect 24400 24284 24452 24336
rect 32404 24284 32456 24336
rect 23112 24216 23164 24268
rect 24952 24259 25004 24268
rect 24952 24225 24961 24259
rect 24961 24225 24995 24259
rect 24995 24225 25004 24259
rect 24952 24216 25004 24225
rect 27068 24259 27120 24268
rect 22560 24080 22612 24132
rect 22652 24123 22704 24132
rect 22652 24089 22661 24123
rect 22661 24089 22695 24123
rect 22695 24089 22704 24123
rect 22652 24080 22704 24089
rect 23204 24080 23256 24132
rect 21180 24012 21232 24064
rect 22192 24055 22244 24064
rect 22192 24021 22201 24055
rect 22201 24021 22235 24055
rect 22235 24021 22244 24055
rect 22192 24012 22244 24021
rect 22284 24012 22336 24064
rect 22744 24012 22796 24064
rect 25044 24148 25096 24200
rect 25964 24148 26016 24200
rect 27068 24225 27077 24259
rect 27077 24225 27111 24259
rect 27111 24225 27120 24259
rect 27068 24216 27120 24225
rect 28448 24259 28500 24268
rect 28448 24225 28457 24259
rect 28457 24225 28491 24259
rect 28491 24225 28500 24259
rect 28448 24216 28500 24225
rect 28724 24216 28776 24268
rect 29552 24216 29604 24268
rect 30932 24216 30984 24268
rect 31024 24216 31076 24268
rect 34152 24216 34204 24268
rect 26884 24148 26936 24200
rect 26976 24191 27028 24200
rect 26976 24157 26985 24191
rect 26985 24157 27019 24191
rect 27019 24157 27028 24191
rect 28356 24191 28408 24200
rect 26976 24148 27028 24157
rect 28356 24157 28365 24191
rect 28365 24157 28399 24191
rect 28399 24157 28408 24191
rect 28356 24148 28408 24157
rect 30288 24148 30340 24200
rect 30656 24191 30708 24200
rect 30656 24157 30665 24191
rect 30665 24157 30699 24191
rect 30699 24157 30708 24191
rect 30656 24148 30708 24157
rect 31116 24148 31168 24200
rect 31852 24148 31904 24200
rect 32036 24191 32088 24200
rect 32036 24157 32045 24191
rect 32045 24157 32079 24191
rect 32079 24157 32088 24191
rect 32036 24148 32088 24157
rect 32496 24191 32548 24200
rect 32496 24157 32505 24191
rect 32505 24157 32539 24191
rect 32539 24157 32548 24191
rect 32496 24148 32548 24157
rect 26700 24080 26752 24132
rect 28724 24080 28776 24132
rect 32680 24123 32732 24132
rect 32680 24089 32689 24123
rect 32689 24089 32723 24123
rect 32723 24089 32732 24123
rect 32680 24080 32732 24089
rect 34336 24123 34388 24132
rect 34336 24089 34345 24123
rect 34345 24089 34379 24123
rect 34379 24089 34388 24123
rect 34336 24080 34388 24089
rect 28172 24055 28224 24064
rect 28172 24021 28181 24055
rect 28181 24021 28215 24055
rect 28215 24021 28224 24055
rect 28172 24012 28224 24021
rect 28448 24012 28500 24064
rect 30196 24012 30248 24064
rect 31852 24012 31904 24064
rect 32220 24012 32272 24064
rect 9390 23910 9442 23962
rect 9454 23910 9506 23962
rect 9518 23910 9570 23962
rect 9582 23910 9634 23962
rect 9646 23910 9698 23962
rect 17831 23910 17883 23962
rect 17895 23910 17947 23962
rect 17959 23910 18011 23962
rect 18023 23910 18075 23962
rect 18087 23910 18139 23962
rect 26272 23910 26324 23962
rect 26336 23910 26388 23962
rect 26400 23910 26452 23962
rect 26464 23910 26516 23962
rect 26528 23910 26580 23962
rect 34713 23910 34765 23962
rect 34777 23910 34829 23962
rect 34841 23910 34893 23962
rect 34905 23910 34957 23962
rect 34969 23910 35021 23962
rect 8944 23808 8996 23860
rect 22192 23808 22244 23860
rect 22376 23808 22428 23860
rect 22652 23808 22704 23860
rect 23296 23808 23348 23860
rect 23848 23808 23900 23860
rect 27620 23808 27672 23860
rect 29736 23808 29788 23860
rect 31760 23808 31812 23860
rect 32404 23808 32456 23860
rect 17500 23740 17552 23792
rect 17684 23740 17736 23792
rect 16028 23647 16080 23656
rect 16028 23613 16037 23647
rect 16037 23613 16071 23647
rect 16071 23613 16080 23647
rect 16028 23604 16080 23613
rect 17224 23715 17276 23724
rect 17224 23681 17233 23715
rect 17233 23681 17267 23715
rect 17267 23681 17276 23715
rect 17224 23672 17276 23681
rect 17960 23672 18012 23724
rect 18328 23672 18380 23724
rect 19064 23715 19116 23724
rect 16856 23604 16908 23656
rect 17316 23647 17368 23656
rect 17316 23613 17325 23647
rect 17325 23613 17359 23647
rect 17359 23613 17368 23647
rect 17316 23604 17368 23613
rect 18604 23604 18656 23656
rect 17500 23536 17552 23588
rect 19064 23681 19073 23715
rect 19073 23681 19107 23715
rect 19107 23681 19116 23715
rect 19064 23672 19116 23681
rect 22284 23740 22336 23792
rect 23388 23740 23440 23792
rect 22468 23672 22520 23724
rect 24308 23740 24360 23792
rect 26884 23740 26936 23792
rect 28540 23740 28592 23792
rect 22652 23604 22704 23656
rect 16120 23468 16172 23520
rect 20720 23536 20772 23588
rect 24400 23672 24452 23724
rect 25688 23715 25740 23724
rect 25688 23681 25697 23715
rect 25697 23681 25731 23715
rect 25731 23681 25740 23715
rect 25688 23672 25740 23681
rect 25964 23672 26016 23724
rect 26976 23672 27028 23724
rect 29000 23672 29052 23724
rect 31484 23672 31536 23724
rect 26608 23604 26660 23656
rect 27068 23604 27120 23656
rect 28448 23604 28500 23656
rect 28816 23604 28868 23656
rect 29092 23604 29144 23656
rect 30104 23604 30156 23656
rect 20260 23468 20312 23520
rect 20536 23468 20588 23520
rect 27528 23536 27580 23588
rect 28632 23536 28684 23588
rect 30288 23536 30340 23588
rect 30656 23604 30708 23656
rect 31392 23604 31444 23656
rect 34428 23740 34480 23792
rect 32496 23647 32548 23656
rect 32496 23613 32505 23647
rect 32505 23613 32539 23647
rect 32539 23613 32548 23647
rect 32496 23604 32548 23613
rect 32680 23647 32732 23656
rect 32680 23613 32689 23647
rect 32689 23613 32723 23647
rect 32723 23613 32732 23647
rect 32680 23604 32732 23613
rect 22376 23468 22428 23520
rect 23020 23511 23072 23520
rect 23020 23477 23029 23511
rect 23029 23477 23063 23511
rect 23063 23477 23072 23511
rect 23020 23468 23072 23477
rect 25044 23468 25096 23520
rect 25412 23511 25464 23520
rect 25412 23477 25421 23511
rect 25421 23477 25455 23511
rect 25455 23477 25464 23511
rect 25412 23468 25464 23477
rect 28356 23468 28408 23520
rect 28908 23468 28960 23520
rect 30840 23511 30892 23520
rect 30840 23477 30849 23511
rect 30849 23477 30883 23511
rect 30883 23477 30892 23511
rect 30840 23468 30892 23477
rect 30932 23468 30984 23520
rect 32036 23536 32088 23588
rect 32864 23536 32916 23588
rect 32312 23468 32364 23520
rect 5170 23366 5222 23418
rect 5234 23366 5286 23418
rect 5298 23366 5350 23418
rect 5362 23366 5414 23418
rect 5426 23366 5478 23418
rect 13611 23366 13663 23418
rect 13675 23366 13727 23418
rect 13739 23366 13791 23418
rect 13803 23366 13855 23418
rect 13867 23366 13919 23418
rect 22052 23366 22104 23418
rect 22116 23366 22168 23418
rect 22180 23366 22232 23418
rect 22244 23366 22296 23418
rect 22308 23366 22360 23418
rect 30493 23366 30545 23418
rect 30557 23366 30609 23418
rect 30621 23366 30673 23418
rect 30685 23366 30737 23418
rect 30749 23366 30801 23418
rect 16672 23307 16724 23316
rect 16672 23273 16681 23307
rect 16681 23273 16715 23307
rect 16715 23273 16724 23307
rect 16672 23264 16724 23273
rect 18420 23264 18472 23316
rect 18696 23264 18748 23316
rect 21916 23264 21968 23316
rect 17592 23171 17644 23180
rect 17592 23137 17601 23171
rect 17601 23137 17635 23171
rect 17635 23137 17644 23171
rect 17592 23128 17644 23137
rect 18788 23196 18840 23248
rect 22376 23196 22428 23248
rect 22560 23196 22612 23248
rect 16580 23103 16632 23112
rect 16580 23069 16589 23103
rect 16589 23069 16623 23103
rect 16623 23069 16632 23103
rect 16580 23060 16632 23069
rect 16764 23103 16816 23112
rect 16764 23069 16773 23103
rect 16773 23069 16807 23103
rect 16807 23069 16816 23103
rect 16764 23060 16816 23069
rect 17408 23060 17460 23112
rect 19708 23128 19760 23180
rect 20076 23128 20128 23180
rect 28264 23264 28316 23316
rect 26884 23239 26936 23248
rect 26884 23205 26893 23239
rect 26893 23205 26927 23239
rect 26927 23205 26936 23239
rect 26884 23196 26936 23205
rect 18236 22992 18288 23044
rect 19984 23060 20036 23112
rect 20444 23060 20496 23112
rect 20812 23103 20864 23112
rect 20812 23069 20821 23103
rect 20821 23069 20855 23103
rect 20855 23069 20864 23103
rect 20812 23060 20864 23069
rect 23204 23103 23256 23112
rect 23204 23069 23213 23103
rect 23213 23069 23247 23103
rect 23247 23069 23256 23103
rect 23204 23060 23256 23069
rect 23480 23103 23532 23112
rect 23480 23069 23489 23103
rect 23489 23069 23523 23103
rect 23523 23069 23532 23103
rect 23480 23060 23532 23069
rect 24952 23103 25004 23112
rect 20352 22992 20404 23044
rect 24952 23069 24961 23103
rect 24961 23069 24995 23103
rect 24995 23069 25004 23103
rect 24952 23060 25004 23069
rect 25228 23060 25280 23112
rect 29092 23264 29144 23316
rect 31944 23264 31996 23316
rect 29368 23196 29420 23248
rect 31300 23239 31352 23248
rect 31300 23205 31309 23239
rect 31309 23205 31343 23239
rect 31343 23205 31352 23239
rect 31300 23196 31352 23205
rect 28816 23171 28868 23180
rect 28816 23137 28825 23171
rect 28825 23137 28859 23171
rect 28859 23137 28868 23171
rect 28816 23128 28868 23137
rect 28448 23103 28500 23112
rect 28448 23069 28457 23103
rect 28457 23069 28491 23103
rect 28491 23069 28500 23103
rect 28448 23060 28500 23069
rect 25320 22992 25372 23044
rect 25412 22992 25464 23044
rect 27068 22992 27120 23044
rect 27528 22992 27580 23044
rect 27620 22992 27672 23044
rect 28356 22992 28408 23044
rect 29000 23103 29052 23112
rect 29000 23069 29020 23103
rect 29020 23069 29052 23103
rect 29000 23060 29052 23069
rect 18788 22967 18840 22976
rect 18788 22933 18797 22967
rect 18797 22933 18831 22967
rect 18831 22933 18840 22967
rect 18788 22924 18840 22933
rect 19432 22967 19484 22976
rect 19432 22933 19441 22967
rect 19441 22933 19475 22967
rect 19475 22933 19484 22967
rect 19432 22924 19484 22933
rect 22744 22924 22796 22976
rect 24584 22967 24636 22976
rect 24584 22933 24593 22967
rect 24593 22933 24627 22967
rect 24627 22933 24636 22967
rect 24584 22924 24636 22933
rect 28632 22924 28684 22976
rect 29184 22967 29236 22976
rect 29184 22933 29193 22967
rect 29193 22933 29227 22967
rect 29227 22933 29236 22967
rect 29184 22924 29236 22933
rect 31024 23060 31076 23112
rect 34336 23171 34388 23180
rect 34336 23137 34345 23171
rect 34345 23137 34379 23171
rect 34379 23137 34388 23171
rect 34336 23128 34388 23137
rect 32036 23060 32088 23112
rect 32496 23103 32548 23112
rect 32496 23069 32505 23103
rect 32505 23069 32539 23103
rect 32539 23069 32548 23103
rect 32496 23060 32548 23069
rect 32680 23035 32732 23044
rect 30104 22924 30156 22976
rect 30288 22924 30340 22976
rect 30472 22924 30524 22976
rect 31116 22924 31168 22976
rect 32680 23001 32689 23035
rect 32689 23001 32723 23035
rect 32723 23001 32732 23035
rect 32680 22992 32732 23001
rect 34520 22924 34572 22976
rect 9390 22822 9442 22874
rect 9454 22822 9506 22874
rect 9518 22822 9570 22874
rect 9582 22822 9634 22874
rect 9646 22822 9698 22874
rect 17831 22822 17883 22874
rect 17895 22822 17947 22874
rect 17959 22822 18011 22874
rect 18023 22822 18075 22874
rect 18087 22822 18139 22874
rect 26272 22822 26324 22874
rect 26336 22822 26388 22874
rect 26400 22822 26452 22874
rect 26464 22822 26516 22874
rect 26528 22822 26580 22874
rect 34713 22822 34765 22874
rect 34777 22822 34829 22874
rect 34841 22822 34893 22874
rect 34905 22822 34957 22874
rect 34969 22822 35021 22874
rect 17316 22720 17368 22772
rect 19708 22720 19760 22772
rect 23480 22720 23532 22772
rect 16580 22584 16632 22636
rect 17592 22584 17644 22636
rect 19064 22652 19116 22704
rect 19432 22584 19484 22636
rect 20628 22627 20680 22636
rect 20628 22593 20637 22627
rect 20637 22593 20671 22627
rect 20671 22593 20680 22627
rect 20628 22584 20680 22593
rect 20720 22584 20772 22636
rect 20904 22627 20956 22636
rect 20904 22593 20913 22627
rect 20913 22593 20947 22627
rect 20947 22593 20956 22627
rect 20904 22584 20956 22593
rect 20996 22627 21048 22636
rect 20996 22593 21005 22627
rect 21005 22593 21039 22627
rect 21039 22593 21048 22627
rect 24584 22652 24636 22704
rect 20996 22584 21048 22593
rect 23020 22584 23072 22636
rect 24124 22627 24176 22636
rect 24124 22593 24158 22627
rect 24158 22593 24176 22627
rect 24124 22584 24176 22593
rect 17500 22559 17552 22568
rect 17500 22525 17509 22559
rect 17509 22525 17543 22559
rect 17543 22525 17552 22559
rect 17500 22516 17552 22525
rect 21916 22516 21968 22568
rect 23480 22516 23532 22568
rect 16764 22448 16816 22500
rect 16396 22380 16448 22432
rect 20076 22380 20128 22432
rect 23388 22423 23440 22432
rect 23388 22389 23397 22423
rect 23397 22389 23431 22423
rect 23431 22389 23440 22423
rect 25228 22720 25280 22772
rect 26608 22763 26660 22772
rect 26608 22729 26617 22763
rect 26617 22729 26651 22763
rect 26651 22729 26660 22763
rect 26608 22720 26660 22729
rect 26884 22720 26936 22772
rect 24952 22652 25004 22704
rect 25136 22652 25188 22704
rect 25412 22584 25464 22636
rect 26700 22652 26752 22704
rect 29000 22652 29052 22704
rect 30472 22720 30524 22772
rect 31392 22763 31444 22772
rect 29276 22652 29328 22704
rect 30840 22652 30892 22704
rect 31392 22729 31401 22763
rect 31401 22729 31435 22763
rect 31435 22729 31444 22763
rect 31392 22720 31444 22729
rect 27252 22584 27304 22636
rect 27528 22584 27580 22636
rect 28908 22627 28960 22636
rect 28908 22593 28917 22627
rect 28917 22593 28951 22627
rect 28951 22593 28960 22627
rect 28908 22584 28960 22593
rect 25596 22516 25648 22568
rect 30104 22584 30156 22636
rect 32312 22627 32364 22636
rect 32312 22593 32321 22627
rect 32321 22593 32355 22627
rect 32355 22593 32364 22627
rect 32312 22584 32364 22593
rect 33140 22584 33192 22636
rect 34244 22763 34296 22772
rect 34244 22729 34253 22763
rect 34253 22729 34287 22763
rect 34287 22729 34296 22763
rect 34244 22720 34296 22729
rect 34336 22627 34388 22636
rect 34336 22593 34345 22627
rect 34345 22593 34379 22627
rect 34379 22593 34388 22627
rect 34336 22584 34388 22593
rect 25320 22448 25372 22500
rect 29736 22516 29788 22568
rect 29920 22448 29972 22500
rect 31300 22448 31352 22500
rect 25228 22423 25280 22432
rect 23388 22380 23440 22389
rect 25228 22389 25237 22423
rect 25237 22389 25271 22423
rect 25271 22389 25280 22423
rect 25228 22380 25280 22389
rect 27804 22380 27856 22432
rect 28724 22423 28776 22432
rect 28724 22389 28733 22423
rect 28733 22389 28767 22423
rect 28767 22389 28776 22423
rect 28724 22380 28776 22389
rect 5170 22278 5222 22330
rect 5234 22278 5286 22330
rect 5298 22278 5350 22330
rect 5362 22278 5414 22330
rect 5426 22278 5478 22330
rect 13611 22278 13663 22330
rect 13675 22278 13727 22330
rect 13739 22278 13791 22330
rect 13803 22278 13855 22330
rect 13867 22278 13919 22330
rect 22052 22278 22104 22330
rect 22116 22278 22168 22330
rect 22180 22278 22232 22330
rect 22244 22278 22296 22330
rect 22308 22278 22360 22330
rect 30493 22278 30545 22330
rect 30557 22278 30609 22330
rect 30621 22278 30673 22330
rect 30685 22278 30737 22330
rect 30749 22278 30801 22330
rect 21824 22176 21876 22228
rect 24400 22176 24452 22228
rect 28816 22219 28868 22228
rect 28816 22185 28825 22219
rect 28825 22185 28859 22219
rect 28859 22185 28868 22219
rect 28816 22176 28868 22185
rect 16580 22108 16632 22160
rect 18696 22151 18748 22160
rect 16488 22083 16540 22092
rect 16488 22049 16497 22083
rect 16497 22049 16531 22083
rect 16531 22049 16540 22083
rect 16488 22040 16540 22049
rect 17316 22083 17368 22092
rect 17316 22049 17325 22083
rect 17325 22049 17359 22083
rect 17359 22049 17368 22083
rect 17316 22040 17368 22049
rect 16672 21972 16724 22024
rect 18696 22117 18705 22151
rect 18705 22117 18739 22151
rect 18739 22117 18748 22151
rect 18696 22108 18748 22117
rect 20352 22083 20404 22092
rect 20352 22049 20361 22083
rect 20361 22049 20395 22083
rect 20395 22049 20404 22083
rect 20352 22040 20404 22049
rect 23112 22108 23164 22160
rect 18604 22015 18656 22024
rect 18604 21981 18613 22015
rect 18613 21981 18647 22015
rect 18647 21981 18656 22015
rect 18604 21972 18656 21981
rect 19064 21972 19116 22024
rect 17500 21904 17552 21956
rect 18972 21904 19024 21956
rect 21088 22040 21140 22092
rect 22008 22040 22060 22092
rect 20720 21972 20772 22024
rect 21180 21972 21232 22024
rect 21364 21972 21416 22024
rect 21456 21972 21508 22024
rect 23572 22040 23624 22092
rect 23940 22108 23992 22160
rect 24032 22083 24084 22092
rect 22744 22015 22796 22024
rect 20812 21904 20864 21956
rect 20996 21904 21048 21956
rect 22744 21981 22753 22015
rect 22753 21981 22787 22015
rect 22787 21981 22796 22015
rect 22744 21972 22796 21981
rect 22836 21972 22888 22024
rect 24032 22049 24041 22083
rect 24041 22049 24075 22083
rect 24075 22049 24084 22083
rect 24032 22040 24084 22049
rect 24400 22040 24452 22092
rect 27252 22108 27304 22160
rect 28356 22108 28408 22160
rect 29644 22108 29696 22160
rect 24768 22015 24820 22024
rect 24768 21981 24777 22015
rect 24777 21981 24811 22015
rect 24811 21981 24820 22015
rect 24768 21972 24820 21981
rect 25044 22015 25096 22024
rect 25044 21981 25053 22015
rect 25053 21981 25087 22015
rect 25087 21981 25096 22015
rect 25044 21972 25096 21981
rect 28448 22040 28500 22092
rect 30104 22176 30156 22228
rect 31024 22176 31076 22228
rect 32588 22040 32640 22092
rect 27068 21972 27120 22024
rect 27436 21972 27488 22024
rect 19708 21879 19760 21888
rect 19708 21845 19733 21879
rect 19733 21845 19760 21879
rect 19708 21836 19760 21845
rect 20536 21836 20588 21888
rect 21180 21836 21232 21888
rect 21732 21836 21784 21888
rect 22468 21904 22520 21956
rect 22560 21904 22612 21956
rect 23020 21947 23072 21956
rect 23020 21913 23029 21947
rect 23029 21913 23063 21947
rect 23063 21913 23072 21947
rect 23020 21904 23072 21913
rect 25688 21904 25740 21956
rect 26884 21904 26936 21956
rect 27252 21904 27304 21956
rect 27804 22015 27856 22024
rect 27804 21981 27813 22015
rect 27813 21981 27847 22015
rect 27847 21981 27856 22015
rect 27804 21972 27856 21981
rect 28080 21972 28132 22024
rect 29184 21972 29236 22024
rect 31760 22015 31812 22024
rect 31760 21981 31769 22015
rect 31769 21981 31803 22015
rect 31803 21981 31812 22015
rect 31944 22015 31996 22024
rect 31760 21972 31812 21981
rect 31944 21981 31953 22015
rect 31953 21981 31987 22015
rect 31987 21981 31996 22015
rect 31944 21972 31996 21981
rect 32404 21972 32456 22024
rect 32772 22015 32824 22024
rect 32772 21981 32781 22015
rect 32781 21981 32815 22015
rect 32815 21981 32824 22015
rect 32772 21972 32824 21981
rect 27896 21904 27948 21956
rect 22192 21836 22244 21888
rect 22376 21836 22428 21888
rect 23296 21879 23348 21888
rect 23296 21845 23305 21879
rect 23305 21845 23339 21879
rect 23339 21845 23348 21879
rect 23296 21836 23348 21845
rect 24032 21879 24084 21888
rect 24032 21845 24041 21879
rect 24041 21845 24075 21879
rect 24075 21845 24084 21879
rect 24032 21836 24084 21845
rect 25780 21836 25832 21888
rect 27344 21879 27396 21888
rect 27344 21845 27353 21879
rect 27353 21845 27387 21879
rect 27387 21845 27396 21879
rect 27344 21836 27396 21845
rect 27988 21836 28040 21888
rect 29000 21879 29052 21888
rect 29000 21845 29009 21879
rect 29009 21845 29043 21879
rect 29043 21845 29052 21879
rect 29000 21836 29052 21845
rect 30288 21836 30340 21888
rect 32404 21836 32456 21888
rect 9390 21734 9442 21786
rect 9454 21734 9506 21786
rect 9518 21734 9570 21786
rect 9582 21734 9634 21786
rect 9646 21734 9698 21786
rect 17831 21734 17883 21786
rect 17895 21734 17947 21786
rect 17959 21734 18011 21786
rect 18023 21734 18075 21786
rect 18087 21734 18139 21786
rect 26272 21734 26324 21786
rect 26336 21734 26388 21786
rect 26400 21734 26452 21786
rect 26464 21734 26516 21786
rect 26528 21734 26580 21786
rect 34713 21734 34765 21786
rect 34777 21734 34829 21786
rect 34841 21734 34893 21786
rect 34905 21734 34957 21786
rect 34969 21734 35021 21786
rect 17132 21675 17184 21684
rect 17132 21641 17141 21675
rect 17141 21641 17175 21675
rect 17175 21641 17184 21675
rect 17132 21632 17184 21641
rect 17316 21632 17368 21684
rect 19800 21632 19852 21684
rect 21180 21632 21232 21684
rect 21456 21675 21508 21684
rect 21456 21641 21465 21675
rect 21465 21641 21499 21675
rect 21499 21641 21508 21675
rect 21456 21632 21508 21641
rect 23204 21632 23256 21684
rect 27160 21632 27212 21684
rect 33048 21632 33100 21684
rect 16120 21564 16172 21616
rect 20260 21564 20312 21616
rect 21548 21564 21600 21616
rect 25044 21564 25096 21616
rect 16028 21539 16080 21548
rect 16028 21505 16037 21539
rect 16037 21505 16071 21539
rect 16071 21505 16080 21539
rect 16028 21496 16080 21505
rect 17592 21539 17644 21548
rect 17592 21505 17601 21539
rect 17601 21505 17635 21539
rect 17635 21505 17644 21539
rect 17592 21496 17644 21505
rect 18972 21539 19024 21548
rect 18972 21505 19006 21539
rect 19006 21505 19024 21539
rect 18972 21496 19024 21505
rect 15936 21471 15988 21480
rect 15936 21437 15945 21471
rect 15945 21437 15979 21471
rect 15979 21437 15988 21471
rect 15936 21428 15988 21437
rect 16120 21471 16172 21480
rect 16120 21437 16129 21471
rect 16129 21437 16163 21471
rect 16163 21437 16172 21471
rect 16120 21428 16172 21437
rect 16856 21428 16908 21480
rect 17500 21471 17552 21480
rect 17500 21437 17509 21471
rect 17509 21437 17543 21471
rect 17543 21437 17552 21471
rect 17500 21428 17552 21437
rect 16028 21360 16080 21412
rect 16488 21360 16540 21412
rect 17592 21360 17644 21412
rect 16948 21292 17000 21344
rect 19432 21292 19484 21344
rect 20076 21335 20128 21344
rect 20076 21301 20085 21335
rect 20085 21301 20119 21335
rect 20119 21301 20128 21335
rect 20076 21292 20128 21301
rect 20996 21539 21048 21548
rect 20996 21505 21005 21539
rect 21005 21505 21039 21539
rect 21039 21505 21048 21539
rect 20996 21496 21048 21505
rect 21180 21496 21232 21548
rect 21364 21496 21416 21548
rect 22100 21496 22152 21548
rect 21456 21428 21508 21480
rect 22468 21360 22520 21412
rect 23572 21496 23624 21548
rect 25412 21496 25464 21548
rect 25596 21539 25648 21548
rect 25596 21505 25605 21539
rect 25605 21505 25639 21539
rect 25639 21505 25648 21539
rect 25596 21496 25648 21505
rect 26884 21564 26936 21616
rect 27344 21564 27396 21616
rect 27896 21564 27948 21616
rect 28080 21564 28132 21616
rect 29276 21607 29328 21616
rect 29276 21573 29285 21607
rect 29285 21573 29319 21607
rect 29319 21573 29328 21607
rect 29276 21564 29328 21573
rect 23480 21471 23532 21480
rect 23480 21437 23489 21471
rect 23489 21437 23523 21471
rect 23523 21437 23532 21471
rect 23480 21428 23532 21437
rect 27068 21428 27120 21480
rect 23388 21292 23440 21344
rect 24768 21360 24820 21412
rect 23664 21292 23716 21344
rect 25136 21292 25188 21344
rect 26056 21335 26108 21344
rect 26056 21301 26065 21335
rect 26065 21301 26099 21335
rect 26099 21301 26108 21335
rect 26056 21292 26108 21301
rect 26516 21335 26568 21344
rect 26516 21301 26525 21335
rect 26525 21301 26559 21335
rect 26559 21301 26568 21335
rect 26516 21292 26568 21301
rect 26884 21292 26936 21344
rect 27528 21496 27580 21548
rect 28264 21496 28316 21548
rect 28908 21496 28960 21548
rect 30288 21607 30340 21616
rect 30288 21573 30297 21607
rect 30297 21573 30331 21607
rect 30331 21573 30340 21607
rect 30288 21564 30340 21573
rect 31668 21564 31720 21616
rect 31760 21496 31812 21548
rect 32772 21496 32824 21548
rect 33140 21539 33192 21548
rect 33140 21505 33174 21539
rect 33174 21505 33192 21539
rect 33140 21496 33192 21505
rect 29644 21403 29696 21412
rect 29644 21369 29653 21403
rect 29653 21369 29687 21403
rect 29687 21369 29696 21403
rect 29644 21360 29696 21369
rect 30932 21428 30984 21480
rect 31116 21471 31168 21480
rect 31116 21437 31125 21471
rect 31125 21437 31159 21471
rect 31159 21437 31168 21471
rect 31116 21428 31168 21437
rect 27436 21292 27488 21344
rect 29736 21292 29788 21344
rect 31852 21360 31904 21412
rect 30840 21292 30892 21344
rect 31116 21292 31168 21344
rect 31576 21292 31628 21344
rect 33600 21292 33652 21344
rect 5170 21190 5222 21242
rect 5234 21190 5286 21242
rect 5298 21190 5350 21242
rect 5362 21190 5414 21242
rect 5426 21190 5478 21242
rect 13611 21190 13663 21242
rect 13675 21190 13727 21242
rect 13739 21190 13791 21242
rect 13803 21190 13855 21242
rect 13867 21190 13919 21242
rect 22052 21190 22104 21242
rect 22116 21190 22168 21242
rect 22180 21190 22232 21242
rect 22244 21190 22296 21242
rect 22308 21190 22360 21242
rect 30493 21190 30545 21242
rect 30557 21190 30609 21242
rect 30621 21190 30673 21242
rect 30685 21190 30737 21242
rect 30749 21190 30801 21242
rect 15936 21088 15988 21140
rect 16672 21131 16724 21140
rect 16672 21097 16681 21131
rect 16681 21097 16715 21131
rect 16715 21097 16724 21131
rect 16672 21088 16724 21097
rect 19708 21088 19760 21140
rect 22652 21088 22704 21140
rect 23572 21131 23624 21140
rect 23572 21097 23581 21131
rect 23581 21097 23615 21131
rect 23615 21097 23624 21131
rect 23572 21088 23624 21097
rect 16580 20952 16632 21004
rect 18236 20952 18288 21004
rect 16672 20884 16724 20936
rect 17132 20884 17184 20936
rect 18420 20884 18472 20936
rect 25136 21088 25188 21140
rect 29460 21088 29512 21140
rect 18604 20887 18626 20914
rect 18626 20887 18656 20914
rect 18880 20927 18932 20936
rect 18604 20862 18656 20887
rect 18880 20893 18889 20927
rect 18889 20893 18923 20927
rect 18923 20893 18932 20927
rect 18880 20884 18932 20893
rect 18144 20748 18196 20800
rect 19340 20748 19392 20800
rect 19524 20791 19576 20800
rect 19524 20757 19533 20791
rect 19533 20757 19567 20791
rect 19567 20757 19576 20791
rect 19524 20748 19576 20757
rect 20352 20927 20404 20936
rect 20352 20893 20361 20927
rect 20361 20893 20395 20927
rect 20395 20893 20404 20927
rect 20352 20884 20404 20893
rect 20904 20884 20956 20936
rect 21456 20884 21508 20936
rect 21732 20884 21784 20936
rect 19984 20816 20036 20868
rect 22100 20816 22152 20868
rect 23480 20816 23532 20868
rect 24492 21020 24544 21072
rect 24216 20952 24268 21004
rect 24492 20816 24544 20868
rect 25044 20884 25096 20936
rect 28356 20952 28408 21004
rect 28724 20995 28776 21004
rect 28724 20961 28733 20995
rect 28733 20961 28767 20995
rect 28767 20961 28776 20995
rect 28724 20952 28776 20961
rect 29000 20995 29052 21004
rect 29000 20961 29009 20995
rect 29009 20961 29043 20995
rect 29043 20961 29052 20995
rect 29000 20952 29052 20961
rect 29276 21020 29328 21072
rect 29920 21020 29972 21072
rect 30472 20952 30524 21004
rect 31576 21088 31628 21140
rect 28540 20884 28592 20936
rect 29092 20884 29144 20936
rect 29828 20884 29880 20936
rect 30104 20884 30156 20936
rect 32128 21020 32180 21072
rect 30840 20952 30892 21004
rect 31392 20952 31444 21004
rect 31576 20952 31628 21004
rect 32404 20952 32456 21004
rect 31300 20884 31352 20936
rect 32496 20927 32548 20936
rect 24676 20859 24728 20868
rect 24676 20825 24685 20859
rect 24685 20825 24719 20859
rect 24719 20825 24728 20859
rect 24676 20816 24728 20825
rect 26516 20816 26568 20868
rect 27436 20816 27488 20868
rect 30012 20816 30064 20868
rect 32496 20893 32505 20927
rect 32505 20893 32539 20927
rect 32539 20893 32548 20927
rect 32496 20884 32548 20893
rect 25412 20748 25464 20800
rect 25964 20748 26016 20800
rect 26884 20748 26936 20800
rect 27528 20791 27580 20800
rect 27528 20757 27537 20791
rect 27537 20757 27571 20791
rect 27571 20757 27580 20791
rect 27528 20748 27580 20757
rect 31392 20748 31444 20800
rect 34336 20859 34388 20868
rect 34336 20825 34345 20859
rect 34345 20825 34379 20859
rect 34379 20825 34388 20859
rect 34336 20816 34388 20825
rect 31852 20791 31904 20800
rect 31852 20757 31877 20791
rect 31877 20757 31904 20791
rect 31852 20748 31904 20757
rect 32128 20748 32180 20800
rect 32956 20748 33008 20800
rect 9390 20646 9442 20698
rect 9454 20646 9506 20698
rect 9518 20646 9570 20698
rect 9582 20646 9634 20698
rect 9646 20646 9698 20698
rect 17831 20646 17883 20698
rect 17895 20646 17947 20698
rect 17959 20646 18011 20698
rect 18023 20646 18075 20698
rect 18087 20646 18139 20698
rect 26272 20646 26324 20698
rect 26336 20646 26388 20698
rect 26400 20646 26452 20698
rect 26464 20646 26516 20698
rect 26528 20646 26580 20698
rect 34713 20646 34765 20698
rect 34777 20646 34829 20698
rect 34841 20646 34893 20698
rect 34905 20646 34957 20698
rect 34969 20646 35021 20698
rect 16856 20544 16908 20596
rect 18236 20544 18288 20596
rect 20812 20544 20864 20596
rect 21640 20544 21692 20596
rect 23020 20544 23072 20596
rect 23388 20544 23440 20596
rect 24492 20544 24544 20596
rect 25044 20544 25096 20596
rect 25228 20544 25280 20596
rect 26056 20544 26108 20596
rect 26332 20544 26384 20596
rect 26976 20544 27028 20596
rect 30196 20544 30248 20596
rect 16120 20476 16172 20528
rect 16028 20451 16080 20460
rect 16028 20417 16037 20451
rect 16037 20417 16071 20451
rect 16071 20417 16080 20451
rect 16028 20408 16080 20417
rect 16212 20451 16264 20460
rect 16212 20417 16221 20451
rect 16221 20417 16255 20451
rect 16255 20417 16264 20451
rect 16212 20408 16264 20417
rect 16580 20408 16632 20460
rect 17592 20476 17644 20528
rect 19340 20476 19392 20528
rect 22376 20476 22428 20528
rect 22836 20476 22888 20528
rect 26608 20476 26660 20528
rect 19432 20451 19484 20460
rect 19432 20417 19441 20451
rect 19441 20417 19475 20451
rect 19475 20417 19484 20451
rect 19432 20408 19484 20417
rect 16672 20340 16724 20392
rect 19340 20340 19392 20392
rect 16764 20272 16816 20324
rect 17500 20315 17552 20324
rect 17040 20204 17092 20256
rect 17500 20281 17509 20315
rect 17509 20281 17543 20315
rect 17543 20281 17552 20315
rect 17500 20272 17552 20281
rect 18512 20272 18564 20324
rect 20812 20408 20864 20460
rect 21916 20408 21968 20460
rect 22744 20408 22796 20460
rect 23756 20408 23808 20460
rect 25780 20408 25832 20460
rect 25964 20408 26016 20460
rect 26332 20451 26384 20460
rect 26332 20417 26341 20451
rect 26341 20417 26375 20451
rect 26375 20417 26384 20451
rect 26332 20408 26384 20417
rect 26424 20451 26476 20460
rect 26424 20417 26433 20451
rect 26433 20417 26467 20451
rect 26467 20417 26476 20451
rect 27528 20476 27580 20528
rect 29828 20476 29880 20528
rect 32772 20476 32824 20528
rect 26424 20408 26476 20417
rect 27252 20408 27304 20460
rect 28172 20408 28224 20460
rect 28908 20408 28960 20460
rect 29000 20408 29052 20460
rect 31208 20451 31260 20460
rect 31208 20417 31217 20451
rect 31217 20417 31251 20451
rect 31251 20417 31260 20451
rect 31208 20408 31260 20417
rect 31392 20451 31444 20460
rect 31392 20417 31401 20451
rect 31401 20417 31435 20451
rect 31435 20417 31444 20451
rect 31392 20408 31444 20417
rect 32312 20451 32364 20460
rect 32312 20417 32321 20451
rect 32321 20417 32355 20451
rect 32355 20417 32364 20451
rect 32312 20408 32364 20417
rect 33692 20408 33744 20460
rect 34244 20587 34296 20596
rect 34244 20553 34253 20587
rect 34253 20553 34287 20587
rect 34287 20553 34296 20587
rect 34244 20544 34296 20553
rect 34244 20408 34296 20460
rect 21640 20272 21692 20324
rect 23020 20272 23072 20324
rect 21364 20204 21416 20256
rect 23112 20204 23164 20256
rect 23388 20247 23440 20256
rect 23388 20213 23397 20247
rect 23397 20213 23431 20247
rect 23431 20213 23440 20247
rect 23388 20204 23440 20213
rect 26056 20272 26108 20324
rect 26424 20272 26476 20324
rect 28816 20340 28868 20392
rect 28724 20272 28776 20324
rect 28908 20272 28960 20324
rect 29460 20383 29512 20392
rect 29460 20349 29469 20383
rect 29469 20349 29503 20383
rect 29503 20349 29512 20383
rect 30104 20383 30156 20392
rect 29460 20340 29512 20349
rect 30104 20349 30113 20383
rect 30113 20349 30147 20383
rect 30147 20349 30156 20383
rect 30104 20340 30156 20349
rect 31852 20340 31904 20392
rect 31944 20272 31996 20324
rect 26516 20204 26568 20256
rect 28632 20204 28684 20256
rect 31024 20247 31076 20256
rect 31024 20213 31033 20247
rect 31033 20213 31067 20247
rect 31067 20213 31076 20247
rect 31024 20204 31076 20213
rect 33784 20204 33836 20256
rect 5170 20102 5222 20154
rect 5234 20102 5286 20154
rect 5298 20102 5350 20154
rect 5362 20102 5414 20154
rect 5426 20102 5478 20154
rect 13611 20102 13663 20154
rect 13675 20102 13727 20154
rect 13739 20102 13791 20154
rect 13803 20102 13855 20154
rect 13867 20102 13919 20154
rect 22052 20102 22104 20154
rect 22116 20102 22168 20154
rect 22180 20102 22232 20154
rect 22244 20102 22296 20154
rect 22308 20102 22360 20154
rect 30493 20102 30545 20154
rect 30557 20102 30609 20154
rect 30621 20102 30673 20154
rect 30685 20102 30737 20154
rect 30749 20102 30801 20154
rect 1952 19796 2004 19848
rect 2504 19796 2556 19848
rect 18420 20000 18472 20052
rect 16028 19932 16080 19984
rect 21088 20000 21140 20052
rect 22560 20000 22612 20052
rect 27252 20000 27304 20052
rect 31852 20000 31904 20052
rect 31944 20000 31996 20052
rect 33232 20000 33284 20052
rect 21364 19932 21416 19984
rect 16764 19796 16816 19848
rect 16948 19864 17000 19916
rect 19432 19907 19484 19916
rect 17040 19839 17092 19848
rect 17040 19805 17049 19839
rect 17049 19805 17083 19839
rect 17083 19805 17092 19839
rect 17040 19796 17092 19805
rect 17132 19839 17184 19848
rect 17132 19805 17141 19839
rect 17141 19805 17175 19839
rect 17175 19805 17184 19839
rect 17132 19796 17184 19805
rect 19064 19796 19116 19848
rect 19432 19873 19441 19907
rect 19441 19873 19475 19907
rect 19475 19873 19484 19907
rect 19432 19864 19484 19873
rect 20444 19864 20496 19916
rect 22376 19932 22428 19984
rect 21640 19864 21692 19916
rect 20720 19796 20772 19848
rect 21088 19796 21140 19848
rect 21456 19839 21508 19848
rect 21456 19805 21465 19839
rect 21465 19805 21499 19839
rect 21499 19805 21508 19839
rect 21456 19796 21508 19805
rect 21548 19839 21600 19848
rect 21548 19805 21557 19839
rect 21557 19805 21591 19839
rect 21591 19805 21600 19839
rect 21548 19796 21600 19805
rect 21916 19796 21968 19848
rect 23480 19796 23532 19848
rect 23848 19796 23900 19848
rect 26792 19839 26844 19848
rect 26792 19805 26801 19839
rect 26801 19805 26835 19839
rect 26835 19805 26844 19839
rect 26792 19796 26844 19805
rect 27344 19864 27396 19916
rect 29736 19932 29788 19984
rect 33784 19932 33836 19984
rect 18328 19771 18380 19780
rect 18328 19737 18337 19771
rect 18337 19737 18371 19771
rect 18371 19737 18380 19771
rect 18328 19728 18380 19737
rect 1952 19660 2004 19712
rect 16672 19703 16724 19712
rect 16672 19669 16681 19703
rect 16681 19669 16715 19703
rect 16715 19669 16724 19703
rect 16672 19660 16724 19669
rect 18604 19660 18656 19712
rect 19340 19660 19392 19712
rect 20076 19728 20128 19780
rect 22928 19728 22980 19780
rect 23020 19660 23072 19712
rect 23756 19703 23808 19712
rect 23756 19669 23765 19703
rect 23765 19669 23799 19703
rect 23799 19669 23808 19703
rect 23756 19660 23808 19669
rect 24768 19660 24820 19712
rect 25596 19728 25648 19780
rect 27896 19796 27948 19848
rect 29276 19796 29328 19848
rect 29828 19796 29880 19848
rect 25964 19703 26016 19712
rect 25964 19669 25973 19703
rect 25973 19669 26007 19703
rect 26007 19669 26016 19703
rect 25964 19660 26016 19669
rect 28816 19771 28868 19780
rect 28816 19737 28825 19771
rect 28825 19737 28859 19771
rect 28859 19737 28868 19771
rect 28816 19728 28868 19737
rect 28908 19728 28960 19780
rect 30840 19728 30892 19780
rect 33416 19864 33468 19916
rect 31760 19796 31812 19848
rect 34336 19839 34388 19848
rect 27712 19703 27764 19712
rect 27712 19669 27721 19703
rect 27721 19669 27755 19703
rect 27755 19669 27764 19703
rect 27712 19660 27764 19669
rect 27804 19660 27856 19712
rect 29092 19660 29144 19712
rect 30196 19660 30248 19712
rect 31392 19660 31444 19712
rect 32220 19728 32272 19780
rect 34336 19805 34345 19839
rect 34345 19805 34379 19839
rect 34379 19805 34388 19839
rect 34336 19796 34388 19805
rect 32772 19728 32824 19780
rect 32956 19728 33008 19780
rect 33324 19728 33376 19780
rect 33048 19660 33100 19712
rect 9390 19558 9442 19610
rect 9454 19558 9506 19610
rect 9518 19558 9570 19610
rect 9582 19558 9634 19610
rect 9646 19558 9698 19610
rect 17831 19558 17883 19610
rect 17895 19558 17947 19610
rect 17959 19558 18011 19610
rect 18023 19558 18075 19610
rect 18087 19558 18139 19610
rect 26272 19558 26324 19610
rect 26336 19558 26388 19610
rect 26400 19558 26452 19610
rect 26464 19558 26516 19610
rect 26528 19558 26580 19610
rect 34713 19558 34765 19610
rect 34777 19558 34829 19610
rect 34841 19558 34893 19610
rect 34905 19558 34957 19610
rect 34969 19558 35021 19610
rect 1952 19431 2004 19440
rect 1952 19397 1961 19431
rect 1961 19397 1995 19431
rect 1995 19397 2004 19431
rect 1952 19388 2004 19397
rect 15568 19456 15620 19508
rect 16028 19456 16080 19508
rect 18604 19499 18656 19508
rect 18604 19465 18613 19499
rect 18613 19465 18647 19499
rect 18647 19465 18656 19499
rect 18604 19456 18656 19465
rect 20444 19456 20496 19508
rect 21456 19456 21508 19508
rect 22468 19499 22520 19508
rect 16212 19388 16264 19440
rect 22468 19465 22477 19499
rect 22477 19465 22511 19499
rect 22511 19465 22520 19499
rect 22468 19456 22520 19465
rect 22928 19499 22980 19508
rect 22928 19465 22937 19499
rect 22937 19465 22971 19499
rect 22971 19465 22980 19499
rect 22928 19456 22980 19465
rect 23664 19456 23716 19508
rect 24492 19456 24544 19508
rect 25964 19456 26016 19508
rect 26332 19456 26384 19508
rect 30104 19456 30156 19508
rect 31392 19456 31444 19508
rect 1768 19295 1820 19304
rect 1768 19261 1777 19295
rect 1777 19261 1811 19295
rect 1811 19261 1820 19295
rect 1768 19252 1820 19261
rect 2228 19295 2280 19304
rect 2228 19261 2237 19295
rect 2237 19261 2271 19295
rect 2271 19261 2280 19295
rect 2228 19252 2280 19261
rect 15568 19320 15620 19372
rect 16580 19320 16632 19372
rect 16672 19320 16724 19372
rect 18420 19363 18472 19372
rect 18420 19329 18429 19363
rect 18429 19329 18463 19363
rect 18463 19329 18472 19363
rect 18420 19320 18472 19329
rect 19340 19363 19392 19372
rect 19340 19329 19349 19363
rect 19349 19329 19383 19363
rect 19383 19329 19392 19363
rect 19340 19320 19392 19329
rect 20628 19363 20680 19372
rect 20628 19329 20637 19363
rect 20637 19329 20671 19363
rect 20671 19329 20680 19363
rect 20628 19320 20680 19329
rect 20812 19363 20864 19372
rect 20812 19329 20821 19363
rect 20821 19329 20855 19363
rect 20855 19329 20864 19363
rect 20812 19320 20864 19329
rect 23940 19388 23992 19440
rect 24952 19431 25004 19440
rect 24952 19397 24961 19431
rect 24961 19397 24995 19431
rect 24995 19397 25004 19431
rect 24952 19388 25004 19397
rect 25044 19388 25096 19440
rect 16948 19295 17000 19304
rect 16948 19261 16957 19295
rect 16957 19261 16991 19295
rect 16991 19261 17000 19295
rect 16948 19252 17000 19261
rect 18328 19184 18380 19236
rect 18696 19184 18748 19236
rect 22376 19320 22428 19372
rect 23112 19363 23164 19372
rect 23112 19329 23121 19363
rect 23121 19329 23155 19363
rect 23155 19329 23164 19363
rect 23112 19320 23164 19329
rect 23296 19320 23348 19372
rect 24216 19363 24268 19372
rect 24216 19329 24225 19363
rect 24225 19329 24259 19363
rect 24259 19329 24268 19363
rect 24216 19320 24268 19329
rect 24860 19320 24912 19372
rect 26056 19363 26108 19372
rect 26056 19329 26065 19363
rect 26065 19329 26099 19363
rect 26099 19329 26108 19363
rect 26056 19320 26108 19329
rect 26148 19363 26200 19372
rect 26148 19329 26157 19363
rect 26157 19329 26191 19363
rect 26191 19329 26200 19363
rect 26148 19320 26200 19329
rect 26792 19320 26844 19372
rect 27344 19363 27396 19372
rect 27344 19329 27353 19363
rect 27353 19329 27387 19363
rect 27387 19329 27396 19363
rect 27344 19320 27396 19329
rect 21824 19252 21876 19304
rect 23756 19252 23808 19304
rect 25872 19252 25924 19304
rect 21272 19184 21324 19236
rect 23020 19184 23072 19236
rect 25780 19184 25832 19236
rect 18420 19116 18472 19168
rect 20720 19116 20772 19168
rect 22652 19116 22704 19168
rect 23296 19159 23348 19168
rect 23296 19125 23305 19159
rect 23305 19125 23339 19159
rect 23339 19125 23348 19159
rect 23296 19116 23348 19125
rect 25136 19159 25188 19168
rect 25136 19125 25145 19159
rect 25145 19125 25179 19159
rect 25179 19125 25188 19159
rect 25136 19116 25188 19125
rect 25320 19159 25372 19168
rect 25320 19125 25329 19159
rect 25329 19125 25363 19159
rect 25363 19125 25372 19159
rect 25320 19116 25372 19125
rect 26148 19116 26200 19168
rect 27252 19252 27304 19304
rect 26976 19184 27028 19236
rect 27804 19320 27856 19372
rect 27712 19252 27764 19304
rect 29276 19320 29328 19372
rect 29368 19320 29420 19372
rect 28724 19252 28776 19304
rect 28356 19184 28408 19236
rect 29828 19252 29880 19304
rect 32312 19388 32364 19440
rect 31024 19320 31076 19372
rect 31760 19320 31812 19372
rect 32128 19320 32180 19372
rect 31944 19252 31996 19304
rect 32312 19252 32364 19304
rect 34336 19295 34388 19304
rect 34336 19261 34345 19295
rect 34345 19261 34379 19295
rect 34379 19261 34388 19295
rect 34336 19252 34388 19261
rect 27344 19116 27396 19168
rect 29736 19159 29788 19168
rect 29736 19125 29745 19159
rect 29745 19125 29779 19159
rect 29779 19125 29788 19159
rect 29736 19116 29788 19125
rect 30748 19116 30800 19168
rect 31024 19116 31076 19168
rect 31116 19116 31168 19168
rect 31944 19116 31996 19168
rect 5170 19014 5222 19066
rect 5234 19014 5286 19066
rect 5298 19014 5350 19066
rect 5362 19014 5414 19066
rect 5426 19014 5478 19066
rect 13611 19014 13663 19066
rect 13675 19014 13727 19066
rect 13739 19014 13791 19066
rect 13803 19014 13855 19066
rect 13867 19014 13919 19066
rect 22052 19014 22104 19066
rect 22116 19014 22168 19066
rect 22180 19014 22232 19066
rect 22244 19014 22296 19066
rect 22308 19014 22360 19066
rect 30493 19014 30545 19066
rect 30557 19014 30609 19066
rect 30621 19014 30673 19066
rect 30685 19014 30737 19066
rect 30749 19014 30801 19066
rect 1768 18912 1820 18964
rect 16948 18955 17000 18964
rect 16948 18921 16957 18955
rect 16957 18921 16991 18955
rect 16991 18921 17000 18955
rect 16948 18912 17000 18921
rect 16580 18844 16632 18896
rect 2044 18776 2096 18828
rect 2228 18776 2280 18828
rect 1768 18708 1820 18760
rect 16764 18708 16816 18760
rect 17408 18708 17460 18760
rect 18420 18708 18472 18760
rect 18604 18751 18656 18760
rect 18604 18717 18613 18751
rect 18613 18717 18647 18751
rect 18647 18717 18656 18751
rect 18604 18708 18656 18717
rect 19984 18912 20036 18964
rect 20812 18912 20864 18964
rect 21364 18912 21416 18964
rect 22560 18955 22612 18964
rect 22560 18921 22569 18955
rect 22569 18921 22603 18955
rect 22603 18921 22612 18955
rect 22560 18912 22612 18921
rect 22652 18912 22704 18964
rect 25412 18912 25464 18964
rect 28448 18912 28500 18964
rect 29460 18912 29512 18964
rect 30840 18912 30892 18964
rect 33692 18955 33744 18964
rect 33692 18921 33701 18955
rect 33701 18921 33735 18955
rect 33735 18921 33744 18955
rect 33692 18912 33744 18921
rect 21180 18844 21232 18896
rect 23572 18844 23624 18896
rect 23756 18887 23808 18896
rect 23756 18853 23765 18887
rect 23765 18853 23799 18887
rect 23799 18853 23808 18887
rect 23756 18844 23808 18853
rect 24676 18844 24728 18896
rect 27252 18844 27304 18896
rect 19432 18776 19484 18828
rect 18880 18751 18932 18760
rect 18880 18717 18889 18751
rect 18889 18717 18923 18751
rect 18923 18717 18932 18751
rect 18880 18708 18932 18717
rect 20352 18708 20404 18760
rect 24952 18776 25004 18828
rect 20260 18640 20312 18692
rect 21088 18640 21140 18692
rect 21456 18640 21508 18692
rect 22376 18683 22428 18692
rect 22376 18649 22385 18683
rect 22385 18649 22419 18683
rect 22419 18649 22428 18683
rect 22376 18640 22428 18649
rect 18512 18572 18564 18624
rect 21272 18572 21324 18624
rect 21640 18572 21692 18624
rect 22468 18572 22520 18624
rect 25136 18708 25188 18760
rect 26148 18751 26200 18760
rect 24584 18640 24636 18692
rect 26148 18717 26157 18751
rect 26157 18717 26191 18751
rect 26191 18717 26200 18751
rect 26148 18708 26200 18717
rect 26608 18708 26660 18760
rect 27712 18776 27764 18828
rect 26332 18640 26384 18692
rect 27160 18708 27212 18760
rect 27620 18708 27672 18760
rect 28724 18844 28776 18896
rect 32404 18844 32456 18896
rect 28356 18776 28408 18828
rect 28816 18776 28868 18828
rect 29092 18776 29144 18828
rect 28264 18708 28316 18760
rect 29000 18751 29052 18760
rect 29000 18717 29009 18751
rect 29009 18717 29043 18751
rect 29043 18717 29052 18751
rect 29000 18708 29052 18717
rect 26976 18640 27028 18692
rect 28540 18640 28592 18692
rect 29644 18776 29696 18828
rect 30196 18819 30248 18828
rect 30196 18785 30205 18819
rect 30205 18785 30239 18819
rect 30239 18785 30248 18819
rect 30196 18776 30248 18785
rect 32680 18776 32732 18828
rect 24952 18572 25004 18624
rect 27344 18572 27396 18624
rect 28356 18572 28408 18624
rect 31668 18708 31720 18760
rect 31760 18708 31812 18760
rect 33232 18751 33284 18760
rect 33232 18717 33241 18751
rect 33241 18717 33275 18751
rect 33275 18717 33284 18751
rect 33232 18708 33284 18717
rect 30840 18640 30892 18692
rect 30288 18572 30340 18624
rect 33048 18640 33100 18692
rect 33692 18572 33744 18624
rect 9390 18470 9442 18522
rect 9454 18470 9506 18522
rect 9518 18470 9570 18522
rect 9582 18470 9634 18522
rect 9646 18470 9698 18522
rect 17831 18470 17883 18522
rect 17895 18470 17947 18522
rect 17959 18470 18011 18522
rect 18023 18470 18075 18522
rect 18087 18470 18139 18522
rect 26272 18470 26324 18522
rect 26336 18470 26388 18522
rect 26400 18470 26452 18522
rect 26464 18470 26516 18522
rect 26528 18470 26580 18522
rect 34713 18470 34765 18522
rect 34777 18470 34829 18522
rect 34841 18470 34893 18522
rect 34905 18470 34957 18522
rect 34969 18470 35021 18522
rect 17408 18411 17460 18420
rect 17408 18377 17417 18411
rect 17417 18377 17451 18411
rect 17451 18377 17460 18411
rect 17408 18368 17460 18377
rect 18420 18368 18472 18420
rect 19800 18411 19852 18420
rect 19800 18377 19809 18411
rect 19809 18377 19843 18411
rect 19843 18377 19852 18411
rect 19800 18368 19852 18377
rect 20260 18411 20312 18420
rect 20260 18377 20269 18411
rect 20269 18377 20303 18411
rect 20303 18377 20312 18411
rect 20260 18368 20312 18377
rect 21364 18411 21416 18420
rect 1768 18275 1820 18284
rect 1768 18241 1777 18275
rect 1777 18241 1811 18275
rect 1811 18241 1820 18275
rect 1768 18232 1820 18241
rect 17040 18275 17092 18284
rect 17040 18241 17049 18275
rect 17049 18241 17083 18275
rect 17083 18241 17092 18275
rect 17040 18232 17092 18241
rect 19432 18300 19484 18352
rect 18512 18232 18564 18284
rect 21364 18377 21373 18411
rect 21373 18377 21407 18411
rect 21407 18377 21416 18411
rect 21364 18368 21416 18377
rect 24952 18368 25004 18420
rect 26608 18368 26660 18420
rect 27988 18411 28040 18420
rect 21180 18343 21232 18352
rect 21180 18309 21189 18343
rect 21189 18309 21223 18343
rect 21223 18309 21232 18343
rect 21180 18300 21232 18309
rect 27252 18300 27304 18352
rect 27988 18377 27997 18411
rect 27997 18377 28031 18411
rect 28031 18377 28040 18411
rect 27988 18368 28040 18377
rect 31300 18368 31352 18420
rect 29000 18300 29052 18352
rect 1952 18207 2004 18216
rect 1952 18173 1961 18207
rect 1961 18173 1995 18207
rect 1995 18173 2004 18207
rect 1952 18164 2004 18173
rect 2780 18207 2832 18216
rect 2780 18173 2789 18207
rect 2789 18173 2823 18207
rect 2823 18173 2832 18207
rect 2780 18164 2832 18173
rect 17132 18207 17184 18216
rect 17132 18173 17141 18207
rect 17141 18173 17175 18207
rect 17175 18173 17184 18207
rect 17132 18164 17184 18173
rect 21640 18232 21692 18284
rect 22836 18232 22888 18284
rect 23848 18275 23900 18284
rect 23848 18241 23857 18275
rect 23857 18241 23891 18275
rect 23891 18241 23900 18275
rect 23848 18232 23900 18241
rect 23940 18232 23992 18284
rect 24584 18232 24636 18284
rect 25320 18232 25372 18284
rect 27344 18275 27396 18284
rect 27344 18241 27353 18275
rect 27353 18241 27387 18275
rect 27387 18241 27396 18275
rect 27344 18232 27396 18241
rect 27712 18275 27764 18284
rect 20812 18164 20864 18216
rect 21272 18164 21324 18216
rect 21548 18164 21600 18216
rect 21916 18164 21968 18216
rect 25136 18096 25188 18148
rect 27712 18241 27721 18275
rect 27721 18241 27755 18275
rect 27755 18241 27764 18275
rect 27712 18232 27764 18241
rect 28080 18232 28132 18284
rect 28356 18232 28408 18284
rect 30196 18232 30248 18284
rect 30932 18300 30984 18352
rect 31116 18300 31168 18352
rect 32404 18368 32456 18420
rect 27620 18164 27672 18216
rect 28264 18164 28316 18216
rect 28448 18207 28500 18216
rect 28448 18173 28457 18207
rect 28457 18173 28491 18207
rect 28491 18173 28500 18207
rect 28448 18164 28500 18173
rect 30932 18164 30984 18216
rect 31300 18232 31352 18284
rect 32496 18343 32548 18352
rect 32496 18309 32505 18343
rect 32505 18309 32539 18343
rect 32539 18309 32548 18343
rect 32496 18300 32548 18309
rect 31944 18232 31996 18284
rect 32956 18368 33008 18420
rect 33692 18300 33744 18352
rect 32864 18232 32916 18284
rect 31852 18164 31904 18216
rect 33232 18164 33284 18216
rect 33600 18232 33652 18284
rect 22376 18028 22428 18080
rect 26056 18071 26108 18080
rect 26056 18037 26065 18071
rect 26065 18037 26099 18071
rect 26099 18037 26108 18071
rect 26056 18028 26108 18037
rect 28264 18028 28316 18080
rect 31484 18071 31536 18080
rect 31484 18037 31493 18071
rect 31493 18037 31527 18071
rect 31527 18037 31536 18071
rect 31484 18028 31536 18037
rect 31852 18028 31904 18080
rect 33968 18071 34020 18080
rect 33968 18037 33977 18071
rect 33977 18037 34011 18071
rect 34011 18037 34020 18071
rect 33968 18028 34020 18037
rect 5170 17926 5222 17978
rect 5234 17926 5286 17978
rect 5298 17926 5350 17978
rect 5362 17926 5414 17978
rect 5426 17926 5478 17978
rect 13611 17926 13663 17978
rect 13675 17926 13727 17978
rect 13739 17926 13791 17978
rect 13803 17926 13855 17978
rect 13867 17926 13919 17978
rect 22052 17926 22104 17978
rect 22116 17926 22168 17978
rect 22180 17926 22232 17978
rect 22244 17926 22296 17978
rect 22308 17926 22360 17978
rect 30493 17926 30545 17978
rect 30557 17926 30609 17978
rect 30621 17926 30673 17978
rect 30685 17926 30737 17978
rect 30749 17926 30801 17978
rect 1952 17824 2004 17876
rect 20812 17867 20864 17876
rect 20812 17833 20821 17867
rect 20821 17833 20855 17867
rect 20855 17833 20864 17867
rect 20812 17824 20864 17833
rect 26056 17824 26108 17876
rect 28356 17867 28408 17876
rect 28356 17833 28365 17867
rect 28365 17833 28399 17867
rect 28399 17833 28408 17867
rect 28356 17824 28408 17833
rect 28448 17824 28500 17876
rect 29828 17824 29880 17876
rect 31208 17824 31260 17876
rect 19432 17731 19484 17740
rect 19432 17697 19441 17731
rect 19441 17697 19475 17731
rect 19475 17697 19484 17731
rect 19432 17688 19484 17697
rect 2136 17620 2188 17672
rect 21548 17663 21600 17672
rect 21548 17629 21557 17663
rect 21557 17629 21591 17663
rect 21591 17629 21600 17663
rect 21548 17620 21600 17629
rect 23664 17663 23716 17672
rect 23664 17629 23673 17663
rect 23673 17629 23707 17663
rect 23707 17629 23716 17663
rect 23664 17620 23716 17629
rect 19340 17552 19392 17604
rect 21640 17552 21692 17604
rect 22560 17484 22612 17536
rect 23480 17527 23532 17536
rect 23480 17493 23489 17527
rect 23489 17493 23523 17527
rect 23523 17493 23532 17527
rect 23480 17484 23532 17493
rect 27160 17620 27212 17672
rect 28448 17620 28500 17672
rect 29460 17756 29512 17808
rect 29736 17756 29788 17808
rect 30932 17756 30984 17808
rect 31852 17756 31904 17808
rect 31024 17688 31076 17740
rect 34336 17731 34388 17740
rect 34336 17697 34345 17731
rect 34345 17697 34379 17731
rect 34379 17697 34388 17731
rect 34336 17688 34388 17697
rect 25320 17552 25372 17604
rect 26700 17595 26752 17604
rect 26700 17561 26734 17595
rect 26734 17561 26752 17595
rect 26700 17552 26752 17561
rect 28264 17552 28316 17604
rect 28908 17620 28960 17672
rect 24952 17484 25004 17536
rect 25688 17484 25740 17536
rect 26148 17484 26200 17536
rect 27896 17484 27948 17536
rect 31208 17620 31260 17672
rect 31852 17620 31904 17672
rect 32220 17620 32272 17672
rect 29736 17552 29788 17604
rect 33232 17552 33284 17604
rect 30656 17484 30708 17536
rect 32220 17484 32272 17536
rect 32956 17484 33008 17536
rect 9390 17382 9442 17434
rect 9454 17382 9506 17434
rect 9518 17382 9570 17434
rect 9582 17382 9634 17434
rect 9646 17382 9698 17434
rect 17831 17382 17883 17434
rect 17895 17382 17947 17434
rect 17959 17382 18011 17434
rect 18023 17382 18075 17434
rect 18087 17382 18139 17434
rect 26272 17382 26324 17434
rect 26336 17382 26388 17434
rect 26400 17382 26452 17434
rect 26464 17382 26516 17434
rect 26528 17382 26580 17434
rect 34713 17382 34765 17434
rect 34777 17382 34829 17434
rect 34841 17382 34893 17434
rect 34905 17382 34957 17434
rect 34969 17382 35021 17434
rect 19340 17323 19392 17332
rect 19340 17289 19349 17323
rect 19349 17289 19383 17323
rect 19383 17289 19392 17323
rect 19340 17280 19392 17289
rect 19432 17280 19484 17332
rect 21456 17323 21508 17332
rect 21456 17289 21465 17323
rect 21465 17289 21499 17323
rect 21499 17289 21508 17323
rect 21456 17280 21508 17289
rect 19064 17212 19116 17264
rect 19432 17187 19484 17196
rect 1768 17119 1820 17128
rect 1768 17085 1777 17119
rect 1777 17085 1811 17119
rect 1811 17085 1820 17119
rect 1768 17076 1820 17085
rect 2596 17076 2648 17128
rect 2780 17119 2832 17128
rect 2780 17085 2789 17119
rect 2789 17085 2823 17119
rect 2823 17085 2832 17119
rect 2780 17076 2832 17085
rect 19432 17153 19441 17187
rect 19441 17153 19475 17187
rect 19475 17153 19484 17187
rect 19432 17144 19484 17153
rect 20812 17212 20864 17264
rect 21548 17212 21600 17264
rect 20628 17144 20680 17196
rect 22100 17144 22152 17196
rect 22468 17144 22520 17196
rect 23480 17212 23532 17264
rect 25688 17280 25740 17332
rect 26884 17280 26936 17332
rect 29828 17280 29880 17332
rect 30288 17323 30340 17332
rect 30288 17289 30297 17323
rect 30297 17289 30331 17323
rect 30331 17289 30340 17323
rect 30288 17280 30340 17289
rect 30380 17280 30432 17332
rect 25044 17255 25096 17264
rect 25044 17221 25085 17255
rect 25085 17221 25096 17255
rect 25044 17212 25096 17221
rect 25596 17212 25648 17264
rect 26056 17212 26108 17264
rect 28448 17212 28500 17264
rect 30656 17212 30708 17264
rect 32220 17212 32272 17264
rect 26792 17144 26844 17196
rect 27160 17187 27212 17196
rect 27160 17153 27169 17187
rect 27169 17153 27203 17187
rect 27203 17153 27212 17187
rect 27160 17144 27212 17153
rect 29184 17187 29236 17196
rect 29184 17153 29193 17187
rect 29193 17153 29227 17187
rect 29227 17153 29236 17187
rect 29184 17144 29236 17153
rect 29644 17144 29696 17196
rect 22560 17076 22612 17128
rect 25872 17076 25924 17128
rect 26056 17076 26108 17128
rect 21824 16940 21876 16992
rect 22376 16983 22428 16992
rect 22376 16949 22385 16983
rect 22385 16949 22419 16983
rect 22419 16949 22428 16983
rect 22376 16940 22428 16949
rect 24952 16940 25004 16992
rect 25504 17008 25556 17060
rect 25228 16983 25280 16992
rect 25228 16949 25237 16983
rect 25237 16949 25271 16983
rect 25271 16949 25280 16983
rect 25228 16940 25280 16949
rect 26516 16983 26568 16992
rect 26516 16949 26525 16983
rect 26525 16949 26559 16983
rect 26559 16949 26568 16983
rect 26516 16940 26568 16949
rect 28816 17076 28868 17128
rect 29368 17076 29420 17128
rect 30472 17144 30524 17196
rect 30932 17144 30984 17196
rect 30012 17008 30064 17060
rect 27804 16940 27856 16992
rect 29368 16940 29420 16992
rect 30380 17008 30432 17060
rect 30472 16940 30524 16992
rect 31852 17144 31904 17196
rect 32496 17119 32548 17128
rect 32496 17085 32505 17119
rect 32505 17085 32539 17119
rect 32539 17085 32548 17119
rect 32496 17076 32548 17085
rect 34336 17119 34388 17128
rect 34336 17085 34345 17119
rect 34345 17085 34379 17119
rect 34379 17085 34388 17119
rect 34336 17076 34388 17085
rect 32680 17008 32732 17060
rect 33784 16940 33836 16992
rect 5170 16838 5222 16890
rect 5234 16838 5286 16890
rect 5298 16838 5350 16890
rect 5362 16838 5414 16890
rect 5426 16838 5478 16890
rect 13611 16838 13663 16890
rect 13675 16838 13727 16890
rect 13739 16838 13791 16890
rect 13803 16838 13855 16890
rect 13867 16838 13919 16890
rect 22052 16838 22104 16890
rect 22116 16838 22168 16890
rect 22180 16838 22232 16890
rect 22244 16838 22296 16890
rect 22308 16838 22360 16890
rect 30493 16838 30545 16890
rect 30557 16838 30609 16890
rect 30621 16838 30673 16890
rect 30685 16838 30737 16890
rect 30749 16838 30801 16890
rect 1768 16736 1820 16788
rect 2596 16779 2648 16788
rect 2596 16745 2605 16779
rect 2605 16745 2639 16779
rect 2639 16745 2648 16779
rect 2596 16736 2648 16745
rect 20628 16779 20680 16788
rect 20628 16745 20637 16779
rect 20637 16745 20671 16779
rect 20671 16745 20680 16779
rect 20628 16736 20680 16745
rect 21640 16779 21692 16788
rect 21640 16745 21649 16779
rect 21649 16745 21683 16779
rect 21683 16745 21692 16779
rect 21640 16736 21692 16745
rect 22376 16779 22428 16788
rect 22376 16745 22385 16779
rect 22385 16745 22419 16779
rect 22419 16745 22428 16779
rect 22376 16736 22428 16745
rect 20720 16711 20772 16720
rect 20720 16677 20729 16711
rect 20729 16677 20763 16711
rect 20763 16677 20772 16711
rect 20720 16668 20772 16677
rect 24308 16736 24360 16788
rect 24768 16779 24820 16788
rect 24768 16745 24777 16779
rect 24777 16745 24811 16779
rect 24811 16745 24820 16779
rect 24768 16736 24820 16745
rect 27712 16736 27764 16788
rect 28448 16736 28500 16788
rect 28816 16779 28868 16788
rect 28816 16745 28825 16779
rect 28825 16745 28859 16779
rect 28859 16745 28868 16779
rect 28816 16736 28868 16745
rect 29736 16779 29788 16788
rect 29736 16745 29745 16779
rect 29745 16745 29779 16779
rect 29779 16745 29788 16779
rect 29736 16736 29788 16745
rect 29828 16736 29880 16788
rect 19432 16600 19484 16652
rect 2504 16575 2556 16584
rect 2504 16541 2513 16575
rect 2513 16541 2547 16575
rect 2547 16541 2556 16575
rect 2504 16532 2556 16541
rect 22376 16600 22428 16652
rect 22652 16668 22704 16720
rect 21824 16575 21876 16584
rect 21824 16541 21833 16575
rect 21833 16541 21867 16575
rect 21867 16541 21876 16575
rect 21824 16532 21876 16541
rect 22468 16532 22520 16584
rect 23388 16600 23440 16652
rect 23756 16668 23808 16720
rect 24400 16600 24452 16652
rect 27160 16668 27212 16720
rect 29368 16668 29420 16720
rect 25228 16600 25280 16652
rect 24584 16575 24636 16584
rect 21916 16464 21968 16516
rect 22192 16464 22244 16516
rect 21732 16396 21784 16448
rect 24584 16541 24593 16575
rect 24593 16541 24627 16575
rect 24627 16541 24636 16575
rect 24584 16532 24636 16541
rect 24768 16532 24820 16584
rect 25136 16532 25188 16584
rect 25504 16575 25556 16584
rect 25504 16541 25513 16575
rect 25513 16541 25547 16575
rect 25547 16541 25556 16575
rect 25504 16532 25556 16541
rect 25596 16575 25648 16584
rect 25596 16541 25605 16575
rect 25605 16541 25639 16575
rect 25639 16541 25648 16575
rect 26148 16575 26200 16584
rect 25596 16532 25648 16541
rect 26148 16541 26157 16575
rect 26157 16541 26191 16575
rect 26191 16541 26200 16575
rect 26148 16532 26200 16541
rect 28172 16600 28224 16652
rect 30472 16668 30524 16720
rect 27804 16532 27856 16584
rect 28448 16575 28500 16584
rect 28448 16541 28457 16575
rect 28457 16541 28491 16575
rect 28491 16541 28500 16575
rect 28448 16532 28500 16541
rect 30012 16575 30064 16584
rect 30012 16541 30021 16575
rect 30021 16541 30055 16575
rect 30055 16541 30064 16575
rect 30012 16532 30064 16541
rect 32864 16600 32916 16652
rect 31208 16532 31260 16584
rect 31760 16575 31812 16584
rect 31760 16541 31769 16575
rect 31769 16541 31803 16575
rect 31803 16541 31812 16575
rect 31760 16532 31812 16541
rect 23020 16396 23072 16448
rect 23848 16396 23900 16448
rect 24308 16396 24360 16448
rect 24676 16396 24728 16448
rect 24952 16464 25004 16516
rect 25688 16464 25740 16516
rect 29092 16464 29144 16516
rect 29552 16464 29604 16516
rect 30380 16464 30432 16516
rect 30472 16464 30524 16516
rect 32220 16464 32272 16516
rect 32680 16507 32732 16516
rect 32680 16473 32689 16507
rect 32689 16473 32723 16507
rect 32723 16473 32732 16507
rect 32680 16464 32732 16473
rect 35164 16464 35216 16516
rect 25412 16439 25464 16448
rect 25412 16405 25427 16439
rect 25427 16405 25461 16439
rect 25461 16405 25464 16439
rect 25412 16396 25464 16405
rect 26516 16439 26568 16448
rect 26516 16405 26525 16439
rect 26525 16405 26559 16439
rect 26559 16405 26568 16439
rect 26516 16396 26568 16405
rect 26884 16396 26936 16448
rect 28540 16396 28592 16448
rect 29460 16396 29512 16448
rect 30012 16396 30064 16448
rect 9390 16294 9442 16346
rect 9454 16294 9506 16346
rect 9518 16294 9570 16346
rect 9582 16294 9634 16346
rect 9646 16294 9698 16346
rect 17831 16294 17883 16346
rect 17895 16294 17947 16346
rect 17959 16294 18011 16346
rect 18023 16294 18075 16346
rect 18087 16294 18139 16346
rect 26272 16294 26324 16346
rect 26336 16294 26388 16346
rect 26400 16294 26452 16346
rect 26464 16294 26516 16346
rect 26528 16294 26580 16346
rect 34713 16294 34765 16346
rect 34777 16294 34829 16346
rect 34841 16294 34893 16346
rect 34905 16294 34957 16346
rect 34969 16294 35021 16346
rect 22376 16235 22428 16244
rect 22376 16201 22385 16235
rect 22385 16201 22419 16235
rect 22419 16201 22428 16235
rect 22376 16192 22428 16201
rect 22744 16192 22796 16244
rect 24032 16192 24084 16244
rect 24492 16235 24544 16244
rect 24492 16201 24501 16235
rect 24501 16201 24535 16235
rect 24535 16201 24544 16235
rect 24492 16192 24544 16201
rect 25320 16235 25372 16244
rect 25320 16201 25329 16235
rect 25329 16201 25363 16235
rect 25363 16201 25372 16235
rect 25320 16192 25372 16201
rect 28908 16192 28960 16244
rect 30748 16192 30800 16244
rect 31484 16235 31536 16244
rect 31484 16201 31493 16235
rect 31493 16201 31527 16235
rect 31527 16201 31536 16235
rect 31484 16192 31536 16201
rect 32404 16235 32456 16244
rect 32404 16201 32413 16235
rect 32413 16201 32447 16235
rect 32447 16201 32456 16235
rect 32404 16192 32456 16201
rect 33508 16192 33560 16244
rect 34520 16192 34572 16244
rect 22100 16099 22152 16108
rect 22100 16065 22109 16099
rect 22109 16065 22143 16099
rect 22143 16065 22152 16099
rect 22100 16056 22152 16065
rect 23572 16124 23624 16176
rect 25504 16124 25556 16176
rect 22192 16031 22244 16040
rect 22192 15997 22201 16031
rect 22201 15997 22235 16031
rect 22235 15997 22244 16031
rect 22192 15988 22244 15997
rect 22652 15988 22704 16040
rect 20536 15920 20588 15972
rect 24032 16056 24084 16108
rect 23664 15963 23716 15972
rect 23664 15929 23673 15963
rect 23673 15929 23707 15963
rect 23707 15929 23716 15963
rect 23664 15920 23716 15929
rect 1584 15852 1636 15904
rect 22100 15852 22152 15904
rect 22560 15852 22612 15904
rect 25228 16056 25280 16108
rect 25412 16099 25464 16108
rect 25412 16065 25421 16099
rect 25421 16065 25455 16099
rect 25455 16065 25464 16099
rect 25412 16056 25464 16065
rect 26148 16056 26200 16108
rect 28264 16124 28316 16176
rect 28816 16124 28868 16176
rect 29276 16167 29328 16176
rect 29276 16133 29285 16167
rect 29285 16133 29319 16167
rect 29319 16133 29328 16167
rect 29276 16124 29328 16133
rect 29460 16124 29512 16176
rect 28172 16056 28224 16108
rect 28356 16099 28408 16108
rect 28356 16065 28365 16099
rect 28365 16065 28399 16099
rect 28399 16065 28408 16099
rect 28356 16056 28408 16065
rect 28724 16056 28776 16108
rect 29092 16056 29144 16108
rect 25596 16031 25648 16040
rect 25596 15997 25605 16031
rect 25605 15997 25639 16031
rect 25639 15997 25648 16031
rect 25596 15988 25648 15997
rect 27160 15988 27212 16040
rect 28632 15988 28684 16040
rect 29368 16099 29420 16108
rect 29368 16065 29377 16099
rect 29377 16065 29411 16099
rect 29411 16065 29420 16099
rect 29828 16099 29880 16108
rect 29368 16056 29420 16065
rect 29828 16065 29837 16099
rect 29837 16065 29871 16099
rect 29871 16065 29880 16099
rect 29828 16056 29880 16065
rect 30196 16124 30248 16176
rect 30472 16099 30524 16108
rect 30472 16065 30481 16099
rect 30481 16065 30515 16099
rect 30515 16065 30524 16099
rect 30472 16056 30524 16065
rect 30656 16099 30708 16108
rect 30656 16065 30665 16099
rect 30665 16065 30699 16099
rect 30699 16065 30708 16099
rect 30656 16056 30708 16065
rect 31944 16124 31996 16176
rect 32956 16099 33008 16108
rect 24952 15852 25004 15904
rect 25596 15852 25648 15904
rect 26608 15852 26660 15904
rect 28448 15852 28500 15904
rect 29552 15988 29604 16040
rect 31116 15988 31168 16040
rect 32956 16065 32965 16099
rect 32965 16065 32999 16099
rect 32999 16065 33008 16099
rect 32956 16056 33008 16065
rect 33324 16056 33376 16108
rect 29092 15920 29144 15972
rect 31208 15920 31260 15972
rect 32680 15920 32732 15972
rect 29000 15852 29052 15904
rect 5170 15750 5222 15802
rect 5234 15750 5286 15802
rect 5298 15750 5350 15802
rect 5362 15750 5414 15802
rect 5426 15750 5478 15802
rect 13611 15750 13663 15802
rect 13675 15750 13727 15802
rect 13739 15750 13791 15802
rect 13803 15750 13855 15802
rect 13867 15750 13919 15802
rect 22052 15750 22104 15802
rect 22116 15750 22168 15802
rect 22180 15750 22232 15802
rect 22244 15750 22296 15802
rect 22308 15750 22360 15802
rect 30493 15750 30545 15802
rect 30557 15750 30609 15802
rect 30621 15750 30673 15802
rect 30685 15750 30737 15802
rect 30749 15750 30801 15802
rect 22836 15648 22888 15700
rect 23940 15648 23992 15700
rect 24124 15648 24176 15700
rect 26792 15648 26844 15700
rect 26976 15648 27028 15700
rect 29184 15648 29236 15700
rect 30840 15648 30892 15700
rect 31576 15648 31628 15700
rect 32036 15691 32088 15700
rect 32036 15657 32045 15691
rect 32045 15657 32079 15691
rect 32079 15657 32088 15691
rect 32036 15648 32088 15657
rect 33140 15648 33192 15700
rect 34060 15648 34112 15700
rect 23112 15580 23164 15632
rect 26424 15580 26476 15632
rect 31300 15580 31352 15632
rect 31852 15580 31904 15632
rect 32680 15580 32732 15632
rect 1584 15555 1636 15564
rect 1584 15521 1593 15555
rect 1593 15521 1627 15555
rect 1627 15521 1636 15555
rect 1584 15512 1636 15521
rect 2780 15555 2832 15564
rect 2780 15521 2789 15555
rect 2789 15521 2823 15555
rect 2823 15521 2832 15555
rect 2780 15512 2832 15521
rect 24216 15512 24268 15564
rect 23020 15487 23072 15496
rect 23020 15453 23029 15487
rect 23029 15453 23063 15487
rect 23063 15453 23072 15487
rect 23020 15444 23072 15453
rect 23296 15444 23348 15496
rect 23848 15487 23900 15496
rect 23848 15453 23857 15487
rect 23857 15453 23891 15487
rect 23891 15453 23900 15487
rect 23848 15444 23900 15453
rect 24032 15487 24084 15496
rect 24032 15453 24041 15487
rect 24041 15453 24075 15487
rect 24075 15453 24084 15487
rect 24032 15444 24084 15453
rect 25044 15444 25096 15496
rect 1768 15419 1820 15428
rect 1768 15385 1777 15419
rect 1777 15385 1811 15419
rect 1811 15385 1820 15419
rect 1768 15376 1820 15385
rect 25688 15512 25740 15564
rect 25872 15444 25924 15496
rect 26884 15487 26936 15496
rect 25596 15376 25648 15428
rect 26424 15376 26476 15428
rect 25412 15308 25464 15360
rect 26516 15308 26568 15360
rect 26884 15453 26893 15487
rect 26893 15453 26927 15487
rect 26927 15453 26936 15487
rect 26884 15444 26936 15453
rect 27804 15376 27856 15428
rect 28448 15487 28500 15496
rect 28448 15453 28457 15487
rect 28457 15453 28491 15487
rect 28491 15453 28500 15487
rect 28448 15444 28500 15453
rect 28632 15444 28684 15496
rect 29828 15444 29880 15496
rect 30380 15444 30432 15496
rect 30840 15487 30892 15496
rect 30840 15453 30849 15487
rect 30849 15453 30883 15487
rect 30883 15453 30892 15487
rect 30840 15444 30892 15453
rect 32312 15512 32364 15564
rect 31668 15444 31720 15496
rect 33968 15512 34020 15564
rect 32680 15444 32732 15496
rect 33784 15487 33836 15496
rect 33784 15453 33793 15487
rect 33793 15453 33827 15487
rect 33827 15453 33836 15487
rect 33784 15444 33836 15453
rect 34244 15376 34296 15428
rect 28356 15308 28408 15360
rect 9390 15206 9442 15258
rect 9454 15206 9506 15258
rect 9518 15206 9570 15258
rect 9582 15206 9634 15258
rect 9646 15206 9698 15258
rect 17831 15206 17883 15258
rect 17895 15206 17947 15258
rect 17959 15206 18011 15258
rect 18023 15206 18075 15258
rect 18087 15206 18139 15258
rect 26272 15206 26324 15258
rect 26336 15206 26388 15258
rect 26400 15206 26452 15258
rect 26464 15206 26516 15258
rect 26528 15206 26580 15258
rect 34713 15206 34765 15258
rect 34777 15206 34829 15258
rect 34841 15206 34893 15258
rect 34905 15206 34957 15258
rect 34969 15206 35021 15258
rect 1768 15104 1820 15156
rect 24860 15147 24912 15156
rect 24860 15113 24869 15147
rect 24869 15113 24903 15147
rect 24903 15113 24912 15147
rect 24860 15104 24912 15113
rect 25596 15147 25648 15156
rect 25596 15113 25605 15147
rect 25605 15113 25639 15147
rect 25639 15113 25648 15147
rect 25596 15104 25648 15113
rect 27068 15104 27120 15156
rect 27252 15147 27304 15156
rect 27252 15113 27261 15147
rect 27261 15113 27295 15147
rect 27295 15113 27304 15147
rect 27252 15104 27304 15113
rect 28080 15147 28132 15156
rect 28080 15113 28089 15147
rect 28089 15113 28123 15147
rect 28123 15113 28132 15147
rect 28080 15104 28132 15113
rect 29368 15147 29420 15156
rect 29368 15113 29377 15147
rect 29377 15113 29411 15147
rect 29411 15113 29420 15147
rect 29368 15104 29420 15113
rect 30288 15104 30340 15156
rect 32772 15104 32824 15156
rect 33048 15147 33100 15156
rect 33048 15113 33057 15147
rect 33057 15113 33091 15147
rect 33091 15113 33100 15147
rect 33048 15104 33100 15113
rect 29828 15036 29880 15088
rect 30104 15036 30156 15088
rect 2872 14968 2924 15020
rect 22008 14968 22060 15020
rect 24768 15011 24820 15020
rect 24768 14977 24777 15011
rect 24777 14977 24811 15011
rect 24811 14977 24820 15011
rect 24768 14968 24820 14977
rect 25412 15011 25464 15020
rect 25412 14977 25421 15011
rect 25421 14977 25455 15011
rect 25455 14977 25464 15011
rect 25412 14968 25464 14977
rect 25596 15011 25648 15020
rect 25596 14977 25605 15011
rect 25605 14977 25639 15011
rect 25639 14977 25648 15011
rect 25596 14968 25648 14977
rect 25780 14968 25832 15020
rect 26148 14968 26200 15020
rect 27804 14968 27856 15020
rect 28172 14968 28224 15020
rect 28816 15011 28868 15020
rect 28816 14977 28825 15011
rect 28825 14977 28859 15011
rect 28859 14977 28868 15011
rect 28816 14968 28868 14977
rect 15292 14900 15344 14952
rect 29000 14900 29052 14952
rect 30932 14968 30984 15020
rect 31668 14968 31720 15020
rect 32772 14968 32824 15020
rect 33600 14968 33652 15020
rect 33784 15011 33836 15020
rect 33784 14977 33793 15011
rect 33793 14977 33827 15011
rect 33827 14977 33836 15011
rect 33784 14968 33836 14977
rect 32128 14900 32180 14952
rect 1768 14764 1820 14816
rect 5170 14662 5222 14714
rect 5234 14662 5286 14714
rect 5298 14662 5350 14714
rect 5362 14662 5414 14714
rect 5426 14662 5478 14714
rect 13611 14662 13663 14714
rect 13675 14662 13727 14714
rect 13739 14662 13791 14714
rect 13803 14662 13855 14714
rect 13867 14662 13919 14714
rect 22052 14662 22104 14714
rect 22116 14662 22168 14714
rect 22180 14662 22232 14714
rect 22244 14662 22296 14714
rect 22308 14662 22360 14714
rect 30493 14662 30545 14714
rect 30557 14662 30609 14714
rect 30621 14662 30673 14714
rect 30685 14662 30737 14714
rect 30749 14662 30801 14714
rect 26700 14560 26752 14612
rect 31024 14603 31076 14612
rect 31024 14569 31033 14603
rect 31033 14569 31067 14603
rect 31067 14569 31076 14603
rect 31024 14560 31076 14569
rect 32496 14560 32548 14612
rect 27436 14492 27488 14544
rect 1768 14467 1820 14476
rect 1768 14433 1777 14467
rect 1777 14433 1811 14467
rect 1811 14433 1820 14467
rect 1768 14424 1820 14433
rect 2780 14467 2832 14476
rect 2780 14433 2789 14467
rect 2789 14433 2823 14467
rect 2823 14433 2832 14467
rect 2780 14424 2832 14433
rect 1584 14399 1636 14408
rect 1584 14365 1593 14399
rect 1593 14365 1627 14399
rect 1627 14365 1636 14399
rect 1584 14356 1636 14365
rect 25504 14356 25556 14408
rect 25964 14399 26016 14408
rect 25964 14365 25973 14399
rect 25973 14365 26007 14399
rect 26007 14365 26016 14399
rect 25964 14356 26016 14365
rect 26608 14399 26660 14408
rect 26608 14365 26617 14399
rect 26617 14365 26651 14399
rect 26651 14365 26660 14399
rect 26608 14356 26660 14365
rect 26884 14356 26936 14408
rect 34336 14399 34388 14408
rect 26056 14288 26108 14340
rect 34336 14365 34345 14399
rect 34345 14365 34379 14399
rect 34379 14365 34388 14399
rect 34336 14356 34388 14365
rect 32680 14331 32732 14340
rect 32680 14297 32689 14331
rect 32689 14297 32723 14331
rect 32723 14297 32732 14331
rect 32680 14288 32732 14297
rect 33508 14220 33560 14272
rect 9390 14118 9442 14170
rect 9454 14118 9506 14170
rect 9518 14118 9570 14170
rect 9582 14118 9634 14170
rect 9646 14118 9698 14170
rect 17831 14118 17883 14170
rect 17895 14118 17947 14170
rect 17959 14118 18011 14170
rect 18023 14118 18075 14170
rect 18087 14118 18139 14170
rect 26272 14118 26324 14170
rect 26336 14118 26388 14170
rect 26400 14118 26452 14170
rect 26464 14118 26516 14170
rect 26528 14118 26580 14170
rect 34713 14118 34765 14170
rect 34777 14118 34829 14170
rect 34841 14118 34893 14170
rect 34905 14118 34957 14170
rect 34969 14118 35021 14170
rect 30840 14016 30892 14068
rect 31392 14016 31444 14068
rect 30288 13923 30340 13932
rect 30288 13889 30297 13923
rect 30297 13889 30331 13923
rect 30331 13889 30340 13923
rect 30288 13880 30340 13889
rect 30932 13923 30984 13932
rect 30932 13889 30941 13923
rect 30941 13889 30975 13923
rect 30975 13889 30984 13923
rect 30932 13880 30984 13889
rect 31576 13923 31628 13932
rect 31576 13889 31585 13923
rect 31585 13889 31619 13923
rect 31619 13889 31628 13923
rect 31576 13880 31628 13889
rect 1768 13855 1820 13864
rect 1768 13821 1777 13855
rect 1777 13821 1811 13855
rect 1811 13821 1820 13855
rect 1768 13812 1820 13821
rect 1952 13855 2004 13864
rect 1952 13821 1961 13855
rect 1961 13821 1995 13855
rect 1995 13821 2004 13855
rect 1952 13812 2004 13821
rect 2780 13855 2832 13864
rect 2780 13821 2789 13855
rect 2789 13821 2823 13855
rect 2823 13821 2832 13855
rect 2780 13812 2832 13821
rect 32496 13855 32548 13864
rect 32496 13821 32505 13855
rect 32505 13821 32539 13855
rect 32539 13821 32548 13855
rect 32496 13812 32548 13821
rect 34336 13855 34388 13864
rect 34336 13821 34345 13855
rect 34345 13821 34379 13855
rect 34379 13821 34388 13855
rect 34336 13812 34388 13821
rect 5170 13574 5222 13626
rect 5234 13574 5286 13626
rect 5298 13574 5350 13626
rect 5362 13574 5414 13626
rect 5426 13574 5478 13626
rect 13611 13574 13663 13626
rect 13675 13574 13727 13626
rect 13739 13574 13791 13626
rect 13803 13574 13855 13626
rect 13867 13574 13919 13626
rect 22052 13574 22104 13626
rect 22116 13574 22168 13626
rect 22180 13574 22232 13626
rect 22244 13574 22296 13626
rect 22308 13574 22360 13626
rect 30493 13574 30545 13626
rect 30557 13574 30609 13626
rect 30621 13574 30673 13626
rect 30685 13574 30737 13626
rect 30749 13574 30801 13626
rect 1768 13472 1820 13524
rect 31208 13515 31260 13524
rect 31208 13481 31217 13515
rect 31217 13481 31251 13515
rect 31251 13481 31260 13515
rect 31208 13472 31260 13481
rect 31852 13515 31904 13524
rect 31852 13481 31861 13515
rect 31861 13481 31895 13515
rect 31895 13481 31904 13515
rect 31852 13472 31904 13481
rect 32588 13515 32640 13524
rect 32588 13481 32597 13515
rect 32597 13481 32631 13515
rect 32631 13481 32640 13515
rect 32588 13472 32640 13481
rect 33600 13515 33652 13524
rect 33600 13481 33609 13515
rect 33609 13481 33643 13515
rect 33643 13481 33652 13515
rect 33600 13472 33652 13481
rect 1584 13404 1636 13456
rect 30380 13268 30432 13320
rect 31760 13311 31812 13320
rect 31760 13277 31769 13311
rect 31769 13277 31803 13311
rect 31803 13277 31812 13311
rect 33784 13311 33836 13320
rect 31760 13268 31812 13277
rect 33784 13277 33793 13311
rect 33793 13277 33827 13311
rect 33827 13277 33836 13311
rect 33784 13268 33836 13277
rect 9390 13030 9442 13082
rect 9454 13030 9506 13082
rect 9518 13030 9570 13082
rect 9582 13030 9634 13082
rect 9646 13030 9698 13082
rect 17831 13030 17883 13082
rect 17895 13030 17947 13082
rect 17959 13030 18011 13082
rect 18023 13030 18075 13082
rect 18087 13030 18139 13082
rect 26272 13030 26324 13082
rect 26336 13030 26388 13082
rect 26400 13030 26452 13082
rect 26464 13030 26516 13082
rect 26528 13030 26580 13082
rect 34713 13030 34765 13082
rect 34777 13030 34829 13082
rect 34841 13030 34893 13082
rect 34905 13030 34957 13082
rect 34969 13030 35021 13082
rect 1952 12928 2004 12980
rect 34336 12903 34388 12912
rect 34336 12869 34345 12903
rect 34345 12869 34379 12903
rect 34379 12869 34388 12903
rect 34336 12860 34388 12869
rect 2228 12792 2280 12844
rect 2688 12792 2740 12844
rect 30932 12792 30984 12844
rect 31484 12792 31536 12844
rect 33140 12724 33192 12776
rect 5170 12486 5222 12538
rect 5234 12486 5286 12538
rect 5298 12486 5350 12538
rect 5362 12486 5414 12538
rect 5426 12486 5478 12538
rect 13611 12486 13663 12538
rect 13675 12486 13727 12538
rect 13739 12486 13791 12538
rect 13803 12486 13855 12538
rect 13867 12486 13919 12538
rect 22052 12486 22104 12538
rect 22116 12486 22168 12538
rect 22180 12486 22232 12538
rect 22244 12486 22296 12538
rect 22308 12486 22360 12538
rect 30493 12486 30545 12538
rect 30557 12486 30609 12538
rect 30621 12486 30673 12538
rect 30685 12486 30737 12538
rect 30749 12486 30801 12538
rect 32496 12384 32548 12436
rect 33324 12248 33376 12300
rect 34336 12291 34388 12300
rect 34336 12257 34345 12291
rect 34345 12257 34379 12291
rect 34379 12257 34388 12291
rect 34336 12248 34388 12257
rect 2136 12180 2188 12232
rect 14372 12180 14424 12232
rect 31576 12180 31628 12232
rect 1952 12044 2004 12096
rect 9390 11942 9442 11994
rect 9454 11942 9506 11994
rect 9518 11942 9570 11994
rect 9582 11942 9634 11994
rect 9646 11942 9698 11994
rect 17831 11942 17883 11994
rect 17895 11942 17947 11994
rect 17959 11942 18011 11994
rect 18023 11942 18075 11994
rect 18087 11942 18139 11994
rect 26272 11942 26324 11994
rect 26336 11942 26388 11994
rect 26400 11942 26452 11994
rect 26464 11942 26516 11994
rect 26528 11942 26580 11994
rect 34713 11942 34765 11994
rect 34777 11942 34829 11994
rect 34841 11942 34893 11994
rect 34905 11942 34957 11994
rect 34969 11942 35021 11994
rect 1952 11815 2004 11824
rect 1952 11781 1961 11815
rect 1961 11781 1995 11815
rect 1995 11781 2004 11815
rect 1952 11772 2004 11781
rect 32864 11704 32916 11756
rect 33232 11704 33284 11756
rect 33968 11747 34020 11756
rect 33968 11713 33977 11747
rect 33977 11713 34011 11747
rect 34011 11713 34020 11747
rect 33968 11704 34020 11713
rect 2044 11636 2096 11688
rect 2780 11679 2832 11688
rect 2780 11645 2789 11679
rect 2789 11645 2823 11679
rect 2823 11645 2832 11679
rect 2780 11636 2832 11645
rect 5170 11398 5222 11450
rect 5234 11398 5286 11450
rect 5298 11398 5350 11450
rect 5362 11398 5414 11450
rect 5426 11398 5478 11450
rect 13611 11398 13663 11450
rect 13675 11398 13727 11450
rect 13739 11398 13791 11450
rect 13803 11398 13855 11450
rect 13867 11398 13919 11450
rect 22052 11398 22104 11450
rect 22116 11398 22168 11450
rect 22180 11398 22232 11450
rect 22244 11398 22296 11450
rect 22308 11398 22360 11450
rect 30493 11398 30545 11450
rect 30557 11398 30609 11450
rect 30621 11398 30673 11450
rect 30685 11398 30737 11450
rect 30749 11398 30801 11450
rect 2044 11339 2096 11348
rect 2044 11305 2053 11339
rect 2053 11305 2087 11339
rect 2087 11305 2096 11339
rect 2044 11296 2096 11305
rect 33140 11296 33192 11348
rect 33416 11296 33468 11348
rect 1768 11092 1820 11144
rect 33508 11092 33560 11144
rect 9390 10854 9442 10906
rect 9454 10854 9506 10906
rect 9518 10854 9570 10906
rect 9582 10854 9634 10906
rect 9646 10854 9698 10906
rect 17831 10854 17883 10906
rect 17895 10854 17947 10906
rect 17959 10854 18011 10906
rect 18023 10854 18075 10906
rect 18087 10854 18139 10906
rect 26272 10854 26324 10906
rect 26336 10854 26388 10906
rect 26400 10854 26452 10906
rect 26464 10854 26516 10906
rect 26528 10854 26580 10906
rect 34713 10854 34765 10906
rect 34777 10854 34829 10906
rect 34841 10854 34893 10906
rect 34905 10854 34957 10906
rect 34969 10854 35021 10906
rect 32680 10752 32732 10804
rect 1768 10659 1820 10668
rect 1768 10625 1777 10659
rect 1777 10625 1811 10659
rect 1811 10625 1820 10659
rect 1768 10616 1820 10625
rect 33324 10659 33376 10668
rect 33324 10625 33333 10659
rect 33333 10625 33367 10659
rect 33367 10625 33376 10659
rect 33324 10616 33376 10625
rect 2044 10548 2096 10600
rect 2780 10591 2832 10600
rect 2780 10557 2789 10591
rect 2789 10557 2823 10591
rect 2823 10557 2832 10591
rect 2780 10548 2832 10557
rect 31484 10548 31536 10600
rect 5170 10310 5222 10362
rect 5234 10310 5286 10362
rect 5298 10310 5350 10362
rect 5362 10310 5414 10362
rect 5426 10310 5478 10362
rect 13611 10310 13663 10362
rect 13675 10310 13727 10362
rect 13739 10310 13791 10362
rect 13803 10310 13855 10362
rect 13867 10310 13919 10362
rect 22052 10310 22104 10362
rect 22116 10310 22168 10362
rect 22180 10310 22232 10362
rect 22244 10310 22296 10362
rect 22308 10310 22360 10362
rect 30493 10310 30545 10362
rect 30557 10310 30609 10362
rect 30621 10310 30673 10362
rect 30685 10310 30737 10362
rect 30749 10310 30801 10362
rect 2044 10251 2096 10260
rect 2044 10217 2053 10251
rect 2053 10217 2087 10251
rect 2087 10217 2096 10251
rect 2044 10208 2096 10217
rect 34244 10251 34296 10260
rect 34244 10217 34253 10251
rect 34253 10217 34287 10251
rect 34287 10217 34296 10251
rect 34244 10208 34296 10217
rect 4712 10004 4764 10056
rect 34060 10047 34112 10056
rect 34060 10013 34069 10047
rect 34069 10013 34103 10047
rect 34103 10013 34112 10047
rect 34060 10004 34112 10013
rect 9390 9766 9442 9818
rect 9454 9766 9506 9818
rect 9518 9766 9570 9818
rect 9582 9766 9634 9818
rect 9646 9766 9698 9818
rect 17831 9766 17883 9818
rect 17895 9766 17947 9818
rect 17959 9766 18011 9818
rect 18023 9766 18075 9818
rect 18087 9766 18139 9818
rect 26272 9766 26324 9818
rect 26336 9766 26388 9818
rect 26400 9766 26452 9818
rect 26464 9766 26516 9818
rect 26528 9766 26580 9818
rect 34713 9766 34765 9818
rect 34777 9766 34829 9818
rect 34841 9766 34893 9818
rect 34905 9766 34957 9818
rect 34969 9766 35021 9818
rect 2872 9528 2924 9580
rect 9128 9528 9180 9580
rect 1584 9324 1636 9376
rect 2596 9367 2648 9376
rect 2596 9333 2605 9367
rect 2605 9333 2639 9367
rect 2639 9333 2648 9367
rect 2596 9324 2648 9333
rect 5170 9222 5222 9274
rect 5234 9222 5286 9274
rect 5298 9222 5350 9274
rect 5362 9222 5414 9274
rect 5426 9222 5478 9274
rect 13611 9222 13663 9274
rect 13675 9222 13727 9274
rect 13739 9222 13791 9274
rect 13803 9222 13855 9274
rect 13867 9222 13919 9274
rect 22052 9222 22104 9274
rect 22116 9222 22168 9274
rect 22180 9222 22232 9274
rect 22244 9222 22296 9274
rect 22308 9222 22360 9274
rect 30493 9222 30545 9274
rect 30557 9222 30609 9274
rect 30621 9222 30673 9274
rect 30685 9222 30737 9274
rect 30749 9222 30801 9274
rect 1584 9027 1636 9036
rect 1584 8993 1593 9027
rect 1593 8993 1627 9027
rect 1627 8993 1636 9027
rect 1584 8984 1636 8993
rect 2596 8984 2648 9036
rect 2780 9027 2832 9036
rect 2780 8993 2789 9027
rect 2789 8993 2823 9027
rect 2823 8993 2832 9027
rect 2780 8984 2832 8993
rect 32496 8916 32548 8968
rect 9390 8678 9442 8730
rect 9454 8678 9506 8730
rect 9518 8678 9570 8730
rect 9582 8678 9634 8730
rect 9646 8678 9698 8730
rect 17831 8678 17883 8730
rect 17895 8678 17947 8730
rect 17959 8678 18011 8730
rect 18023 8678 18075 8730
rect 18087 8678 18139 8730
rect 26272 8678 26324 8730
rect 26336 8678 26388 8730
rect 26400 8678 26452 8730
rect 26464 8678 26516 8730
rect 26528 8678 26580 8730
rect 34713 8678 34765 8730
rect 34777 8678 34829 8730
rect 34841 8678 34893 8730
rect 34905 8678 34957 8730
rect 34969 8678 35021 8730
rect 34336 8551 34388 8560
rect 34336 8517 34345 8551
rect 34345 8517 34379 8551
rect 34379 8517 34388 8551
rect 34336 8508 34388 8517
rect 32496 8483 32548 8492
rect 32496 8449 32505 8483
rect 32505 8449 32539 8483
rect 32539 8449 32548 8483
rect 32496 8440 32548 8449
rect 1768 8415 1820 8424
rect 1768 8381 1777 8415
rect 1777 8381 1811 8415
rect 1811 8381 1820 8415
rect 1768 8372 1820 8381
rect 2596 8372 2648 8424
rect 2780 8415 2832 8424
rect 2780 8381 2789 8415
rect 2789 8381 2823 8415
rect 2823 8381 2832 8415
rect 2780 8372 2832 8381
rect 33876 8372 33928 8424
rect 5170 8134 5222 8186
rect 5234 8134 5286 8186
rect 5298 8134 5350 8186
rect 5362 8134 5414 8186
rect 5426 8134 5478 8186
rect 13611 8134 13663 8186
rect 13675 8134 13727 8186
rect 13739 8134 13791 8186
rect 13803 8134 13855 8186
rect 13867 8134 13919 8186
rect 22052 8134 22104 8186
rect 22116 8134 22168 8186
rect 22180 8134 22232 8186
rect 22244 8134 22296 8186
rect 22308 8134 22360 8186
rect 30493 8134 30545 8186
rect 30557 8134 30609 8186
rect 30621 8134 30673 8186
rect 30685 8134 30737 8186
rect 30749 8134 30801 8186
rect 1768 8032 1820 8084
rect 2596 8075 2648 8084
rect 2596 8041 2605 8075
rect 2605 8041 2639 8075
rect 2639 8041 2648 8075
rect 2596 8032 2648 8041
rect 31668 8032 31720 8084
rect 33140 8032 33192 8084
rect 33876 8075 33928 8084
rect 33876 8041 33885 8075
rect 33885 8041 33919 8075
rect 33919 8041 33928 8075
rect 33876 8032 33928 8041
rect 7196 7896 7248 7948
rect 7380 7896 7432 7948
rect 33324 7871 33376 7880
rect 1768 7760 1820 7812
rect 33324 7837 33333 7871
rect 33333 7837 33367 7871
rect 33367 7837 33376 7871
rect 33324 7828 33376 7837
rect 33784 7871 33836 7880
rect 33784 7837 33793 7871
rect 33793 7837 33827 7871
rect 33827 7837 33836 7871
rect 33784 7828 33836 7837
rect 9390 7590 9442 7642
rect 9454 7590 9506 7642
rect 9518 7590 9570 7642
rect 9582 7590 9634 7642
rect 9646 7590 9698 7642
rect 17831 7590 17883 7642
rect 17895 7590 17947 7642
rect 17959 7590 18011 7642
rect 18023 7590 18075 7642
rect 18087 7590 18139 7642
rect 26272 7590 26324 7642
rect 26336 7590 26388 7642
rect 26400 7590 26452 7642
rect 26464 7590 26516 7642
rect 26528 7590 26580 7642
rect 34713 7590 34765 7642
rect 34777 7590 34829 7642
rect 34841 7590 34893 7642
rect 34905 7590 34957 7642
rect 34969 7590 35021 7642
rect 1768 7395 1820 7404
rect 1768 7361 1777 7395
rect 1777 7361 1811 7395
rect 1811 7361 1820 7395
rect 1768 7352 1820 7361
rect 33508 7352 33560 7404
rect 1952 7327 2004 7336
rect 1952 7293 1961 7327
rect 1961 7293 1995 7327
rect 1995 7293 2004 7327
rect 1952 7284 2004 7293
rect 2780 7327 2832 7336
rect 2780 7293 2789 7327
rect 2789 7293 2823 7327
rect 2823 7293 2832 7327
rect 2780 7284 2832 7293
rect 4252 7191 4304 7200
rect 4252 7157 4261 7191
rect 4261 7157 4295 7191
rect 4295 7157 4304 7191
rect 4252 7148 4304 7157
rect 33232 7191 33284 7200
rect 33232 7157 33241 7191
rect 33241 7157 33275 7191
rect 33275 7157 33284 7191
rect 33232 7148 33284 7157
rect 33968 7191 34020 7200
rect 33968 7157 33977 7191
rect 33977 7157 34011 7191
rect 34011 7157 34020 7191
rect 33968 7148 34020 7157
rect 5170 7046 5222 7098
rect 5234 7046 5286 7098
rect 5298 7046 5350 7098
rect 5362 7046 5414 7098
rect 5426 7046 5478 7098
rect 13611 7046 13663 7098
rect 13675 7046 13727 7098
rect 13739 7046 13791 7098
rect 13803 7046 13855 7098
rect 13867 7046 13919 7098
rect 22052 7046 22104 7098
rect 22116 7046 22168 7098
rect 22180 7046 22232 7098
rect 22244 7046 22296 7098
rect 22308 7046 22360 7098
rect 30493 7046 30545 7098
rect 30557 7046 30609 7098
rect 30621 7046 30673 7098
rect 30685 7046 30737 7098
rect 30749 7046 30801 7098
rect 1952 6944 2004 6996
rect 33232 6808 33284 6860
rect 34336 6851 34388 6860
rect 34336 6817 34345 6851
rect 34345 6817 34379 6851
rect 34379 6817 34388 6851
rect 34336 6808 34388 6817
rect 2320 6740 2372 6792
rect 2688 6783 2740 6792
rect 2688 6749 2697 6783
rect 2697 6749 2731 6783
rect 2731 6749 2740 6783
rect 2688 6740 2740 6749
rect 1768 6672 1820 6724
rect 4344 6740 4396 6792
rect 4896 6740 4948 6792
rect 9128 6740 9180 6792
rect 19984 6740 20036 6792
rect 31944 6740 31996 6792
rect 7196 6672 7248 6724
rect 30288 6672 30340 6724
rect 33968 6672 34020 6724
rect 1952 6604 2004 6656
rect 2964 6604 3016 6656
rect 32680 6604 32732 6656
rect 9390 6502 9442 6554
rect 9454 6502 9506 6554
rect 9518 6502 9570 6554
rect 9582 6502 9634 6554
rect 9646 6502 9698 6554
rect 17831 6502 17883 6554
rect 17895 6502 17947 6554
rect 17959 6502 18011 6554
rect 18023 6502 18075 6554
rect 18087 6502 18139 6554
rect 26272 6502 26324 6554
rect 26336 6502 26388 6554
rect 26400 6502 26452 6554
rect 26464 6502 26516 6554
rect 26528 6502 26580 6554
rect 34713 6502 34765 6554
rect 34777 6502 34829 6554
rect 34841 6502 34893 6554
rect 34905 6502 34957 6554
rect 34969 6502 35021 6554
rect 1952 6375 2004 6384
rect 1952 6341 1961 6375
rect 1961 6341 1995 6375
rect 1995 6341 2004 6375
rect 1952 6332 2004 6341
rect 1768 6307 1820 6316
rect 1768 6273 1777 6307
rect 1777 6273 1811 6307
rect 1811 6273 1820 6307
rect 1768 6264 1820 6273
rect 3884 6264 3936 6316
rect 10508 6264 10560 6316
rect 31484 6264 31536 6316
rect 2872 6239 2924 6248
rect 2872 6205 2881 6239
rect 2881 6205 2915 6239
rect 2915 6205 2924 6239
rect 2872 6196 2924 6205
rect 33324 6196 33376 6248
rect 34336 6239 34388 6248
rect 34336 6205 34345 6239
rect 34345 6205 34379 6239
rect 34379 6205 34388 6239
rect 34336 6196 34388 6205
rect 3056 6128 3108 6180
rect 1584 6060 1636 6112
rect 4804 6103 4856 6112
rect 4804 6069 4813 6103
rect 4813 6069 4847 6103
rect 4847 6069 4856 6103
rect 4804 6060 4856 6069
rect 5170 5958 5222 6010
rect 5234 5958 5286 6010
rect 5298 5958 5350 6010
rect 5362 5958 5414 6010
rect 5426 5958 5478 6010
rect 13611 5958 13663 6010
rect 13675 5958 13727 6010
rect 13739 5958 13791 6010
rect 13803 5958 13855 6010
rect 13867 5958 13919 6010
rect 22052 5958 22104 6010
rect 22116 5958 22168 6010
rect 22180 5958 22232 6010
rect 22244 5958 22296 6010
rect 22308 5958 22360 6010
rect 30493 5958 30545 6010
rect 30557 5958 30609 6010
rect 30621 5958 30673 6010
rect 30685 5958 30737 6010
rect 30749 5958 30801 6010
rect 2320 5788 2372 5840
rect 1584 5763 1636 5772
rect 1584 5729 1593 5763
rect 1593 5729 1627 5763
rect 1627 5729 1636 5763
rect 1584 5720 1636 5729
rect 6460 5720 6512 5772
rect 28816 5720 28868 5772
rect 4344 5652 4396 5704
rect 4620 5695 4672 5704
rect 4620 5661 4629 5695
rect 4629 5661 4663 5695
rect 4663 5661 4672 5695
rect 4620 5652 4672 5661
rect 5080 5652 5132 5704
rect 5632 5652 5684 5704
rect 6092 5695 6144 5704
rect 6092 5661 6101 5695
rect 6101 5661 6135 5695
rect 6135 5661 6144 5695
rect 6092 5652 6144 5661
rect 6552 5695 6604 5704
rect 6552 5661 6561 5695
rect 6561 5661 6595 5695
rect 6595 5661 6604 5695
rect 6552 5652 6604 5661
rect 7380 5695 7432 5704
rect 7380 5661 7389 5695
rect 7389 5661 7423 5695
rect 7423 5661 7432 5695
rect 7380 5652 7432 5661
rect 31300 5652 31352 5704
rect 31852 5652 31904 5704
rect 32036 5695 32088 5704
rect 32036 5661 32045 5695
rect 32045 5661 32079 5695
rect 32079 5661 32088 5695
rect 32036 5652 32088 5661
rect 3424 5627 3476 5636
rect 3424 5593 3433 5627
rect 3433 5593 3467 5627
rect 3467 5593 3476 5627
rect 3424 5584 3476 5593
rect 4160 5584 4212 5636
rect 32128 5584 32180 5636
rect 34612 5584 34664 5636
rect 4712 5559 4764 5568
rect 4712 5525 4721 5559
rect 4721 5525 4755 5559
rect 4755 5525 4764 5559
rect 4712 5516 4764 5525
rect 6736 5516 6788 5568
rect 9390 5414 9442 5466
rect 9454 5414 9506 5466
rect 9518 5414 9570 5466
rect 9582 5414 9634 5466
rect 9646 5414 9698 5466
rect 17831 5414 17883 5466
rect 17895 5414 17947 5466
rect 17959 5414 18011 5466
rect 18023 5414 18075 5466
rect 18087 5414 18139 5466
rect 26272 5414 26324 5466
rect 26336 5414 26388 5466
rect 26400 5414 26452 5466
rect 26464 5414 26516 5466
rect 26528 5414 26580 5466
rect 34713 5414 34765 5466
rect 34777 5414 34829 5466
rect 34841 5414 34893 5466
rect 34905 5414 34957 5466
rect 34969 5414 35021 5466
rect 4712 5312 4764 5364
rect 34060 5244 34112 5296
rect 6460 5176 6512 5228
rect 7196 5219 7248 5228
rect 1768 5151 1820 5160
rect 1768 5117 1777 5151
rect 1777 5117 1811 5151
rect 1811 5117 1820 5151
rect 1768 5108 1820 5117
rect 2780 5151 2832 5160
rect 2780 5117 2789 5151
rect 2789 5117 2823 5151
rect 2823 5117 2832 5151
rect 2780 5108 2832 5117
rect 4896 5108 4948 5160
rect 7196 5185 7205 5219
rect 7205 5185 7239 5219
rect 7239 5185 7248 5219
rect 7196 5176 7248 5185
rect 28080 5176 28132 5228
rect 32036 5176 32088 5228
rect 4436 5040 4488 5092
rect 13176 5108 13228 5160
rect 33048 5151 33100 5160
rect 33048 5117 33057 5151
rect 33057 5117 33091 5151
rect 33091 5117 33100 5151
rect 33048 5108 33100 5117
rect 1860 4972 1912 5024
rect 31024 4972 31076 5024
rect 31208 5015 31260 5024
rect 31208 4981 31217 5015
rect 31217 4981 31251 5015
rect 31251 4981 31260 5015
rect 31208 4972 31260 4981
rect 5170 4870 5222 4922
rect 5234 4870 5286 4922
rect 5298 4870 5350 4922
rect 5362 4870 5414 4922
rect 5426 4870 5478 4922
rect 13611 4870 13663 4922
rect 13675 4870 13727 4922
rect 13739 4870 13791 4922
rect 13803 4870 13855 4922
rect 13867 4870 13919 4922
rect 22052 4870 22104 4922
rect 22116 4870 22168 4922
rect 22180 4870 22232 4922
rect 22244 4870 22296 4922
rect 22308 4870 22360 4922
rect 30493 4870 30545 4922
rect 30557 4870 30609 4922
rect 30621 4870 30673 4922
rect 30685 4870 30737 4922
rect 30749 4870 30801 4922
rect 6092 4700 6144 4752
rect 1860 4632 1912 4684
rect 2780 4675 2832 4684
rect 2780 4641 2789 4675
rect 2789 4641 2823 4675
rect 2823 4641 2832 4675
rect 2780 4632 2832 4641
rect 4804 4632 4856 4684
rect 4896 4675 4948 4684
rect 4896 4641 4905 4675
rect 4905 4641 4939 4675
rect 4939 4641 4948 4675
rect 4896 4632 4948 4641
rect 5080 4632 5132 4684
rect 6460 4607 6512 4616
rect 6460 4573 6469 4607
rect 6469 4573 6503 4607
rect 6503 4573 6512 4607
rect 6460 4564 6512 4573
rect 8024 4632 8076 4684
rect 31852 4632 31904 4684
rect 32680 4675 32732 4684
rect 32680 4641 32689 4675
rect 32689 4641 32723 4675
rect 32723 4641 32732 4675
rect 32680 4632 32732 4641
rect 7196 4564 7248 4616
rect 8392 4607 8444 4616
rect 8392 4573 8401 4607
rect 8401 4573 8435 4607
rect 8435 4573 8444 4607
rect 8392 4564 8444 4573
rect 19984 4607 20036 4616
rect 19984 4573 19993 4607
rect 19993 4573 20027 4607
rect 20027 4573 20036 4607
rect 19984 4564 20036 4573
rect 28080 4564 28132 4616
rect 5540 4496 5592 4548
rect 5816 4496 5868 4548
rect 30840 4496 30892 4548
rect 34336 4539 34388 4548
rect 6920 4428 6972 4480
rect 19800 4428 19852 4480
rect 34336 4505 34345 4539
rect 34345 4505 34379 4539
rect 34379 4505 34388 4539
rect 34336 4496 34388 4505
rect 34520 4428 34572 4480
rect 9390 4326 9442 4378
rect 9454 4326 9506 4378
rect 9518 4326 9570 4378
rect 9582 4326 9634 4378
rect 9646 4326 9698 4378
rect 17831 4326 17883 4378
rect 17895 4326 17947 4378
rect 17959 4326 18011 4378
rect 18023 4326 18075 4378
rect 18087 4326 18139 4378
rect 26272 4326 26324 4378
rect 26336 4326 26388 4378
rect 26400 4326 26452 4378
rect 26464 4326 26516 4378
rect 26528 4326 26580 4378
rect 34713 4326 34765 4378
rect 34777 4326 34829 4378
rect 34841 4326 34893 4378
rect 34905 4326 34957 4378
rect 34969 4326 35021 4378
rect 19800 4199 19852 4208
rect 1768 4088 1820 4140
rect 3976 4088 4028 4140
rect 4160 4020 4212 4072
rect 4344 4088 4396 4140
rect 5632 4131 5684 4140
rect 5632 4097 5641 4131
rect 5641 4097 5675 4131
rect 5675 4097 5684 4131
rect 5632 4088 5684 4097
rect 6552 4131 6604 4140
rect 6552 4097 6561 4131
rect 6561 4097 6595 4131
rect 6595 4097 6604 4131
rect 19800 4165 19809 4199
rect 19809 4165 19843 4199
rect 19843 4165 19852 4199
rect 19800 4156 19852 4165
rect 6552 4088 6604 4097
rect 5540 4020 5592 4072
rect 8024 4131 8076 4140
rect 8024 4097 8033 4131
rect 8033 4097 8067 4131
rect 8067 4097 8076 4131
rect 9128 4131 9180 4140
rect 8024 4088 8076 4097
rect 9128 4097 9137 4131
rect 9137 4097 9171 4131
rect 9171 4097 9180 4131
rect 9128 4088 9180 4097
rect 28816 4131 28868 4140
rect 28816 4097 28825 4131
rect 28825 4097 28859 4131
rect 28859 4097 28868 4131
rect 28816 4088 28868 4097
rect 31300 4088 31352 4140
rect 13084 4063 13136 4072
rect 13084 4029 13093 4063
rect 13093 4029 13127 4063
rect 13127 4029 13136 4063
rect 13084 4020 13136 4029
rect 13268 4063 13320 4072
rect 13268 4029 13277 4063
rect 13277 4029 13311 4063
rect 13311 4029 13320 4063
rect 13268 4020 13320 4029
rect 13452 4020 13504 4072
rect 20260 4020 20312 4072
rect 20628 4063 20680 4072
rect 20628 4029 20637 4063
rect 20637 4029 20671 4063
rect 20671 4029 20680 4063
rect 20628 4020 20680 4029
rect 27896 4020 27948 4072
rect 30104 4063 30156 4072
rect 30104 4029 30113 4063
rect 30113 4029 30147 4063
rect 30147 4029 30156 4063
rect 30104 4020 30156 4029
rect 31852 4020 31904 4072
rect 32680 4063 32732 4072
rect 32680 4029 32689 4063
rect 32689 4029 32723 4063
rect 32723 4029 32732 4063
rect 32680 4020 32732 4029
rect 35440 4020 35492 4072
rect 6460 3952 6512 4004
rect 6552 3952 6604 4004
rect 15660 3952 15712 4004
rect 27712 3952 27764 4004
rect 33140 3952 33192 4004
rect 4344 3884 4396 3936
rect 5724 3927 5776 3936
rect 5724 3893 5733 3927
rect 5733 3893 5767 3927
rect 5767 3893 5776 3927
rect 5724 3884 5776 3893
rect 6092 3884 6144 3936
rect 7196 3884 7248 3936
rect 9220 3927 9272 3936
rect 9220 3893 9229 3927
rect 9229 3893 9263 3927
rect 9263 3893 9272 3927
rect 9220 3884 9272 3893
rect 15568 3884 15620 3936
rect 16856 3884 16908 3936
rect 20076 3884 20128 3936
rect 27620 3884 27672 3936
rect 31668 3884 31720 3936
rect 5170 3782 5222 3834
rect 5234 3782 5286 3834
rect 5298 3782 5350 3834
rect 5362 3782 5414 3834
rect 5426 3782 5478 3834
rect 13611 3782 13663 3834
rect 13675 3782 13727 3834
rect 13739 3782 13791 3834
rect 13803 3782 13855 3834
rect 13867 3782 13919 3834
rect 22052 3782 22104 3834
rect 22116 3782 22168 3834
rect 22180 3782 22232 3834
rect 22244 3782 22296 3834
rect 22308 3782 22360 3834
rect 30493 3782 30545 3834
rect 30557 3782 30609 3834
rect 30621 3782 30673 3834
rect 30685 3782 30737 3834
rect 30749 3782 30801 3834
rect 13084 3723 13136 3732
rect 13084 3689 13093 3723
rect 13093 3689 13127 3723
rect 13127 3689 13136 3723
rect 13084 3680 13136 3689
rect 8392 3612 8444 3664
rect 10508 3612 10560 3664
rect 20076 3680 20128 3732
rect 20260 3723 20312 3732
rect 20260 3689 20269 3723
rect 20269 3689 20303 3723
rect 20303 3689 20312 3723
rect 20260 3680 20312 3689
rect 23756 3680 23808 3732
rect 27712 3680 27764 3732
rect 27896 3723 27948 3732
rect 27896 3689 27905 3723
rect 27905 3689 27939 3723
rect 27939 3689 27948 3723
rect 27896 3680 27948 3689
rect 30104 3680 30156 3732
rect 14372 3612 14424 3664
rect 2780 3587 2832 3596
rect 2780 3553 2789 3587
rect 2789 3553 2823 3587
rect 2823 3553 2832 3587
rect 2780 3544 2832 3553
rect 6092 3587 6144 3596
rect 6092 3553 6101 3587
rect 6101 3553 6135 3587
rect 6135 3553 6144 3587
rect 6092 3544 6144 3553
rect 6460 3587 6512 3596
rect 6460 3553 6469 3587
rect 6469 3553 6503 3587
rect 6503 3553 6512 3587
rect 6460 3544 6512 3553
rect 15568 3587 15620 3596
rect 15568 3553 15577 3587
rect 15577 3553 15611 3587
rect 15611 3553 15620 3587
rect 15568 3544 15620 3553
rect 16120 3587 16172 3596
rect 16120 3553 16129 3587
rect 16129 3553 16163 3587
rect 16163 3553 16172 3587
rect 16120 3544 16172 3553
rect 21272 3587 21324 3596
rect 21272 3553 21281 3587
rect 21281 3553 21315 3587
rect 21315 3553 21324 3587
rect 21272 3544 21324 3553
rect 4160 3519 4212 3528
rect 4160 3485 4169 3519
rect 4169 3485 4203 3519
rect 4203 3485 4212 3519
rect 4160 3476 4212 3485
rect 4804 3519 4856 3528
rect 4804 3485 4813 3519
rect 4813 3485 4847 3519
rect 4847 3485 4856 3519
rect 4804 3476 4856 3485
rect 9312 3519 9364 3528
rect 2964 3408 3016 3460
rect 7012 3408 7064 3460
rect 9312 3485 9321 3519
rect 9321 3485 9355 3519
rect 9355 3485 9364 3519
rect 9312 3476 9364 3485
rect 10048 3519 10100 3528
rect 10048 3485 10057 3519
rect 10057 3485 10091 3519
rect 10091 3485 10100 3519
rect 10048 3476 10100 3485
rect 10508 3519 10560 3528
rect 10508 3485 10517 3519
rect 10517 3485 10551 3519
rect 10551 3485 10560 3519
rect 10508 3476 10560 3485
rect 14280 3476 14332 3528
rect 14372 3519 14424 3528
rect 14372 3485 14381 3519
rect 14381 3485 14415 3519
rect 14415 3485 14424 3519
rect 14372 3476 14424 3485
rect 19432 3476 19484 3528
rect 20720 3519 20772 3528
rect 20720 3485 20729 3519
rect 20729 3485 20763 3519
rect 20763 3485 20772 3519
rect 20720 3476 20772 3485
rect 23756 3476 23808 3528
rect 24768 3519 24820 3528
rect 24768 3485 24777 3519
rect 24777 3485 24811 3519
rect 24811 3485 24820 3519
rect 24768 3476 24820 3485
rect 31944 3680 31996 3732
rect 34060 3723 34112 3732
rect 34060 3689 34069 3723
rect 34069 3689 34103 3723
rect 34103 3689 34112 3723
rect 34060 3680 34112 3689
rect 9128 3408 9180 3460
rect 15752 3451 15804 3460
rect 9772 3340 9824 3392
rect 14464 3383 14516 3392
rect 14464 3349 14473 3383
rect 14473 3349 14507 3383
rect 14507 3349 14516 3383
rect 14464 3340 14516 3349
rect 15752 3417 15761 3451
rect 15761 3417 15795 3451
rect 15795 3417 15804 3451
rect 15752 3408 15804 3417
rect 22100 3408 22152 3460
rect 27712 3408 27764 3460
rect 28448 3476 28500 3528
rect 29644 3476 29696 3528
rect 31760 3612 31812 3664
rect 33140 3612 33192 3664
rect 31208 3544 31260 3596
rect 31300 3544 31352 3596
rect 33784 3544 33836 3596
rect 30380 3476 30432 3528
rect 33508 3519 33560 3528
rect 33508 3485 33517 3519
rect 33517 3485 33551 3519
rect 33551 3485 33560 3519
rect 33508 3476 33560 3485
rect 31024 3408 31076 3460
rect 35900 3408 35952 3460
rect 24032 3340 24084 3392
rect 32496 3340 32548 3392
rect 9390 3238 9442 3290
rect 9454 3238 9506 3290
rect 9518 3238 9570 3290
rect 9582 3238 9634 3290
rect 9646 3238 9698 3290
rect 17831 3238 17883 3290
rect 17895 3238 17947 3290
rect 17959 3238 18011 3290
rect 18023 3238 18075 3290
rect 18087 3238 18139 3290
rect 26272 3238 26324 3290
rect 26336 3238 26388 3290
rect 26400 3238 26452 3290
rect 26464 3238 26516 3290
rect 26528 3238 26580 3290
rect 34713 3238 34765 3290
rect 34777 3238 34829 3290
rect 34841 3238 34893 3290
rect 34905 3238 34957 3290
rect 34969 3238 35021 3290
rect 6920 3136 6972 3188
rect 8024 3136 8076 3188
rect 13268 3179 13320 3188
rect 4344 3111 4396 3120
rect 4344 3077 4353 3111
rect 4353 3077 4387 3111
rect 4387 3077 4396 3111
rect 4344 3068 4396 3077
rect 7196 3111 7248 3120
rect 7196 3077 7205 3111
rect 7205 3077 7239 3111
rect 7239 3077 7248 3111
rect 7196 3068 7248 3077
rect 9772 3068 9824 3120
rect 13268 3145 13277 3179
rect 13277 3145 13311 3179
rect 13311 3145 13320 3179
rect 13268 3136 13320 3145
rect 19340 3136 19392 3188
rect 22100 3179 22152 3188
rect 22100 3145 22109 3179
rect 22109 3145 22143 3179
rect 22143 3145 22152 3179
rect 22100 3136 22152 3145
rect 14464 3111 14516 3120
rect 14464 3077 14473 3111
rect 14473 3077 14507 3111
rect 14507 3077 14516 3111
rect 14464 3068 14516 3077
rect 7012 3043 7064 3052
rect 7012 3009 7021 3043
rect 7021 3009 7055 3043
rect 7055 3009 7064 3043
rect 7012 3000 7064 3009
rect 13176 3043 13228 3052
rect 13176 3009 13185 3043
rect 13185 3009 13219 3043
rect 13219 3009 13228 3043
rect 13176 3000 13228 3009
rect 14280 3043 14332 3052
rect 14280 3009 14289 3043
rect 14289 3009 14323 3043
rect 14323 3009 14332 3043
rect 14280 3000 14332 3009
rect 3056 2932 3108 2984
rect 3240 2975 3292 2984
rect 3240 2941 3249 2975
rect 3249 2941 3283 2975
rect 3283 2941 3292 2975
rect 3240 2932 3292 2941
rect 4804 2932 4856 2984
rect 5080 2975 5132 2984
rect 5080 2941 5089 2975
rect 5089 2941 5123 2975
rect 5123 2941 5132 2975
rect 5080 2932 5132 2941
rect 8392 2975 8444 2984
rect 8392 2941 8401 2975
rect 8401 2941 8435 2975
rect 8435 2941 8444 2975
rect 8392 2932 8444 2941
rect 10048 2932 10100 2984
rect 10324 2975 10376 2984
rect 10324 2941 10333 2975
rect 10333 2941 10367 2975
rect 10367 2941 10376 2975
rect 10324 2932 10376 2941
rect 3884 2864 3936 2916
rect 4896 2864 4948 2916
rect 14832 2975 14884 2984
rect 14832 2941 14841 2975
rect 14841 2941 14875 2975
rect 14875 2941 14884 2975
rect 14832 2932 14884 2941
rect 23756 3068 23808 3120
rect 16856 3043 16908 3052
rect 16856 3009 16865 3043
rect 16865 3009 16899 3043
rect 16899 3009 16908 3043
rect 16856 3000 16908 3009
rect 19432 3043 19484 3052
rect 19432 3009 19441 3043
rect 19441 3009 19475 3043
rect 19475 3009 19484 3043
rect 19432 3000 19484 3009
rect 21916 3000 21968 3052
rect 24768 3136 24820 3188
rect 32680 3136 32732 3188
rect 24032 3111 24084 3120
rect 24032 3077 24041 3111
rect 24041 3077 24075 3111
rect 24075 3077 24084 3111
rect 24032 3068 24084 3077
rect 27620 3068 27672 3120
rect 28540 3068 28592 3120
rect 29920 3068 29972 3120
rect 31300 3068 31352 3120
rect 32496 3111 32548 3120
rect 32496 3077 32505 3111
rect 32505 3077 32539 3111
rect 32539 3077 32548 3111
rect 32496 3068 32548 3077
rect 17040 2975 17092 2984
rect 17040 2941 17049 2975
rect 17049 2941 17083 2975
rect 17083 2941 17092 2975
rect 17040 2932 17092 2941
rect 17408 2975 17460 2984
rect 17408 2941 17417 2975
rect 17417 2941 17451 2975
rect 17451 2941 17460 2975
rect 17408 2932 17460 2941
rect 19616 2975 19668 2984
rect 19616 2941 19625 2975
rect 19625 2941 19659 2975
rect 19659 2941 19668 2975
rect 19616 2932 19668 2941
rect 19984 2975 20036 2984
rect 19984 2941 19993 2975
rect 19993 2941 20027 2975
rect 20027 2941 20036 2975
rect 19984 2932 20036 2941
rect 24492 2975 24544 2984
rect 24492 2941 24501 2975
rect 24501 2941 24535 2975
rect 24535 2941 24544 2975
rect 24492 2932 24544 2941
rect 28448 3000 28500 3052
rect 29644 3043 29696 3052
rect 29644 3009 29653 3043
rect 29653 3009 29687 3043
rect 29687 3009 29696 3043
rect 29644 3000 29696 3009
rect 29092 2932 29144 2984
rect 29920 2932 29972 2984
rect 30288 2975 30340 2984
rect 30288 2941 30297 2975
rect 30297 2941 30331 2975
rect 30331 2941 30340 2975
rect 30288 2932 30340 2941
rect 33508 2932 33560 2984
rect 28540 2864 28592 2916
rect 664 2796 716 2848
rect 6828 2796 6880 2848
rect 30196 2796 30248 2848
rect 32220 2864 32272 2916
rect 32772 2796 32824 2848
rect 5170 2694 5222 2746
rect 5234 2694 5286 2746
rect 5298 2694 5350 2746
rect 5362 2694 5414 2746
rect 5426 2694 5478 2746
rect 13611 2694 13663 2746
rect 13675 2694 13727 2746
rect 13739 2694 13791 2746
rect 13803 2694 13855 2746
rect 13867 2694 13919 2746
rect 22052 2694 22104 2746
rect 22116 2694 22168 2746
rect 22180 2694 22232 2746
rect 22244 2694 22296 2746
rect 22308 2694 22360 2746
rect 30493 2694 30545 2746
rect 30557 2694 30609 2746
rect 30621 2694 30673 2746
rect 30685 2694 30737 2746
rect 30749 2694 30801 2746
rect 15752 2635 15804 2644
rect 15752 2601 15761 2635
rect 15761 2601 15795 2635
rect 15795 2601 15804 2635
rect 15752 2592 15804 2601
rect 17040 2635 17092 2644
rect 17040 2601 17049 2635
rect 17049 2601 17083 2635
rect 17083 2601 17092 2635
rect 17040 2592 17092 2601
rect 19064 2592 19116 2644
rect 19616 2592 19668 2644
rect 20720 2592 20772 2644
rect 30840 2592 30892 2644
rect 4252 2524 4304 2576
rect 2596 2499 2648 2508
rect 2596 2465 2605 2499
rect 2605 2465 2639 2499
rect 2639 2465 2648 2499
rect 2596 2456 2648 2465
rect 4160 2499 4212 2508
rect 4160 2465 4169 2499
rect 4169 2465 4203 2499
rect 4203 2465 4212 2499
rect 4160 2456 4212 2465
rect 4528 2456 4580 2508
rect 7380 2524 7432 2576
rect 32128 2524 32180 2576
rect 6736 2499 6788 2508
rect 6736 2465 6745 2499
rect 6745 2465 6779 2499
rect 6779 2465 6788 2499
rect 6736 2456 6788 2465
rect 6828 2456 6880 2508
rect 9312 2456 9364 2508
rect 9772 2499 9824 2508
rect 9772 2465 9781 2499
rect 9781 2465 9815 2499
rect 9815 2465 9824 2499
rect 9772 2456 9824 2465
rect 15660 2431 15712 2440
rect 15660 2397 15669 2431
rect 15669 2397 15703 2431
rect 15703 2397 15712 2431
rect 15660 2388 15712 2397
rect 18236 2388 18288 2440
rect 19340 2388 19392 2440
rect 29092 2456 29144 2508
rect 30380 2456 30432 2508
rect 30932 2499 30984 2508
rect 30932 2465 30941 2499
rect 30941 2465 30975 2499
rect 30975 2465 30984 2499
rect 30932 2456 30984 2465
rect 31668 2456 31720 2508
rect 32864 2499 32916 2508
rect 32864 2465 32873 2499
rect 32873 2465 32907 2499
rect 32907 2465 32916 2499
rect 32864 2456 32916 2465
rect 27712 2431 27764 2440
rect 27712 2397 27721 2431
rect 27721 2397 27755 2431
rect 27755 2397 27764 2431
rect 27712 2388 27764 2397
rect 28540 2388 28592 2440
rect 29000 2431 29052 2440
rect 29000 2397 29009 2431
rect 29009 2397 29043 2431
rect 29043 2397 29052 2431
rect 29000 2388 29052 2397
rect 5724 2320 5776 2372
rect 9312 2363 9364 2372
rect 9312 2329 9321 2363
rect 9321 2329 9355 2363
rect 9355 2329 9364 2363
rect 9312 2320 9364 2329
rect 5816 2252 5868 2304
rect 30196 2320 30248 2372
rect 33416 2252 33468 2304
rect 9390 2150 9442 2202
rect 9454 2150 9506 2202
rect 9518 2150 9570 2202
rect 9582 2150 9634 2202
rect 9646 2150 9698 2202
rect 17831 2150 17883 2202
rect 17895 2150 17947 2202
rect 17959 2150 18011 2202
rect 18023 2150 18075 2202
rect 18087 2150 18139 2202
rect 26272 2150 26324 2202
rect 26336 2150 26388 2202
rect 26400 2150 26452 2202
rect 26464 2150 26516 2202
rect 26528 2150 26580 2202
rect 34713 2150 34765 2202
rect 34777 2150 34829 2202
rect 34841 2150 34893 2202
rect 34905 2150 34957 2202
rect 34969 2150 35021 2202
rect 34520 1096 34572 1148
rect 34796 1096 34848 1148
<< metal2 >>
rect -10 41200 102 41800
rect 634 41200 746 41800
rect 1278 41200 1390 41800
rect 1922 41200 2034 41800
rect 2566 41200 2678 41800
rect 2778 41576 2834 41585
rect 2778 41511 2834 41520
rect 676 38282 704 41200
rect 1320 39370 1348 41200
rect 1308 39364 1360 39370
rect 1308 39306 1360 39312
rect 2792 38894 2820 41511
rect 3210 41200 3322 41800
rect 4498 41200 4610 41800
rect 5142 41200 5254 41800
rect 5786 41200 5898 41800
rect 6430 41200 6542 41800
rect 7074 41200 7186 41800
rect 7718 41200 7830 41800
rect 8362 41200 8474 41800
rect 9006 41200 9118 41800
rect 9650 41200 9762 41800
rect 10938 41200 11050 41800
rect 11582 41200 11694 41800
rect 12226 41200 12338 41800
rect 12870 41200 12982 41800
rect 13514 41200 13626 41800
rect 14158 41200 14270 41800
rect 14802 41200 14914 41800
rect 15446 41200 15558 41800
rect 16090 41200 16202 41800
rect 17378 41200 17490 41800
rect 18022 41200 18134 41800
rect 18666 41200 18778 41800
rect 19310 41200 19422 41800
rect 19954 41200 20066 41800
rect 20598 41200 20710 41800
rect 21242 41200 21354 41800
rect 21886 41200 21998 41800
rect 22530 41200 22642 41800
rect 23818 41200 23930 41800
rect 24462 41200 24574 41800
rect 25106 41200 25218 41800
rect 25750 41200 25862 41800
rect 26394 41200 26506 41800
rect 27038 41200 27150 41800
rect 27682 41200 27794 41800
rect 28326 41200 28438 41800
rect 28970 41200 29082 41800
rect 30258 41200 30370 41800
rect 30902 41200 31014 41800
rect 31546 41200 31658 41800
rect 32190 41200 32302 41800
rect 32834 41200 32946 41800
rect 33478 41200 33590 41800
rect 34122 41200 34234 41800
rect 34766 41200 34878 41800
rect 35410 41200 35522 41800
rect 3252 39386 3280 41200
rect 3422 40896 3478 40905
rect 3422 40831 3478 40840
rect 3252 39358 3372 39386
rect 3240 39296 3292 39302
rect 3240 39238 3292 39244
rect 2780 38888 2832 38894
rect 2780 38830 2832 38836
rect 664 38276 716 38282
rect 664 38218 716 38224
rect 3252 37942 3280 39238
rect 3240 37936 3292 37942
rect 3240 37878 3292 37884
rect 1676 37868 1728 37874
rect 1676 37810 1728 37816
rect 2964 37868 3016 37874
rect 2964 37810 3016 37816
rect 1688 33114 1716 37810
rect 2042 37496 2098 37505
rect 2042 37431 2098 37440
rect 2056 37330 2084 37431
rect 2044 37324 2096 37330
rect 2044 37266 2096 37272
rect 2976 37262 3004 37810
rect 3056 37800 3108 37806
rect 3056 37742 3108 37748
rect 3068 37466 3096 37742
rect 3056 37460 3108 37466
rect 3056 37402 3108 37408
rect 3344 37330 3372 39358
rect 3436 37806 3464 40831
rect 5170 39740 5478 39749
rect 5170 39738 5176 39740
rect 5232 39738 5256 39740
rect 5312 39738 5336 39740
rect 5392 39738 5416 39740
rect 5472 39738 5478 39740
rect 5232 39686 5234 39738
rect 5414 39686 5416 39738
rect 5170 39684 5176 39686
rect 5232 39684 5256 39686
rect 5312 39684 5336 39686
rect 5392 39684 5416 39686
rect 5472 39684 5478 39686
rect 5170 39675 5478 39684
rect 3884 39432 3936 39438
rect 3884 39374 3936 39380
rect 4160 39432 4212 39438
rect 4160 39374 4212 39380
rect 3516 39092 3568 39098
rect 3516 39034 3568 39040
rect 3528 38865 3556 39034
rect 3514 38856 3570 38865
rect 3514 38791 3570 38800
rect 3896 38758 3924 39374
rect 4172 38962 4200 39374
rect 5080 39024 5132 39030
rect 5080 38966 5132 38972
rect 4160 38956 4212 38962
rect 4160 38898 4212 38904
rect 3976 38820 4028 38826
rect 3976 38762 4028 38768
rect 3884 38752 3936 38758
rect 3884 38694 3936 38700
rect 3424 37800 3476 37806
rect 3424 37742 3476 37748
rect 3332 37324 3384 37330
rect 3332 37266 3384 37272
rect 2964 37256 3016 37262
rect 2964 37198 3016 37204
rect 2778 36816 2834 36825
rect 2778 36751 2834 36760
rect 2792 36718 2820 36751
rect 2780 36712 2832 36718
rect 2780 36654 2832 36660
rect 3240 36236 3292 36242
rect 3240 36178 3292 36184
rect 1768 36168 1820 36174
rect 1768 36110 1820 36116
rect 2044 36168 2096 36174
rect 2044 36110 2096 36116
rect 2870 36136 2926 36145
rect 1780 34610 1808 36110
rect 2056 35630 2084 36110
rect 2870 36071 2926 36080
rect 2884 35894 2912 36071
rect 2884 35866 3004 35894
rect 2504 35692 2556 35698
rect 2504 35634 2556 35640
rect 2044 35624 2096 35630
rect 2044 35566 2096 35572
rect 1768 34604 1820 34610
rect 1768 34546 1820 34552
rect 1952 34536 2004 34542
rect 1952 34478 2004 34484
rect 1964 34202 1992 34478
rect 1952 34196 2004 34202
rect 1952 34138 2004 34144
rect 1676 33108 1728 33114
rect 1676 33050 1728 33056
rect 1768 31816 1820 31822
rect 1768 31758 1820 31764
rect 1780 31346 1808 31758
rect 1768 31340 1820 31346
rect 1768 31282 1820 31288
rect 2056 26234 2084 35566
rect 2516 35018 2544 35634
rect 2778 35456 2834 35465
rect 2778 35391 2834 35400
rect 2792 35154 2820 35391
rect 2780 35148 2832 35154
rect 2780 35090 2832 35096
rect 2136 35012 2188 35018
rect 2136 34954 2188 34960
rect 2504 35012 2556 35018
rect 2504 34954 2556 34960
rect 2148 33658 2176 34954
rect 2516 33998 2544 34954
rect 2872 34944 2924 34950
rect 2872 34886 2924 34892
rect 2780 34536 2832 34542
rect 2780 34478 2832 34484
rect 2792 34105 2820 34478
rect 2778 34096 2834 34105
rect 2778 34031 2834 34040
rect 2504 33992 2556 33998
rect 2504 33934 2556 33940
rect 2136 33652 2188 33658
rect 2136 33594 2188 33600
rect 2884 33522 2912 34886
rect 2320 33516 2372 33522
rect 2320 33458 2372 33464
rect 2872 33516 2924 33522
rect 2872 33458 2924 33464
rect 2136 31272 2188 31278
rect 2136 31214 2188 31220
rect 2148 30938 2176 31214
rect 2136 30932 2188 30938
rect 2136 30874 2188 30880
rect 2136 30728 2188 30734
rect 2136 30670 2188 30676
rect 2148 26994 2176 30670
rect 2136 26988 2188 26994
rect 2136 26930 2188 26936
rect 1964 26206 2084 26234
rect 1584 25696 1636 25702
rect 1584 25638 1636 25644
rect 1596 25362 1624 25638
rect 1584 25356 1636 25362
rect 1584 25298 1636 25304
rect 1768 25220 1820 25226
rect 1768 25162 1820 25168
rect 1780 24954 1808 25162
rect 1768 24948 1820 24954
rect 1768 24890 1820 24896
rect 1964 19854 1992 26206
rect 2044 24812 2096 24818
rect 2044 24754 2096 24760
rect 1952 19848 2004 19854
rect 1952 19790 2004 19796
rect 1952 19712 2004 19718
rect 1952 19654 2004 19660
rect 1964 19446 1992 19654
rect 1952 19440 2004 19446
rect 1952 19382 2004 19388
rect 1768 19304 1820 19310
rect 1768 19246 1820 19252
rect 1780 18970 1808 19246
rect 1768 18964 1820 18970
rect 1768 18906 1820 18912
rect 2056 18834 2084 24754
rect 2044 18828 2096 18834
rect 2044 18770 2096 18776
rect 1768 18760 1820 18766
rect 1768 18702 1820 18708
rect 1780 18290 1808 18702
rect 1768 18284 1820 18290
rect 1768 18226 1820 18232
rect 1952 18216 2004 18222
rect 1952 18158 2004 18164
rect 1964 17882 1992 18158
rect 1952 17876 2004 17882
rect 1952 17818 2004 17824
rect 2148 17678 2176 26930
rect 2228 19304 2280 19310
rect 2228 19246 2280 19252
rect 2240 19145 2268 19246
rect 2226 19136 2282 19145
rect 2226 19071 2282 19080
rect 2228 18828 2280 18834
rect 2228 18770 2280 18776
rect 2136 17672 2188 17678
rect 2136 17614 2188 17620
rect 1768 17128 1820 17134
rect 1768 17070 1820 17076
rect 1780 16794 1808 17070
rect 1768 16788 1820 16794
rect 1768 16730 1820 16736
rect 1584 15904 1636 15910
rect 1584 15846 1636 15852
rect 1596 15570 1624 15846
rect 1584 15564 1636 15570
rect 1584 15506 1636 15512
rect 1768 15428 1820 15434
rect 1768 15370 1820 15376
rect 1780 15162 1808 15370
rect 1768 15156 1820 15162
rect 1768 15098 1820 15104
rect 1768 14816 1820 14822
rect 1768 14758 1820 14764
rect 1780 14482 1808 14758
rect 1768 14476 1820 14482
rect 1768 14418 1820 14424
rect 1584 14408 1636 14414
rect 1584 14350 1636 14356
rect 1596 13462 1624 14350
rect 1768 13864 1820 13870
rect 1768 13806 1820 13812
rect 1952 13864 2004 13870
rect 1952 13806 2004 13812
rect 1780 13530 1808 13806
rect 1768 13524 1820 13530
rect 1768 13466 1820 13472
rect 1584 13456 1636 13462
rect 1584 13398 1636 13404
rect 1964 12986 1992 13806
rect 1952 12980 2004 12986
rect 1952 12922 2004 12928
rect 2148 12238 2176 17614
rect 2240 12850 2268 18770
rect 2228 12844 2280 12850
rect 2228 12786 2280 12792
rect 2136 12232 2188 12238
rect 2136 12174 2188 12180
rect 1952 12096 2004 12102
rect 1952 12038 2004 12044
rect 1964 11830 1992 12038
rect 1952 11824 2004 11830
rect 1952 11766 2004 11772
rect 2044 11688 2096 11694
rect 2044 11630 2096 11636
rect 2056 11354 2084 11630
rect 2044 11348 2096 11354
rect 2044 11290 2096 11296
rect 1768 11144 1820 11150
rect 1768 11086 1820 11092
rect 1780 10674 1808 11086
rect 1768 10668 1820 10674
rect 1768 10610 1820 10616
rect 2044 10600 2096 10606
rect 2044 10542 2096 10548
rect 2056 10266 2084 10542
rect 2044 10260 2096 10266
rect 2044 10202 2096 10208
rect 1584 9376 1636 9382
rect 1584 9318 1636 9324
rect 1596 9042 1624 9318
rect 1584 9036 1636 9042
rect 1584 8978 1636 8984
rect 1768 8424 1820 8430
rect 1768 8366 1820 8372
rect 1780 8090 1808 8366
rect 1768 8084 1820 8090
rect 1768 8026 1820 8032
rect 1768 7812 1820 7818
rect 1768 7754 1820 7760
rect 1780 7410 1808 7754
rect 1768 7404 1820 7410
rect 1768 7346 1820 7352
rect 1952 7336 2004 7342
rect 1952 7278 2004 7284
rect 1964 7002 1992 7278
rect 1952 6996 2004 7002
rect 1952 6938 2004 6944
rect 2332 6798 2360 33458
rect 2976 32910 3004 35866
rect 3056 33924 3108 33930
rect 3056 33866 3108 33872
rect 2964 32904 3016 32910
rect 2964 32846 3016 32852
rect 2778 31376 2834 31385
rect 2778 31311 2834 31320
rect 2792 31278 2820 31311
rect 2780 31272 2832 31278
rect 2780 31214 2832 31220
rect 2780 25356 2832 25362
rect 2780 25298 2832 25304
rect 2792 25265 2820 25298
rect 2778 25256 2834 25265
rect 2778 25191 2834 25200
rect 3068 24818 3096 33866
rect 3252 33590 3280 36178
rect 3896 35630 3924 38694
rect 3988 37398 4016 38762
rect 4160 38344 4212 38350
rect 4160 38286 4212 38292
rect 4896 38344 4948 38350
rect 4896 38286 4948 38292
rect 4068 38208 4120 38214
rect 4068 38150 4120 38156
rect 3976 37392 4028 37398
rect 3976 37334 4028 37340
rect 3976 37256 4028 37262
rect 3976 37198 4028 37204
rect 3988 36786 4016 37198
rect 4080 37194 4108 38150
rect 4068 37188 4120 37194
rect 4068 37130 4120 37136
rect 4172 37126 4200 38286
rect 4436 38276 4488 38282
rect 4436 38218 4488 38224
rect 4160 37120 4212 37126
rect 4160 37062 4212 37068
rect 3976 36780 4028 36786
rect 3976 36722 4028 36728
rect 3988 36174 4016 36722
rect 4448 36718 4476 38218
rect 4908 37942 4936 38286
rect 4896 37936 4948 37942
rect 4896 37878 4948 37884
rect 4804 37868 4856 37874
rect 4804 37810 4856 37816
rect 4620 37188 4672 37194
rect 4620 37130 4672 37136
rect 4436 36712 4488 36718
rect 4436 36654 4488 36660
rect 3976 36168 4028 36174
rect 3976 36110 4028 36116
rect 3988 35698 4016 36110
rect 4632 35894 4660 37130
rect 4816 36242 4844 37810
rect 4804 36236 4856 36242
rect 4804 36178 4856 36184
rect 4804 36100 4856 36106
rect 4804 36042 4856 36048
rect 4448 35866 4660 35894
rect 3976 35692 4028 35698
rect 3976 35634 4028 35640
rect 3884 35624 3936 35630
rect 3884 35566 3936 35572
rect 3240 33584 3292 33590
rect 3240 33526 3292 33532
rect 3514 32056 3570 32065
rect 3514 31991 3570 32000
rect 3528 27334 3556 31991
rect 3516 27328 3568 27334
rect 3516 27270 3568 27276
rect 3056 24812 3108 24818
rect 3056 24754 3108 24760
rect 2504 19848 2556 19854
rect 2504 19790 2556 19796
rect 2516 16590 2544 19790
rect 2778 18456 2834 18465
rect 2778 18391 2834 18400
rect 2792 18222 2820 18391
rect 2780 18216 2832 18222
rect 2780 18158 2832 18164
rect 2596 17128 2648 17134
rect 2780 17128 2832 17134
rect 2596 17070 2648 17076
rect 2778 17096 2780 17105
rect 2832 17096 2834 17105
rect 2608 16794 2636 17070
rect 2778 17031 2834 17040
rect 2596 16788 2648 16794
rect 2596 16730 2648 16736
rect 2504 16584 2556 16590
rect 2556 16546 2912 16574
rect 2504 16526 2556 16532
rect 2778 15736 2834 15745
rect 2778 15671 2834 15680
rect 2792 15570 2820 15671
rect 2780 15564 2832 15570
rect 2780 15506 2832 15512
rect 2884 15026 2912 16546
rect 2872 15020 2924 15026
rect 2872 14962 2924 14968
rect 2780 14476 2832 14482
rect 2780 14418 2832 14424
rect 2792 14385 2820 14418
rect 2778 14376 2834 14385
rect 2778 14311 2834 14320
rect 2780 13864 2832 13870
rect 2780 13806 2832 13812
rect 2792 13705 2820 13806
rect 2778 13696 2834 13705
rect 2778 13631 2834 13640
rect 2688 12844 2740 12850
rect 2688 12786 2740 12792
rect 2596 9376 2648 9382
rect 2596 9318 2648 9324
rect 2608 9042 2636 9318
rect 2596 9036 2648 9042
rect 2596 8978 2648 8984
rect 2596 8424 2648 8430
rect 2596 8366 2648 8372
rect 2608 8090 2636 8366
rect 2596 8084 2648 8090
rect 2596 8026 2648 8032
rect 2700 6798 2728 12786
rect 2780 11688 2832 11694
rect 2778 11656 2780 11665
rect 2832 11656 2834 11665
rect 2778 11591 2834 11600
rect 2778 10976 2834 10985
rect 2778 10911 2834 10920
rect 2792 10606 2820 10911
rect 2780 10600 2832 10606
rect 2780 10542 2832 10548
rect 2884 9586 2912 14962
rect 2872 9580 2924 9586
rect 2872 9522 2924 9528
rect 2780 9036 2832 9042
rect 2780 8978 2832 8984
rect 2792 8945 2820 8978
rect 2778 8936 2834 8945
rect 2778 8871 2834 8880
rect 2780 8424 2832 8430
rect 2780 8366 2832 8372
rect 2792 8265 2820 8366
rect 2778 8256 2834 8265
rect 2778 8191 2834 8200
rect 2778 7576 2834 7585
rect 2778 7511 2834 7520
rect 2792 7342 2820 7511
rect 2780 7336 2832 7342
rect 2780 7278 2832 7284
rect 2320 6792 2372 6798
rect 2320 6734 2372 6740
rect 2688 6792 2740 6798
rect 2688 6734 2740 6740
rect 1768 6724 1820 6730
rect 1768 6666 1820 6672
rect 1780 6322 1808 6666
rect 1952 6656 2004 6662
rect 1952 6598 2004 6604
rect 1964 6390 1992 6598
rect 1952 6384 2004 6390
rect 1952 6326 2004 6332
rect 1768 6316 1820 6322
rect 1768 6258 1820 6264
rect 1584 6112 1636 6118
rect 1584 6054 1636 6060
rect 1596 5778 1624 6054
rect 2332 5846 2360 6734
rect 2964 6656 3016 6662
rect 2964 6598 3016 6604
rect 2872 6248 2924 6254
rect 2872 6190 2924 6196
rect 2320 5840 2372 5846
rect 2320 5782 2372 5788
rect 1584 5772 1636 5778
rect 1584 5714 1636 5720
rect 1768 5160 1820 5166
rect 1768 5102 1820 5108
rect 2780 5160 2832 5166
rect 2780 5102 2832 5108
rect 1780 4146 1808 5102
rect 1860 5024 1912 5030
rect 1860 4966 1912 4972
rect 1872 4690 1900 4966
rect 2792 4865 2820 5102
rect 2778 4856 2834 4865
rect 2778 4791 2834 4800
rect 1860 4684 1912 4690
rect 1860 4626 1912 4632
rect 2780 4684 2832 4690
rect 2780 4626 2832 4632
rect 2792 4185 2820 4626
rect 2778 4176 2834 4185
rect 1768 4140 1820 4146
rect 2778 4111 2834 4120
rect 1768 4082 1820 4088
rect 2780 3596 2832 3602
rect 2780 3538 2832 3544
rect 664 2848 716 2854
rect 664 2790 716 2796
rect 676 800 704 2790
rect 2596 2508 2648 2514
rect 2596 2450 2648 2456
rect 2608 800 2636 2450
rect 2792 2145 2820 3538
rect 2884 3505 2912 6190
rect 2870 3496 2926 3505
rect 2976 3466 3004 6598
rect 3896 6322 3924 35566
rect 3988 35086 4016 35634
rect 3976 35080 4028 35086
rect 3976 35022 4028 35028
rect 4448 34066 4476 35866
rect 4712 35012 4764 35018
rect 4712 34954 4764 34960
rect 4436 34060 4488 34066
rect 4436 34002 4488 34008
rect 4252 7200 4304 7206
rect 4252 7142 4304 7148
rect 3884 6316 3936 6322
rect 3884 6258 3936 6264
rect 3056 6180 3108 6186
rect 3056 6122 3108 6128
rect 2870 3431 2926 3440
rect 2964 3460 3016 3466
rect 2964 3402 3016 3408
rect 3068 2990 3096 6122
rect 3424 5636 3476 5642
rect 3424 5578 3476 5584
rect 4160 5636 4212 5642
rect 4160 5578 4212 5584
rect 3436 5545 3464 5578
rect 3422 5536 3478 5545
rect 3422 5471 3478 5480
rect 3976 4140 4028 4146
rect 3976 4082 4028 4088
rect 3056 2984 3108 2990
rect 3056 2926 3108 2932
rect 3240 2984 3292 2990
rect 3240 2926 3292 2932
rect 2778 2136 2834 2145
rect 2778 2071 2834 2080
rect 3252 800 3280 2926
rect 3884 2916 3936 2922
rect 3884 2858 3936 2864
rect 3896 800 3924 2858
rect 3988 2825 4016 4082
rect 4172 4078 4200 5578
rect 4160 4072 4212 4078
rect 4160 4014 4212 4020
rect 4160 3528 4212 3534
rect 4160 3470 4212 3476
rect 3974 2816 4030 2825
rect 3974 2751 4030 2760
rect 4172 2514 4200 3470
rect 4264 2582 4292 7142
rect 4448 6914 4476 34002
rect 4724 10062 4752 34954
rect 4816 16574 4844 36042
rect 4908 33930 4936 37878
rect 5092 36718 5120 38966
rect 5828 38894 5856 41200
rect 7116 39506 7144 41200
rect 7104 39500 7156 39506
rect 7104 39442 7156 39448
rect 6736 39364 6788 39370
rect 6736 39306 6788 39312
rect 5540 38888 5592 38894
rect 5540 38830 5592 38836
rect 5816 38888 5868 38894
rect 5816 38830 5868 38836
rect 5170 38652 5478 38661
rect 5170 38650 5176 38652
rect 5232 38650 5256 38652
rect 5312 38650 5336 38652
rect 5392 38650 5416 38652
rect 5472 38650 5478 38652
rect 5232 38598 5234 38650
rect 5414 38598 5416 38650
rect 5170 38596 5176 38598
rect 5232 38596 5256 38598
rect 5312 38596 5336 38598
rect 5392 38596 5416 38598
rect 5472 38596 5478 38598
rect 5170 38587 5478 38596
rect 5552 38010 5580 38830
rect 6748 38554 6776 39306
rect 7288 39296 7340 39302
rect 7288 39238 7340 39244
rect 6736 38548 6788 38554
rect 6736 38490 6788 38496
rect 7196 38276 7248 38282
rect 7196 38218 7248 38224
rect 7208 38010 7236 38218
rect 5540 38004 5592 38010
rect 5540 37946 5592 37952
rect 7196 38004 7248 38010
rect 7196 37946 7248 37952
rect 6368 37868 6420 37874
rect 6368 37810 6420 37816
rect 5724 37664 5776 37670
rect 5724 37606 5776 37612
rect 5170 37564 5478 37573
rect 5170 37562 5176 37564
rect 5232 37562 5256 37564
rect 5312 37562 5336 37564
rect 5392 37562 5416 37564
rect 5472 37562 5478 37564
rect 5232 37510 5234 37562
rect 5414 37510 5416 37562
rect 5170 37508 5176 37510
rect 5232 37508 5256 37510
rect 5312 37508 5336 37510
rect 5392 37508 5416 37510
rect 5472 37508 5478 37510
rect 5170 37499 5478 37508
rect 5540 37256 5592 37262
rect 5540 37198 5592 37204
rect 5552 36922 5580 37198
rect 5540 36916 5592 36922
rect 5540 36858 5592 36864
rect 5736 36786 5764 37606
rect 6380 37466 6408 37810
rect 6368 37460 6420 37466
rect 6368 37402 6420 37408
rect 6736 37256 6788 37262
rect 6788 37204 6868 37210
rect 6736 37198 6868 37204
rect 6748 37182 6868 37198
rect 6840 37126 6868 37182
rect 6828 37120 6880 37126
rect 6828 37062 6880 37068
rect 7300 36922 7328 39238
rect 7760 38418 7788 41200
rect 8116 38752 8168 38758
rect 8116 38694 8168 38700
rect 7748 38412 7800 38418
rect 7748 38354 7800 38360
rect 7472 38208 7524 38214
rect 7472 38150 7524 38156
rect 7484 37262 7512 38150
rect 8128 37942 8156 38694
rect 8404 37942 8432 41200
rect 9048 38894 9076 41200
rect 13611 39740 13919 39749
rect 13611 39738 13617 39740
rect 13673 39738 13697 39740
rect 13753 39738 13777 39740
rect 13833 39738 13857 39740
rect 13913 39738 13919 39740
rect 13673 39686 13675 39738
rect 13855 39686 13857 39738
rect 13611 39684 13617 39686
rect 13673 39684 13697 39686
rect 13753 39684 13777 39686
rect 13833 39684 13857 39686
rect 13913 39684 13919 39686
rect 13611 39675 13919 39684
rect 14844 39506 14872 41200
rect 14832 39500 14884 39506
rect 14832 39442 14884 39448
rect 9312 39432 9364 39438
rect 13728 39432 13780 39438
rect 9312 39374 9364 39380
rect 13726 39400 13728 39409
rect 14004 39432 14056 39438
rect 13780 39400 13782 39409
rect 8576 38888 8628 38894
rect 8576 38830 8628 38836
rect 9036 38888 9088 38894
rect 9036 38830 9088 38836
rect 8588 38554 8616 38830
rect 8576 38548 8628 38554
rect 8576 38490 8628 38496
rect 9128 38344 9180 38350
rect 9128 38286 9180 38292
rect 9140 38010 9168 38286
rect 9128 38004 9180 38010
rect 9128 37946 9180 37952
rect 8116 37936 8168 37942
rect 8116 37878 8168 37884
rect 8392 37936 8444 37942
rect 8392 37878 8444 37884
rect 7380 37256 7432 37262
rect 7380 37198 7432 37204
rect 7472 37256 7524 37262
rect 7472 37198 7524 37204
rect 7288 36916 7340 36922
rect 7288 36858 7340 36864
rect 7392 36786 7420 37198
rect 5540 36780 5592 36786
rect 5540 36722 5592 36728
rect 5724 36780 5776 36786
rect 5724 36722 5776 36728
rect 6552 36780 6604 36786
rect 6552 36722 6604 36728
rect 7380 36780 7432 36786
rect 7380 36722 7432 36728
rect 4988 36712 5040 36718
rect 4988 36654 5040 36660
rect 5080 36712 5132 36718
rect 5080 36654 5132 36660
rect 5000 35894 5028 36654
rect 5170 36476 5478 36485
rect 5170 36474 5176 36476
rect 5232 36474 5256 36476
rect 5312 36474 5336 36476
rect 5392 36474 5416 36476
rect 5472 36474 5478 36476
rect 5232 36422 5234 36474
rect 5414 36422 5416 36474
rect 5170 36420 5176 36422
rect 5232 36420 5256 36422
rect 5312 36420 5336 36422
rect 5392 36420 5416 36422
rect 5472 36420 5478 36422
rect 5170 36411 5478 36420
rect 5000 35866 5120 35894
rect 4896 33924 4948 33930
rect 4896 33866 4948 33872
rect 4816 16546 5028 16574
rect 4712 10056 4764 10062
rect 4712 9998 4764 10004
rect 4724 6914 4752 9998
rect 4356 6886 4476 6914
rect 4632 6886 4752 6914
rect 4356 6798 4384 6886
rect 4344 6792 4396 6798
rect 4344 6734 4396 6740
rect 4356 5710 4384 6734
rect 4632 5710 4660 6886
rect 4896 6792 4948 6798
rect 4896 6734 4948 6740
rect 4804 6112 4856 6118
rect 4804 6054 4856 6060
rect 4344 5704 4396 5710
rect 4344 5646 4396 5652
rect 4620 5704 4672 5710
rect 4620 5646 4672 5652
rect 4356 4146 4384 5646
rect 4712 5568 4764 5574
rect 4712 5510 4764 5516
rect 4724 5370 4752 5510
rect 4712 5364 4764 5370
rect 4712 5306 4764 5312
rect 4436 5092 4488 5098
rect 4436 5034 4488 5040
rect 4344 4140 4396 4146
rect 4344 4082 4396 4088
rect 4344 3936 4396 3942
rect 4344 3878 4396 3884
rect 4356 3126 4384 3878
rect 4344 3120 4396 3126
rect 4344 3062 4396 3068
rect 4252 2576 4304 2582
rect 4252 2518 4304 2524
rect 4160 2508 4212 2514
rect 4160 2450 4212 2456
rect 4066 1456 4122 1465
rect 4448 1442 4476 5034
rect 4816 4690 4844 6054
rect 4908 5166 4936 6734
rect 5000 5522 5028 16546
rect 5092 5710 5120 35866
rect 5170 35388 5478 35397
rect 5170 35386 5176 35388
rect 5232 35386 5256 35388
rect 5312 35386 5336 35388
rect 5392 35386 5416 35388
rect 5472 35386 5478 35388
rect 5232 35334 5234 35386
rect 5414 35334 5416 35386
rect 5170 35332 5176 35334
rect 5232 35332 5256 35334
rect 5312 35332 5336 35334
rect 5392 35332 5416 35334
rect 5472 35332 5478 35334
rect 5170 35323 5478 35332
rect 5552 35018 5580 36722
rect 6564 36038 6592 36722
rect 6552 36032 6604 36038
rect 6552 35974 6604 35980
rect 6552 35624 6604 35630
rect 6552 35566 6604 35572
rect 5540 35012 5592 35018
rect 5540 34954 5592 34960
rect 5170 34300 5478 34309
rect 5170 34298 5176 34300
rect 5232 34298 5256 34300
rect 5312 34298 5336 34300
rect 5392 34298 5416 34300
rect 5472 34298 5478 34300
rect 5232 34246 5234 34298
rect 5414 34246 5416 34298
rect 5170 34244 5176 34246
rect 5232 34244 5256 34246
rect 5312 34244 5336 34246
rect 5392 34244 5416 34246
rect 5472 34244 5478 34246
rect 5170 34235 5478 34244
rect 6564 34066 6592 35566
rect 6552 34060 6604 34066
rect 6552 34002 6604 34008
rect 5170 33212 5478 33221
rect 5170 33210 5176 33212
rect 5232 33210 5256 33212
rect 5312 33210 5336 33212
rect 5392 33210 5416 33212
rect 5472 33210 5478 33212
rect 5232 33158 5234 33210
rect 5414 33158 5416 33210
rect 5170 33156 5176 33158
rect 5232 33156 5256 33158
rect 5312 33156 5336 33158
rect 5392 33156 5416 33158
rect 5472 33156 5478 33158
rect 5170 33147 5478 33156
rect 5170 32124 5478 32133
rect 5170 32122 5176 32124
rect 5232 32122 5256 32124
rect 5312 32122 5336 32124
rect 5392 32122 5416 32124
rect 5472 32122 5478 32124
rect 5232 32070 5234 32122
rect 5414 32070 5416 32122
rect 5170 32068 5176 32070
rect 5232 32068 5256 32070
rect 5312 32068 5336 32070
rect 5392 32068 5416 32070
rect 5472 32068 5478 32070
rect 5170 32059 5478 32068
rect 5170 31036 5478 31045
rect 5170 31034 5176 31036
rect 5232 31034 5256 31036
rect 5312 31034 5336 31036
rect 5392 31034 5416 31036
rect 5472 31034 5478 31036
rect 5232 30982 5234 31034
rect 5414 30982 5416 31034
rect 5170 30980 5176 30982
rect 5232 30980 5256 30982
rect 5312 30980 5336 30982
rect 5392 30980 5416 30982
rect 5472 30980 5478 30982
rect 5170 30971 5478 30980
rect 5170 29948 5478 29957
rect 5170 29946 5176 29948
rect 5232 29946 5256 29948
rect 5312 29946 5336 29948
rect 5392 29946 5416 29948
rect 5472 29946 5478 29948
rect 5232 29894 5234 29946
rect 5414 29894 5416 29946
rect 5170 29892 5176 29894
rect 5232 29892 5256 29894
rect 5312 29892 5336 29894
rect 5392 29892 5416 29894
rect 5472 29892 5478 29894
rect 5170 29883 5478 29892
rect 5170 28860 5478 28869
rect 5170 28858 5176 28860
rect 5232 28858 5256 28860
rect 5312 28858 5336 28860
rect 5392 28858 5416 28860
rect 5472 28858 5478 28860
rect 5232 28806 5234 28858
rect 5414 28806 5416 28858
rect 5170 28804 5176 28806
rect 5232 28804 5256 28806
rect 5312 28804 5336 28806
rect 5392 28804 5416 28806
rect 5472 28804 5478 28806
rect 5170 28795 5478 28804
rect 5170 27772 5478 27781
rect 5170 27770 5176 27772
rect 5232 27770 5256 27772
rect 5312 27770 5336 27772
rect 5392 27770 5416 27772
rect 5472 27770 5478 27772
rect 5232 27718 5234 27770
rect 5414 27718 5416 27770
rect 5170 27716 5176 27718
rect 5232 27716 5256 27718
rect 5312 27716 5336 27718
rect 5392 27716 5416 27718
rect 5472 27716 5478 27718
rect 5170 27707 5478 27716
rect 6564 26994 6592 34002
rect 6644 27396 6696 27402
rect 6644 27338 6696 27344
rect 6656 27130 6684 27338
rect 6644 27124 6696 27130
rect 6644 27066 6696 27072
rect 6552 26988 6604 26994
rect 6552 26930 6604 26936
rect 5170 26684 5478 26693
rect 5170 26682 5176 26684
rect 5232 26682 5256 26684
rect 5312 26682 5336 26684
rect 5392 26682 5416 26684
rect 5472 26682 5478 26684
rect 5232 26630 5234 26682
rect 5414 26630 5416 26682
rect 5170 26628 5176 26630
rect 5232 26628 5256 26630
rect 5312 26628 5336 26630
rect 5392 26628 5416 26630
rect 5472 26628 5478 26630
rect 5170 26619 5478 26628
rect 5170 25596 5478 25605
rect 5170 25594 5176 25596
rect 5232 25594 5256 25596
rect 5312 25594 5336 25596
rect 5392 25594 5416 25596
rect 5472 25594 5478 25596
rect 5232 25542 5234 25594
rect 5414 25542 5416 25594
rect 5170 25540 5176 25542
rect 5232 25540 5256 25542
rect 5312 25540 5336 25542
rect 5392 25540 5416 25542
rect 5472 25540 5478 25542
rect 5170 25531 5478 25540
rect 5170 24508 5478 24517
rect 5170 24506 5176 24508
rect 5232 24506 5256 24508
rect 5312 24506 5336 24508
rect 5392 24506 5416 24508
rect 5472 24506 5478 24508
rect 5232 24454 5234 24506
rect 5414 24454 5416 24506
rect 5170 24452 5176 24454
rect 5232 24452 5256 24454
rect 5312 24452 5336 24454
rect 5392 24452 5416 24454
rect 5472 24452 5478 24454
rect 5170 24443 5478 24452
rect 5170 23420 5478 23429
rect 5170 23418 5176 23420
rect 5232 23418 5256 23420
rect 5312 23418 5336 23420
rect 5392 23418 5416 23420
rect 5472 23418 5478 23420
rect 5232 23366 5234 23418
rect 5414 23366 5416 23418
rect 5170 23364 5176 23366
rect 5232 23364 5256 23366
rect 5312 23364 5336 23366
rect 5392 23364 5416 23366
rect 5472 23364 5478 23366
rect 5170 23355 5478 23364
rect 5170 22332 5478 22341
rect 5170 22330 5176 22332
rect 5232 22330 5256 22332
rect 5312 22330 5336 22332
rect 5392 22330 5416 22332
rect 5472 22330 5478 22332
rect 5232 22278 5234 22330
rect 5414 22278 5416 22330
rect 5170 22276 5176 22278
rect 5232 22276 5256 22278
rect 5312 22276 5336 22278
rect 5392 22276 5416 22278
rect 5472 22276 5478 22278
rect 5170 22267 5478 22276
rect 5170 21244 5478 21253
rect 5170 21242 5176 21244
rect 5232 21242 5256 21244
rect 5312 21242 5336 21244
rect 5392 21242 5416 21244
rect 5472 21242 5478 21244
rect 5232 21190 5234 21242
rect 5414 21190 5416 21242
rect 5170 21188 5176 21190
rect 5232 21188 5256 21190
rect 5312 21188 5336 21190
rect 5392 21188 5416 21190
rect 5472 21188 5478 21190
rect 5170 21179 5478 21188
rect 5170 20156 5478 20165
rect 5170 20154 5176 20156
rect 5232 20154 5256 20156
rect 5312 20154 5336 20156
rect 5392 20154 5416 20156
rect 5472 20154 5478 20156
rect 5232 20102 5234 20154
rect 5414 20102 5416 20154
rect 5170 20100 5176 20102
rect 5232 20100 5256 20102
rect 5312 20100 5336 20102
rect 5392 20100 5416 20102
rect 5472 20100 5478 20102
rect 5170 20091 5478 20100
rect 5170 19068 5478 19077
rect 5170 19066 5176 19068
rect 5232 19066 5256 19068
rect 5312 19066 5336 19068
rect 5392 19066 5416 19068
rect 5472 19066 5478 19068
rect 5232 19014 5234 19066
rect 5414 19014 5416 19066
rect 5170 19012 5176 19014
rect 5232 19012 5256 19014
rect 5312 19012 5336 19014
rect 5392 19012 5416 19014
rect 5472 19012 5478 19014
rect 5170 19003 5478 19012
rect 5170 17980 5478 17989
rect 5170 17978 5176 17980
rect 5232 17978 5256 17980
rect 5312 17978 5336 17980
rect 5392 17978 5416 17980
rect 5472 17978 5478 17980
rect 5232 17926 5234 17978
rect 5414 17926 5416 17978
rect 5170 17924 5176 17926
rect 5232 17924 5256 17926
rect 5312 17924 5336 17926
rect 5392 17924 5416 17926
rect 5472 17924 5478 17926
rect 5170 17915 5478 17924
rect 5170 16892 5478 16901
rect 5170 16890 5176 16892
rect 5232 16890 5256 16892
rect 5312 16890 5336 16892
rect 5392 16890 5416 16892
rect 5472 16890 5478 16892
rect 5232 16838 5234 16890
rect 5414 16838 5416 16890
rect 5170 16836 5176 16838
rect 5232 16836 5256 16838
rect 5312 16836 5336 16838
rect 5392 16836 5416 16838
rect 5472 16836 5478 16838
rect 5170 16827 5478 16836
rect 5170 15804 5478 15813
rect 5170 15802 5176 15804
rect 5232 15802 5256 15804
rect 5312 15802 5336 15804
rect 5392 15802 5416 15804
rect 5472 15802 5478 15804
rect 5232 15750 5234 15802
rect 5414 15750 5416 15802
rect 5170 15748 5176 15750
rect 5232 15748 5256 15750
rect 5312 15748 5336 15750
rect 5392 15748 5416 15750
rect 5472 15748 5478 15750
rect 5170 15739 5478 15748
rect 5170 14716 5478 14725
rect 5170 14714 5176 14716
rect 5232 14714 5256 14716
rect 5312 14714 5336 14716
rect 5392 14714 5416 14716
rect 5472 14714 5478 14716
rect 5232 14662 5234 14714
rect 5414 14662 5416 14714
rect 5170 14660 5176 14662
rect 5232 14660 5256 14662
rect 5312 14660 5336 14662
rect 5392 14660 5416 14662
rect 5472 14660 5478 14662
rect 5170 14651 5478 14660
rect 5170 13628 5478 13637
rect 5170 13626 5176 13628
rect 5232 13626 5256 13628
rect 5312 13626 5336 13628
rect 5392 13626 5416 13628
rect 5472 13626 5478 13628
rect 5232 13574 5234 13626
rect 5414 13574 5416 13626
rect 5170 13572 5176 13574
rect 5232 13572 5256 13574
rect 5312 13572 5336 13574
rect 5392 13572 5416 13574
rect 5472 13572 5478 13574
rect 5170 13563 5478 13572
rect 5170 12540 5478 12549
rect 5170 12538 5176 12540
rect 5232 12538 5256 12540
rect 5312 12538 5336 12540
rect 5392 12538 5416 12540
rect 5472 12538 5478 12540
rect 5232 12486 5234 12538
rect 5414 12486 5416 12538
rect 5170 12484 5176 12486
rect 5232 12484 5256 12486
rect 5312 12484 5336 12486
rect 5392 12484 5416 12486
rect 5472 12484 5478 12486
rect 5170 12475 5478 12484
rect 5170 11452 5478 11461
rect 5170 11450 5176 11452
rect 5232 11450 5256 11452
rect 5312 11450 5336 11452
rect 5392 11450 5416 11452
rect 5472 11450 5478 11452
rect 5232 11398 5234 11450
rect 5414 11398 5416 11450
rect 5170 11396 5176 11398
rect 5232 11396 5256 11398
rect 5312 11396 5336 11398
rect 5392 11396 5416 11398
rect 5472 11396 5478 11398
rect 5170 11387 5478 11396
rect 5170 10364 5478 10373
rect 5170 10362 5176 10364
rect 5232 10362 5256 10364
rect 5312 10362 5336 10364
rect 5392 10362 5416 10364
rect 5472 10362 5478 10364
rect 5232 10310 5234 10362
rect 5414 10310 5416 10362
rect 5170 10308 5176 10310
rect 5232 10308 5256 10310
rect 5312 10308 5336 10310
rect 5392 10308 5416 10310
rect 5472 10308 5478 10310
rect 5170 10299 5478 10308
rect 5170 9276 5478 9285
rect 5170 9274 5176 9276
rect 5232 9274 5256 9276
rect 5312 9274 5336 9276
rect 5392 9274 5416 9276
rect 5472 9274 5478 9276
rect 5232 9222 5234 9274
rect 5414 9222 5416 9274
rect 5170 9220 5176 9222
rect 5232 9220 5256 9222
rect 5312 9220 5336 9222
rect 5392 9220 5416 9222
rect 5472 9220 5478 9222
rect 5170 9211 5478 9220
rect 5170 8188 5478 8197
rect 5170 8186 5176 8188
rect 5232 8186 5256 8188
rect 5312 8186 5336 8188
rect 5392 8186 5416 8188
rect 5472 8186 5478 8188
rect 5232 8134 5234 8186
rect 5414 8134 5416 8186
rect 5170 8132 5176 8134
rect 5232 8132 5256 8134
rect 5312 8132 5336 8134
rect 5392 8132 5416 8134
rect 5472 8132 5478 8134
rect 5170 8123 5478 8132
rect 7392 7954 7420 36722
rect 9140 36174 9168 37946
rect 9324 37806 9352 39374
rect 14004 39374 14056 39380
rect 13726 39335 13782 39344
rect 13452 39296 13504 39302
rect 13452 39238 13504 39244
rect 9390 39196 9698 39205
rect 9390 39194 9396 39196
rect 9452 39194 9476 39196
rect 9532 39194 9556 39196
rect 9612 39194 9636 39196
rect 9692 39194 9698 39196
rect 9452 39142 9454 39194
rect 9634 39142 9636 39194
rect 9390 39140 9396 39142
rect 9452 39140 9476 39142
rect 9532 39140 9556 39142
rect 9612 39140 9636 39142
rect 9692 39140 9698 39142
rect 9390 39131 9698 39140
rect 9390 38108 9698 38117
rect 9390 38106 9396 38108
rect 9452 38106 9476 38108
rect 9532 38106 9556 38108
rect 9612 38106 9636 38108
rect 9692 38106 9698 38108
rect 9452 38054 9454 38106
rect 9634 38054 9636 38106
rect 9390 38052 9396 38054
rect 9452 38052 9476 38054
rect 9532 38052 9556 38054
rect 9612 38052 9636 38054
rect 9692 38052 9698 38054
rect 9390 38043 9698 38052
rect 9312 37800 9364 37806
rect 9312 37742 9364 37748
rect 9390 37020 9698 37029
rect 9390 37018 9396 37020
rect 9452 37018 9476 37020
rect 9532 37018 9556 37020
rect 9612 37018 9636 37020
rect 9692 37018 9698 37020
rect 9452 36966 9454 37018
rect 9634 36966 9636 37018
rect 9390 36964 9396 36966
rect 9452 36964 9476 36966
rect 9532 36964 9556 36966
rect 9612 36964 9636 36966
rect 9692 36964 9698 36966
rect 9390 36955 9698 36964
rect 9128 36168 9180 36174
rect 9128 36110 9180 36116
rect 9390 35932 9698 35941
rect 9390 35930 9396 35932
rect 9452 35930 9476 35932
rect 9532 35930 9556 35932
rect 9612 35930 9636 35932
rect 9692 35930 9698 35932
rect 9452 35878 9454 35930
rect 9634 35878 9636 35930
rect 9390 35876 9396 35878
rect 9452 35876 9476 35878
rect 9532 35876 9556 35878
rect 9612 35876 9636 35878
rect 9692 35876 9698 35878
rect 9390 35867 9698 35876
rect 9390 34844 9698 34853
rect 9390 34842 9396 34844
rect 9452 34842 9476 34844
rect 9532 34842 9556 34844
rect 9612 34842 9636 34844
rect 9692 34842 9698 34844
rect 9452 34790 9454 34842
rect 9634 34790 9636 34842
rect 9390 34788 9396 34790
rect 9452 34788 9476 34790
rect 9532 34788 9556 34790
rect 9612 34788 9636 34790
rect 9692 34788 9698 34790
rect 9390 34779 9698 34788
rect 9390 33756 9698 33765
rect 9390 33754 9396 33756
rect 9452 33754 9476 33756
rect 9532 33754 9556 33756
rect 9612 33754 9636 33756
rect 9692 33754 9698 33756
rect 9452 33702 9454 33754
rect 9634 33702 9636 33754
rect 9390 33700 9396 33702
rect 9452 33700 9476 33702
rect 9532 33700 9556 33702
rect 9612 33700 9636 33702
rect 9692 33700 9698 33702
rect 9390 33691 9698 33700
rect 13464 33046 13492 39238
rect 14016 38962 14044 39374
rect 14464 39364 14516 39370
rect 14464 39306 14516 39312
rect 14004 38956 14056 38962
rect 14004 38898 14056 38904
rect 14372 38820 14424 38826
rect 14372 38762 14424 38768
rect 13611 38652 13919 38661
rect 13611 38650 13617 38652
rect 13673 38650 13697 38652
rect 13753 38650 13777 38652
rect 13833 38650 13857 38652
rect 13913 38650 13919 38652
rect 13673 38598 13675 38650
rect 13855 38598 13857 38650
rect 13611 38596 13617 38598
rect 13673 38596 13697 38598
rect 13753 38596 13777 38598
rect 13833 38596 13857 38598
rect 13913 38596 13919 38598
rect 13611 38587 13919 38596
rect 14384 38350 14412 38762
rect 14476 38554 14504 39306
rect 16132 38894 16160 41200
rect 16856 39432 16908 39438
rect 16856 39374 16908 39380
rect 17316 39432 17368 39438
rect 17316 39374 17368 39380
rect 16580 39296 16632 39302
rect 16580 39238 16632 39244
rect 15200 38888 15252 38894
rect 15200 38830 15252 38836
rect 16120 38888 16172 38894
rect 16120 38830 16172 38836
rect 15212 38554 15240 38830
rect 15660 38820 15712 38826
rect 15660 38762 15712 38768
rect 14464 38548 14516 38554
rect 14464 38490 14516 38496
rect 15200 38548 15252 38554
rect 15200 38490 15252 38496
rect 14280 38344 14332 38350
rect 14280 38286 14332 38292
rect 14372 38344 14424 38350
rect 14372 38286 14424 38292
rect 13611 37564 13919 37573
rect 13611 37562 13617 37564
rect 13673 37562 13697 37564
rect 13753 37562 13777 37564
rect 13833 37562 13857 37564
rect 13913 37562 13919 37564
rect 13673 37510 13675 37562
rect 13855 37510 13857 37562
rect 13611 37508 13617 37510
rect 13673 37508 13697 37510
rect 13753 37508 13777 37510
rect 13833 37508 13857 37510
rect 13913 37508 13919 37510
rect 13611 37499 13919 37508
rect 14292 37466 14320 38286
rect 15672 37874 15700 38762
rect 16028 38480 16080 38486
rect 16028 38422 16080 38428
rect 15660 37868 15712 37874
rect 15660 37810 15712 37816
rect 16040 37670 16068 38422
rect 16592 38418 16620 39238
rect 16672 38752 16724 38758
rect 16672 38694 16724 38700
rect 16580 38412 16632 38418
rect 16580 38354 16632 38360
rect 16396 37868 16448 37874
rect 16396 37810 16448 37816
rect 16028 37664 16080 37670
rect 16028 37606 16080 37612
rect 16120 37664 16172 37670
rect 16120 37606 16172 37612
rect 14280 37460 14332 37466
rect 14280 37402 14332 37408
rect 15292 37460 15344 37466
rect 15292 37402 15344 37408
rect 14292 37126 14320 37402
rect 14280 37120 14332 37126
rect 14280 37062 14332 37068
rect 13611 36476 13919 36485
rect 13611 36474 13617 36476
rect 13673 36474 13697 36476
rect 13753 36474 13777 36476
rect 13833 36474 13857 36476
rect 13913 36474 13919 36476
rect 13673 36422 13675 36474
rect 13855 36422 13857 36474
rect 13611 36420 13617 36422
rect 13673 36420 13697 36422
rect 13753 36420 13777 36422
rect 13833 36420 13857 36422
rect 13913 36420 13919 36422
rect 13611 36411 13919 36420
rect 13611 35388 13919 35397
rect 13611 35386 13617 35388
rect 13673 35386 13697 35388
rect 13753 35386 13777 35388
rect 13833 35386 13857 35388
rect 13913 35386 13919 35388
rect 13673 35334 13675 35386
rect 13855 35334 13857 35386
rect 13611 35332 13617 35334
rect 13673 35332 13697 35334
rect 13753 35332 13777 35334
rect 13833 35332 13857 35334
rect 13913 35332 13919 35334
rect 13611 35323 13919 35332
rect 13611 34300 13919 34309
rect 13611 34298 13617 34300
rect 13673 34298 13697 34300
rect 13753 34298 13777 34300
rect 13833 34298 13857 34300
rect 13913 34298 13919 34300
rect 13673 34246 13675 34298
rect 13855 34246 13857 34298
rect 13611 34244 13617 34246
rect 13673 34244 13697 34246
rect 13753 34244 13777 34246
rect 13833 34244 13857 34246
rect 13913 34244 13919 34246
rect 13611 34235 13919 34244
rect 13611 33212 13919 33221
rect 13611 33210 13617 33212
rect 13673 33210 13697 33212
rect 13753 33210 13777 33212
rect 13833 33210 13857 33212
rect 13913 33210 13919 33212
rect 13673 33158 13675 33210
rect 13855 33158 13857 33210
rect 13611 33156 13617 33158
rect 13673 33156 13697 33158
rect 13753 33156 13777 33158
rect 13833 33156 13857 33158
rect 13913 33156 13919 33158
rect 13611 33147 13919 33156
rect 13452 33040 13504 33046
rect 13452 32982 13504 32988
rect 9390 32668 9698 32677
rect 9390 32666 9396 32668
rect 9452 32666 9476 32668
rect 9532 32666 9556 32668
rect 9612 32666 9636 32668
rect 9692 32666 9698 32668
rect 9452 32614 9454 32666
rect 9634 32614 9636 32666
rect 9390 32612 9396 32614
rect 9452 32612 9476 32614
rect 9532 32612 9556 32614
rect 9612 32612 9636 32614
rect 9692 32612 9698 32614
rect 9390 32603 9698 32612
rect 13611 32124 13919 32133
rect 13611 32122 13617 32124
rect 13673 32122 13697 32124
rect 13753 32122 13777 32124
rect 13833 32122 13857 32124
rect 13913 32122 13919 32124
rect 13673 32070 13675 32122
rect 13855 32070 13857 32122
rect 13611 32068 13617 32070
rect 13673 32068 13697 32070
rect 13753 32068 13777 32070
rect 13833 32068 13857 32070
rect 13913 32068 13919 32070
rect 13611 32059 13919 32068
rect 9390 31580 9698 31589
rect 9390 31578 9396 31580
rect 9452 31578 9476 31580
rect 9532 31578 9556 31580
rect 9612 31578 9636 31580
rect 9692 31578 9698 31580
rect 9452 31526 9454 31578
rect 9634 31526 9636 31578
rect 9390 31524 9396 31526
rect 9452 31524 9476 31526
rect 9532 31524 9556 31526
rect 9612 31524 9636 31526
rect 9692 31524 9698 31526
rect 9390 31515 9698 31524
rect 13611 31036 13919 31045
rect 13611 31034 13617 31036
rect 13673 31034 13697 31036
rect 13753 31034 13777 31036
rect 13833 31034 13857 31036
rect 13913 31034 13919 31036
rect 13673 30982 13675 31034
rect 13855 30982 13857 31034
rect 13611 30980 13617 30982
rect 13673 30980 13697 30982
rect 13753 30980 13777 30982
rect 13833 30980 13857 30982
rect 13913 30980 13919 30982
rect 13611 30971 13919 30980
rect 9390 30492 9698 30501
rect 9390 30490 9396 30492
rect 9452 30490 9476 30492
rect 9532 30490 9556 30492
rect 9612 30490 9636 30492
rect 9692 30490 9698 30492
rect 9452 30438 9454 30490
rect 9634 30438 9636 30490
rect 9390 30436 9396 30438
rect 9452 30436 9476 30438
rect 9532 30436 9556 30438
rect 9612 30436 9636 30438
rect 9692 30436 9698 30438
rect 9390 30427 9698 30436
rect 13611 29948 13919 29957
rect 13611 29946 13617 29948
rect 13673 29946 13697 29948
rect 13753 29946 13777 29948
rect 13833 29946 13857 29948
rect 13913 29946 13919 29948
rect 13673 29894 13675 29946
rect 13855 29894 13857 29946
rect 13611 29892 13617 29894
rect 13673 29892 13697 29894
rect 13753 29892 13777 29894
rect 13833 29892 13857 29894
rect 13913 29892 13919 29894
rect 13611 29883 13919 29892
rect 9390 29404 9698 29413
rect 9390 29402 9396 29404
rect 9452 29402 9476 29404
rect 9532 29402 9556 29404
rect 9612 29402 9636 29404
rect 9692 29402 9698 29404
rect 9452 29350 9454 29402
rect 9634 29350 9636 29402
rect 9390 29348 9396 29350
rect 9452 29348 9476 29350
rect 9532 29348 9556 29350
rect 9612 29348 9636 29350
rect 9692 29348 9698 29350
rect 9390 29339 9698 29348
rect 13611 28860 13919 28869
rect 13611 28858 13617 28860
rect 13673 28858 13697 28860
rect 13753 28858 13777 28860
rect 13833 28858 13857 28860
rect 13913 28858 13919 28860
rect 13673 28806 13675 28858
rect 13855 28806 13857 28858
rect 13611 28804 13617 28806
rect 13673 28804 13697 28806
rect 13753 28804 13777 28806
rect 13833 28804 13857 28806
rect 13913 28804 13919 28806
rect 13611 28795 13919 28804
rect 9390 28316 9698 28325
rect 9390 28314 9396 28316
rect 9452 28314 9476 28316
rect 9532 28314 9556 28316
rect 9612 28314 9636 28316
rect 9692 28314 9698 28316
rect 9452 28262 9454 28314
rect 9634 28262 9636 28314
rect 9390 28260 9396 28262
rect 9452 28260 9476 28262
rect 9532 28260 9556 28262
rect 9612 28260 9636 28262
rect 9692 28260 9698 28262
rect 9390 28251 9698 28260
rect 13611 27772 13919 27781
rect 13611 27770 13617 27772
rect 13673 27770 13697 27772
rect 13753 27770 13777 27772
rect 13833 27770 13857 27772
rect 13913 27770 13919 27772
rect 13673 27718 13675 27770
rect 13855 27718 13857 27770
rect 13611 27716 13617 27718
rect 13673 27716 13697 27718
rect 13753 27716 13777 27718
rect 13833 27716 13857 27718
rect 13913 27716 13919 27718
rect 13611 27707 13919 27716
rect 7656 27532 7708 27538
rect 7656 27474 7708 27480
rect 7668 27130 7696 27474
rect 9390 27228 9698 27237
rect 9390 27226 9396 27228
rect 9452 27226 9476 27228
rect 9532 27226 9556 27228
rect 9612 27226 9636 27228
rect 9692 27226 9698 27228
rect 9452 27174 9454 27226
rect 9634 27174 9636 27226
rect 9390 27172 9396 27174
rect 9452 27172 9476 27174
rect 9532 27172 9556 27174
rect 9612 27172 9636 27174
rect 9692 27172 9698 27174
rect 9390 27163 9698 27172
rect 7656 27124 7708 27130
rect 7656 27066 7708 27072
rect 8944 26988 8996 26994
rect 8944 26930 8996 26936
rect 8956 23866 8984 26930
rect 13611 26684 13919 26693
rect 13611 26682 13617 26684
rect 13673 26682 13697 26684
rect 13753 26682 13777 26684
rect 13833 26682 13857 26684
rect 13913 26682 13919 26684
rect 13673 26630 13675 26682
rect 13855 26630 13857 26682
rect 13611 26628 13617 26630
rect 13673 26628 13697 26630
rect 13753 26628 13777 26630
rect 13833 26628 13857 26630
rect 13913 26628 13919 26630
rect 13611 26619 13919 26628
rect 9390 26140 9698 26149
rect 9390 26138 9396 26140
rect 9452 26138 9476 26140
rect 9532 26138 9556 26140
rect 9612 26138 9636 26140
rect 9692 26138 9698 26140
rect 9452 26086 9454 26138
rect 9634 26086 9636 26138
rect 9390 26084 9396 26086
rect 9452 26084 9476 26086
rect 9532 26084 9556 26086
rect 9612 26084 9636 26086
rect 9692 26084 9698 26086
rect 9390 26075 9698 26084
rect 13611 25596 13919 25605
rect 13611 25594 13617 25596
rect 13673 25594 13697 25596
rect 13753 25594 13777 25596
rect 13833 25594 13857 25596
rect 13913 25594 13919 25596
rect 13673 25542 13675 25594
rect 13855 25542 13857 25594
rect 13611 25540 13617 25542
rect 13673 25540 13697 25542
rect 13753 25540 13777 25542
rect 13833 25540 13857 25542
rect 13913 25540 13919 25542
rect 13611 25531 13919 25540
rect 15304 25294 15332 37402
rect 16132 34406 16160 37606
rect 16120 34400 16172 34406
rect 16120 34342 16172 34348
rect 16212 33584 16264 33590
rect 16212 33526 16264 33532
rect 16028 32768 16080 32774
rect 16028 32710 16080 32716
rect 16040 27470 16068 32710
rect 16224 29850 16252 33526
rect 16304 32564 16356 32570
rect 16304 32506 16356 32512
rect 16212 29844 16264 29850
rect 16212 29786 16264 29792
rect 16316 28558 16344 32506
rect 16304 28552 16356 28558
rect 16118 28520 16174 28529
rect 16304 28494 16356 28500
rect 16118 28455 16174 28464
rect 16132 28082 16160 28455
rect 16120 28076 16172 28082
rect 16120 28018 16172 28024
rect 16304 27872 16356 27878
rect 16304 27814 16356 27820
rect 16028 27464 16080 27470
rect 16028 27406 16080 27412
rect 16316 26994 16344 27814
rect 16304 26988 16356 26994
rect 16304 26930 16356 26936
rect 16120 26784 16172 26790
rect 16120 26726 16172 26732
rect 16132 26518 16160 26726
rect 16120 26512 16172 26518
rect 16120 26454 16172 26460
rect 16028 26308 16080 26314
rect 16028 26250 16080 26256
rect 15292 25288 15344 25294
rect 15292 25230 15344 25236
rect 9390 25052 9698 25061
rect 9390 25050 9396 25052
rect 9452 25050 9476 25052
rect 9532 25050 9556 25052
rect 9612 25050 9636 25052
rect 9692 25050 9698 25052
rect 9452 24998 9454 25050
rect 9634 24998 9636 25050
rect 9390 24996 9396 24998
rect 9452 24996 9476 24998
rect 9532 24996 9556 24998
rect 9612 24996 9636 24998
rect 9692 24996 9698 24998
rect 9390 24987 9698 24996
rect 13611 24508 13919 24517
rect 13611 24506 13617 24508
rect 13673 24506 13697 24508
rect 13753 24506 13777 24508
rect 13833 24506 13857 24508
rect 13913 24506 13919 24508
rect 13673 24454 13675 24506
rect 13855 24454 13857 24506
rect 13611 24452 13617 24454
rect 13673 24452 13697 24454
rect 13753 24452 13777 24454
rect 13833 24452 13857 24454
rect 13913 24452 13919 24454
rect 13611 24443 13919 24452
rect 9390 23964 9698 23973
rect 9390 23962 9396 23964
rect 9452 23962 9476 23964
rect 9532 23962 9556 23964
rect 9612 23962 9636 23964
rect 9692 23962 9698 23964
rect 9452 23910 9454 23962
rect 9634 23910 9636 23962
rect 9390 23908 9396 23910
rect 9452 23908 9476 23910
rect 9532 23908 9556 23910
rect 9612 23908 9636 23910
rect 9692 23908 9698 23910
rect 9390 23899 9698 23908
rect 8944 23860 8996 23866
rect 8944 23802 8996 23808
rect 13611 23420 13919 23429
rect 13611 23418 13617 23420
rect 13673 23418 13697 23420
rect 13753 23418 13777 23420
rect 13833 23418 13857 23420
rect 13913 23418 13919 23420
rect 13673 23366 13675 23418
rect 13855 23366 13857 23418
rect 13611 23364 13617 23366
rect 13673 23364 13697 23366
rect 13753 23364 13777 23366
rect 13833 23364 13857 23366
rect 13913 23364 13919 23366
rect 13611 23355 13919 23364
rect 9390 22876 9698 22885
rect 9390 22874 9396 22876
rect 9452 22874 9476 22876
rect 9532 22874 9556 22876
rect 9612 22874 9636 22876
rect 9692 22874 9698 22876
rect 9452 22822 9454 22874
rect 9634 22822 9636 22874
rect 9390 22820 9396 22822
rect 9452 22820 9476 22822
rect 9532 22820 9556 22822
rect 9612 22820 9636 22822
rect 9692 22820 9698 22822
rect 9390 22811 9698 22820
rect 13611 22332 13919 22341
rect 13611 22330 13617 22332
rect 13673 22330 13697 22332
rect 13753 22330 13777 22332
rect 13833 22330 13857 22332
rect 13913 22330 13919 22332
rect 13673 22278 13675 22330
rect 13855 22278 13857 22330
rect 13611 22276 13617 22278
rect 13673 22276 13697 22278
rect 13753 22276 13777 22278
rect 13833 22276 13857 22278
rect 13913 22276 13919 22278
rect 13611 22267 13919 22276
rect 9390 21788 9698 21797
rect 9390 21786 9396 21788
rect 9452 21786 9476 21788
rect 9532 21786 9556 21788
rect 9612 21786 9636 21788
rect 9692 21786 9698 21788
rect 9452 21734 9454 21786
rect 9634 21734 9636 21786
rect 9390 21732 9396 21734
rect 9452 21732 9476 21734
rect 9532 21732 9556 21734
rect 9612 21732 9636 21734
rect 9692 21732 9698 21734
rect 9390 21723 9698 21732
rect 13611 21244 13919 21253
rect 13611 21242 13617 21244
rect 13673 21242 13697 21244
rect 13753 21242 13777 21244
rect 13833 21242 13857 21244
rect 13913 21242 13919 21244
rect 13673 21190 13675 21242
rect 13855 21190 13857 21242
rect 13611 21188 13617 21190
rect 13673 21188 13697 21190
rect 13753 21188 13777 21190
rect 13833 21188 13857 21190
rect 13913 21188 13919 21190
rect 13611 21179 13919 21188
rect 9390 20700 9698 20709
rect 9390 20698 9396 20700
rect 9452 20698 9476 20700
rect 9532 20698 9556 20700
rect 9612 20698 9636 20700
rect 9692 20698 9698 20700
rect 9452 20646 9454 20698
rect 9634 20646 9636 20698
rect 9390 20644 9396 20646
rect 9452 20644 9476 20646
rect 9532 20644 9556 20646
rect 9612 20644 9636 20646
rect 9692 20644 9698 20646
rect 9390 20635 9698 20644
rect 13611 20156 13919 20165
rect 13611 20154 13617 20156
rect 13673 20154 13697 20156
rect 13753 20154 13777 20156
rect 13833 20154 13857 20156
rect 13913 20154 13919 20156
rect 13673 20102 13675 20154
rect 13855 20102 13857 20154
rect 13611 20100 13617 20102
rect 13673 20100 13697 20102
rect 13753 20100 13777 20102
rect 13833 20100 13857 20102
rect 13913 20100 13919 20102
rect 13611 20091 13919 20100
rect 9390 19612 9698 19621
rect 9390 19610 9396 19612
rect 9452 19610 9476 19612
rect 9532 19610 9556 19612
rect 9612 19610 9636 19612
rect 9692 19610 9698 19612
rect 9452 19558 9454 19610
rect 9634 19558 9636 19610
rect 9390 19556 9396 19558
rect 9452 19556 9476 19558
rect 9532 19556 9556 19558
rect 9612 19556 9636 19558
rect 9692 19556 9698 19558
rect 9390 19547 9698 19556
rect 13611 19068 13919 19077
rect 13611 19066 13617 19068
rect 13673 19066 13697 19068
rect 13753 19066 13777 19068
rect 13833 19066 13857 19068
rect 13913 19066 13919 19068
rect 13673 19014 13675 19066
rect 13855 19014 13857 19066
rect 13611 19012 13617 19014
rect 13673 19012 13697 19014
rect 13753 19012 13777 19014
rect 13833 19012 13857 19014
rect 13913 19012 13919 19014
rect 13611 19003 13919 19012
rect 9390 18524 9698 18533
rect 9390 18522 9396 18524
rect 9452 18522 9476 18524
rect 9532 18522 9556 18524
rect 9612 18522 9636 18524
rect 9692 18522 9698 18524
rect 9452 18470 9454 18522
rect 9634 18470 9636 18522
rect 9390 18468 9396 18470
rect 9452 18468 9476 18470
rect 9532 18468 9556 18470
rect 9612 18468 9636 18470
rect 9692 18468 9698 18470
rect 9390 18459 9698 18468
rect 13611 17980 13919 17989
rect 13611 17978 13617 17980
rect 13673 17978 13697 17980
rect 13753 17978 13777 17980
rect 13833 17978 13857 17980
rect 13913 17978 13919 17980
rect 13673 17926 13675 17978
rect 13855 17926 13857 17978
rect 13611 17924 13617 17926
rect 13673 17924 13697 17926
rect 13753 17924 13777 17926
rect 13833 17924 13857 17926
rect 13913 17924 13919 17926
rect 13611 17915 13919 17924
rect 9390 17436 9698 17445
rect 9390 17434 9396 17436
rect 9452 17434 9476 17436
rect 9532 17434 9556 17436
rect 9612 17434 9636 17436
rect 9692 17434 9698 17436
rect 9452 17382 9454 17434
rect 9634 17382 9636 17434
rect 9390 17380 9396 17382
rect 9452 17380 9476 17382
rect 9532 17380 9556 17382
rect 9612 17380 9636 17382
rect 9692 17380 9698 17382
rect 9390 17371 9698 17380
rect 13611 16892 13919 16901
rect 13611 16890 13617 16892
rect 13673 16890 13697 16892
rect 13753 16890 13777 16892
rect 13833 16890 13857 16892
rect 13913 16890 13919 16892
rect 13673 16838 13675 16890
rect 13855 16838 13857 16890
rect 13611 16836 13617 16838
rect 13673 16836 13697 16838
rect 13753 16836 13777 16838
rect 13833 16836 13857 16838
rect 13913 16836 13919 16838
rect 13611 16827 13919 16836
rect 9390 16348 9698 16357
rect 9390 16346 9396 16348
rect 9452 16346 9476 16348
rect 9532 16346 9556 16348
rect 9612 16346 9636 16348
rect 9692 16346 9698 16348
rect 9452 16294 9454 16346
rect 9634 16294 9636 16346
rect 9390 16292 9396 16294
rect 9452 16292 9476 16294
rect 9532 16292 9556 16294
rect 9612 16292 9636 16294
rect 9692 16292 9698 16294
rect 9390 16283 9698 16292
rect 13611 15804 13919 15813
rect 13611 15802 13617 15804
rect 13673 15802 13697 15804
rect 13753 15802 13777 15804
rect 13833 15802 13857 15804
rect 13913 15802 13919 15804
rect 13673 15750 13675 15802
rect 13855 15750 13857 15802
rect 13611 15748 13617 15750
rect 13673 15748 13697 15750
rect 13753 15748 13777 15750
rect 13833 15748 13857 15750
rect 13913 15748 13919 15750
rect 13611 15739 13919 15748
rect 9390 15260 9698 15269
rect 9390 15258 9396 15260
rect 9452 15258 9476 15260
rect 9532 15258 9556 15260
rect 9612 15258 9636 15260
rect 9692 15258 9698 15260
rect 9452 15206 9454 15258
rect 9634 15206 9636 15258
rect 9390 15204 9396 15206
rect 9452 15204 9476 15206
rect 9532 15204 9556 15206
rect 9612 15204 9636 15206
rect 9692 15204 9698 15206
rect 9390 15195 9698 15204
rect 15304 14958 15332 25230
rect 16040 24818 16068 26250
rect 16028 24812 16080 24818
rect 16028 24754 16080 24760
rect 16040 24274 16068 24754
rect 16028 24268 16080 24274
rect 16028 24210 16080 24216
rect 15752 24200 15804 24206
rect 15750 24168 15752 24177
rect 15804 24168 15806 24177
rect 15750 24103 15806 24112
rect 16040 23662 16068 24210
rect 16028 23656 16080 23662
rect 16028 23598 16080 23604
rect 16120 23520 16172 23526
rect 16120 23462 16172 23468
rect 16132 21622 16160 23462
rect 16408 22438 16436 37810
rect 16580 37732 16632 37738
rect 16580 37674 16632 37680
rect 16592 35698 16620 37674
rect 16580 35692 16632 35698
rect 16580 35634 16632 35640
rect 16684 35154 16712 38694
rect 16868 38282 16896 39374
rect 17040 39296 17092 39302
rect 17040 39238 17092 39244
rect 17052 39030 17080 39238
rect 17040 39024 17092 39030
rect 17040 38966 17092 38972
rect 16856 38276 16908 38282
rect 16856 38218 16908 38224
rect 17132 37868 17184 37874
rect 17132 37810 17184 37816
rect 16672 35148 16724 35154
rect 16672 35090 16724 35096
rect 17144 34746 17172 37810
rect 17328 36786 17356 39374
rect 17420 38418 17448 41200
rect 18064 40066 18092 41200
rect 18064 40038 18276 40066
rect 17831 39196 18139 39205
rect 17831 39194 17837 39196
rect 17893 39194 17917 39196
rect 17973 39194 17997 39196
rect 18053 39194 18077 39196
rect 18133 39194 18139 39196
rect 17893 39142 17895 39194
rect 18075 39142 18077 39194
rect 17831 39140 17837 39142
rect 17893 39140 17917 39142
rect 17973 39140 17997 39142
rect 18053 39140 18077 39142
rect 18133 39140 18139 39142
rect 17831 39131 18139 39140
rect 18248 38894 18276 40038
rect 18708 39438 18736 41200
rect 18972 39636 19024 39642
rect 18972 39578 19024 39584
rect 18696 39432 18748 39438
rect 18696 39374 18748 39380
rect 18328 39296 18380 39302
rect 18328 39238 18380 39244
rect 17684 38888 17736 38894
rect 17684 38830 17736 38836
rect 18236 38888 18288 38894
rect 18236 38830 18288 38836
rect 17408 38412 17460 38418
rect 17408 38354 17460 38360
rect 17696 37874 17724 38830
rect 18236 38208 18288 38214
rect 18236 38150 18288 38156
rect 17831 38108 18139 38117
rect 17831 38106 17837 38108
rect 17893 38106 17917 38108
rect 17973 38106 17997 38108
rect 18053 38106 18077 38108
rect 18133 38106 18139 38108
rect 17893 38054 17895 38106
rect 18075 38054 18077 38106
rect 17831 38052 17837 38054
rect 17893 38052 17917 38054
rect 17973 38052 17997 38054
rect 18053 38052 18077 38054
rect 18133 38052 18139 38054
rect 17831 38043 18139 38052
rect 17684 37868 17736 37874
rect 17684 37810 17736 37816
rect 17408 37256 17460 37262
rect 17408 37198 17460 37204
rect 17316 36780 17368 36786
rect 17316 36722 17368 36728
rect 17420 36106 17448 37198
rect 17500 37120 17552 37126
rect 17500 37062 17552 37068
rect 17408 36100 17460 36106
rect 17408 36042 17460 36048
rect 17132 34740 17184 34746
rect 17132 34682 17184 34688
rect 17408 32496 17460 32502
rect 17408 32438 17460 32444
rect 17420 32026 17448 32438
rect 17408 32020 17460 32026
rect 17408 31962 17460 31968
rect 17512 31686 17540 37062
rect 17831 37020 18139 37029
rect 17831 37018 17837 37020
rect 17893 37018 17917 37020
rect 17973 37018 17997 37020
rect 18053 37018 18077 37020
rect 18133 37018 18139 37020
rect 17893 36966 17895 37018
rect 18075 36966 18077 37018
rect 17831 36964 17837 36966
rect 17893 36964 17917 36966
rect 17973 36964 17997 36966
rect 18053 36964 18077 36966
rect 18133 36964 18139 36966
rect 17831 36955 18139 36964
rect 17590 36816 17646 36825
rect 18248 36786 18276 38150
rect 17590 36751 17592 36760
rect 17644 36751 17646 36760
rect 18236 36780 18288 36786
rect 17592 36722 17644 36728
rect 18236 36722 18288 36728
rect 17684 36576 17736 36582
rect 17684 36518 17736 36524
rect 17696 35698 17724 36518
rect 18236 36032 18288 36038
rect 18236 35974 18288 35980
rect 17831 35932 18139 35941
rect 17831 35930 17837 35932
rect 17893 35930 17917 35932
rect 17973 35930 17997 35932
rect 18053 35930 18077 35932
rect 18133 35930 18139 35932
rect 17893 35878 17895 35930
rect 18075 35878 18077 35930
rect 17831 35876 17837 35878
rect 17893 35876 17917 35878
rect 17973 35876 17997 35878
rect 18053 35876 18077 35878
rect 18133 35876 18139 35878
rect 17831 35867 18139 35876
rect 18248 35766 18276 35974
rect 18236 35760 18288 35766
rect 18236 35702 18288 35708
rect 17684 35692 17736 35698
rect 17684 35634 17736 35640
rect 17592 35488 17644 35494
rect 17592 35430 17644 35436
rect 17604 34649 17632 35430
rect 18340 35086 18368 39238
rect 18604 38344 18656 38350
rect 18604 38286 18656 38292
rect 18616 37942 18644 38286
rect 18696 38004 18748 38010
rect 18696 37946 18748 37952
rect 18604 37936 18656 37942
rect 18604 37878 18656 37884
rect 18616 37262 18644 37878
rect 18708 37806 18736 37946
rect 18984 37874 19012 39578
rect 19156 39432 19208 39438
rect 19156 39374 19208 39380
rect 19168 38962 19196 39374
rect 19156 38956 19208 38962
rect 19156 38898 19208 38904
rect 19996 38894 20024 41200
rect 20352 40044 20404 40050
rect 20352 39986 20404 39992
rect 20260 39432 20312 39438
rect 20260 39374 20312 39380
rect 19340 38888 19392 38894
rect 19340 38830 19392 38836
rect 19984 38888 20036 38894
rect 19984 38830 20036 38836
rect 19352 38554 19380 38830
rect 19340 38548 19392 38554
rect 19340 38490 19392 38496
rect 20272 38418 20300 39374
rect 20260 38412 20312 38418
rect 20260 38354 20312 38360
rect 20168 38276 20220 38282
rect 20168 38218 20220 38224
rect 20180 38010 20208 38218
rect 20168 38004 20220 38010
rect 20168 37946 20220 37952
rect 18972 37868 19024 37874
rect 18972 37810 19024 37816
rect 18696 37800 18748 37806
rect 18696 37742 18748 37748
rect 18604 37256 18656 37262
rect 18604 37198 18656 37204
rect 18708 36786 18736 37742
rect 20364 37466 20392 39986
rect 20536 38820 20588 38826
rect 20536 38762 20588 38768
rect 20444 37868 20496 37874
rect 20444 37810 20496 37816
rect 20352 37460 20404 37466
rect 20352 37402 20404 37408
rect 19248 37392 19300 37398
rect 19432 37392 19484 37398
rect 19300 37340 19432 37346
rect 19248 37334 19484 37340
rect 19156 37324 19208 37330
rect 19260 37318 19472 37334
rect 19156 37266 19208 37272
rect 18880 37256 18932 37262
rect 18878 37224 18880 37233
rect 18932 37224 18934 37233
rect 18878 37159 18934 37168
rect 19064 37120 19116 37126
rect 19064 37062 19116 37068
rect 18696 36780 18748 36786
rect 18696 36722 18748 36728
rect 18972 36576 19024 36582
rect 18972 36518 19024 36524
rect 18420 36168 18472 36174
rect 18420 36110 18472 36116
rect 18432 35290 18460 36110
rect 18420 35284 18472 35290
rect 18420 35226 18472 35232
rect 18328 35080 18380 35086
rect 18328 35022 18380 35028
rect 18328 34944 18380 34950
rect 18328 34886 18380 34892
rect 17831 34844 18139 34853
rect 17831 34842 17837 34844
rect 17893 34842 17917 34844
rect 17973 34842 17997 34844
rect 18053 34842 18077 34844
rect 18133 34842 18139 34844
rect 17893 34790 17895 34842
rect 18075 34790 18077 34842
rect 17831 34788 17837 34790
rect 17893 34788 17917 34790
rect 17973 34788 17997 34790
rect 18053 34788 18077 34790
rect 18133 34788 18139 34790
rect 17831 34779 18139 34788
rect 18236 34672 18288 34678
rect 17590 34640 17646 34649
rect 18236 34614 18288 34620
rect 17590 34575 17646 34584
rect 17831 33756 18139 33765
rect 17831 33754 17837 33756
rect 17893 33754 17917 33756
rect 17973 33754 17997 33756
rect 18053 33754 18077 33756
rect 18133 33754 18139 33756
rect 17893 33702 17895 33754
rect 18075 33702 18077 33754
rect 17831 33700 17837 33702
rect 17893 33700 17917 33702
rect 17973 33700 17997 33702
rect 18053 33700 18077 33702
rect 18133 33700 18139 33702
rect 17831 33691 18139 33700
rect 18248 33522 18276 34614
rect 18340 33998 18368 34886
rect 18696 34604 18748 34610
rect 18696 34546 18748 34552
rect 18708 34202 18736 34546
rect 18696 34196 18748 34202
rect 18696 34138 18748 34144
rect 18328 33992 18380 33998
rect 18328 33934 18380 33940
rect 18420 33856 18472 33862
rect 18420 33798 18472 33804
rect 18432 33522 18460 33798
rect 18984 33522 19012 36518
rect 19076 33658 19104 37062
rect 19064 33652 19116 33658
rect 19064 33594 19116 33600
rect 18236 33516 18288 33522
rect 18236 33458 18288 33464
rect 18420 33516 18472 33522
rect 18420 33458 18472 33464
rect 18972 33516 19024 33522
rect 18972 33458 19024 33464
rect 17831 32668 18139 32677
rect 17831 32666 17837 32668
rect 17893 32666 17917 32668
rect 17973 32666 17997 32668
rect 18053 32666 18077 32668
rect 18133 32666 18139 32668
rect 17893 32614 17895 32666
rect 18075 32614 18077 32666
rect 17831 32612 17837 32614
rect 17893 32612 17917 32614
rect 17973 32612 17997 32614
rect 18053 32612 18077 32614
rect 18133 32612 18139 32614
rect 17831 32603 18139 32612
rect 18248 32434 18276 33458
rect 18420 32972 18472 32978
rect 18420 32914 18472 32920
rect 18236 32428 18288 32434
rect 18236 32370 18288 32376
rect 17592 32020 17644 32026
rect 17592 31962 17644 31968
rect 17500 31680 17552 31686
rect 17500 31622 17552 31628
rect 17604 31346 17632 31962
rect 17684 31952 17736 31958
rect 17684 31894 17736 31900
rect 17592 31340 17644 31346
rect 17592 31282 17644 31288
rect 17500 30048 17552 30054
rect 17500 29990 17552 29996
rect 17512 29782 17540 29990
rect 17500 29776 17552 29782
rect 17500 29718 17552 29724
rect 16856 29640 16908 29646
rect 16856 29582 16908 29588
rect 16672 29504 16724 29510
rect 16672 29446 16724 29452
rect 16684 29306 16712 29446
rect 16672 29300 16724 29306
rect 16672 29242 16724 29248
rect 16868 29209 16896 29582
rect 17592 29572 17644 29578
rect 17592 29514 17644 29520
rect 16854 29200 16910 29209
rect 17604 29170 17632 29514
rect 16854 29135 16910 29144
rect 17592 29164 17644 29170
rect 17592 29106 17644 29112
rect 17590 28928 17646 28937
rect 17590 28863 17646 28872
rect 17604 28558 17632 28863
rect 17592 28552 17644 28558
rect 17592 28494 17644 28500
rect 17132 28484 17184 28490
rect 17132 28426 17184 28432
rect 16764 28416 16816 28422
rect 16764 28358 16816 28364
rect 16776 28218 16804 28358
rect 16764 28212 16816 28218
rect 16764 28154 16816 28160
rect 17144 28082 17172 28426
rect 17696 28150 17724 31894
rect 18248 31754 18276 32370
rect 18432 31754 18460 32914
rect 18880 32904 18932 32910
rect 18880 32846 18932 32852
rect 18892 32570 18920 32846
rect 18880 32564 18932 32570
rect 18880 32506 18932 32512
rect 19064 32224 19116 32230
rect 19064 32166 19116 32172
rect 19076 31822 19104 32166
rect 19064 31816 19116 31822
rect 19064 31758 19116 31764
rect 18248 31726 18460 31754
rect 17831 31580 18139 31589
rect 17831 31578 17837 31580
rect 17893 31578 17917 31580
rect 17973 31578 17997 31580
rect 18053 31578 18077 31580
rect 18133 31578 18139 31580
rect 17893 31526 17895 31578
rect 18075 31526 18077 31578
rect 17831 31524 17837 31526
rect 17893 31524 17917 31526
rect 17973 31524 17997 31526
rect 18053 31524 18077 31526
rect 18133 31524 18139 31526
rect 17831 31515 18139 31524
rect 18236 31272 18288 31278
rect 18432 31226 18460 31726
rect 18512 31748 18564 31754
rect 18512 31690 18564 31696
rect 18288 31220 18460 31226
rect 18236 31214 18460 31220
rect 18248 31198 18460 31214
rect 17776 30932 17828 30938
rect 17776 30874 17828 30880
rect 17788 30734 17816 30874
rect 17776 30728 17828 30734
rect 17776 30670 17828 30676
rect 17831 30492 18139 30501
rect 17831 30490 17837 30492
rect 17893 30490 17917 30492
rect 17973 30490 17997 30492
rect 18053 30490 18077 30492
rect 18133 30490 18139 30492
rect 17893 30438 17895 30490
rect 18075 30438 18077 30490
rect 17831 30436 17837 30438
rect 17893 30436 17917 30438
rect 17973 30436 17997 30438
rect 18053 30436 18077 30438
rect 18133 30436 18139 30438
rect 17831 30427 18139 30436
rect 18248 30274 18276 31198
rect 18420 30864 18472 30870
rect 18420 30806 18472 30812
rect 18156 30258 18276 30274
rect 18144 30252 18276 30258
rect 18196 30246 18276 30252
rect 18144 30194 18196 30200
rect 17866 29744 17922 29753
rect 17866 29679 17922 29688
rect 17880 29646 17908 29679
rect 18432 29646 18460 30806
rect 18524 30802 18552 31690
rect 18604 31340 18656 31346
rect 18604 31282 18656 31288
rect 18616 31142 18644 31282
rect 18604 31136 18656 31142
rect 18604 31078 18656 31084
rect 18512 30796 18564 30802
rect 18512 30738 18564 30744
rect 18524 30666 18552 30738
rect 18512 30660 18564 30666
rect 18512 30602 18564 30608
rect 18512 30048 18564 30054
rect 18512 29990 18564 29996
rect 17868 29640 17920 29646
rect 17868 29582 17920 29588
rect 18420 29640 18472 29646
rect 18420 29582 18472 29588
rect 17831 29404 18139 29413
rect 17831 29402 17837 29404
rect 17893 29402 17917 29404
rect 17973 29402 17997 29404
rect 18053 29402 18077 29404
rect 18133 29402 18139 29404
rect 17893 29350 17895 29402
rect 18075 29350 18077 29402
rect 17831 29348 17837 29350
rect 17893 29348 17917 29350
rect 17973 29348 17997 29350
rect 18053 29348 18077 29350
rect 18133 29348 18139 29350
rect 17831 29339 18139 29348
rect 18420 29232 18472 29238
rect 18326 29200 18382 29209
rect 18144 29164 18196 29170
rect 18420 29174 18472 29180
rect 18326 29135 18382 29144
rect 18144 29106 18196 29112
rect 18156 28558 18184 29106
rect 18340 28665 18368 29135
rect 18326 28656 18382 28665
rect 18326 28591 18382 28600
rect 18144 28552 18196 28558
rect 18196 28512 18276 28540
rect 18144 28494 18196 28500
rect 17831 28316 18139 28325
rect 17831 28314 17837 28316
rect 17893 28314 17917 28316
rect 17973 28314 17997 28316
rect 18053 28314 18077 28316
rect 18133 28314 18139 28316
rect 17893 28262 17895 28314
rect 18075 28262 18077 28314
rect 17831 28260 17837 28262
rect 17893 28260 17917 28262
rect 17973 28260 17997 28262
rect 18053 28260 18077 28262
rect 18133 28260 18139 28262
rect 17831 28251 18139 28260
rect 17684 28144 17736 28150
rect 17604 28104 17684 28132
rect 17040 28076 17092 28082
rect 17040 28018 17092 28024
rect 17132 28076 17184 28082
rect 17132 28018 17184 28024
rect 17052 27674 17080 28018
rect 17408 27872 17460 27878
rect 17408 27814 17460 27820
rect 17040 27668 17092 27674
rect 17040 27610 17092 27616
rect 17040 27532 17092 27538
rect 17040 27474 17092 27480
rect 16764 27056 16816 27062
rect 16764 26998 16816 27004
rect 16776 26382 16804 26998
rect 17052 26994 17080 27474
rect 17420 27470 17448 27814
rect 17604 27606 17632 28104
rect 17736 28104 17908 28132
rect 17684 28086 17736 28092
rect 17592 27600 17644 27606
rect 17592 27542 17644 27548
rect 17880 27538 17908 28104
rect 18248 27946 18276 28512
rect 18432 28150 18460 29174
rect 18524 28506 18552 29990
rect 18616 29696 18644 31078
rect 19076 30734 19104 31758
rect 19168 31686 19196 37266
rect 20456 37262 20484 37810
rect 20444 37256 20496 37262
rect 20444 37198 20496 37204
rect 19340 36780 19392 36786
rect 19340 36722 19392 36728
rect 19352 36310 19380 36722
rect 20456 36718 20484 37198
rect 20548 36786 20576 38762
rect 20640 38418 20668 41200
rect 22052 39740 22360 39749
rect 22052 39738 22058 39740
rect 22114 39738 22138 39740
rect 22194 39738 22218 39740
rect 22274 39738 22298 39740
rect 22354 39738 22360 39740
rect 22114 39686 22116 39738
rect 22296 39686 22298 39738
rect 22052 39684 22058 39686
rect 22114 39684 22138 39686
rect 22194 39684 22218 39686
rect 22274 39684 22298 39686
rect 22354 39684 22360 39686
rect 22052 39675 22360 39684
rect 21456 39432 21508 39438
rect 21456 39374 21508 39380
rect 22100 39432 22152 39438
rect 22100 39374 22152 39380
rect 21468 39001 21496 39374
rect 21454 38992 21510 39001
rect 21454 38927 21510 38936
rect 22112 38842 22140 39374
rect 22192 39296 22244 39302
rect 22192 39238 22244 39244
rect 22204 39030 22232 39238
rect 22192 39024 22244 39030
rect 22192 38966 22244 38972
rect 22572 38894 22600 41200
rect 23940 39840 23992 39846
rect 23940 39782 23992 39788
rect 23952 39642 23980 39782
rect 23940 39636 23992 39642
rect 23940 39578 23992 39584
rect 23388 39432 23440 39438
rect 23388 39374 23440 39380
rect 23848 39432 23900 39438
rect 23848 39374 23900 39380
rect 23400 39098 23428 39374
rect 23388 39092 23440 39098
rect 23388 39034 23440 39040
rect 21928 38814 22140 38842
rect 22376 38888 22428 38894
rect 22376 38830 22428 38836
rect 22560 38888 22612 38894
rect 22560 38830 22612 38836
rect 20628 38412 20680 38418
rect 20628 38354 20680 38360
rect 21362 38312 21418 38321
rect 21362 38247 21418 38256
rect 21180 37664 21232 37670
rect 21180 37606 21232 37612
rect 20720 37120 20772 37126
rect 20720 37062 20772 37068
rect 20732 36922 20760 37062
rect 20720 36916 20772 36922
rect 20720 36858 20772 36864
rect 20536 36780 20588 36786
rect 20536 36722 20588 36728
rect 20444 36712 20496 36718
rect 20628 36712 20680 36718
rect 20444 36654 20496 36660
rect 20626 36680 20628 36689
rect 20680 36680 20682 36689
rect 20626 36615 20682 36624
rect 20536 36576 20588 36582
rect 20536 36518 20588 36524
rect 19340 36304 19392 36310
rect 19340 36246 19392 36252
rect 19800 36168 19852 36174
rect 19800 36110 19852 36116
rect 19812 35601 19840 36110
rect 19892 36032 19944 36038
rect 19892 35974 19944 35980
rect 20168 36032 20220 36038
rect 20168 35974 20220 35980
rect 19798 35592 19854 35601
rect 19798 35527 19854 35536
rect 19248 35488 19300 35494
rect 19248 35430 19300 35436
rect 19524 35488 19576 35494
rect 19524 35430 19576 35436
rect 19260 34610 19288 35430
rect 19338 35184 19394 35193
rect 19338 35119 19394 35128
rect 19352 34678 19380 35119
rect 19536 35086 19564 35430
rect 19524 35080 19576 35086
rect 19524 35022 19576 35028
rect 19800 34944 19852 34950
rect 19800 34886 19852 34892
rect 19340 34672 19392 34678
rect 19340 34614 19392 34620
rect 19248 34604 19300 34610
rect 19248 34546 19300 34552
rect 19260 32978 19288 34546
rect 19812 33998 19840 34886
rect 19800 33992 19852 33998
rect 19800 33934 19852 33940
rect 19800 33856 19852 33862
rect 19800 33798 19852 33804
rect 19524 33312 19576 33318
rect 19524 33254 19576 33260
rect 19432 33040 19484 33046
rect 19430 33008 19432 33017
rect 19484 33008 19486 33017
rect 19248 32972 19300 32978
rect 19430 32943 19486 32952
rect 19248 32914 19300 32920
rect 19260 31958 19288 32914
rect 19340 32224 19392 32230
rect 19340 32166 19392 32172
rect 19248 31952 19300 31958
rect 19248 31894 19300 31900
rect 19156 31680 19208 31686
rect 19156 31622 19208 31628
rect 19248 31136 19300 31142
rect 19248 31078 19300 31084
rect 19260 30802 19288 31078
rect 19352 30870 19380 32166
rect 19536 31890 19564 33254
rect 19708 33108 19760 33114
rect 19708 33050 19760 33056
rect 19616 32360 19668 32366
rect 19616 32302 19668 32308
rect 19524 31884 19576 31890
rect 19524 31826 19576 31832
rect 19536 30938 19564 31826
rect 19628 31822 19656 32302
rect 19616 31816 19668 31822
rect 19616 31758 19668 31764
rect 19524 30932 19576 30938
rect 19524 30874 19576 30880
rect 19340 30864 19392 30870
rect 19340 30806 19392 30812
rect 19248 30796 19300 30802
rect 19248 30738 19300 30744
rect 19064 30728 19116 30734
rect 19064 30670 19116 30676
rect 19432 30728 19484 30734
rect 19432 30670 19484 30676
rect 18972 30592 19024 30598
rect 18972 30534 19024 30540
rect 18984 30326 19012 30534
rect 18972 30320 19024 30326
rect 18972 30262 19024 30268
rect 18788 30048 18840 30054
rect 18788 29990 18840 29996
rect 18696 29708 18748 29714
rect 18616 29668 18696 29696
rect 18696 29650 18748 29656
rect 18694 29608 18750 29617
rect 18694 29543 18696 29552
rect 18748 29543 18750 29552
rect 18696 29514 18748 29520
rect 18604 29504 18656 29510
rect 18602 29472 18604 29481
rect 18656 29472 18658 29481
rect 18602 29407 18658 29416
rect 18800 28694 18828 29990
rect 18972 29640 19024 29646
rect 18972 29582 19024 29588
rect 18984 29102 19012 29582
rect 18972 29096 19024 29102
rect 18972 29038 19024 29044
rect 18972 28960 19024 28966
rect 18970 28928 18972 28937
rect 19024 28928 19026 28937
rect 18970 28863 19026 28872
rect 18788 28688 18840 28694
rect 18788 28630 18840 28636
rect 18970 28656 19026 28665
rect 18970 28591 19026 28600
rect 18984 28558 19012 28591
rect 18972 28552 19024 28558
rect 18524 28478 18828 28506
rect 18972 28494 19024 28500
rect 18604 28416 18656 28422
rect 18604 28358 18656 28364
rect 18420 28144 18472 28150
rect 18420 28086 18472 28092
rect 18236 27940 18288 27946
rect 18236 27882 18288 27888
rect 18420 27872 18472 27878
rect 18420 27814 18472 27820
rect 18512 27872 18564 27878
rect 18512 27814 18564 27820
rect 17868 27532 17920 27538
rect 17868 27474 17920 27480
rect 17408 27464 17460 27470
rect 17408 27406 17460 27412
rect 18328 27464 18380 27470
rect 18328 27406 18380 27412
rect 17408 27328 17460 27334
rect 17408 27270 17460 27276
rect 18236 27328 18288 27334
rect 18236 27270 18288 27276
rect 17040 26988 17092 26994
rect 17040 26930 17092 26936
rect 16948 26920 17000 26926
rect 16948 26862 17000 26868
rect 16960 26586 16988 26862
rect 17040 26784 17092 26790
rect 17040 26726 17092 26732
rect 16948 26580 17000 26586
rect 16948 26522 17000 26528
rect 17052 26382 17080 26726
rect 16764 26376 16816 26382
rect 16764 26318 16816 26324
rect 17040 26376 17092 26382
rect 17040 26318 17092 26324
rect 17316 26376 17368 26382
rect 17316 26318 17368 26324
rect 17328 25378 17356 26318
rect 17420 26314 17448 27270
rect 17831 27228 18139 27237
rect 17831 27226 17837 27228
rect 17893 27226 17917 27228
rect 17973 27226 17997 27228
rect 18053 27226 18077 27228
rect 18133 27226 18139 27228
rect 17893 27174 17895 27226
rect 18075 27174 18077 27226
rect 17831 27172 17837 27174
rect 17893 27172 17917 27174
rect 17973 27172 17997 27174
rect 18053 27172 18077 27174
rect 18133 27172 18139 27174
rect 17831 27163 18139 27172
rect 18248 27062 18276 27270
rect 18340 27130 18368 27406
rect 18328 27124 18380 27130
rect 18328 27066 18380 27072
rect 18236 27056 18288 27062
rect 17512 26994 18092 27010
rect 18236 26998 18288 27004
rect 17512 26988 18104 26994
rect 17512 26982 18052 26988
rect 17512 26382 17540 26982
rect 18052 26930 18104 26936
rect 18432 26926 18460 27814
rect 18524 27606 18552 27814
rect 18512 27600 18564 27606
rect 18512 27542 18564 27548
rect 18524 26994 18552 27542
rect 18616 27470 18644 28358
rect 18694 27568 18750 27577
rect 18694 27503 18750 27512
rect 18604 27464 18656 27470
rect 18604 27406 18656 27412
rect 18512 26988 18564 26994
rect 18512 26930 18564 26936
rect 18144 26920 18196 26926
rect 18144 26862 18196 26868
rect 18420 26920 18472 26926
rect 18420 26862 18472 26868
rect 17868 26784 17920 26790
rect 17868 26726 17920 26732
rect 17880 26466 17908 26726
rect 17604 26450 17908 26466
rect 17604 26444 17920 26450
rect 17604 26438 17868 26444
rect 17500 26376 17552 26382
rect 17500 26318 17552 26324
rect 17408 26308 17460 26314
rect 17408 26250 17460 26256
rect 17420 25838 17448 26250
rect 17604 25906 17632 26438
rect 17868 26386 17920 26392
rect 18156 26382 18184 26862
rect 18236 26852 18288 26858
rect 18236 26794 18288 26800
rect 17684 26376 17736 26382
rect 17684 26318 17736 26324
rect 18144 26376 18196 26382
rect 18144 26318 18196 26324
rect 17696 25906 17724 26318
rect 17831 26140 18139 26149
rect 17831 26138 17837 26140
rect 17893 26138 17917 26140
rect 17973 26138 17997 26140
rect 18053 26138 18077 26140
rect 18133 26138 18139 26140
rect 17893 26086 17895 26138
rect 18075 26086 18077 26138
rect 17831 26084 17837 26086
rect 17893 26084 17917 26086
rect 17973 26084 17997 26086
rect 18053 26084 18077 26086
rect 18133 26084 18139 26086
rect 17831 26075 18139 26084
rect 18248 25974 18276 26794
rect 18604 26376 18656 26382
rect 18604 26318 18656 26324
rect 18328 26308 18380 26314
rect 18328 26250 18380 26256
rect 18144 25968 18196 25974
rect 18144 25910 18196 25916
rect 18236 25968 18288 25974
rect 18236 25910 18288 25916
rect 17592 25900 17644 25906
rect 17592 25842 17644 25848
rect 17684 25900 17736 25906
rect 17684 25842 17736 25848
rect 17408 25832 17460 25838
rect 17408 25774 17460 25780
rect 17408 25696 17460 25702
rect 17408 25638 17460 25644
rect 17052 25350 17356 25378
rect 17052 25294 17080 25350
rect 16580 25288 16632 25294
rect 16580 25230 16632 25236
rect 17040 25288 17092 25294
rect 17040 25230 17092 25236
rect 17132 25288 17184 25294
rect 17132 25230 17184 25236
rect 16592 24954 16620 25230
rect 16856 25220 16908 25226
rect 16856 25162 16908 25168
rect 16580 24948 16632 24954
rect 16580 24890 16632 24896
rect 16592 23118 16620 24890
rect 16868 24410 16896 25162
rect 16856 24404 16908 24410
rect 16856 24346 16908 24352
rect 16764 24268 16816 24274
rect 16764 24210 16816 24216
rect 16672 24064 16724 24070
rect 16672 24006 16724 24012
rect 16684 23322 16712 24006
rect 16672 23316 16724 23322
rect 16672 23258 16724 23264
rect 16776 23118 16804 24210
rect 16868 23662 16896 24346
rect 17144 24177 17172 25230
rect 17328 24954 17356 25350
rect 17420 25294 17448 25638
rect 17408 25288 17460 25294
rect 17408 25230 17460 25236
rect 18050 25256 18106 25265
rect 18156 25242 18184 25910
rect 18340 25906 18368 26250
rect 18420 26240 18472 26246
rect 18420 26182 18472 26188
rect 18328 25900 18380 25906
rect 18328 25842 18380 25848
rect 18432 25362 18460 26182
rect 18616 25906 18644 26318
rect 18604 25900 18656 25906
rect 18604 25842 18656 25848
rect 18420 25356 18472 25362
rect 18420 25298 18472 25304
rect 18156 25214 18368 25242
rect 18050 25191 18052 25200
rect 18104 25191 18106 25200
rect 18052 25162 18104 25168
rect 17592 25152 17644 25158
rect 17592 25094 17644 25100
rect 17316 24948 17368 24954
rect 17316 24890 17368 24896
rect 17408 24880 17460 24886
rect 17408 24822 17460 24828
rect 17500 24880 17552 24886
rect 17500 24822 17552 24828
rect 17224 24812 17276 24818
rect 17224 24754 17276 24760
rect 17236 24410 17264 24754
rect 17316 24608 17368 24614
rect 17316 24550 17368 24556
rect 17224 24404 17276 24410
rect 17224 24346 17276 24352
rect 17130 24168 17186 24177
rect 17328 24138 17356 24550
rect 17130 24103 17186 24112
rect 17316 24132 17368 24138
rect 17144 23712 17172 24103
rect 17316 24074 17368 24080
rect 17328 23746 17356 24074
rect 17420 24070 17448 24822
rect 17512 24206 17540 24822
rect 17500 24200 17552 24206
rect 17500 24142 17552 24148
rect 17408 24064 17460 24070
rect 17408 24006 17460 24012
rect 17512 23798 17540 24142
rect 17500 23792 17552 23798
rect 17224 23724 17276 23730
rect 17144 23684 17224 23712
rect 17328 23718 17448 23746
rect 17500 23734 17552 23740
rect 17224 23666 17276 23672
rect 16856 23656 16908 23662
rect 16856 23598 16908 23604
rect 17316 23656 17368 23662
rect 17316 23598 17368 23604
rect 16580 23112 16632 23118
rect 16580 23054 16632 23060
rect 16764 23112 16816 23118
rect 16764 23054 16816 23060
rect 16592 22642 16620 23054
rect 16580 22636 16632 22642
rect 16580 22578 16632 22584
rect 16396 22432 16448 22438
rect 16396 22374 16448 22380
rect 16592 22166 16620 22578
rect 16776 22506 16804 23054
rect 17328 22778 17356 23598
rect 17420 23118 17448 23718
rect 17500 23588 17552 23594
rect 17500 23530 17552 23536
rect 17408 23112 17460 23118
rect 17408 23054 17460 23060
rect 17316 22772 17368 22778
rect 17316 22714 17368 22720
rect 17512 22574 17540 23530
rect 17604 23186 17632 25094
rect 17831 25052 18139 25061
rect 17831 25050 17837 25052
rect 17893 25050 17917 25052
rect 17973 25050 17997 25052
rect 18053 25050 18077 25052
rect 18133 25050 18139 25052
rect 17893 24998 17895 25050
rect 18075 24998 18077 25050
rect 17831 24996 17837 24998
rect 17893 24996 17917 24998
rect 17973 24996 17997 24998
rect 18053 24996 18077 24998
rect 18133 24996 18139 24998
rect 17831 24987 18139 24996
rect 18340 24818 18368 25214
rect 18604 25220 18656 25226
rect 18708 25208 18736 27503
rect 18800 27062 18828 28478
rect 19076 28422 19104 30670
rect 19248 30184 19300 30190
rect 19248 30126 19300 30132
rect 19156 30116 19208 30122
rect 19156 30058 19208 30064
rect 19168 29170 19196 30058
rect 19260 30054 19288 30126
rect 19248 30048 19300 30054
rect 19444 30036 19472 30670
rect 19616 30320 19668 30326
rect 19614 30288 19616 30297
rect 19668 30288 19670 30297
rect 19614 30223 19670 30232
rect 19614 30152 19670 30161
rect 19614 30087 19670 30096
rect 19524 30048 19576 30054
rect 19444 30008 19524 30036
rect 19248 29990 19300 29996
rect 19524 29990 19576 29996
rect 19536 29714 19564 29990
rect 19628 29782 19656 30087
rect 19616 29776 19668 29782
rect 19616 29718 19668 29724
rect 19524 29708 19576 29714
rect 19524 29650 19576 29656
rect 19246 29608 19302 29617
rect 19246 29543 19248 29552
rect 19300 29543 19302 29552
rect 19248 29514 19300 29520
rect 19340 29504 19392 29510
rect 19340 29446 19392 29452
rect 19156 29164 19208 29170
rect 19156 29106 19208 29112
rect 19248 29164 19300 29170
rect 19248 29106 19300 29112
rect 19064 28416 19116 28422
rect 19064 28358 19116 28364
rect 19168 28150 19196 29106
rect 19260 28626 19288 29106
rect 19248 28620 19300 28626
rect 19248 28562 19300 28568
rect 19352 28506 19380 29446
rect 19536 28558 19564 29650
rect 19260 28478 19380 28506
rect 19524 28552 19576 28558
rect 19524 28494 19576 28500
rect 19156 28144 19208 28150
rect 19156 28086 19208 28092
rect 19064 28076 19116 28082
rect 19064 28018 19116 28024
rect 19076 27538 19104 28018
rect 19064 27532 19116 27538
rect 19064 27474 19116 27480
rect 19156 27464 19208 27470
rect 19156 27406 19208 27412
rect 18788 27056 18840 27062
rect 18788 26998 18840 27004
rect 19062 26888 19118 26897
rect 19062 26823 19118 26832
rect 19076 26586 19104 26823
rect 19064 26580 19116 26586
rect 19064 26522 19116 26528
rect 18972 26512 19024 26518
rect 18970 26480 18972 26489
rect 19024 26480 19026 26489
rect 18788 26444 18840 26450
rect 18970 26415 19026 26424
rect 18788 26386 18840 26392
rect 18800 25906 18828 26386
rect 18880 26376 18932 26382
rect 18880 26318 18932 26324
rect 18788 25900 18840 25906
rect 18788 25842 18840 25848
rect 18800 25294 18828 25842
rect 18892 25498 18920 26318
rect 18880 25492 18932 25498
rect 18880 25434 18932 25440
rect 18788 25288 18840 25294
rect 18788 25230 18840 25236
rect 18656 25180 18736 25208
rect 18604 25162 18656 25168
rect 18328 24812 18380 24818
rect 18328 24754 18380 24760
rect 18340 24698 18368 24754
rect 18248 24670 18368 24698
rect 18604 24744 18656 24750
rect 18604 24686 18656 24692
rect 17684 24608 17736 24614
rect 17684 24550 17736 24556
rect 17696 23798 17724 24550
rect 17831 23964 18139 23973
rect 17831 23962 17837 23964
rect 17893 23962 17917 23964
rect 17973 23962 17997 23964
rect 18053 23962 18077 23964
rect 18133 23962 18139 23964
rect 17893 23910 17895 23962
rect 18075 23910 18077 23962
rect 17831 23908 17837 23910
rect 17893 23908 17917 23910
rect 17973 23908 17997 23910
rect 18053 23908 18077 23910
rect 18133 23908 18139 23910
rect 17831 23899 18139 23908
rect 17684 23792 17736 23798
rect 17684 23734 17736 23740
rect 17958 23760 18014 23769
rect 17958 23695 17960 23704
rect 18012 23695 18014 23704
rect 17960 23666 18012 23672
rect 17592 23180 17644 23186
rect 17592 23122 17644 23128
rect 18248 23050 18276 24670
rect 18328 24608 18380 24614
rect 18328 24550 18380 24556
rect 18340 23730 18368 24550
rect 18420 24404 18472 24410
rect 18420 24346 18472 24352
rect 18328 23724 18380 23730
rect 18328 23666 18380 23672
rect 18432 23322 18460 24346
rect 18616 24206 18644 24686
rect 18604 24200 18656 24206
rect 18604 24142 18656 24148
rect 18616 23662 18644 24142
rect 18604 23656 18656 23662
rect 18604 23598 18656 23604
rect 18420 23316 18472 23322
rect 18420 23258 18472 23264
rect 18616 23304 18644 23598
rect 18696 23316 18748 23322
rect 18616 23276 18696 23304
rect 18236 23044 18288 23050
rect 18236 22986 18288 22992
rect 17831 22876 18139 22885
rect 17831 22874 17837 22876
rect 17893 22874 17917 22876
rect 17973 22874 17997 22876
rect 18053 22874 18077 22876
rect 18133 22874 18139 22876
rect 17893 22822 17895 22874
rect 18075 22822 18077 22874
rect 17831 22820 17837 22822
rect 17893 22820 17917 22822
rect 17973 22820 17997 22822
rect 18053 22820 18077 22822
rect 18133 22820 18139 22822
rect 17831 22811 18139 22820
rect 17592 22636 17644 22642
rect 17592 22578 17644 22584
rect 17500 22568 17552 22574
rect 17500 22510 17552 22516
rect 16764 22500 16816 22506
rect 16764 22442 16816 22448
rect 16580 22160 16632 22166
rect 16580 22102 16632 22108
rect 16488 22092 16540 22098
rect 16488 22034 16540 22040
rect 16120 21616 16172 21622
rect 16120 21558 16172 21564
rect 16028 21548 16080 21554
rect 16028 21490 16080 21496
rect 15936 21480 15988 21486
rect 15936 21422 15988 21428
rect 15948 21146 15976 21422
rect 16040 21418 16068 21490
rect 16132 21486 16160 21558
rect 16120 21480 16172 21486
rect 16120 21422 16172 21428
rect 16028 21412 16080 21418
rect 16028 21354 16080 21360
rect 15936 21140 15988 21146
rect 15936 21082 15988 21088
rect 16132 20534 16160 21422
rect 16500 21418 16528 22034
rect 16488 21412 16540 21418
rect 16488 21354 16540 21360
rect 16592 21010 16620 22102
rect 17316 22092 17368 22098
rect 17316 22034 17368 22040
rect 16672 22024 16724 22030
rect 16672 21966 16724 21972
rect 16684 21146 16712 21966
rect 17328 21690 17356 22034
rect 17500 21956 17552 21962
rect 17500 21898 17552 21904
rect 17132 21684 17184 21690
rect 17132 21626 17184 21632
rect 17316 21684 17368 21690
rect 17316 21626 17368 21632
rect 16856 21480 16908 21486
rect 16856 21422 16908 21428
rect 16672 21140 16724 21146
rect 16672 21082 16724 21088
rect 16580 21004 16632 21010
rect 16580 20946 16632 20952
rect 16120 20528 16172 20534
rect 16120 20470 16172 20476
rect 16592 20466 16620 20946
rect 16672 20936 16724 20942
rect 16672 20878 16724 20884
rect 16028 20460 16080 20466
rect 16028 20402 16080 20408
rect 16212 20460 16264 20466
rect 16212 20402 16264 20408
rect 16580 20460 16632 20466
rect 16580 20402 16632 20408
rect 16040 19990 16068 20402
rect 16028 19984 16080 19990
rect 16028 19926 16080 19932
rect 16040 19514 16068 19926
rect 15568 19508 15620 19514
rect 15568 19450 15620 19456
rect 16028 19508 16080 19514
rect 16028 19450 16080 19456
rect 15580 19378 15608 19450
rect 16224 19446 16252 20402
rect 16212 19440 16264 19446
rect 16212 19382 16264 19388
rect 16592 19378 16620 20402
rect 16684 20398 16712 20878
rect 16868 20602 16896 21422
rect 16948 21344 17000 21350
rect 16948 21286 17000 21292
rect 16856 20596 16908 20602
rect 16856 20538 16908 20544
rect 16672 20392 16724 20398
rect 16672 20334 16724 20340
rect 16764 20324 16816 20330
rect 16764 20266 16816 20272
rect 16776 19854 16804 20266
rect 16960 19922 16988 21286
rect 17144 20942 17172 21626
rect 17512 21486 17540 21898
rect 17604 21554 17632 22578
rect 17831 21788 18139 21797
rect 17831 21786 17837 21788
rect 17893 21786 17917 21788
rect 17973 21786 17997 21788
rect 18053 21786 18077 21788
rect 18133 21786 18139 21788
rect 17893 21734 17895 21786
rect 18075 21734 18077 21786
rect 17831 21732 17837 21734
rect 17893 21732 17917 21734
rect 17973 21732 17997 21734
rect 18053 21732 18077 21734
rect 18133 21732 18139 21734
rect 17831 21723 18139 21732
rect 17592 21548 17644 21554
rect 18248 21536 18276 22986
rect 18616 22030 18644 23276
rect 18696 23258 18748 23264
rect 18800 23254 18828 25230
rect 19064 25220 19116 25226
rect 19064 25162 19116 25168
rect 18880 25152 18932 25158
rect 18880 25094 18932 25100
rect 18892 24818 18920 25094
rect 19076 24818 19104 25162
rect 18880 24812 18932 24818
rect 18880 24754 18932 24760
rect 19064 24812 19116 24818
rect 19064 24754 19116 24760
rect 18880 24200 18932 24206
rect 18880 24142 18932 24148
rect 19064 24200 19116 24206
rect 19064 24142 19116 24148
rect 18788 23248 18840 23254
rect 18788 23190 18840 23196
rect 18800 22982 18828 23190
rect 18788 22976 18840 22982
rect 18788 22918 18840 22924
rect 18696 22160 18748 22166
rect 18696 22102 18748 22108
rect 18604 22024 18656 22030
rect 18604 21966 18656 21972
rect 17592 21490 17644 21496
rect 18156 21508 18368 21536
rect 17500 21480 17552 21486
rect 17500 21422 17552 21428
rect 17132 20936 17184 20942
rect 17132 20878 17184 20884
rect 17512 20330 17540 21422
rect 17592 21412 17644 21418
rect 17592 21354 17644 21360
rect 17604 20534 17632 21354
rect 18156 20806 18184 21508
rect 18236 21004 18288 21010
rect 18236 20946 18288 20952
rect 18144 20800 18196 20806
rect 18144 20742 18196 20748
rect 17831 20700 18139 20709
rect 17831 20698 17837 20700
rect 17893 20698 17917 20700
rect 17973 20698 17997 20700
rect 18053 20698 18077 20700
rect 18133 20698 18139 20700
rect 17893 20646 17895 20698
rect 18075 20646 18077 20698
rect 17831 20644 17837 20646
rect 17893 20644 17917 20646
rect 17973 20644 17997 20646
rect 18053 20644 18077 20646
rect 18133 20644 18139 20646
rect 17831 20635 18139 20644
rect 18248 20602 18276 20946
rect 18236 20596 18288 20602
rect 18236 20538 18288 20544
rect 17592 20528 17644 20534
rect 17592 20470 17644 20476
rect 18340 20346 18368 21508
rect 18420 20936 18472 20942
rect 18472 20896 18552 20924
rect 18616 20920 18644 21966
rect 18420 20878 18472 20884
rect 17500 20324 17552 20330
rect 18340 20318 18460 20346
rect 18524 20330 18552 20896
rect 18604 20914 18656 20920
rect 18604 20856 18656 20862
rect 17500 20266 17552 20272
rect 17040 20256 17092 20262
rect 17040 20198 17092 20204
rect 16948 19916 17000 19922
rect 16948 19858 17000 19864
rect 17052 19854 17080 20198
rect 18432 20058 18460 20318
rect 18512 20324 18564 20330
rect 18512 20266 18564 20272
rect 18420 20052 18472 20058
rect 18420 19994 18472 20000
rect 16764 19848 16816 19854
rect 16764 19790 16816 19796
rect 17040 19848 17092 19854
rect 17040 19790 17092 19796
rect 17132 19848 17184 19854
rect 17132 19790 17184 19796
rect 16672 19712 16724 19718
rect 16672 19654 16724 19660
rect 16684 19378 16712 19654
rect 15568 19372 15620 19378
rect 15568 19314 15620 19320
rect 16580 19372 16632 19378
rect 16580 19314 16632 19320
rect 16672 19372 16724 19378
rect 16672 19314 16724 19320
rect 16592 18902 16620 19314
rect 16580 18896 16632 18902
rect 16580 18838 16632 18844
rect 16776 18766 16804 19790
rect 16948 19304 17000 19310
rect 16948 19246 17000 19252
rect 16960 18970 16988 19246
rect 16948 18964 17000 18970
rect 16948 18906 17000 18912
rect 16764 18760 16816 18766
rect 16764 18702 16816 18708
rect 17052 18290 17080 19790
rect 17040 18284 17092 18290
rect 17040 18226 17092 18232
rect 17144 18222 17172 19790
rect 18328 19780 18380 19786
rect 18328 19722 18380 19728
rect 17831 19612 18139 19621
rect 17831 19610 17837 19612
rect 17893 19610 17917 19612
rect 17973 19610 17997 19612
rect 18053 19610 18077 19612
rect 18133 19610 18139 19612
rect 17893 19558 17895 19610
rect 18075 19558 18077 19610
rect 17831 19556 17837 19558
rect 17893 19556 17917 19558
rect 17973 19556 17997 19558
rect 18053 19556 18077 19558
rect 18133 19556 18139 19558
rect 17831 19547 18139 19556
rect 18340 19242 18368 19722
rect 18432 19378 18460 19994
rect 18616 19718 18644 20856
rect 18604 19712 18656 19718
rect 18604 19654 18656 19660
rect 18616 19514 18644 19654
rect 18604 19508 18656 19514
rect 18604 19450 18656 19456
rect 18420 19372 18472 19378
rect 18420 19314 18472 19320
rect 18328 19236 18380 19242
rect 18328 19178 18380 19184
rect 18420 19168 18472 19174
rect 18420 19110 18472 19116
rect 18432 18766 18460 19110
rect 18616 18766 18644 19450
rect 18708 19242 18736 22102
rect 18892 20942 18920 24142
rect 19076 23730 19104 24142
rect 19064 23724 19116 23730
rect 19064 23666 19116 23672
rect 19076 22710 19104 23666
rect 19064 22704 19116 22710
rect 19064 22646 19116 22652
rect 19064 22024 19116 22030
rect 19064 21966 19116 21972
rect 18972 21956 19024 21962
rect 18972 21898 19024 21904
rect 18984 21554 19012 21898
rect 18972 21548 19024 21554
rect 18972 21490 19024 21496
rect 18880 20936 18932 20942
rect 18880 20878 18932 20884
rect 18696 19236 18748 19242
rect 18696 19178 18748 19184
rect 18892 18766 18920 20878
rect 19076 19854 19104 21966
rect 19064 19848 19116 19854
rect 19064 19790 19116 19796
rect 17408 18760 17460 18766
rect 17408 18702 17460 18708
rect 18420 18760 18472 18766
rect 18420 18702 18472 18708
rect 18604 18760 18656 18766
rect 18604 18702 18656 18708
rect 18880 18760 18932 18766
rect 18880 18702 18932 18708
rect 17420 18426 17448 18702
rect 17831 18524 18139 18533
rect 17831 18522 17837 18524
rect 17893 18522 17917 18524
rect 17973 18522 17997 18524
rect 18053 18522 18077 18524
rect 18133 18522 18139 18524
rect 17893 18470 17895 18522
rect 18075 18470 18077 18522
rect 17831 18468 17837 18470
rect 17893 18468 17917 18470
rect 17973 18468 17997 18470
rect 18053 18468 18077 18470
rect 18133 18468 18139 18470
rect 17831 18459 18139 18468
rect 18432 18426 18460 18702
rect 18512 18624 18564 18630
rect 18512 18566 18564 18572
rect 17408 18420 17460 18426
rect 17408 18362 17460 18368
rect 18420 18420 18472 18426
rect 18420 18362 18472 18368
rect 18524 18290 18552 18566
rect 18512 18284 18564 18290
rect 18512 18226 18564 18232
rect 17132 18216 17184 18222
rect 17132 18158 17184 18164
rect 17831 17436 18139 17445
rect 17831 17434 17837 17436
rect 17893 17434 17917 17436
rect 17973 17434 17997 17436
rect 18053 17434 18077 17436
rect 18133 17434 18139 17436
rect 17893 17382 17895 17434
rect 18075 17382 18077 17434
rect 17831 17380 17837 17382
rect 17893 17380 17917 17382
rect 17973 17380 17997 17382
rect 18053 17380 18077 17382
rect 18133 17380 18139 17382
rect 17831 17371 18139 17380
rect 19076 17270 19104 19790
rect 19064 17264 19116 17270
rect 19064 17206 19116 17212
rect 17831 16348 18139 16357
rect 17831 16346 17837 16348
rect 17893 16346 17917 16348
rect 17973 16346 17997 16348
rect 18053 16346 18077 16348
rect 18133 16346 18139 16348
rect 17893 16294 17895 16346
rect 18075 16294 18077 16346
rect 17831 16292 17837 16294
rect 17893 16292 17917 16294
rect 17973 16292 17997 16294
rect 18053 16292 18077 16294
rect 18133 16292 18139 16294
rect 17831 16283 18139 16292
rect 17831 15260 18139 15269
rect 17831 15258 17837 15260
rect 17893 15258 17917 15260
rect 17973 15258 17997 15260
rect 18053 15258 18077 15260
rect 18133 15258 18139 15260
rect 17893 15206 17895 15258
rect 18075 15206 18077 15258
rect 17831 15204 17837 15206
rect 17893 15204 17917 15206
rect 17973 15204 17997 15206
rect 18053 15204 18077 15206
rect 18133 15204 18139 15206
rect 17831 15195 18139 15204
rect 15292 14952 15344 14958
rect 15292 14894 15344 14900
rect 13611 14716 13919 14725
rect 13611 14714 13617 14716
rect 13673 14714 13697 14716
rect 13753 14714 13777 14716
rect 13833 14714 13857 14716
rect 13913 14714 13919 14716
rect 13673 14662 13675 14714
rect 13855 14662 13857 14714
rect 13611 14660 13617 14662
rect 13673 14660 13697 14662
rect 13753 14660 13777 14662
rect 13833 14660 13857 14662
rect 13913 14660 13919 14662
rect 13611 14651 13919 14660
rect 9390 14172 9698 14181
rect 9390 14170 9396 14172
rect 9452 14170 9476 14172
rect 9532 14170 9556 14172
rect 9612 14170 9636 14172
rect 9692 14170 9698 14172
rect 9452 14118 9454 14170
rect 9634 14118 9636 14170
rect 9390 14116 9396 14118
rect 9452 14116 9476 14118
rect 9532 14116 9556 14118
rect 9612 14116 9636 14118
rect 9692 14116 9698 14118
rect 9390 14107 9698 14116
rect 17831 14172 18139 14181
rect 17831 14170 17837 14172
rect 17893 14170 17917 14172
rect 17973 14170 17997 14172
rect 18053 14170 18077 14172
rect 18133 14170 18139 14172
rect 17893 14118 17895 14170
rect 18075 14118 18077 14170
rect 17831 14116 17837 14118
rect 17893 14116 17917 14118
rect 17973 14116 17997 14118
rect 18053 14116 18077 14118
rect 18133 14116 18139 14118
rect 17831 14107 18139 14116
rect 13611 13628 13919 13637
rect 13611 13626 13617 13628
rect 13673 13626 13697 13628
rect 13753 13626 13777 13628
rect 13833 13626 13857 13628
rect 13913 13626 13919 13628
rect 13673 13574 13675 13626
rect 13855 13574 13857 13626
rect 13611 13572 13617 13574
rect 13673 13572 13697 13574
rect 13753 13572 13777 13574
rect 13833 13572 13857 13574
rect 13913 13572 13919 13574
rect 13611 13563 13919 13572
rect 9390 13084 9698 13093
rect 9390 13082 9396 13084
rect 9452 13082 9476 13084
rect 9532 13082 9556 13084
rect 9612 13082 9636 13084
rect 9692 13082 9698 13084
rect 9452 13030 9454 13082
rect 9634 13030 9636 13082
rect 9390 13028 9396 13030
rect 9452 13028 9476 13030
rect 9532 13028 9556 13030
rect 9612 13028 9636 13030
rect 9692 13028 9698 13030
rect 9390 13019 9698 13028
rect 17831 13084 18139 13093
rect 17831 13082 17837 13084
rect 17893 13082 17917 13084
rect 17973 13082 17997 13084
rect 18053 13082 18077 13084
rect 18133 13082 18139 13084
rect 17893 13030 17895 13082
rect 18075 13030 18077 13082
rect 17831 13028 17837 13030
rect 17893 13028 17917 13030
rect 17973 13028 17997 13030
rect 18053 13028 18077 13030
rect 18133 13028 18139 13030
rect 17831 13019 18139 13028
rect 13611 12540 13919 12549
rect 13611 12538 13617 12540
rect 13673 12538 13697 12540
rect 13753 12538 13777 12540
rect 13833 12538 13857 12540
rect 13913 12538 13919 12540
rect 13673 12486 13675 12538
rect 13855 12486 13857 12538
rect 13611 12484 13617 12486
rect 13673 12484 13697 12486
rect 13753 12484 13777 12486
rect 13833 12484 13857 12486
rect 13913 12484 13919 12486
rect 13611 12475 13919 12484
rect 14372 12232 14424 12238
rect 14372 12174 14424 12180
rect 9390 11996 9698 12005
rect 9390 11994 9396 11996
rect 9452 11994 9476 11996
rect 9532 11994 9556 11996
rect 9612 11994 9636 11996
rect 9692 11994 9698 11996
rect 9452 11942 9454 11994
rect 9634 11942 9636 11994
rect 9390 11940 9396 11942
rect 9452 11940 9476 11942
rect 9532 11940 9556 11942
rect 9612 11940 9636 11942
rect 9692 11940 9698 11942
rect 9390 11931 9698 11940
rect 13611 11452 13919 11461
rect 13611 11450 13617 11452
rect 13673 11450 13697 11452
rect 13753 11450 13777 11452
rect 13833 11450 13857 11452
rect 13913 11450 13919 11452
rect 13673 11398 13675 11450
rect 13855 11398 13857 11450
rect 13611 11396 13617 11398
rect 13673 11396 13697 11398
rect 13753 11396 13777 11398
rect 13833 11396 13857 11398
rect 13913 11396 13919 11398
rect 13611 11387 13919 11396
rect 9390 10908 9698 10917
rect 9390 10906 9396 10908
rect 9452 10906 9476 10908
rect 9532 10906 9556 10908
rect 9612 10906 9636 10908
rect 9692 10906 9698 10908
rect 9452 10854 9454 10906
rect 9634 10854 9636 10906
rect 9390 10852 9396 10854
rect 9452 10852 9476 10854
rect 9532 10852 9556 10854
rect 9612 10852 9636 10854
rect 9692 10852 9698 10854
rect 9390 10843 9698 10852
rect 13611 10364 13919 10373
rect 13611 10362 13617 10364
rect 13673 10362 13697 10364
rect 13753 10362 13777 10364
rect 13833 10362 13857 10364
rect 13913 10362 13919 10364
rect 13673 10310 13675 10362
rect 13855 10310 13857 10362
rect 13611 10308 13617 10310
rect 13673 10308 13697 10310
rect 13753 10308 13777 10310
rect 13833 10308 13857 10310
rect 13913 10308 13919 10310
rect 13611 10299 13919 10308
rect 9390 9820 9698 9829
rect 9390 9818 9396 9820
rect 9452 9818 9476 9820
rect 9532 9818 9556 9820
rect 9612 9818 9636 9820
rect 9692 9818 9698 9820
rect 9452 9766 9454 9818
rect 9634 9766 9636 9818
rect 9390 9764 9396 9766
rect 9452 9764 9476 9766
rect 9532 9764 9556 9766
rect 9612 9764 9636 9766
rect 9692 9764 9698 9766
rect 9390 9755 9698 9764
rect 9128 9580 9180 9586
rect 9128 9522 9180 9528
rect 7196 7948 7248 7954
rect 7196 7890 7248 7896
rect 7380 7948 7432 7954
rect 7380 7890 7432 7896
rect 5170 7100 5478 7109
rect 5170 7098 5176 7100
rect 5232 7098 5256 7100
rect 5312 7098 5336 7100
rect 5392 7098 5416 7100
rect 5472 7098 5478 7100
rect 5232 7046 5234 7098
rect 5414 7046 5416 7098
rect 5170 7044 5176 7046
rect 5232 7044 5256 7046
rect 5312 7044 5336 7046
rect 5392 7044 5416 7046
rect 5472 7044 5478 7046
rect 5170 7035 5478 7044
rect 7208 6730 7236 7890
rect 9140 6798 9168 9522
rect 13611 9276 13919 9285
rect 13611 9274 13617 9276
rect 13673 9274 13697 9276
rect 13753 9274 13777 9276
rect 13833 9274 13857 9276
rect 13913 9274 13919 9276
rect 13673 9222 13675 9274
rect 13855 9222 13857 9274
rect 13611 9220 13617 9222
rect 13673 9220 13697 9222
rect 13753 9220 13777 9222
rect 13833 9220 13857 9222
rect 13913 9220 13919 9222
rect 13611 9211 13919 9220
rect 9390 8732 9698 8741
rect 9390 8730 9396 8732
rect 9452 8730 9476 8732
rect 9532 8730 9556 8732
rect 9612 8730 9636 8732
rect 9692 8730 9698 8732
rect 9452 8678 9454 8730
rect 9634 8678 9636 8730
rect 9390 8676 9396 8678
rect 9452 8676 9476 8678
rect 9532 8676 9556 8678
rect 9612 8676 9636 8678
rect 9692 8676 9698 8678
rect 9390 8667 9698 8676
rect 13611 8188 13919 8197
rect 13611 8186 13617 8188
rect 13673 8186 13697 8188
rect 13753 8186 13777 8188
rect 13833 8186 13857 8188
rect 13913 8186 13919 8188
rect 13673 8134 13675 8186
rect 13855 8134 13857 8186
rect 13611 8132 13617 8134
rect 13673 8132 13697 8134
rect 13753 8132 13777 8134
rect 13833 8132 13857 8134
rect 13913 8132 13919 8134
rect 13611 8123 13919 8132
rect 9390 7644 9698 7653
rect 9390 7642 9396 7644
rect 9452 7642 9476 7644
rect 9532 7642 9556 7644
rect 9612 7642 9636 7644
rect 9692 7642 9698 7644
rect 9452 7590 9454 7642
rect 9634 7590 9636 7642
rect 9390 7588 9396 7590
rect 9452 7588 9476 7590
rect 9532 7588 9556 7590
rect 9612 7588 9636 7590
rect 9692 7588 9698 7590
rect 9390 7579 9698 7588
rect 13611 7100 13919 7109
rect 13611 7098 13617 7100
rect 13673 7098 13697 7100
rect 13753 7098 13777 7100
rect 13833 7098 13857 7100
rect 13913 7098 13919 7100
rect 13673 7046 13675 7098
rect 13855 7046 13857 7098
rect 13611 7044 13617 7046
rect 13673 7044 13697 7046
rect 13753 7044 13777 7046
rect 13833 7044 13857 7046
rect 13913 7044 13919 7046
rect 13611 7035 13919 7044
rect 9128 6792 9180 6798
rect 9128 6734 9180 6740
rect 7196 6724 7248 6730
rect 7196 6666 7248 6672
rect 5170 6012 5478 6021
rect 5170 6010 5176 6012
rect 5232 6010 5256 6012
rect 5312 6010 5336 6012
rect 5392 6010 5416 6012
rect 5472 6010 5478 6012
rect 5232 5958 5234 6010
rect 5414 5958 5416 6010
rect 5170 5956 5176 5958
rect 5232 5956 5256 5958
rect 5312 5956 5336 5958
rect 5392 5956 5416 5958
rect 5472 5956 5478 5958
rect 5170 5947 5478 5956
rect 6460 5772 6512 5778
rect 6460 5714 6512 5720
rect 5080 5704 5132 5710
rect 5080 5646 5132 5652
rect 5632 5704 5684 5710
rect 5632 5646 5684 5652
rect 6092 5704 6144 5710
rect 6092 5646 6144 5652
rect 5000 5494 5120 5522
rect 4896 5160 4948 5166
rect 4896 5102 4948 5108
rect 5092 4690 5120 5494
rect 5170 4924 5478 4933
rect 5170 4922 5176 4924
rect 5232 4922 5256 4924
rect 5312 4922 5336 4924
rect 5392 4922 5416 4924
rect 5472 4922 5478 4924
rect 5232 4870 5234 4922
rect 5414 4870 5416 4922
rect 5170 4868 5176 4870
rect 5232 4868 5256 4870
rect 5312 4868 5336 4870
rect 5392 4868 5416 4870
rect 5472 4868 5478 4870
rect 5170 4859 5478 4868
rect 4804 4684 4856 4690
rect 4804 4626 4856 4632
rect 4896 4684 4948 4690
rect 4896 4626 4948 4632
rect 5080 4684 5132 4690
rect 5080 4626 5132 4632
rect 4804 3528 4856 3534
rect 4804 3470 4856 3476
rect 4816 2990 4844 3470
rect 4804 2984 4856 2990
rect 4804 2926 4856 2932
rect 4908 2922 4936 4626
rect 5540 4548 5592 4554
rect 5540 4490 5592 4496
rect 5552 4078 5580 4490
rect 5644 4146 5672 5646
rect 6104 4758 6132 5646
rect 6472 5234 6500 5714
rect 6552 5704 6604 5710
rect 6552 5646 6604 5652
rect 6460 5228 6512 5234
rect 6460 5170 6512 5176
rect 6092 4752 6144 4758
rect 6092 4694 6144 4700
rect 6460 4616 6512 4622
rect 6460 4558 6512 4564
rect 5816 4548 5868 4554
rect 5816 4490 5868 4496
rect 5632 4140 5684 4146
rect 5632 4082 5684 4088
rect 5540 4072 5592 4078
rect 5540 4014 5592 4020
rect 5724 3936 5776 3942
rect 5724 3878 5776 3884
rect 5170 3836 5478 3845
rect 5170 3834 5176 3836
rect 5232 3834 5256 3836
rect 5312 3834 5336 3836
rect 5392 3834 5416 3836
rect 5472 3834 5478 3836
rect 5232 3782 5234 3834
rect 5414 3782 5416 3834
rect 5170 3780 5176 3782
rect 5232 3780 5256 3782
rect 5312 3780 5336 3782
rect 5392 3780 5416 3782
rect 5472 3780 5478 3782
rect 5170 3771 5478 3780
rect 5080 2984 5132 2990
rect 5080 2926 5132 2932
rect 4896 2916 4948 2922
rect 4896 2858 4948 2864
rect 4528 2508 4580 2514
rect 4528 2450 4580 2456
rect 4122 1414 4476 1442
rect 4066 1391 4122 1400
rect 4540 800 4568 2450
rect 5092 1714 5120 2926
rect 5170 2748 5478 2757
rect 5170 2746 5176 2748
rect 5232 2746 5256 2748
rect 5312 2746 5336 2748
rect 5392 2746 5416 2748
rect 5472 2746 5478 2748
rect 5232 2694 5234 2746
rect 5414 2694 5416 2746
rect 5170 2692 5176 2694
rect 5232 2692 5256 2694
rect 5312 2692 5336 2694
rect 5392 2692 5416 2694
rect 5472 2692 5478 2694
rect 5170 2683 5478 2692
rect 5736 2378 5764 3878
rect 5724 2372 5776 2378
rect 5724 2314 5776 2320
rect 5828 2310 5856 4490
rect 6472 4010 6500 4558
rect 6564 4146 6592 5646
rect 6736 5568 6788 5574
rect 6736 5510 6788 5516
rect 6552 4140 6604 4146
rect 6552 4082 6604 4088
rect 6564 4010 6592 4082
rect 6460 4004 6512 4010
rect 6460 3946 6512 3952
rect 6552 4004 6604 4010
rect 6552 3946 6604 3952
rect 6092 3936 6144 3942
rect 6092 3878 6144 3884
rect 6104 3602 6132 3878
rect 6092 3596 6144 3602
rect 6092 3538 6144 3544
rect 6460 3596 6512 3602
rect 6460 3538 6512 3544
rect 5816 2304 5868 2310
rect 5816 2246 5868 2252
rect 5092 1686 5212 1714
rect 5184 800 5212 1686
rect 6472 800 6500 3538
rect 6748 2514 6776 5510
rect 7208 5234 7236 6666
rect 9390 6556 9698 6565
rect 9390 6554 9396 6556
rect 9452 6554 9476 6556
rect 9532 6554 9556 6556
rect 9612 6554 9636 6556
rect 9692 6554 9698 6556
rect 9452 6502 9454 6554
rect 9634 6502 9636 6554
rect 9390 6500 9396 6502
rect 9452 6500 9476 6502
rect 9532 6500 9556 6502
rect 9612 6500 9636 6502
rect 9692 6500 9698 6502
rect 9390 6491 9698 6500
rect 10508 6316 10560 6322
rect 10508 6258 10560 6264
rect 7380 5704 7432 5710
rect 7380 5646 7432 5652
rect 7196 5228 7248 5234
rect 7196 5170 7248 5176
rect 7208 4622 7236 5170
rect 7196 4616 7248 4622
rect 7196 4558 7248 4564
rect 6920 4480 6972 4486
rect 6920 4422 6972 4428
rect 6932 3194 6960 4422
rect 7196 3936 7248 3942
rect 7196 3878 7248 3884
rect 7012 3460 7064 3466
rect 7012 3402 7064 3408
rect 6920 3188 6972 3194
rect 6920 3130 6972 3136
rect 7024 3058 7052 3402
rect 7208 3126 7236 3878
rect 7196 3120 7248 3126
rect 7196 3062 7248 3068
rect 7012 3052 7064 3058
rect 7012 2994 7064 3000
rect 6828 2848 6880 2854
rect 6828 2790 6880 2796
rect 6840 2514 6868 2790
rect 7392 2582 7420 5646
rect 9390 5468 9698 5477
rect 9390 5466 9396 5468
rect 9452 5466 9476 5468
rect 9532 5466 9556 5468
rect 9612 5466 9636 5468
rect 9692 5466 9698 5468
rect 9452 5414 9454 5466
rect 9634 5414 9636 5466
rect 9390 5412 9396 5414
rect 9452 5412 9476 5414
rect 9532 5412 9556 5414
rect 9612 5412 9636 5414
rect 9692 5412 9698 5414
rect 9390 5403 9698 5412
rect 8024 4684 8076 4690
rect 8024 4626 8076 4632
rect 8036 4146 8064 4626
rect 8392 4616 8444 4622
rect 8392 4558 8444 4564
rect 8024 4140 8076 4146
rect 8024 4082 8076 4088
rect 8036 3194 8064 4082
rect 8404 3670 8432 4558
rect 9390 4380 9698 4389
rect 9390 4378 9396 4380
rect 9452 4378 9476 4380
rect 9532 4378 9556 4380
rect 9612 4378 9636 4380
rect 9692 4378 9698 4380
rect 9452 4326 9454 4378
rect 9634 4326 9636 4378
rect 9390 4324 9396 4326
rect 9452 4324 9476 4326
rect 9532 4324 9556 4326
rect 9612 4324 9636 4326
rect 9692 4324 9698 4326
rect 9390 4315 9698 4324
rect 9128 4140 9180 4146
rect 9128 4082 9180 4088
rect 8392 3664 8444 3670
rect 8392 3606 8444 3612
rect 9140 3466 9168 4082
rect 9220 3936 9272 3942
rect 9220 3878 9272 3884
rect 9128 3460 9180 3466
rect 9128 3402 9180 3408
rect 8024 3188 8076 3194
rect 8024 3130 8076 3136
rect 8392 2984 8444 2990
rect 8392 2926 8444 2932
rect 7380 2576 7432 2582
rect 7380 2518 7432 2524
rect 6736 2508 6788 2514
rect 6736 2450 6788 2456
rect 6828 2508 6880 2514
rect 6828 2450 6880 2456
rect 8404 800 8432 2926
rect 9232 2394 9260 3878
rect 10520 3670 10548 6258
rect 13611 6012 13919 6021
rect 13611 6010 13617 6012
rect 13673 6010 13697 6012
rect 13753 6010 13777 6012
rect 13833 6010 13857 6012
rect 13913 6010 13919 6012
rect 13673 5958 13675 6010
rect 13855 5958 13857 6010
rect 13611 5956 13617 5958
rect 13673 5956 13697 5958
rect 13753 5956 13777 5958
rect 13833 5956 13857 5958
rect 13913 5956 13919 5958
rect 13611 5947 13919 5956
rect 13176 5160 13228 5166
rect 13176 5102 13228 5108
rect 13084 4072 13136 4078
rect 13084 4014 13136 4020
rect 13096 3738 13124 4014
rect 13084 3732 13136 3738
rect 13084 3674 13136 3680
rect 10508 3664 10560 3670
rect 10508 3606 10560 3612
rect 10520 3534 10548 3606
rect 9312 3528 9364 3534
rect 9312 3470 9364 3476
rect 10048 3528 10100 3534
rect 10048 3470 10100 3476
rect 10508 3528 10560 3534
rect 10508 3470 10560 3476
rect 9324 2514 9352 3470
rect 9772 3392 9824 3398
rect 9772 3334 9824 3340
rect 9390 3292 9698 3301
rect 9390 3290 9396 3292
rect 9452 3290 9476 3292
rect 9532 3290 9556 3292
rect 9612 3290 9636 3292
rect 9692 3290 9698 3292
rect 9452 3238 9454 3290
rect 9634 3238 9636 3290
rect 9390 3236 9396 3238
rect 9452 3236 9476 3238
rect 9532 3236 9556 3238
rect 9612 3236 9636 3238
rect 9692 3236 9698 3238
rect 9390 3227 9698 3236
rect 9784 3126 9812 3334
rect 9772 3120 9824 3126
rect 9772 3062 9824 3068
rect 10060 2990 10088 3470
rect 13188 3058 13216 5102
rect 13611 4924 13919 4933
rect 13611 4922 13617 4924
rect 13673 4922 13697 4924
rect 13753 4922 13777 4924
rect 13833 4922 13857 4924
rect 13913 4922 13919 4924
rect 13673 4870 13675 4922
rect 13855 4870 13857 4922
rect 13611 4868 13617 4870
rect 13673 4868 13697 4870
rect 13753 4868 13777 4870
rect 13833 4868 13857 4870
rect 13913 4868 13919 4870
rect 13611 4859 13919 4868
rect 13268 4072 13320 4078
rect 13268 4014 13320 4020
rect 13452 4072 13504 4078
rect 13452 4014 13504 4020
rect 13280 3194 13308 4014
rect 13268 3188 13320 3194
rect 13268 3130 13320 3136
rect 13176 3052 13228 3058
rect 13176 2994 13228 3000
rect 10048 2984 10100 2990
rect 10048 2926 10100 2932
rect 10324 2984 10376 2990
rect 10324 2926 10376 2932
rect 9312 2508 9364 2514
rect 9312 2450 9364 2456
rect 9772 2508 9824 2514
rect 9772 2450 9824 2456
rect 9232 2378 9352 2394
rect 9232 2372 9364 2378
rect 9232 2366 9312 2372
rect 9312 2314 9364 2320
rect 9390 2204 9698 2213
rect 9390 2202 9396 2204
rect 9452 2202 9476 2204
rect 9532 2202 9556 2204
rect 9612 2202 9636 2204
rect 9692 2202 9698 2204
rect 9452 2150 9454 2202
rect 9634 2150 9636 2202
rect 9390 2148 9396 2150
rect 9452 2148 9476 2150
rect 9532 2148 9556 2150
rect 9612 2148 9636 2150
rect 9692 2148 9698 2150
rect 9390 2139 9698 2148
rect 9784 1306 9812 2450
rect 9692 1278 9812 1306
rect 9692 800 9720 1278
rect 10336 800 10364 2926
rect 13464 2258 13492 4014
rect 13611 3836 13919 3845
rect 13611 3834 13617 3836
rect 13673 3834 13697 3836
rect 13753 3834 13777 3836
rect 13833 3834 13857 3836
rect 13913 3834 13919 3836
rect 13673 3782 13675 3834
rect 13855 3782 13857 3834
rect 13611 3780 13617 3782
rect 13673 3780 13697 3782
rect 13753 3780 13777 3782
rect 13833 3780 13857 3782
rect 13913 3780 13919 3782
rect 13611 3771 13919 3780
rect 14384 3670 14412 12174
rect 17831 11996 18139 12005
rect 17831 11994 17837 11996
rect 17893 11994 17917 11996
rect 17973 11994 17997 11996
rect 18053 11994 18077 11996
rect 18133 11994 18139 11996
rect 17893 11942 17895 11994
rect 18075 11942 18077 11994
rect 17831 11940 17837 11942
rect 17893 11940 17917 11942
rect 17973 11940 17997 11942
rect 18053 11940 18077 11942
rect 18133 11940 18139 11942
rect 17831 11931 18139 11940
rect 17831 10908 18139 10917
rect 17831 10906 17837 10908
rect 17893 10906 17917 10908
rect 17973 10906 17997 10908
rect 18053 10906 18077 10908
rect 18133 10906 18139 10908
rect 17893 10854 17895 10906
rect 18075 10854 18077 10906
rect 17831 10852 17837 10854
rect 17893 10852 17917 10854
rect 17973 10852 17997 10854
rect 18053 10852 18077 10854
rect 18133 10852 18139 10854
rect 17831 10843 18139 10852
rect 17831 9820 18139 9829
rect 17831 9818 17837 9820
rect 17893 9818 17917 9820
rect 17973 9818 17997 9820
rect 18053 9818 18077 9820
rect 18133 9818 18139 9820
rect 17893 9766 17895 9818
rect 18075 9766 18077 9818
rect 17831 9764 17837 9766
rect 17893 9764 17917 9766
rect 17973 9764 17997 9766
rect 18053 9764 18077 9766
rect 18133 9764 18139 9766
rect 17831 9755 18139 9764
rect 17831 8732 18139 8741
rect 17831 8730 17837 8732
rect 17893 8730 17917 8732
rect 17973 8730 17997 8732
rect 18053 8730 18077 8732
rect 18133 8730 18139 8732
rect 17893 8678 17895 8730
rect 18075 8678 18077 8730
rect 17831 8676 17837 8678
rect 17893 8676 17917 8678
rect 17973 8676 17997 8678
rect 18053 8676 18077 8678
rect 18133 8676 18139 8678
rect 17831 8667 18139 8676
rect 17831 7644 18139 7653
rect 17831 7642 17837 7644
rect 17893 7642 17917 7644
rect 17973 7642 17997 7644
rect 18053 7642 18077 7644
rect 18133 7642 18139 7644
rect 17893 7590 17895 7642
rect 18075 7590 18077 7642
rect 17831 7588 17837 7590
rect 17893 7588 17917 7590
rect 17973 7588 17997 7590
rect 18053 7588 18077 7590
rect 18133 7588 18139 7590
rect 17831 7579 18139 7588
rect 19168 6914 19196 27406
rect 19260 26353 19288 28478
rect 19432 27464 19484 27470
rect 19432 27406 19484 27412
rect 19340 27328 19392 27334
rect 19340 27270 19392 27276
rect 19352 26382 19380 27270
rect 19444 26994 19472 27406
rect 19524 27396 19576 27402
rect 19524 27338 19576 27344
rect 19432 26988 19484 26994
rect 19432 26930 19484 26936
rect 19432 26512 19484 26518
rect 19536 26500 19564 27338
rect 19720 27062 19748 33050
rect 19812 32910 19840 33798
rect 19800 32904 19852 32910
rect 19800 32846 19852 32852
rect 19904 31226 19932 35974
rect 19984 35488 20036 35494
rect 19984 35430 20036 35436
rect 19996 34678 20024 35430
rect 19984 34672 20036 34678
rect 19984 34614 20036 34620
rect 20076 33856 20128 33862
rect 20076 33798 20128 33804
rect 19982 33688 20038 33697
rect 19982 33623 19984 33632
rect 20036 33623 20038 33632
rect 19984 33594 20036 33600
rect 20088 31754 20116 33798
rect 20180 32774 20208 35974
rect 20260 35012 20312 35018
rect 20260 34954 20312 34960
rect 20272 34746 20300 34954
rect 20444 34944 20496 34950
rect 20444 34886 20496 34892
rect 20260 34740 20312 34746
rect 20260 34682 20312 34688
rect 20272 33522 20300 34682
rect 20352 33992 20404 33998
rect 20352 33934 20404 33940
rect 20364 33658 20392 33934
rect 20352 33652 20404 33658
rect 20352 33594 20404 33600
rect 20456 33522 20484 34886
rect 20548 34474 20576 36518
rect 20628 36168 20680 36174
rect 20628 36110 20680 36116
rect 20640 35737 20668 36110
rect 21088 36032 21140 36038
rect 21088 35974 21140 35980
rect 20626 35728 20682 35737
rect 20626 35663 20682 35672
rect 20720 35692 20772 35698
rect 20720 35634 20772 35640
rect 20996 35692 21048 35698
rect 20996 35634 21048 35640
rect 20628 35624 20680 35630
rect 20628 35566 20680 35572
rect 20640 35290 20668 35566
rect 20628 35284 20680 35290
rect 20628 35226 20680 35232
rect 20640 34950 20668 35226
rect 20628 34944 20680 34950
rect 20628 34886 20680 34892
rect 20640 34746 20668 34886
rect 20732 34746 20760 35634
rect 21008 35086 21036 35634
rect 20996 35080 21048 35086
rect 20996 35022 21048 35028
rect 20812 34944 20864 34950
rect 20812 34886 20864 34892
rect 20628 34740 20680 34746
rect 20628 34682 20680 34688
rect 20720 34740 20772 34746
rect 20720 34682 20772 34688
rect 20536 34468 20588 34474
rect 20536 34410 20588 34416
rect 20824 34134 20852 34886
rect 20996 34536 21048 34542
rect 20996 34478 21048 34484
rect 20812 34128 20864 34134
rect 20812 34070 20864 34076
rect 21008 33998 21036 34478
rect 20996 33992 21048 33998
rect 20996 33934 21048 33940
rect 21100 33930 21128 35974
rect 21192 33969 21220 37606
rect 21376 37466 21404 38247
rect 21456 37664 21508 37670
rect 21456 37606 21508 37612
rect 21364 37460 21416 37466
rect 21364 37402 21416 37408
rect 21468 37330 21496 37606
rect 21456 37324 21508 37330
rect 21456 37266 21508 37272
rect 21928 37262 21956 38814
rect 22052 38652 22360 38661
rect 22052 38650 22058 38652
rect 22114 38650 22138 38652
rect 22194 38650 22218 38652
rect 22274 38650 22298 38652
rect 22354 38650 22360 38652
rect 22114 38598 22116 38650
rect 22296 38598 22298 38650
rect 22052 38596 22058 38598
rect 22114 38596 22138 38598
rect 22194 38596 22218 38598
rect 22274 38596 22298 38598
rect 22354 38596 22360 38598
rect 22052 38587 22360 38596
rect 22388 38554 22416 38830
rect 23860 38758 23888 39374
rect 24400 39364 24452 39370
rect 24400 39306 24452 39312
rect 24412 38962 24440 39306
rect 24584 39296 24636 39302
rect 24584 39238 24636 39244
rect 24596 39030 24624 39238
rect 24584 39024 24636 39030
rect 24584 38966 24636 38972
rect 24400 38956 24452 38962
rect 24400 38898 24452 38904
rect 25148 38894 25176 41200
rect 25228 39636 25280 39642
rect 25228 39578 25280 39584
rect 25136 38888 25188 38894
rect 25136 38830 25188 38836
rect 23848 38752 23900 38758
rect 23848 38694 23900 38700
rect 22376 38548 22428 38554
rect 22376 38490 22428 38496
rect 23480 38004 23532 38010
rect 23480 37946 23532 37952
rect 22192 37936 22244 37942
rect 22192 37878 22244 37884
rect 22204 37738 22232 37878
rect 23492 37874 23520 37946
rect 23754 37904 23810 37913
rect 23480 37868 23532 37874
rect 23754 37839 23810 37848
rect 23480 37810 23532 37816
rect 22192 37732 22244 37738
rect 22192 37674 22244 37680
rect 22052 37564 22360 37573
rect 22052 37562 22058 37564
rect 22114 37562 22138 37564
rect 22194 37562 22218 37564
rect 22274 37562 22298 37564
rect 22354 37562 22360 37564
rect 22114 37510 22116 37562
rect 22296 37510 22298 37562
rect 22052 37508 22058 37510
rect 22114 37508 22138 37510
rect 22194 37508 22218 37510
rect 22274 37508 22298 37510
rect 22354 37508 22360 37510
rect 22052 37499 22360 37508
rect 21916 37256 21968 37262
rect 21916 37198 21968 37204
rect 22468 37256 22520 37262
rect 22468 37198 22520 37204
rect 22744 37256 22796 37262
rect 22744 37198 22796 37204
rect 22376 36780 22428 36786
rect 22376 36722 22428 36728
rect 22052 36476 22360 36485
rect 22052 36474 22058 36476
rect 22114 36474 22138 36476
rect 22194 36474 22218 36476
rect 22274 36474 22298 36476
rect 22354 36474 22360 36476
rect 22114 36422 22116 36474
rect 22296 36422 22298 36474
rect 22052 36420 22058 36422
rect 22114 36420 22138 36422
rect 22194 36420 22218 36422
rect 22274 36420 22298 36422
rect 22354 36420 22360 36422
rect 22052 36411 22360 36420
rect 21272 36168 21324 36174
rect 21272 36110 21324 36116
rect 21916 36168 21968 36174
rect 21916 36110 21968 36116
rect 21284 35834 21312 36110
rect 21272 35828 21324 35834
rect 21272 35770 21324 35776
rect 21272 35692 21324 35698
rect 21272 35634 21324 35640
rect 21284 34610 21312 35634
rect 21364 35216 21416 35222
rect 21364 35158 21416 35164
rect 21272 34604 21324 34610
rect 21272 34546 21324 34552
rect 21272 34400 21324 34406
rect 21272 34342 21324 34348
rect 21178 33960 21234 33969
rect 21088 33924 21140 33930
rect 21284 33930 21312 34342
rect 21178 33895 21234 33904
rect 21272 33924 21324 33930
rect 21088 33866 21140 33872
rect 21272 33866 21324 33872
rect 21270 33552 21326 33561
rect 20260 33516 20312 33522
rect 20260 33458 20312 33464
rect 20444 33516 20496 33522
rect 20444 33458 20496 33464
rect 20628 33516 20680 33522
rect 21270 33487 21272 33496
rect 20628 33458 20680 33464
rect 21324 33487 21326 33496
rect 21272 33458 21324 33464
rect 20640 33114 20668 33458
rect 20628 33108 20680 33114
rect 20628 33050 20680 33056
rect 20626 33008 20682 33017
rect 20626 32943 20628 32952
rect 20680 32943 20682 32952
rect 20628 32914 20680 32920
rect 20168 32768 20220 32774
rect 20168 32710 20220 32716
rect 20628 32768 20680 32774
rect 20628 32710 20680 32716
rect 20904 32768 20956 32774
rect 20904 32710 20956 32716
rect 20640 32570 20668 32710
rect 20628 32564 20680 32570
rect 20628 32506 20680 32512
rect 20444 32428 20496 32434
rect 20444 32370 20496 32376
rect 20352 31884 20404 31890
rect 20352 31826 20404 31832
rect 20088 31726 20300 31754
rect 19904 31198 20116 31226
rect 19892 31136 19944 31142
rect 19892 31078 19944 31084
rect 19904 30666 19932 31078
rect 19984 30864 20036 30870
rect 19984 30806 20036 30812
rect 19892 30660 19944 30666
rect 19892 30602 19944 30608
rect 19800 30592 19852 30598
rect 19800 30534 19852 30540
rect 19812 29782 19840 30534
rect 19800 29776 19852 29782
rect 19800 29718 19852 29724
rect 19996 29646 20024 30806
rect 19984 29640 20036 29646
rect 19984 29582 20036 29588
rect 20088 29238 20116 31198
rect 20168 30592 20220 30598
rect 20168 30534 20220 30540
rect 20180 29782 20208 30534
rect 20168 29776 20220 29782
rect 20168 29718 20220 29724
rect 20272 29510 20300 31726
rect 20364 30802 20392 31826
rect 20456 31822 20484 32370
rect 20916 32366 20944 32710
rect 21272 32496 21324 32502
rect 21272 32438 21324 32444
rect 21088 32428 21140 32434
rect 21088 32370 21140 32376
rect 20904 32360 20956 32366
rect 20904 32302 20956 32308
rect 20720 32224 20772 32230
rect 20720 32166 20772 32172
rect 20444 31816 20496 31822
rect 20444 31758 20496 31764
rect 20352 30796 20404 30802
rect 20352 30738 20404 30744
rect 20260 29504 20312 29510
rect 20260 29446 20312 29452
rect 20456 29238 20484 31758
rect 20628 31748 20680 31754
rect 20628 31690 20680 31696
rect 20640 31385 20668 31690
rect 20732 31414 20760 32166
rect 20812 31748 20864 31754
rect 20812 31690 20864 31696
rect 20824 31482 20852 31690
rect 20812 31476 20864 31482
rect 20812 31418 20864 31424
rect 21100 31414 21128 32370
rect 21284 32026 21312 32438
rect 21272 32020 21324 32026
rect 21272 31962 21324 31968
rect 21376 31906 21404 35158
rect 21456 35148 21508 35154
rect 21456 35090 21508 35096
rect 21468 35057 21496 35090
rect 21454 35048 21510 35057
rect 21454 34983 21510 34992
rect 21640 34944 21692 34950
rect 21640 34886 21692 34892
rect 21456 34604 21508 34610
rect 21456 34546 21508 34552
rect 21468 33658 21496 34546
rect 21548 34400 21600 34406
rect 21548 34342 21600 34348
rect 21560 34202 21588 34342
rect 21548 34196 21600 34202
rect 21548 34138 21600 34144
rect 21456 33652 21508 33658
rect 21508 33612 21588 33640
rect 21456 33594 21508 33600
rect 21560 32910 21588 33612
rect 21652 33454 21680 34886
rect 21732 34604 21784 34610
rect 21732 34546 21784 34552
rect 21744 33810 21772 34546
rect 21824 34468 21876 34474
rect 21824 34410 21876 34416
rect 21836 34202 21864 34410
rect 21824 34196 21876 34202
rect 21824 34138 21876 34144
rect 21744 33782 21864 33810
rect 21730 33688 21786 33697
rect 21730 33623 21732 33632
rect 21784 33623 21786 33632
rect 21732 33594 21784 33600
rect 21836 33522 21864 33782
rect 21824 33516 21876 33522
rect 21824 33458 21876 33464
rect 21640 33448 21692 33454
rect 21640 33390 21692 33396
rect 21928 33114 21956 36110
rect 22282 35864 22338 35873
rect 22388 35834 22416 36722
rect 22480 36417 22508 37198
rect 22560 36576 22612 36582
rect 22560 36518 22612 36524
rect 22466 36408 22522 36417
rect 22466 36343 22522 36352
rect 22468 36032 22520 36038
rect 22468 35974 22520 35980
rect 22282 35799 22338 35808
rect 22376 35828 22428 35834
rect 22296 35476 22324 35799
rect 22376 35770 22428 35776
rect 22296 35448 22416 35476
rect 22052 35388 22360 35397
rect 22052 35386 22058 35388
rect 22114 35386 22138 35388
rect 22194 35386 22218 35388
rect 22274 35386 22298 35388
rect 22354 35386 22360 35388
rect 22114 35334 22116 35386
rect 22296 35334 22298 35386
rect 22052 35332 22058 35334
rect 22114 35332 22138 35334
rect 22194 35332 22218 35334
rect 22274 35332 22298 35334
rect 22354 35332 22360 35334
rect 22052 35323 22360 35332
rect 22388 35290 22416 35448
rect 22376 35284 22428 35290
rect 22376 35226 22428 35232
rect 22192 35080 22244 35086
rect 22192 35022 22244 35028
rect 22204 34950 22232 35022
rect 22376 35012 22428 35018
rect 22376 34954 22428 34960
rect 22192 34944 22244 34950
rect 22192 34886 22244 34892
rect 22052 34300 22360 34309
rect 22052 34298 22058 34300
rect 22114 34298 22138 34300
rect 22194 34298 22218 34300
rect 22274 34298 22298 34300
rect 22354 34298 22360 34300
rect 22114 34246 22116 34298
rect 22296 34246 22298 34298
rect 22052 34244 22058 34246
rect 22114 34244 22138 34246
rect 22194 34244 22218 34246
rect 22274 34244 22298 34246
rect 22354 34244 22360 34246
rect 22052 34235 22360 34244
rect 22388 34202 22416 34954
rect 22008 34196 22060 34202
rect 22008 34138 22060 34144
rect 22376 34196 22428 34202
rect 22376 34138 22428 34144
rect 22020 33930 22048 34138
rect 22008 33924 22060 33930
rect 22008 33866 22060 33872
rect 22052 33212 22360 33221
rect 22052 33210 22058 33212
rect 22114 33210 22138 33212
rect 22194 33210 22218 33212
rect 22274 33210 22298 33212
rect 22354 33210 22360 33212
rect 22114 33158 22116 33210
rect 22296 33158 22298 33210
rect 22052 33156 22058 33158
rect 22114 33156 22138 33158
rect 22194 33156 22218 33158
rect 22274 33156 22298 33158
rect 22354 33156 22360 33158
rect 22052 33147 22360 33156
rect 21916 33108 21968 33114
rect 21916 33050 21968 33056
rect 21548 32904 21600 32910
rect 21548 32846 21600 32852
rect 22388 32842 22416 34138
rect 22480 33590 22508 35974
rect 22572 34610 22600 36518
rect 22756 36378 22784 37198
rect 23492 37097 23520 37810
rect 23768 37670 23796 37839
rect 23756 37664 23808 37670
rect 23756 37606 23808 37612
rect 23572 37120 23624 37126
rect 23478 37088 23534 37097
rect 23572 37062 23624 37068
rect 23478 37023 23534 37032
rect 22928 36780 22980 36786
rect 22928 36722 22980 36728
rect 22940 36378 22968 36722
rect 23388 36576 23440 36582
rect 23388 36518 23440 36524
rect 22744 36372 22796 36378
rect 22744 36314 22796 36320
rect 22928 36372 22980 36378
rect 22928 36314 22980 36320
rect 22756 36258 22784 36314
rect 23294 36272 23350 36281
rect 22756 36230 22876 36258
rect 22652 36168 22704 36174
rect 22652 36110 22704 36116
rect 22744 36168 22796 36174
rect 22744 36110 22796 36116
rect 22664 34746 22692 36110
rect 22756 35698 22784 36110
rect 22744 35692 22796 35698
rect 22744 35634 22796 35640
rect 22756 35154 22784 35634
rect 22744 35148 22796 35154
rect 22744 35090 22796 35096
rect 22742 35048 22798 35057
rect 22742 34983 22798 34992
rect 22756 34950 22784 34983
rect 22744 34944 22796 34950
rect 22744 34886 22796 34892
rect 22652 34740 22704 34746
rect 22652 34682 22704 34688
rect 22560 34604 22612 34610
rect 22560 34546 22612 34552
rect 22664 34134 22692 34682
rect 22652 34128 22704 34134
rect 22652 34070 22704 34076
rect 22468 33584 22520 33590
rect 22468 33526 22520 33532
rect 22848 33266 22876 36230
rect 23294 36207 23350 36216
rect 23308 36174 23336 36207
rect 23296 36168 23348 36174
rect 23296 36110 23348 36116
rect 22928 35624 22980 35630
rect 22928 35566 22980 35572
rect 22940 35290 22968 35566
rect 23112 35488 23164 35494
rect 23112 35430 23164 35436
rect 22928 35284 22980 35290
rect 22928 35226 22980 35232
rect 22940 33862 22968 35226
rect 23124 35222 23152 35430
rect 23308 35290 23336 36110
rect 23400 35714 23428 36518
rect 23584 36174 23612 37062
rect 23664 36576 23716 36582
rect 23664 36518 23716 36524
rect 23572 36168 23624 36174
rect 23572 36110 23624 36116
rect 23400 35686 23520 35714
rect 23388 35624 23440 35630
rect 23388 35566 23440 35572
rect 23296 35284 23348 35290
rect 23296 35226 23348 35232
rect 23112 35216 23164 35222
rect 23112 35158 23164 35164
rect 23020 34400 23072 34406
rect 23020 34342 23072 34348
rect 23032 34066 23060 34342
rect 23020 34060 23072 34066
rect 23020 34002 23072 34008
rect 23124 33930 23152 35158
rect 23296 35080 23348 35086
rect 23296 35022 23348 35028
rect 23308 34746 23336 35022
rect 23296 34740 23348 34746
rect 23296 34682 23348 34688
rect 23400 34610 23428 35566
rect 23388 34604 23440 34610
rect 23388 34546 23440 34552
rect 23492 34241 23520 35686
rect 23572 35012 23624 35018
rect 23572 34954 23624 34960
rect 23478 34232 23534 34241
rect 23478 34167 23534 34176
rect 23584 33930 23612 34954
rect 23676 34678 23704 36518
rect 23664 34672 23716 34678
rect 23664 34614 23716 34620
rect 23756 34468 23808 34474
rect 23860 34456 23888 38694
rect 25044 38480 25096 38486
rect 25044 38422 25096 38428
rect 24860 38344 24912 38350
rect 24860 38286 24912 38292
rect 24308 38208 24360 38214
rect 24308 38150 24360 38156
rect 24492 38208 24544 38214
rect 24492 38150 24544 38156
rect 24320 37738 24348 38150
rect 24504 38010 24532 38150
rect 24492 38004 24544 38010
rect 24492 37946 24544 37952
rect 24400 37868 24452 37874
rect 24400 37810 24452 37816
rect 24308 37732 24360 37738
rect 24308 37674 24360 37680
rect 24124 37664 24176 37670
rect 24124 37606 24176 37612
rect 24030 37496 24086 37505
rect 24030 37431 24086 37440
rect 24044 37262 24072 37431
rect 24032 37256 24084 37262
rect 24032 37198 24084 37204
rect 24136 35057 24164 37606
rect 24412 37466 24440 37810
rect 24872 37466 24900 38286
rect 25056 37874 25084 38422
rect 25136 38276 25188 38282
rect 25136 38218 25188 38224
rect 25148 37942 25176 38218
rect 25136 37936 25188 37942
rect 25136 37878 25188 37884
rect 25044 37868 25096 37874
rect 25044 37810 25096 37816
rect 25056 37777 25084 37810
rect 25042 37768 25098 37777
rect 25042 37703 25098 37712
rect 24400 37460 24452 37466
rect 24400 37402 24452 37408
rect 24860 37460 24912 37466
rect 24860 37402 24912 37408
rect 24676 37256 24728 37262
rect 24676 37198 24728 37204
rect 24688 37097 24716 37198
rect 24768 37120 24820 37126
rect 24674 37088 24730 37097
rect 24768 37062 24820 37068
rect 24674 37023 24730 37032
rect 24492 36780 24544 36786
rect 24492 36722 24544 36728
rect 24308 36576 24360 36582
rect 24308 36518 24360 36524
rect 24320 35766 24348 36518
rect 24504 35873 24532 36722
rect 24676 36032 24728 36038
rect 24676 35974 24728 35980
rect 24490 35864 24546 35873
rect 24490 35799 24546 35808
rect 24308 35760 24360 35766
rect 24308 35702 24360 35708
rect 24584 35148 24636 35154
rect 24584 35090 24636 35096
rect 24122 35048 24178 35057
rect 24122 34983 24178 34992
rect 24596 34746 24624 35090
rect 23940 34740 23992 34746
rect 23940 34682 23992 34688
rect 24584 34740 24636 34746
rect 24584 34682 24636 34688
rect 23952 34610 23980 34682
rect 24216 34672 24268 34678
rect 24216 34614 24268 34620
rect 23940 34604 23992 34610
rect 23940 34546 23992 34552
rect 23808 34428 23888 34456
rect 23756 34410 23808 34416
rect 24228 33998 24256 34614
rect 24400 34604 24452 34610
rect 24400 34546 24452 34552
rect 24216 33992 24268 33998
rect 24216 33934 24268 33940
rect 23112 33924 23164 33930
rect 23112 33866 23164 33872
rect 23572 33924 23624 33930
rect 23572 33866 23624 33872
rect 22928 33856 22980 33862
rect 22928 33798 22980 33804
rect 23848 33856 23900 33862
rect 23848 33798 23900 33804
rect 22940 33504 22968 33798
rect 23662 33552 23718 33561
rect 22940 33476 23336 33504
rect 23662 33487 23718 33496
rect 23308 33318 23336 33476
rect 23296 33312 23348 33318
rect 22848 33238 22968 33266
rect 23296 33254 23348 33260
rect 23480 33312 23532 33318
rect 23480 33254 23532 33260
rect 22836 32904 22888 32910
rect 22836 32846 22888 32852
rect 22376 32836 22428 32842
rect 22376 32778 22428 32784
rect 22468 32836 22520 32842
rect 22468 32778 22520 32784
rect 22480 32366 22508 32778
rect 22848 32774 22876 32846
rect 22836 32768 22888 32774
rect 22836 32710 22888 32716
rect 22468 32360 22520 32366
rect 22652 32360 22704 32366
rect 22468 32302 22520 32308
rect 22650 32328 22652 32337
rect 22704 32328 22706 32337
rect 22650 32263 22706 32272
rect 21456 32224 21508 32230
rect 21456 32166 21508 32172
rect 21284 31878 21404 31906
rect 20720 31408 20772 31414
rect 20626 31376 20682 31385
rect 20536 31340 20588 31346
rect 20720 31350 20772 31356
rect 21088 31408 21140 31414
rect 21088 31350 21140 31356
rect 20626 31311 20682 31320
rect 20536 31282 20588 31288
rect 20548 29306 20576 31282
rect 21100 30938 21128 31350
rect 21088 30932 21140 30938
rect 21088 30874 21140 30880
rect 21284 29306 21312 31878
rect 21364 31204 21416 31210
rect 21364 31146 21416 31152
rect 21376 30666 21404 31146
rect 21468 30734 21496 32166
rect 22052 32124 22360 32133
rect 22052 32122 22058 32124
rect 22114 32122 22138 32124
rect 22194 32122 22218 32124
rect 22274 32122 22298 32124
rect 22354 32122 22360 32124
rect 22114 32070 22116 32122
rect 22296 32070 22298 32122
rect 22052 32068 22058 32070
rect 22114 32068 22138 32070
rect 22194 32068 22218 32070
rect 22274 32068 22298 32070
rect 22354 32068 22360 32070
rect 22052 32059 22360 32068
rect 22664 31890 22692 32263
rect 22940 31929 22968 33238
rect 23388 32836 23440 32842
rect 23388 32778 23440 32784
rect 23296 32768 23348 32774
rect 23296 32710 23348 32716
rect 23020 32564 23072 32570
rect 23020 32506 23072 32512
rect 23112 32564 23164 32570
rect 23112 32506 23164 32512
rect 22742 31920 22798 31929
rect 22652 31884 22704 31890
rect 22742 31855 22798 31864
rect 22926 31920 22982 31929
rect 22926 31855 22982 31864
rect 22652 31826 22704 31832
rect 22376 31816 22428 31822
rect 22376 31758 22428 31764
rect 22192 31680 22244 31686
rect 22112 31628 22192 31634
rect 22112 31622 22244 31628
rect 22112 31606 22232 31622
rect 22112 31482 22140 31606
rect 22100 31476 22152 31482
rect 22100 31418 22152 31424
rect 21916 31136 21968 31142
rect 21916 31078 21968 31084
rect 21928 30938 21956 31078
rect 22052 31036 22360 31045
rect 22052 31034 22058 31036
rect 22114 31034 22138 31036
rect 22194 31034 22218 31036
rect 22274 31034 22298 31036
rect 22354 31034 22360 31036
rect 22114 30982 22116 31034
rect 22296 30982 22298 31034
rect 22052 30980 22058 30982
rect 22114 30980 22138 30982
rect 22194 30980 22218 30982
rect 22274 30980 22298 30982
rect 22354 30980 22360 30982
rect 22052 30971 22360 30980
rect 21916 30932 21968 30938
rect 21916 30874 21968 30880
rect 21456 30728 21508 30734
rect 21456 30670 21508 30676
rect 21364 30660 21416 30666
rect 21364 30602 21416 30608
rect 21376 30394 21404 30602
rect 21364 30388 21416 30394
rect 21364 30330 21416 30336
rect 21916 30320 21968 30326
rect 21914 30288 21916 30297
rect 21968 30288 21970 30297
rect 21914 30223 21970 30232
rect 22052 29948 22360 29957
rect 22052 29946 22058 29948
rect 22114 29946 22138 29948
rect 22194 29946 22218 29948
rect 22274 29946 22298 29948
rect 22354 29946 22360 29948
rect 22114 29894 22116 29946
rect 22296 29894 22298 29946
rect 22052 29892 22058 29894
rect 22114 29892 22138 29894
rect 22194 29892 22218 29894
rect 22274 29892 22298 29894
rect 22354 29892 22360 29894
rect 22052 29883 22360 29892
rect 21824 29776 21876 29782
rect 21824 29718 21876 29724
rect 20536 29300 20588 29306
rect 20536 29242 20588 29248
rect 20628 29300 20680 29306
rect 20628 29242 20680 29248
rect 21272 29300 21324 29306
rect 21272 29242 21324 29248
rect 20076 29232 20128 29238
rect 20076 29174 20128 29180
rect 20444 29232 20496 29238
rect 20444 29174 20496 29180
rect 20640 28218 20668 29242
rect 21180 29232 21232 29238
rect 21180 29174 21232 29180
rect 20812 28484 20864 28490
rect 20812 28426 20864 28432
rect 20168 28212 20220 28218
rect 20168 28154 20220 28160
rect 20628 28212 20680 28218
rect 20628 28154 20680 28160
rect 20180 27946 20208 28154
rect 20444 28144 20496 28150
rect 20442 28112 20444 28121
rect 20496 28112 20498 28121
rect 20442 28047 20498 28056
rect 20168 27940 20220 27946
rect 20168 27882 20220 27888
rect 20444 27328 20496 27334
rect 20444 27270 20496 27276
rect 19708 27056 19760 27062
rect 19708 26998 19760 27004
rect 20456 26858 20484 27270
rect 20444 26852 20496 26858
rect 20444 26794 20496 26800
rect 19484 26472 19564 26500
rect 19432 26454 19484 26460
rect 20824 26382 20852 28426
rect 21192 28422 21220 29174
rect 21836 29034 21864 29718
rect 22284 29572 22336 29578
rect 22284 29514 22336 29520
rect 22006 29200 22062 29209
rect 22006 29135 22008 29144
rect 22060 29135 22062 29144
rect 22008 29106 22060 29112
rect 22296 29073 22324 29514
rect 22282 29064 22338 29073
rect 21824 29028 21876 29034
rect 22282 28999 22338 29008
rect 21824 28970 21876 28976
rect 21272 28960 21324 28966
rect 21272 28902 21324 28908
rect 21284 28762 21312 28902
rect 22052 28860 22360 28869
rect 22052 28858 22058 28860
rect 22114 28858 22138 28860
rect 22194 28858 22218 28860
rect 22274 28858 22298 28860
rect 22354 28858 22360 28860
rect 22114 28806 22116 28858
rect 22296 28806 22298 28858
rect 22052 28804 22058 28806
rect 22114 28804 22138 28806
rect 22194 28804 22218 28806
rect 22274 28804 22298 28806
rect 22354 28804 22360 28806
rect 22052 28795 22360 28804
rect 22388 28762 22416 31758
rect 22468 31748 22520 31754
rect 22468 31690 22520 31696
rect 22480 31482 22508 31690
rect 22560 31680 22612 31686
rect 22560 31622 22612 31628
rect 22468 31476 22520 31482
rect 22468 31418 22520 31424
rect 22572 30802 22600 31622
rect 22664 31346 22692 31826
rect 22756 31634 22784 31855
rect 22928 31816 22980 31822
rect 22928 31758 22980 31764
rect 22756 31606 22876 31634
rect 22652 31340 22704 31346
rect 22652 31282 22704 31288
rect 22652 30932 22704 30938
rect 22652 30874 22704 30880
rect 22560 30796 22612 30802
rect 22560 30738 22612 30744
rect 22664 30394 22692 30874
rect 22848 30410 22876 31606
rect 22940 30734 22968 31758
rect 22928 30728 22980 30734
rect 22928 30670 22980 30676
rect 23032 30598 23060 32506
rect 23124 32026 23152 32506
rect 23112 32020 23164 32026
rect 23112 31962 23164 31968
rect 23308 31754 23336 32710
rect 23296 31748 23348 31754
rect 23296 31690 23348 31696
rect 23308 30870 23336 31690
rect 23400 31686 23428 32778
rect 23388 31680 23440 31686
rect 23388 31622 23440 31628
rect 23296 30864 23348 30870
rect 23296 30806 23348 30812
rect 23020 30592 23072 30598
rect 23020 30534 23072 30540
rect 22652 30388 22704 30394
rect 22848 30382 23152 30410
rect 23308 30394 23336 30806
rect 22652 30330 22704 30336
rect 22468 30320 22520 30326
rect 22468 30262 22520 30268
rect 22480 29209 22508 30262
rect 22836 30252 22888 30258
rect 22836 30194 22888 30200
rect 22744 30048 22796 30054
rect 22744 29990 22796 29996
rect 22652 29640 22704 29646
rect 22652 29582 22704 29588
rect 22466 29200 22522 29209
rect 22466 29135 22522 29144
rect 22560 29164 22612 29170
rect 22560 29106 22612 29112
rect 21272 28756 21324 28762
rect 21272 28698 21324 28704
rect 22376 28756 22428 28762
rect 22376 28698 22428 28704
rect 22572 28490 22600 29106
rect 22100 28484 22152 28490
rect 22100 28426 22152 28432
rect 22560 28484 22612 28490
rect 22560 28426 22612 28432
rect 21180 28416 21232 28422
rect 21180 28358 21232 28364
rect 22112 28098 22140 28426
rect 22020 28082 22140 28098
rect 22468 28144 22520 28150
rect 22468 28086 22520 28092
rect 22008 28076 22140 28082
rect 22060 28070 22140 28076
rect 22008 28018 22060 28024
rect 22376 27872 22428 27878
rect 22376 27814 22428 27820
rect 22052 27772 22360 27781
rect 22052 27770 22058 27772
rect 22114 27770 22138 27772
rect 22194 27770 22218 27772
rect 22274 27770 22298 27772
rect 22354 27770 22360 27772
rect 22114 27718 22116 27770
rect 22296 27718 22298 27770
rect 22052 27716 22058 27718
rect 22114 27716 22138 27718
rect 22194 27716 22218 27718
rect 22274 27716 22298 27718
rect 22354 27716 22360 27718
rect 22052 27707 22360 27716
rect 21916 27396 21968 27402
rect 21916 27338 21968 27344
rect 21456 26988 21508 26994
rect 21456 26930 21508 26936
rect 21272 26784 21324 26790
rect 21272 26726 21324 26732
rect 19340 26376 19392 26382
rect 19246 26344 19302 26353
rect 19340 26318 19392 26324
rect 20812 26376 20864 26382
rect 20812 26318 20864 26324
rect 19246 26279 19302 26288
rect 20536 26308 20588 26314
rect 19260 23769 19288 26279
rect 20536 26250 20588 26256
rect 20074 25936 20130 25945
rect 19432 25900 19484 25906
rect 20074 25871 20130 25880
rect 19432 25842 19484 25848
rect 19340 25764 19392 25770
rect 19340 25706 19392 25712
rect 19352 24857 19380 25706
rect 19444 25498 19472 25842
rect 19616 25696 19668 25702
rect 19616 25638 19668 25644
rect 19432 25492 19484 25498
rect 19432 25434 19484 25440
rect 19628 25294 19656 25638
rect 20088 25294 20116 25871
rect 20444 25764 20496 25770
rect 20444 25706 20496 25712
rect 19616 25288 19668 25294
rect 19616 25230 19668 25236
rect 19892 25288 19944 25294
rect 19892 25230 19944 25236
rect 20076 25288 20128 25294
rect 20076 25230 20128 25236
rect 19628 24954 19656 25230
rect 19616 24948 19668 24954
rect 19616 24890 19668 24896
rect 19904 24886 19932 25230
rect 19892 24880 19944 24886
rect 19338 24848 19394 24857
rect 19892 24822 19944 24828
rect 19338 24783 19394 24792
rect 20088 24410 20116 25230
rect 20076 24404 20128 24410
rect 20076 24346 20128 24352
rect 19246 23760 19302 23769
rect 19246 23695 19302 23704
rect 20260 23520 20312 23526
rect 20260 23462 20312 23468
rect 19708 23180 19760 23186
rect 19708 23122 19760 23128
rect 20076 23180 20128 23186
rect 20076 23122 20128 23128
rect 19432 22976 19484 22982
rect 19432 22918 19484 22924
rect 19444 22642 19472 22918
rect 19720 22778 19748 23122
rect 19984 23112 20036 23118
rect 19984 23054 20036 23060
rect 19708 22772 19760 22778
rect 19708 22714 19760 22720
rect 19432 22636 19484 22642
rect 19432 22578 19484 22584
rect 19708 21888 19760 21894
rect 19708 21830 19760 21836
rect 19432 21344 19484 21350
rect 19432 21286 19484 21292
rect 19340 20800 19392 20806
rect 19340 20742 19392 20748
rect 19352 20534 19380 20742
rect 19340 20528 19392 20534
rect 19340 20470 19392 20476
rect 19444 20466 19472 21286
rect 19720 21146 19748 21830
rect 19800 21684 19852 21690
rect 19800 21626 19852 21632
rect 19708 21140 19760 21146
rect 19708 21082 19760 21088
rect 19524 20800 19576 20806
rect 19524 20742 19576 20748
rect 19432 20460 19484 20466
rect 19432 20402 19484 20408
rect 19340 20392 19392 20398
rect 19340 20334 19392 20340
rect 19352 19718 19380 20334
rect 19444 19922 19472 20402
rect 19432 19916 19484 19922
rect 19432 19858 19484 19864
rect 19340 19712 19392 19718
rect 19340 19654 19392 19660
rect 19352 19378 19380 19654
rect 19340 19372 19392 19378
rect 19340 19314 19392 19320
rect 19444 18834 19472 19858
rect 19432 18828 19484 18834
rect 19432 18770 19484 18776
rect 19444 18358 19472 18770
rect 19536 18737 19564 20742
rect 19522 18728 19578 18737
rect 19522 18663 19578 18672
rect 19812 18426 19840 21626
rect 19996 20874 20024 23054
rect 20088 22438 20116 23122
rect 20076 22432 20128 22438
rect 20076 22374 20128 22380
rect 20272 21622 20300 23462
rect 20456 23118 20484 25706
rect 20548 24750 20576 26250
rect 20720 25968 20772 25974
rect 20720 25910 20772 25916
rect 20628 25424 20680 25430
rect 20626 25392 20628 25401
rect 20680 25392 20682 25401
rect 20626 25327 20682 25336
rect 20732 25294 20760 25910
rect 20720 25288 20772 25294
rect 20720 25230 20772 25236
rect 20720 24880 20772 24886
rect 20720 24822 20772 24828
rect 20536 24744 20588 24750
rect 20536 24686 20588 24692
rect 20548 23526 20576 24686
rect 20628 24608 20680 24614
rect 20628 24550 20680 24556
rect 20536 23520 20588 23526
rect 20536 23462 20588 23468
rect 20444 23112 20496 23118
rect 20444 23054 20496 23060
rect 20352 23044 20404 23050
rect 20352 22986 20404 22992
rect 20364 22098 20392 22986
rect 20640 22642 20668 24550
rect 20732 23594 20760 24822
rect 20720 23588 20772 23594
rect 20720 23530 20772 23536
rect 20824 23118 20852 26318
rect 20904 25696 20956 25702
rect 20904 25638 20956 25644
rect 21180 25696 21232 25702
rect 21180 25638 21232 25644
rect 20812 23112 20864 23118
rect 20812 23054 20864 23060
rect 20628 22636 20680 22642
rect 20628 22578 20680 22584
rect 20720 22636 20772 22642
rect 20720 22578 20772 22584
rect 20352 22092 20404 22098
rect 20352 22034 20404 22040
rect 20732 22030 20760 22578
rect 20824 22094 20852 23054
rect 20916 22642 20944 25638
rect 21192 24993 21220 25638
rect 21284 25226 21312 26726
rect 21272 25220 21324 25226
rect 21272 25162 21324 25168
rect 21178 24984 21234 24993
rect 21178 24919 21234 24928
rect 21468 24818 21496 26930
rect 21928 25786 21956 27338
rect 22052 26684 22360 26693
rect 22052 26682 22058 26684
rect 22114 26682 22138 26684
rect 22194 26682 22218 26684
rect 22274 26682 22298 26684
rect 22354 26682 22360 26684
rect 22114 26630 22116 26682
rect 22296 26630 22298 26682
rect 22052 26628 22058 26630
rect 22114 26628 22138 26630
rect 22194 26628 22218 26630
rect 22274 26628 22298 26630
rect 22354 26628 22360 26630
rect 22052 26619 22360 26628
rect 22388 25906 22416 27814
rect 22480 27470 22508 28086
rect 22468 27464 22520 27470
rect 22468 27406 22520 27412
rect 22480 27062 22508 27406
rect 22468 27056 22520 27062
rect 22468 26998 22520 27004
rect 22480 26450 22508 26998
rect 22468 26444 22520 26450
rect 22468 26386 22520 26392
rect 22480 25906 22508 26386
rect 22572 26330 22600 28426
rect 22664 27606 22692 29582
rect 22756 29578 22784 29990
rect 22848 29646 22876 30194
rect 23020 30048 23072 30054
rect 23020 29990 23072 29996
rect 22928 29844 22980 29850
rect 22928 29786 22980 29792
rect 22836 29640 22888 29646
rect 22940 29617 22968 29786
rect 22836 29582 22888 29588
rect 22926 29608 22982 29617
rect 22744 29572 22796 29578
rect 22744 29514 22796 29520
rect 22848 29170 22876 29582
rect 22926 29543 22982 29552
rect 22836 29164 22888 29170
rect 22836 29106 22888 29112
rect 23032 29102 23060 29990
rect 23020 29096 23072 29102
rect 23020 29038 23072 29044
rect 23124 28914 23152 30382
rect 23296 30388 23348 30394
rect 23296 30330 23348 30336
rect 23400 29714 23428 31622
rect 23492 31414 23520 33254
rect 23676 32842 23704 33487
rect 23664 32836 23716 32842
rect 23584 32796 23664 32824
rect 23584 31890 23612 32796
rect 23664 32778 23716 32784
rect 23860 32502 23888 33798
rect 24032 33516 24084 33522
rect 24032 33458 24084 33464
rect 24044 33114 24072 33458
rect 24032 33108 24084 33114
rect 24032 33050 24084 33056
rect 24124 32836 24176 32842
rect 24124 32778 24176 32784
rect 23848 32496 23900 32502
rect 23848 32438 23900 32444
rect 23940 32428 23992 32434
rect 23940 32370 23992 32376
rect 23848 32360 23900 32366
rect 23848 32302 23900 32308
rect 23572 31884 23624 31890
rect 23572 31826 23624 31832
rect 23860 31822 23888 32302
rect 23952 32026 23980 32370
rect 24032 32224 24084 32230
rect 24032 32166 24084 32172
rect 23940 32020 23992 32026
rect 23940 31962 23992 31968
rect 23848 31816 23900 31822
rect 23848 31758 23900 31764
rect 23860 31686 23888 31758
rect 23848 31680 23900 31686
rect 23900 31640 23980 31668
rect 23848 31622 23900 31628
rect 23480 31408 23532 31414
rect 23480 31350 23532 31356
rect 23848 31204 23900 31210
rect 23848 31146 23900 31152
rect 23572 31136 23624 31142
rect 23572 31078 23624 31084
rect 23756 31136 23808 31142
rect 23756 31078 23808 31084
rect 23388 29708 23440 29714
rect 23388 29650 23440 29656
rect 23584 29646 23612 31078
rect 23572 29640 23624 29646
rect 23572 29582 23624 29588
rect 23204 29572 23256 29578
rect 23204 29514 23256 29520
rect 23216 29102 23244 29514
rect 23572 29300 23624 29306
rect 23572 29242 23624 29248
rect 23478 29200 23534 29209
rect 23478 29135 23480 29144
rect 23532 29135 23534 29144
rect 23480 29106 23532 29112
rect 23204 29096 23256 29102
rect 23204 29038 23256 29044
rect 23032 28886 23152 28914
rect 22744 28688 22796 28694
rect 22744 28630 22796 28636
rect 22652 27600 22704 27606
rect 22652 27542 22704 27548
rect 22664 27062 22692 27542
rect 22652 27056 22704 27062
rect 22652 26998 22704 27004
rect 22572 26302 22692 26330
rect 22376 25900 22428 25906
rect 22376 25842 22428 25848
rect 22468 25900 22520 25906
rect 22468 25842 22520 25848
rect 21928 25770 22048 25786
rect 21928 25764 22060 25770
rect 21928 25758 22008 25764
rect 22008 25706 22060 25712
rect 22052 25596 22360 25605
rect 22052 25594 22058 25596
rect 22114 25594 22138 25596
rect 22194 25594 22218 25596
rect 22274 25594 22298 25596
rect 22354 25594 22360 25596
rect 22114 25542 22116 25594
rect 22296 25542 22298 25594
rect 22052 25540 22058 25542
rect 22114 25540 22138 25542
rect 22194 25540 22218 25542
rect 22274 25540 22298 25542
rect 22354 25540 22360 25542
rect 22052 25531 22360 25540
rect 22468 25356 22520 25362
rect 22468 25298 22520 25304
rect 21916 25288 21968 25294
rect 21916 25230 21968 25236
rect 21928 24818 21956 25230
rect 21180 24812 21232 24818
rect 21180 24754 21232 24760
rect 21456 24812 21508 24818
rect 21456 24754 21508 24760
rect 21916 24812 21968 24818
rect 21916 24754 21968 24760
rect 20996 24744 21048 24750
rect 20996 24686 21048 24692
rect 21008 24410 21036 24686
rect 20996 24404 21048 24410
rect 20996 24346 21048 24352
rect 21192 24274 21220 24754
rect 21180 24268 21232 24274
rect 21232 24228 21312 24256
rect 21180 24210 21232 24216
rect 21180 24064 21232 24070
rect 21180 24006 21232 24012
rect 20904 22636 20956 22642
rect 20904 22578 20956 22584
rect 20996 22636 21048 22642
rect 20996 22578 21048 22584
rect 20824 22066 20944 22094
rect 20720 22024 20772 22030
rect 20534 21992 20590 22001
rect 20720 21966 20772 21972
rect 20534 21927 20590 21936
rect 20812 21956 20864 21962
rect 20548 21894 20576 21927
rect 20812 21898 20864 21904
rect 20536 21888 20588 21894
rect 20536 21830 20588 21836
rect 20260 21616 20312 21622
rect 20260 21558 20312 21564
rect 20076 21344 20128 21350
rect 20076 21286 20128 21292
rect 19984 20868 20036 20874
rect 19984 20810 20036 20816
rect 19996 18970 20024 20810
rect 20088 19786 20116 21286
rect 20352 20936 20404 20942
rect 20352 20878 20404 20884
rect 20076 19780 20128 19786
rect 20076 19722 20128 19728
rect 19984 18964 20036 18970
rect 19984 18906 20036 18912
rect 20364 18766 20392 20878
rect 20444 19916 20496 19922
rect 20444 19858 20496 19864
rect 20456 19514 20484 19858
rect 20444 19508 20496 19514
rect 20444 19450 20496 19456
rect 20352 18760 20404 18766
rect 20352 18702 20404 18708
rect 20260 18692 20312 18698
rect 20260 18634 20312 18640
rect 20272 18426 20300 18634
rect 19800 18420 19852 18426
rect 19800 18362 19852 18368
rect 20260 18420 20312 18426
rect 20260 18362 20312 18368
rect 19432 18352 19484 18358
rect 19432 18294 19484 18300
rect 19444 17746 19472 18294
rect 19432 17740 19484 17746
rect 19432 17682 19484 17688
rect 19340 17604 19392 17610
rect 19340 17546 19392 17552
rect 19352 17338 19380 17546
rect 19444 17338 19472 17682
rect 19340 17332 19392 17338
rect 19340 17274 19392 17280
rect 19432 17332 19484 17338
rect 19432 17274 19484 17280
rect 19432 17196 19484 17202
rect 19432 17138 19484 17144
rect 19444 16658 19472 17138
rect 19432 16652 19484 16658
rect 19432 16594 19484 16600
rect 20548 15978 20576 21830
rect 20824 20602 20852 21898
rect 20916 20942 20944 22066
rect 21008 21962 21036 22578
rect 21088 22092 21140 22098
rect 21088 22034 21140 22040
rect 20996 21956 21048 21962
rect 20996 21898 21048 21904
rect 20994 21584 21050 21593
rect 20994 21519 20996 21528
rect 21048 21519 21050 21528
rect 20996 21490 21048 21496
rect 20904 20936 20956 20942
rect 20904 20878 20956 20884
rect 20812 20596 20864 20602
rect 20812 20538 20864 20544
rect 20812 20460 20864 20466
rect 20812 20402 20864 20408
rect 20720 19848 20772 19854
rect 20720 19790 20772 19796
rect 20628 19372 20680 19378
rect 20732 19360 20760 19790
rect 20824 19378 20852 20402
rect 21100 20058 21128 22034
rect 21192 22030 21220 24006
rect 21180 22024 21232 22030
rect 21180 21966 21232 21972
rect 21180 21888 21232 21894
rect 21180 21830 21232 21836
rect 21192 21690 21220 21830
rect 21180 21684 21232 21690
rect 21180 21626 21232 21632
rect 21192 21554 21220 21626
rect 21180 21548 21232 21554
rect 21180 21490 21232 21496
rect 21088 20052 21140 20058
rect 21088 19994 21140 20000
rect 21088 19848 21140 19854
rect 21088 19790 21140 19796
rect 20680 19332 20760 19360
rect 20812 19372 20864 19378
rect 20628 19314 20680 19320
rect 20812 19314 20864 19320
rect 20720 19168 20772 19174
rect 20720 19110 20772 19116
rect 20628 17196 20680 17202
rect 20628 17138 20680 17144
rect 20640 16794 20668 17138
rect 20628 16788 20680 16794
rect 20628 16730 20680 16736
rect 20732 16726 20760 19110
rect 20824 18970 20852 19314
rect 20812 18964 20864 18970
rect 20812 18906 20864 18912
rect 21100 18698 21128 19790
rect 21284 19242 21312 24228
rect 21732 24200 21784 24206
rect 21928 24154 21956 24754
rect 22376 24744 22428 24750
rect 22480 24732 22508 25298
rect 22560 24880 22612 24886
rect 22664 24868 22692 26302
rect 22612 24840 22692 24868
rect 22560 24822 22612 24828
rect 22428 24704 22508 24732
rect 22376 24686 22428 24692
rect 22052 24508 22360 24517
rect 22052 24506 22058 24508
rect 22114 24506 22138 24508
rect 22194 24506 22218 24508
rect 22274 24506 22298 24508
rect 22354 24506 22360 24508
rect 22114 24454 22116 24506
rect 22296 24454 22298 24506
rect 22052 24452 22058 24454
rect 22114 24452 22138 24454
rect 22194 24452 22218 24454
rect 22274 24452 22298 24454
rect 22354 24452 22360 24454
rect 22052 24443 22360 24452
rect 22480 24410 22508 24704
rect 22376 24404 22428 24410
rect 22376 24346 22428 24352
rect 22468 24404 22520 24410
rect 22468 24346 22520 24352
rect 22282 24304 22338 24313
rect 22282 24239 22338 24248
rect 22296 24206 22324 24239
rect 21784 24148 21956 24154
rect 21732 24142 21956 24148
rect 22284 24200 22336 24206
rect 22284 24142 22336 24148
rect 21744 24126 21956 24142
rect 21928 23322 21956 24126
rect 22192 24064 22244 24070
rect 22192 24006 22244 24012
rect 22284 24064 22336 24070
rect 22284 24006 22336 24012
rect 22204 23866 22232 24006
rect 22192 23860 22244 23866
rect 22192 23802 22244 23808
rect 22296 23798 22324 24006
rect 22388 23866 22416 24346
rect 22664 24290 22692 24840
rect 22756 24818 22784 28630
rect 22928 28416 22980 28422
rect 22928 28358 22980 28364
rect 22836 27872 22888 27878
rect 22836 27814 22888 27820
rect 22848 27674 22876 27814
rect 22940 27674 22968 28358
rect 22836 27668 22888 27674
rect 22836 27610 22888 27616
rect 22928 27668 22980 27674
rect 22928 27610 22980 27616
rect 23032 27554 23060 28886
rect 23216 28626 23244 29038
rect 23388 28960 23440 28966
rect 23388 28902 23440 28908
rect 23480 28960 23532 28966
rect 23480 28902 23532 28908
rect 23204 28620 23256 28626
rect 23204 28562 23256 28568
rect 23112 28484 23164 28490
rect 23112 28426 23164 28432
rect 22940 27526 23060 27554
rect 22836 27328 22888 27334
rect 22836 27270 22888 27276
rect 22848 25362 22876 27270
rect 22836 25356 22888 25362
rect 22836 25298 22888 25304
rect 22940 25242 22968 27526
rect 23020 27056 23072 27062
rect 23020 26998 23072 27004
rect 23032 26926 23060 26998
rect 23020 26920 23072 26926
rect 23020 26862 23072 26868
rect 23020 26240 23072 26246
rect 23020 26182 23072 26188
rect 23032 25974 23060 26182
rect 23020 25968 23072 25974
rect 23020 25910 23072 25916
rect 22848 25214 22968 25242
rect 23020 25288 23072 25294
rect 23020 25230 23072 25236
rect 22744 24812 22796 24818
rect 22744 24754 22796 24760
rect 22468 24268 22520 24274
rect 22664 24262 22784 24290
rect 22468 24210 22520 24216
rect 22376 23860 22428 23866
rect 22376 23802 22428 23808
rect 22284 23792 22336 23798
rect 22284 23734 22336 23740
rect 22480 23730 22508 24210
rect 22560 24132 22612 24138
rect 22560 24074 22612 24080
rect 22652 24132 22704 24138
rect 22652 24074 22704 24080
rect 22468 23724 22520 23730
rect 22468 23666 22520 23672
rect 22376 23520 22428 23526
rect 22428 23468 22508 23474
rect 22376 23462 22508 23468
rect 22388 23446 22508 23462
rect 22052 23420 22360 23429
rect 22052 23418 22058 23420
rect 22114 23418 22138 23420
rect 22194 23418 22218 23420
rect 22274 23418 22298 23420
rect 22354 23418 22360 23420
rect 22114 23366 22116 23418
rect 22296 23366 22298 23418
rect 22052 23364 22058 23366
rect 22114 23364 22138 23366
rect 22194 23364 22218 23366
rect 22274 23364 22298 23366
rect 22354 23364 22360 23366
rect 22052 23355 22360 23364
rect 21916 23316 21968 23322
rect 21916 23258 21968 23264
rect 21928 22574 21956 23258
rect 22376 23248 22428 23254
rect 22376 23190 22428 23196
rect 21916 22568 21968 22574
rect 21916 22510 21968 22516
rect 21824 22228 21876 22234
rect 21824 22170 21876 22176
rect 21364 22024 21416 22030
rect 21364 21966 21416 21972
rect 21456 22024 21508 22030
rect 21456 21966 21508 21972
rect 21376 21554 21404 21966
rect 21468 21690 21496 21966
rect 21732 21888 21784 21894
rect 21732 21830 21784 21836
rect 21456 21684 21508 21690
rect 21456 21626 21508 21632
rect 21548 21616 21600 21622
rect 21548 21558 21600 21564
rect 21364 21548 21416 21554
rect 21364 21490 21416 21496
rect 21456 21480 21508 21486
rect 21362 21448 21418 21457
rect 21456 21422 21508 21428
rect 21362 21383 21418 21392
rect 21376 20262 21404 21383
rect 21468 20942 21496 21422
rect 21456 20936 21508 20942
rect 21456 20878 21508 20884
rect 21364 20256 21416 20262
rect 21364 20198 21416 20204
rect 21376 19990 21404 20198
rect 21364 19984 21416 19990
rect 21364 19926 21416 19932
rect 21560 19854 21588 21558
rect 21744 20942 21772 21830
rect 21732 20936 21784 20942
rect 21732 20878 21784 20884
rect 21640 20596 21692 20602
rect 21640 20538 21692 20544
rect 21652 20330 21680 20538
rect 21640 20324 21692 20330
rect 21640 20266 21692 20272
rect 21652 19922 21680 20266
rect 21640 19916 21692 19922
rect 21640 19858 21692 19864
rect 21456 19848 21508 19854
rect 21456 19790 21508 19796
rect 21548 19848 21600 19854
rect 21548 19790 21600 19796
rect 21468 19514 21496 19790
rect 21456 19508 21508 19514
rect 21456 19450 21508 19456
rect 21272 19236 21324 19242
rect 21272 19178 21324 19184
rect 21180 18896 21232 18902
rect 21180 18838 21232 18844
rect 21088 18692 21140 18698
rect 21088 18634 21140 18640
rect 21192 18358 21220 18838
rect 21284 18630 21312 19178
rect 21364 18964 21416 18970
rect 21364 18906 21416 18912
rect 21272 18624 21324 18630
rect 21272 18566 21324 18572
rect 21180 18352 21232 18358
rect 21180 18294 21232 18300
rect 21284 18222 21312 18566
rect 21376 18426 21404 18906
rect 21456 18692 21508 18698
rect 21456 18634 21508 18640
rect 21364 18420 21416 18426
rect 21364 18362 21416 18368
rect 20812 18216 20864 18222
rect 20812 18158 20864 18164
rect 21272 18216 21324 18222
rect 21272 18158 21324 18164
rect 20824 17882 20852 18158
rect 20812 17876 20864 17882
rect 20812 17818 20864 17824
rect 20824 17270 20852 17818
rect 21468 17338 21496 18634
rect 21640 18624 21692 18630
rect 21640 18566 21692 18572
rect 21652 18290 21680 18566
rect 21640 18284 21692 18290
rect 21640 18226 21692 18232
rect 21548 18216 21600 18222
rect 21548 18158 21600 18164
rect 21560 17678 21588 18158
rect 21548 17672 21600 17678
rect 21548 17614 21600 17620
rect 21456 17332 21508 17338
rect 21456 17274 21508 17280
rect 21560 17270 21588 17614
rect 21640 17604 21692 17610
rect 21640 17546 21692 17552
rect 20812 17264 20864 17270
rect 20812 17206 20864 17212
rect 21548 17264 21600 17270
rect 21548 17206 21600 17212
rect 21652 16794 21680 17546
rect 21640 16788 21692 16794
rect 21640 16730 21692 16736
rect 20720 16720 20772 16726
rect 20720 16662 20772 16668
rect 21744 16454 21772 20878
rect 21836 19310 21864 22170
rect 21928 20466 21956 22510
rect 22052 22332 22360 22341
rect 22052 22330 22058 22332
rect 22114 22330 22138 22332
rect 22194 22330 22218 22332
rect 22274 22330 22298 22332
rect 22354 22330 22360 22332
rect 22114 22278 22116 22330
rect 22296 22278 22298 22330
rect 22052 22276 22058 22278
rect 22114 22276 22138 22278
rect 22194 22276 22218 22278
rect 22274 22276 22298 22278
rect 22354 22276 22360 22278
rect 22052 22267 22360 22276
rect 22008 22092 22060 22098
rect 22008 22034 22060 22040
rect 22020 21536 22048 22034
rect 22388 21894 22416 23190
rect 22480 21962 22508 23446
rect 22572 23254 22600 24074
rect 22664 23866 22692 24074
rect 22756 24070 22784 24262
rect 22744 24064 22796 24070
rect 22744 24006 22796 24012
rect 22652 23860 22704 23866
rect 22652 23802 22704 23808
rect 22664 23662 22692 23802
rect 22652 23656 22704 23662
rect 22652 23598 22704 23604
rect 22848 23497 22876 25214
rect 22928 25152 22980 25158
rect 22928 25094 22980 25100
rect 22940 24410 22968 25094
rect 23032 24954 23060 25230
rect 23020 24948 23072 24954
rect 23020 24890 23072 24896
rect 23124 24410 23152 28426
rect 23216 28150 23244 28562
rect 23296 28212 23348 28218
rect 23296 28154 23348 28160
rect 23204 28144 23256 28150
rect 23204 28086 23256 28092
rect 23308 27470 23336 28154
rect 23400 28014 23428 28902
rect 23492 28529 23520 28902
rect 23478 28520 23534 28529
rect 23478 28455 23534 28464
rect 23480 28416 23532 28422
rect 23480 28358 23532 28364
rect 23388 28008 23440 28014
rect 23388 27950 23440 27956
rect 23296 27464 23348 27470
rect 23296 27406 23348 27412
rect 23204 27396 23256 27402
rect 23204 27338 23256 27344
rect 23216 26382 23244 27338
rect 23308 27062 23336 27406
rect 23296 27056 23348 27062
rect 23296 26998 23348 27004
rect 23308 26874 23336 26998
rect 23308 26846 23428 26874
rect 23400 26790 23428 26846
rect 23388 26784 23440 26790
rect 23388 26726 23440 26732
rect 23492 26382 23520 28358
rect 23584 28218 23612 29242
rect 23572 28212 23624 28218
rect 23572 28154 23624 28160
rect 23584 27962 23612 28154
rect 23584 27934 23704 27962
rect 23572 27872 23624 27878
rect 23572 27814 23624 27820
rect 23584 26994 23612 27814
rect 23676 27282 23704 27934
rect 23768 27418 23796 31078
rect 23860 30666 23888 31146
rect 23952 30666 23980 31640
rect 24044 30734 24072 32166
rect 24136 31793 24164 32778
rect 24216 31884 24268 31890
rect 24216 31826 24268 31832
rect 24122 31784 24178 31793
rect 24122 31719 24178 31728
rect 24032 30728 24084 30734
rect 24032 30670 24084 30676
rect 23848 30660 23900 30666
rect 23848 30602 23900 30608
rect 23940 30660 23992 30666
rect 23940 30602 23992 30608
rect 23848 30184 23900 30190
rect 23848 30126 23900 30132
rect 23860 29510 23888 30126
rect 23848 29504 23900 29510
rect 23848 29446 23900 29452
rect 23860 27538 23888 29446
rect 24136 29322 24164 31719
rect 23952 29294 24164 29322
rect 23848 27532 23900 27538
rect 23848 27474 23900 27480
rect 23768 27390 23888 27418
rect 23756 27328 23808 27334
rect 23676 27276 23756 27282
rect 23676 27270 23808 27276
rect 23676 27254 23796 27270
rect 23572 26988 23624 26994
rect 23572 26930 23624 26936
rect 23768 26926 23796 27254
rect 23756 26920 23808 26926
rect 23756 26862 23808 26868
rect 23860 26450 23888 27390
rect 23848 26444 23900 26450
rect 23848 26386 23900 26392
rect 23204 26376 23256 26382
rect 23480 26376 23532 26382
rect 23204 26318 23256 26324
rect 23386 26344 23442 26353
rect 23296 26308 23348 26314
rect 23480 26318 23532 26324
rect 23386 26279 23388 26288
rect 23296 26250 23348 26256
rect 23440 26279 23442 26288
rect 23388 26250 23440 26256
rect 23308 25498 23336 26250
rect 23860 25974 23888 26386
rect 23848 25968 23900 25974
rect 23848 25910 23900 25916
rect 23296 25492 23348 25498
rect 23296 25434 23348 25440
rect 23388 25288 23440 25294
rect 23388 25230 23440 25236
rect 23296 25220 23348 25226
rect 23296 25162 23348 25168
rect 23204 24948 23256 24954
rect 23204 24890 23256 24896
rect 22928 24404 22980 24410
rect 22928 24346 22980 24352
rect 23112 24404 23164 24410
rect 23112 24346 23164 24352
rect 22940 24290 22968 24346
rect 22940 24274 23152 24290
rect 22940 24268 23164 24274
rect 22940 24262 23112 24268
rect 23112 24210 23164 24216
rect 23216 24138 23244 24890
rect 23204 24132 23256 24138
rect 23204 24074 23256 24080
rect 23308 23866 23336 25162
rect 23296 23860 23348 23866
rect 23296 23802 23348 23808
rect 23400 23798 23428 25230
rect 23572 25152 23624 25158
rect 23572 25094 23624 25100
rect 23388 23792 23440 23798
rect 23388 23734 23440 23740
rect 23020 23520 23072 23526
rect 22834 23488 22890 23497
rect 23020 23462 23072 23468
rect 22834 23423 22890 23432
rect 22560 23248 22612 23254
rect 22560 23190 22612 23196
rect 22744 22976 22796 22982
rect 22744 22918 22796 22924
rect 22756 22030 22784 22918
rect 23032 22642 23060 23462
rect 23204 23112 23256 23118
rect 23204 23054 23256 23060
rect 23020 22636 23072 22642
rect 23020 22578 23072 22584
rect 23112 22160 23164 22166
rect 23112 22102 23164 22108
rect 22744 22024 22796 22030
rect 22744 21966 22796 21972
rect 22836 22024 22888 22030
rect 22836 21966 22888 21972
rect 22468 21956 22520 21962
rect 22468 21898 22520 21904
rect 22560 21956 22612 21962
rect 22560 21898 22612 21904
rect 22192 21888 22244 21894
rect 22192 21830 22244 21836
rect 22376 21888 22428 21894
rect 22376 21830 22428 21836
rect 22100 21548 22152 21554
rect 22020 21508 22100 21536
rect 22100 21490 22152 21496
rect 22006 21448 22062 21457
rect 22204 21400 22232 21830
rect 22062 21392 22232 21400
rect 22006 21383 22232 21392
rect 22020 21372 22232 21383
rect 22468 21412 22520 21418
rect 22468 21354 22520 21360
rect 22052 21244 22360 21253
rect 22052 21242 22058 21244
rect 22114 21242 22138 21244
rect 22194 21242 22218 21244
rect 22274 21242 22298 21244
rect 22354 21242 22360 21244
rect 22114 21190 22116 21242
rect 22296 21190 22298 21242
rect 22052 21188 22058 21190
rect 22114 21188 22138 21190
rect 22194 21188 22218 21190
rect 22274 21188 22298 21190
rect 22354 21188 22360 21190
rect 22052 21179 22360 21188
rect 22098 20904 22154 20913
rect 22098 20839 22100 20848
rect 22152 20839 22154 20848
rect 22100 20810 22152 20816
rect 22376 20528 22428 20534
rect 22376 20470 22428 20476
rect 21916 20460 21968 20466
rect 21916 20402 21968 20408
rect 22052 20156 22360 20165
rect 22052 20154 22058 20156
rect 22114 20154 22138 20156
rect 22194 20154 22218 20156
rect 22274 20154 22298 20156
rect 22354 20154 22360 20156
rect 22114 20102 22116 20154
rect 22296 20102 22298 20154
rect 22052 20100 22058 20102
rect 22114 20100 22138 20102
rect 22194 20100 22218 20102
rect 22274 20100 22298 20102
rect 22354 20100 22360 20102
rect 22052 20091 22360 20100
rect 22388 19990 22416 20470
rect 22376 19984 22428 19990
rect 22376 19926 22428 19932
rect 21916 19848 21968 19854
rect 21916 19790 21968 19796
rect 21824 19304 21876 19310
rect 21824 19246 21876 19252
rect 21928 18222 21956 19790
rect 22480 19514 22508 21354
rect 22572 20058 22600 21898
rect 22652 21140 22704 21146
rect 22652 21082 22704 21088
rect 22560 20052 22612 20058
rect 22560 19994 22612 20000
rect 22468 19508 22520 19514
rect 22468 19450 22520 19456
rect 22376 19372 22428 19378
rect 22376 19314 22428 19320
rect 22052 19068 22360 19077
rect 22052 19066 22058 19068
rect 22114 19066 22138 19068
rect 22194 19066 22218 19068
rect 22274 19066 22298 19068
rect 22354 19066 22360 19068
rect 22114 19014 22116 19066
rect 22296 19014 22298 19066
rect 22052 19012 22058 19014
rect 22114 19012 22138 19014
rect 22194 19012 22218 19014
rect 22274 19012 22298 19014
rect 22354 19012 22360 19014
rect 22052 19003 22360 19012
rect 22388 18698 22416 19314
rect 22664 19174 22692 21082
rect 22848 20534 22876 21966
rect 23020 21956 23072 21962
rect 23020 21898 23072 21904
rect 23032 20602 23060 21898
rect 23020 20596 23072 20602
rect 23020 20538 23072 20544
rect 22836 20528 22888 20534
rect 22836 20470 22888 20476
rect 22744 20460 22796 20466
rect 22744 20402 22796 20408
rect 22652 19168 22704 19174
rect 22652 19110 22704 19116
rect 22664 18970 22692 19110
rect 22560 18964 22612 18970
rect 22560 18906 22612 18912
rect 22652 18964 22704 18970
rect 22652 18906 22704 18912
rect 22376 18692 22428 18698
rect 22376 18634 22428 18640
rect 21916 18216 21968 18222
rect 21916 18158 21968 18164
rect 22388 18086 22416 18634
rect 22468 18624 22520 18630
rect 22468 18566 22520 18572
rect 22376 18080 22428 18086
rect 22376 18022 22428 18028
rect 22052 17980 22360 17989
rect 22052 17978 22058 17980
rect 22114 17978 22138 17980
rect 22194 17978 22218 17980
rect 22274 17978 22298 17980
rect 22354 17978 22360 17980
rect 22114 17926 22116 17978
rect 22296 17926 22298 17978
rect 22052 17924 22058 17926
rect 22114 17924 22138 17926
rect 22194 17924 22218 17926
rect 22274 17924 22298 17926
rect 22354 17924 22360 17926
rect 22052 17915 22360 17924
rect 22100 17196 22152 17202
rect 22100 17138 22152 17144
rect 21824 16992 21876 16998
rect 22112 16980 22140 17138
rect 22388 17082 22416 18022
rect 22480 17202 22508 18566
rect 22572 17542 22600 18906
rect 22560 17536 22612 17542
rect 22560 17478 22612 17484
rect 22468 17196 22520 17202
rect 22468 17138 22520 17144
rect 22572 17134 22600 17478
rect 22560 17128 22612 17134
rect 22388 17054 22508 17082
rect 22560 17070 22612 17076
rect 21824 16934 21876 16940
rect 21928 16952 22140 16980
rect 22376 16992 22428 16998
rect 21836 16590 21864 16934
rect 21824 16584 21876 16590
rect 21824 16526 21876 16532
rect 21928 16522 21956 16952
rect 22376 16934 22428 16940
rect 22052 16892 22360 16901
rect 22052 16890 22058 16892
rect 22114 16890 22138 16892
rect 22194 16890 22218 16892
rect 22274 16890 22298 16892
rect 22354 16890 22360 16892
rect 22114 16838 22116 16890
rect 22296 16838 22298 16890
rect 22052 16836 22058 16838
rect 22114 16836 22138 16838
rect 22194 16836 22218 16838
rect 22274 16836 22298 16838
rect 22354 16836 22360 16838
rect 22052 16827 22360 16836
rect 22388 16794 22416 16934
rect 22376 16788 22428 16794
rect 22376 16730 22428 16736
rect 22376 16652 22428 16658
rect 22376 16594 22428 16600
rect 21916 16516 21968 16522
rect 21916 16458 21968 16464
rect 22192 16516 22244 16522
rect 22192 16458 22244 16464
rect 21732 16448 21784 16454
rect 21732 16390 21784 16396
rect 22100 16108 22152 16114
rect 22100 16050 22152 16056
rect 20536 15972 20588 15978
rect 20536 15914 20588 15920
rect 22112 15910 22140 16050
rect 22204 16046 22232 16458
rect 22388 16250 22416 16594
rect 22480 16590 22508 17054
rect 22468 16584 22520 16590
rect 22468 16526 22520 16532
rect 22376 16244 22428 16250
rect 22376 16186 22428 16192
rect 22192 16040 22244 16046
rect 22192 15982 22244 15988
rect 22572 15910 22600 17070
rect 22652 16720 22704 16726
rect 22652 16662 22704 16668
rect 22664 16046 22692 16662
rect 22756 16250 22784 20402
rect 23020 20324 23072 20330
rect 23020 20266 23072 20272
rect 22928 19780 22980 19786
rect 22928 19722 22980 19728
rect 22940 19514 22968 19722
rect 23032 19718 23060 20266
rect 23124 20262 23152 22102
rect 23216 21690 23244 23054
rect 23400 22438 23428 23734
rect 23480 23112 23532 23118
rect 23480 23054 23532 23060
rect 23492 22778 23520 23054
rect 23480 22772 23532 22778
rect 23480 22714 23532 22720
rect 23480 22568 23532 22574
rect 23480 22510 23532 22516
rect 23388 22432 23440 22438
rect 23388 22374 23440 22380
rect 23296 21888 23348 21894
rect 23296 21830 23348 21836
rect 23204 21684 23256 21690
rect 23204 21626 23256 21632
rect 23308 21593 23336 21830
rect 23294 21584 23350 21593
rect 23294 21519 23350 21528
rect 23492 21486 23520 22510
rect 23584 22098 23612 25094
rect 23848 24608 23900 24614
rect 23848 24550 23900 24556
rect 23860 23866 23888 24550
rect 23952 24290 23980 29294
rect 24124 29232 24176 29238
rect 24124 29174 24176 29180
rect 24032 28552 24084 28558
rect 24032 28494 24084 28500
rect 24044 24410 24072 28494
rect 24136 28082 24164 29174
rect 24228 28121 24256 31826
rect 24412 31754 24440 34546
rect 24596 33998 24624 34682
rect 24688 33998 24716 35974
rect 24780 34105 24808 37062
rect 25136 36780 25188 36786
rect 25136 36722 25188 36728
rect 24860 36576 24912 36582
rect 24860 36518 24912 36524
rect 24872 35086 24900 36518
rect 24950 36272 25006 36281
rect 24950 36207 25006 36216
rect 24860 35080 24912 35086
rect 24860 35022 24912 35028
rect 24860 34944 24912 34950
rect 24860 34886 24912 34892
rect 24766 34096 24822 34105
rect 24766 34031 24822 34040
rect 24584 33992 24636 33998
rect 24584 33934 24636 33940
rect 24676 33992 24728 33998
rect 24676 33934 24728 33940
rect 24492 33448 24544 33454
rect 24596 33436 24624 33934
rect 24544 33408 24624 33436
rect 24492 33390 24544 33396
rect 24596 32337 24624 33408
rect 24582 32328 24638 32337
rect 24582 32263 24638 32272
rect 24492 32020 24544 32026
rect 24492 31962 24544 31968
rect 24400 31748 24452 31754
rect 24400 31690 24452 31696
rect 24412 31210 24440 31690
rect 24400 31204 24452 31210
rect 24400 31146 24452 31152
rect 24504 30802 24532 31962
rect 24596 31278 24624 32263
rect 24676 32224 24728 32230
rect 24676 32166 24728 32172
rect 24688 31890 24716 32166
rect 24676 31884 24728 31890
rect 24676 31826 24728 31832
rect 24872 31414 24900 34886
rect 24964 32910 24992 36207
rect 25148 35834 25176 36722
rect 25240 36310 25268 39578
rect 25792 38486 25820 41200
rect 26056 39432 26108 39438
rect 26056 39374 26108 39380
rect 25780 38480 25832 38486
rect 25780 38422 25832 38428
rect 26068 38418 26096 39374
rect 26272 39196 26580 39205
rect 26272 39194 26278 39196
rect 26334 39194 26358 39196
rect 26414 39194 26438 39196
rect 26494 39194 26518 39196
rect 26574 39194 26580 39196
rect 26334 39142 26336 39194
rect 26516 39142 26518 39194
rect 26272 39140 26278 39142
rect 26334 39140 26358 39142
rect 26414 39140 26438 39142
rect 26494 39140 26518 39142
rect 26574 39140 26580 39142
rect 26272 39131 26580 39140
rect 26976 39024 27028 39030
rect 26976 38966 27028 38972
rect 26988 38758 27016 38966
rect 27080 38758 27108 41200
rect 28264 39364 28316 39370
rect 28264 39306 28316 39312
rect 28276 39030 28304 39306
rect 28264 39024 28316 39030
rect 27618 38992 27674 39001
rect 28264 38966 28316 38972
rect 27618 38927 27674 38936
rect 27344 38888 27396 38894
rect 27344 38830 27396 38836
rect 26976 38752 27028 38758
rect 26976 38694 27028 38700
rect 27068 38752 27120 38758
rect 27068 38694 27120 38700
rect 26424 38480 26476 38486
rect 26424 38422 26476 38428
rect 26056 38412 26108 38418
rect 26056 38354 26108 38360
rect 26436 38321 26464 38422
rect 26422 38312 26478 38321
rect 26422 38247 26478 38256
rect 26272 38108 26580 38117
rect 26272 38106 26278 38108
rect 26334 38106 26358 38108
rect 26414 38106 26438 38108
rect 26494 38106 26518 38108
rect 26574 38106 26580 38108
rect 26334 38054 26336 38106
rect 26516 38054 26518 38106
rect 26272 38052 26278 38054
rect 26334 38052 26358 38054
rect 26414 38052 26438 38054
rect 26494 38052 26518 38054
rect 26574 38052 26580 38054
rect 26272 38043 26580 38052
rect 25320 37936 25372 37942
rect 25318 37904 25320 37913
rect 25372 37904 25374 37913
rect 25318 37839 25374 37848
rect 25320 37800 25372 37806
rect 25320 37742 25372 37748
rect 25332 37262 25360 37742
rect 25780 37664 25832 37670
rect 25780 37606 25832 37612
rect 25964 37664 26016 37670
rect 25964 37606 26016 37612
rect 25792 37466 25820 37606
rect 25688 37460 25740 37466
rect 25688 37402 25740 37408
rect 25780 37460 25832 37466
rect 25780 37402 25832 37408
rect 25700 37369 25728 37402
rect 25686 37360 25742 37369
rect 25686 37295 25742 37304
rect 25320 37256 25372 37262
rect 25320 37198 25372 37204
rect 25412 37120 25464 37126
rect 25412 37062 25464 37068
rect 25320 36712 25372 36718
rect 25320 36654 25372 36660
rect 25332 36310 25360 36654
rect 25228 36304 25280 36310
rect 25228 36246 25280 36252
rect 25320 36304 25372 36310
rect 25320 36246 25372 36252
rect 25318 36136 25374 36145
rect 25318 36071 25374 36080
rect 25136 35828 25188 35834
rect 25136 35770 25188 35776
rect 25228 35692 25280 35698
rect 25228 35634 25280 35640
rect 25136 35624 25188 35630
rect 25136 35566 25188 35572
rect 25044 34468 25096 34474
rect 25044 34410 25096 34416
rect 25056 33930 25084 34410
rect 25044 33924 25096 33930
rect 25044 33866 25096 33872
rect 24952 32904 25004 32910
rect 24952 32846 25004 32852
rect 24952 32496 25004 32502
rect 25148 32473 25176 35566
rect 25240 32502 25268 35634
rect 25228 32496 25280 32502
rect 24952 32438 25004 32444
rect 25134 32464 25190 32473
rect 24860 31408 24912 31414
rect 24860 31350 24912 31356
rect 24584 31272 24636 31278
rect 24584 31214 24636 31220
rect 24492 30796 24544 30802
rect 24492 30738 24544 30744
rect 24596 30258 24624 31214
rect 24768 31136 24820 31142
rect 24768 31078 24820 31084
rect 24676 30728 24728 30734
rect 24676 30670 24728 30676
rect 24584 30252 24636 30258
rect 24584 30194 24636 30200
rect 24688 29306 24716 30670
rect 24780 29646 24808 31078
rect 24860 30388 24912 30394
rect 24860 30330 24912 30336
rect 24872 30258 24900 30330
rect 24860 30252 24912 30258
rect 24860 30194 24912 30200
rect 24860 29708 24912 29714
rect 24860 29650 24912 29656
rect 24768 29640 24820 29646
rect 24768 29582 24820 29588
rect 24676 29300 24728 29306
rect 24676 29242 24728 29248
rect 24872 28558 24900 29650
rect 24964 29646 24992 32438
rect 25228 32438 25280 32444
rect 25134 32399 25190 32408
rect 25148 31929 25176 32399
rect 25134 31920 25190 31929
rect 25134 31855 25190 31864
rect 25044 31680 25096 31686
rect 25044 31622 25096 31628
rect 25056 29714 25084 31622
rect 25136 31476 25188 31482
rect 25136 31418 25188 31424
rect 25148 30938 25176 31418
rect 25136 30932 25188 30938
rect 25136 30874 25188 30880
rect 25332 30326 25360 36071
rect 25424 34746 25452 37062
rect 25872 36780 25924 36786
rect 25872 36722 25924 36728
rect 25688 36576 25740 36582
rect 25688 36518 25740 36524
rect 25504 35488 25556 35494
rect 25504 35430 25556 35436
rect 25412 34740 25464 34746
rect 25412 34682 25464 34688
rect 25516 32881 25544 35430
rect 25700 33590 25728 36518
rect 25780 36168 25832 36174
rect 25780 36110 25832 36116
rect 25792 35766 25820 36110
rect 25780 35760 25832 35766
rect 25780 35702 25832 35708
rect 25792 34932 25820 35702
rect 25884 35290 25912 36722
rect 25872 35284 25924 35290
rect 25872 35226 25924 35232
rect 25872 34944 25924 34950
rect 25792 34904 25872 34932
rect 25872 34886 25924 34892
rect 25780 34604 25832 34610
rect 25780 34546 25832 34552
rect 25792 33590 25820 34546
rect 25688 33584 25740 33590
rect 25688 33526 25740 33532
rect 25780 33584 25832 33590
rect 25780 33526 25832 33532
rect 25502 32872 25558 32881
rect 25412 32836 25464 32842
rect 25502 32807 25558 32816
rect 25596 32836 25648 32842
rect 25412 32778 25464 32784
rect 25596 32778 25648 32784
rect 25320 30320 25372 30326
rect 25320 30262 25372 30268
rect 25044 29708 25096 29714
rect 25044 29650 25096 29656
rect 24952 29640 25004 29646
rect 24952 29582 25004 29588
rect 24584 28552 24636 28558
rect 24584 28494 24636 28500
rect 24860 28552 24912 28558
rect 24860 28494 24912 28500
rect 24400 28484 24452 28490
rect 24400 28426 24452 28432
rect 24214 28112 24270 28121
rect 24124 28076 24176 28082
rect 24214 28047 24270 28056
rect 24124 28018 24176 28024
rect 24124 27532 24176 27538
rect 24124 27474 24176 27480
rect 24136 26790 24164 27474
rect 24124 26784 24176 26790
rect 24124 26726 24176 26732
rect 24228 25294 24256 28047
rect 24412 26858 24440 28426
rect 24492 28416 24544 28422
rect 24492 28358 24544 28364
rect 24504 27946 24532 28358
rect 24492 27940 24544 27946
rect 24492 27882 24544 27888
rect 24596 26994 24624 28494
rect 24964 27878 24992 29582
rect 25332 29510 25360 30262
rect 25424 29510 25452 32778
rect 25608 32570 25636 32778
rect 25596 32564 25648 32570
rect 25596 32506 25648 32512
rect 25700 32366 25728 33526
rect 25688 32360 25740 32366
rect 25688 32302 25740 32308
rect 25792 32298 25820 33526
rect 25884 32298 25912 34886
rect 25976 33930 26004 37606
rect 26988 37262 27016 38694
rect 27160 37868 27212 37874
rect 27160 37810 27212 37816
rect 27172 37777 27200 37810
rect 27158 37768 27214 37777
rect 27356 37738 27384 38830
rect 27632 38350 27660 38927
rect 28368 38826 28396 41200
rect 28448 39432 28500 39438
rect 28448 39374 28500 39380
rect 28632 39432 28684 39438
rect 28632 39374 28684 39380
rect 28356 38820 28408 38826
rect 28356 38762 28408 38768
rect 28460 38758 28488 39374
rect 28540 39296 28592 39302
rect 28644 39250 28672 39374
rect 28592 39244 28672 39250
rect 28540 39238 28672 39244
rect 28552 39222 28672 39238
rect 28448 38752 28500 38758
rect 28448 38694 28500 38700
rect 27436 38344 27488 38350
rect 27436 38286 27488 38292
rect 27620 38344 27672 38350
rect 27620 38286 27672 38292
rect 27448 37874 27476 38286
rect 28080 38208 28132 38214
rect 28080 38150 28132 38156
rect 28356 38208 28408 38214
rect 28356 38150 28408 38156
rect 27436 37868 27488 37874
rect 27436 37810 27488 37816
rect 27528 37800 27580 37806
rect 27528 37742 27580 37748
rect 27620 37800 27672 37806
rect 27620 37742 27672 37748
rect 27158 37703 27214 37712
rect 27344 37732 27396 37738
rect 27344 37674 27396 37680
rect 26056 37256 26108 37262
rect 26056 37198 26108 37204
rect 26976 37256 27028 37262
rect 26976 37198 27028 37204
rect 26068 36378 26096 37198
rect 26976 37120 27028 37126
rect 26976 37062 27028 37068
rect 27160 37120 27212 37126
rect 27160 37062 27212 37068
rect 26272 37020 26580 37029
rect 26272 37018 26278 37020
rect 26334 37018 26358 37020
rect 26414 37018 26438 37020
rect 26494 37018 26518 37020
rect 26574 37018 26580 37020
rect 26334 36966 26336 37018
rect 26516 36966 26518 37018
rect 26272 36964 26278 36966
rect 26334 36964 26358 36966
rect 26414 36964 26438 36966
rect 26494 36964 26518 36966
rect 26574 36964 26580 36966
rect 26272 36955 26580 36964
rect 26424 36780 26476 36786
rect 26424 36722 26476 36728
rect 26516 36780 26568 36786
rect 26516 36722 26568 36728
rect 26148 36576 26200 36582
rect 26148 36518 26200 36524
rect 26056 36372 26108 36378
rect 26056 36314 26108 36320
rect 26056 35488 26108 35494
rect 26056 35430 26108 35436
rect 25964 33924 26016 33930
rect 25964 33866 26016 33872
rect 26068 33436 26096 35430
rect 25976 33408 26096 33436
rect 25780 32292 25832 32298
rect 25780 32234 25832 32240
rect 25872 32292 25924 32298
rect 25872 32234 25924 32240
rect 25504 32020 25556 32026
rect 25504 31962 25556 31968
rect 25780 32020 25832 32026
rect 25832 31980 25912 32008
rect 25780 31962 25832 31968
rect 25516 31890 25544 31962
rect 25778 31920 25834 31929
rect 25504 31884 25556 31890
rect 25778 31855 25834 31864
rect 25504 31826 25556 31832
rect 25688 31816 25740 31822
rect 25688 31758 25740 31764
rect 25596 30388 25648 30394
rect 25596 30330 25648 30336
rect 25608 29646 25636 30330
rect 25700 30326 25728 31758
rect 25688 30320 25740 30326
rect 25688 30262 25740 30268
rect 25792 30122 25820 31855
rect 25884 31142 25912 31980
rect 25872 31136 25924 31142
rect 25872 31078 25924 31084
rect 25780 30116 25832 30122
rect 25780 30058 25832 30064
rect 25884 29646 25912 31078
rect 25976 29782 26004 33408
rect 26160 33114 26188 36518
rect 26436 36360 26464 36722
rect 26528 36582 26556 36722
rect 26516 36576 26568 36582
rect 26516 36518 26568 36524
rect 26436 36332 26740 36360
rect 26608 36236 26660 36242
rect 26608 36178 26660 36184
rect 26272 35932 26580 35941
rect 26272 35930 26278 35932
rect 26334 35930 26358 35932
rect 26414 35930 26438 35932
rect 26494 35930 26518 35932
rect 26574 35930 26580 35932
rect 26334 35878 26336 35930
rect 26516 35878 26518 35930
rect 26272 35876 26278 35878
rect 26334 35876 26358 35878
rect 26414 35876 26438 35878
rect 26494 35876 26518 35878
rect 26574 35876 26580 35878
rect 26272 35867 26580 35876
rect 26620 35698 26648 36178
rect 26608 35692 26660 35698
rect 26608 35634 26660 35640
rect 26516 35488 26568 35494
rect 26516 35430 26568 35436
rect 26528 35086 26556 35430
rect 26516 35080 26568 35086
rect 26568 35040 26648 35068
rect 26516 35022 26568 35028
rect 26272 34844 26580 34853
rect 26272 34842 26278 34844
rect 26334 34842 26358 34844
rect 26414 34842 26438 34844
rect 26494 34842 26518 34844
rect 26574 34842 26580 34844
rect 26334 34790 26336 34842
rect 26516 34790 26518 34842
rect 26272 34788 26278 34790
rect 26334 34788 26358 34790
rect 26414 34788 26438 34790
rect 26494 34788 26518 34790
rect 26574 34788 26580 34790
rect 26272 34779 26580 34788
rect 26424 34536 26476 34542
rect 26424 34478 26476 34484
rect 26436 34066 26464 34478
rect 26620 34202 26648 35040
rect 26608 34196 26660 34202
rect 26608 34138 26660 34144
rect 26424 34060 26476 34066
rect 26424 34002 26476 34008
rect 26272 33756 26580 33765
rect 26272 33754 26278 33756
rect 26334 33754 26358 33756
rect 26414 33754 26438 33756
rect 26494 33754 26518 33756
rect 26574 33754 26580 33756
rect 26334 33702 26336 33754
rect 26516 33702 26518 33754
rect 26272 33700 26278 33702
rect 26334 33700 26358 33702
rect 26414 33700 26438 33702
rect 26494 33700 26518 33702
rect 26574 33700 26580 33702
rect 26272 33691 26580 33700
rect 26712 33561 26740 36332
rect 26884 36032 26936 36038
rect 26884 35974 26936 35980
rect 26792 35624 26844 35630
rect 26792 35566 26844 35572
rect 26698 33552 26754 33561
rect 26698 33487 26700 33496
rect 26752 33487 26754 33496
rect 26700 33458 26752 33464
rect 26804 33402 26832 35566
rect 26620 33374 26832 33402
rect 26620 33318 26648 33374
rect 26608 33312 26660 33318
rect 26608 33254 26660 33260
rect 26700 33312 26752 33318
rect 26700 33254 26752 33260
rect 26148 33108 26200 33114
rect 26148 33050 26200 33056
rect 26608 32904 26660 32910
rect 26608 32846 26660 32852
rect 26272 32668 26580 32677
rect 26272 32666 26278 32668
rect 26334 32666 26358 32668
rect 26414 32666 26438 32668
rect 26494 32666 26518 32668
rect 26574 32666 26580 32668
rect 26334 32614 26336 32666
rect 26516 32614 26518 32666
rect 26272 32612 26278 32614
rect 26334 32612 26358 32614
rect 26414 32612 26438 32614
rect 26494 32612 26518 32614
rect 26574 32612 26580 32614
rect 26272 32603 26580 32612
rect 26056 32564 26108 32570
rect 26056 32506 26108 32512
rect 26148 32564 26200 32570
rect 26148 32506 26200 32512
rect 26068 32298 26096 32506
rect 26056 32292 26108 32298
rect 26056 32234 26108 32240
rect 26068 30326 26096 32234
rect 26160 32026 26188 32506
rect 26148 32020 26200 32026
rect 26148 31962 26200 31968
rect 26620 31822 26648 32846
rect 26608 31816 26660 31822
rect 26608 31758 26660 31764
rect 26272 31580 26580 31589
rect 26272 31578 26278 31580
rect 26334 31578 26358 31580
rect 26414 31578 26438 31580
rect 26494 31578 26518 31580
rect 26574 31578 26580 31580
rect 26334 31526 26336 31578
rect 26516 31526 26518 31578
rect 26272 31524 26278 31526
rect 26334 31524 26358 31526
rect 26414 31524 26438 31526
rect 26494 31524 26518 31526
rect 26574 31524 26580 31526
rect 26272 31515 26580 31524
rect 26424 31340 26476 31346
rect 26424 31282 26476 31288
rect 26436 30802 26464 31282
rect 26424 30796 26476 30802
rect 26424 30738 26476 30744
rect 26272 30492 26580 30501
rect 26272 30490 26278 30492
rect 26334 30490 26358 30492
rect 26414 30490 26438 30492
rect 26494 30490 26518 30492
rect 26574 30490 26580 30492
rect 26334 30438 26336 30490
rect 26516 30438 26518 30490
rect 26272 30436 26278 30438
rect 26334 30436 26358 30438
rect 26414 30436 26438 30438
rect 26494 30436 26518 30438
rect 26574 30436 26580 30438
rect 26272 30427 26580 30436
rect 26056 30320 26108 30326
rect 26056 30262 26108 30268
rect 26056 30184 26108 30190
rect 26056 30126 26108 30132
rect 25964 29776 26016 29782
rect 25964 29718 26016 29724
rect 25596 29640 25648 29646
rect 25596 29582 25648 29588
rect 25872 29640 25924 29646
rect 25872 29582 25924 29588
rect 25964 29640 26016 29646
rect 25964 29582 26016 29588
rect 25320 29504 25372 29510
rect 25042 29472 25098 29481
rect 25320 29446 25372 29452
rect 25412 29504 25464 29510
rect 25412 29446 25464 29452
rect 25042 29407 25098 29416
rect 25056 28150 25084 29407
rect 25044 28144 25096 28150
rect 25044 28086 25096 28092
rect 25608 27946 25636 29582
rect 25976 29510 26004 29582
rect 25964 29504 26016 29510
rect 25964 29446 26016 29452
rect 25976 28762 26004 29446
rect 25964 28756 26016 28762
rect 25964 28698 26016 28704
rect 25596 27940 25648 27946
rect 25596 27882 25648 27888
rect 24952 27872 25004 27878
rect 24952 27814 25004 27820
rect 25608 27690 25636 27882
rect 25424 27662 25636 27690
rect 25872 27668 25924 27674
rect 24676 27464 24728 27470
rect 24676 27406 24728 27412
rect 24768 27464 24820 27470
rect 24768 27406 24820 27412
rect 24584 26988 24636 26994
rect 24584 26930 24636 26936
rect 24400 26852 24452 26858
rect 24400 26794 24452 26800
rect 24584 26784 24636 26790
rect 24584 26726 24636 26732
rect 24400 26512 24452 26518
rect 24400 26454 24452 26460
rect 24308 25832 24360 25838
rect 24308 25774 24360 25780
rect 24216 25288 24268 25294
rect 24216 25230 24268 25236
rect 24320 24818 24348 25774
rect 24412 25770 24440 26454
rect 24596 25906 24624 26726
rect 24584 25900 24636 25906
rect 24584 25842 24636 25848
rect 24400 25764 24452 25770
rect 24400 25706 24452 25712
rect 24492 25696 24544 25702
rect 24492 25638 24544 25644
rect 24398 24984 24454 24993
rect 24398 24919 24454 24928
rect 24308 24812 24360 24818
rect 24308 24754 24360 24760
rect 24032 24404 24084 24410
rect 24032 24346 24084 24352
rect 23952 24262 24072 24290
rect 23848 23860 23900 23866
rect 23848 23802 23900 23808
rect 23940 22160 23992 22166
rect 23940 22102 23992 22108
rect 23572 22092 23624 22098
rect 23572 22034 23624 22040
rect 23572 21548 23624 21554
rect 23572 21490 23624 21496
rect 23480 21480 23532 21486
rect 23480 21422 23532 21428
rect 23388 21344 23440 21350
rect 23388 21286 23440 21292
rect 23400 20602 23428 21286
rect 23492 20874 23520 21422
rect 23584 21146 23612 21490
rect 23664 21344 23716 21350
rect 23664 21286 23716 21292
rect 23572 21140 23624 21146
rect 23572 21082 23624 21088
rect 23480 20868 23532 20874
rect 23480 20810 23532 20816
rect 23388 20596 23440 20602
rect 23388 20538 23440 20544
rect 23112 20256 23164 20262
rect 23112 20198 23164 20204
rect 23388 20256 23440 20262
rect 23388 20198 23440 20204
rect 23020 19712 23072 19718
rect 23020 19654 23072 19660
rect 22928 19508 22980 19514
rect 22928 19450 22980 19456
rect 23032 19242 23060 19654
rect 23112 19372 23164 19378
rect 23112 19314 23164 19320
rect 23296 19372 23348 19378
rect 23296 19314 23348 19320
rect 23020 19236 23072 19242
rect 23020 19178 23072 19184
rect 22836 18284 22888 18290
rect 22836 18226 22888 18232
rect 22744 16244 22796 16250
rect 22744 16186 22796 16192
rect 22652 16040 22704 16046
rect 22652 15982 22704 15988
rect 22100 15904 22152 15910
rect 22100 15846 22152 15852
rect 22560 15904 22612 15910
rect 22560 15846 22612 15852
rect 22052 15804 22360 15813
rect 22052 15802 22058 15804
rect 22114 15802 22138 15804
rect 22194 15802 22218 15804
rect 22274 15802 22298 15804
rect 22354 15802 22360 15804
rect 22114 15750 22116 15802
rect 22296 15750 22298 15802
rect 22052 15748 22058 15750
rect 22114 15748 22138 15750
rect 22194 15748 22218 15750
rect 22274 15748 22298 15750
rect 22354 15748 22360 15750
rect 22052 15739 22360 15748
rect 22848 15706 22876 18226
rect 23020 16448 23072 16454
rect 23020 16390 23072 16396
rect 22836 15700 22888 15706
rect 22836 15642 22888 15648
rect 23032 15502 23060 16390
rect 23124 15638 23152 19314
rect 23308 19174 23336 19314
rect 23296 19168 23348 19174
rect 23296 19110 23348 19116
rect 23112 15632 23164 15638
rect 23112 15574 23164 15580
rect 23308 15502 23336 19110
rect 23400 16658 23428 20198
rect 23492 19854 23520 20810
rect 23480 19848 23532 19854
rect 23480 19790 23532 19796
rect 23676 19514 23704 21286
rect 23756 20460 23808 20466
rect 23756 20402 23808 20408
rect 23768 19718 23796 20402
rect 23848 19848 23900 19854
rect 23848 19790 23900 19796
rect 23756 19712 23808 19718
rect 23756 19654 23808 19660
rect 23664 19508 23716 19514
rect 23664 19450 23716 19456
rect 23768 19310 23796 19654
rect 23756 19304 23808 19310
rect 23756 19246 23808 19252
rect 23572 18896 23624 18902
rect 23572 18838 23624 18844
rect 23756 18896 23808 18902
rect 23756 18838 23808 18844
rect 23480 17536 23532 17542
rect 23480 17478 23532 17484
rect 23492 17270 23520 17478
rect 23480 17264 23532 17270
rect 23480 17206 23532 17212
rect 23388 16652 23440 16658
rect 23388 16594 23440 16600
rect 23584 16182 23612 18838
rect 23664 17672 23716 17678
rect 23664 17614 23716 17620
rect 23572 16176 23624 16182
rect 23572 16118 23624 16124
rect 23020 15496 23072 15502
rect 23020 15438 23072 15444
rect 23296 15496 23348 15502
rect 23584 15473 23612 16118
rect 23676 15978 23704 17614
rect 23768 16726 23796 18838
rect 23860 18290 23888 19790
rect 23952 19446 23980 22102
rect 24044 22098 24072 24262
rect 24320 23798 24348 24754
rect 24412 24342 24440 24919
rect 24400 24336 24452 24342
rect 24400 24278 24452 24284
rect 24308 23792 24360 23798
rect 24308 23734 24360 23740
rect 24400 23724 24452 23730
rect 24400 23666 24452 23672
rect 24124 22636 24176 22642
rect 24124 22578 24176 22584
rect 24032 22092 24084 22098
rect 24032 22034 24084 22040
rect 24032 21888 24084 21894
rect 24032 21830 24084 21836
rect 23940 19440 23992 19446
rect 23940 19382 23992 19388
rect 23848 18284 23900 18290
rect 23848 18226 23900 18232
rect 23940 18284 23992 18290
rect 23940 18226 23992 18232
rect 23756 16720 23808 16726
rect 23756 16662 23808 16668
rect 23848 16448 23900 16454
rect 23848 16390 23900 16396
rect 23664 15972 23716 15978
rect 23664 15914 23716 15920
rect 23860 15502 23888 16390
rect 23952 15706 23980 18226
rect 24044 16250 24072 21830
rect 24032 16244 24084 16250
rect 24032 16186 24084 16192
rect 24032 16108 24084 16114
rect 24032 16050 24084 16056
rect 23940 15700 23992 15706
rect 23940 15642 23992 15648
rect 24044 15502 24072 16050
rect 24136 15706 24164 22578
rect 24412 22234 24440 23666
rect 24400 22228 24452 22234
rect 24400 22170 24452 22176
rect 24400 22092 24452 22098
rect 24400 22034 24452 22040
rect 24216 21004 24268 21010
rect 24216 20946 24268 20952
rect 24228 20913 24256 20946
rect 24214 20904 24270 20913
rect 24214 20839 24270 20848
rect 24216 19372 24268 19378
rect 24216 19314 24268 19320
rect 24124 15700 24176 15706
rect 24124 15642 24176 15648
rect 24228 15570 24256 19314
rect 24308 16788 24360 16794
rect 24308 16730 24360 16736
rect 24320 16454 24348 16730
rect 24412 16658 24440 22034
rect 24504 21078 24532 25638
rect 24584 25220 24636 25226
rect 24584 25162 24636 25168
rect 24596 24313 24624 25162
rect 24688 24886 24716 27406
rect 24780 26518 24808 27406
rect 24860 27396 24912 27402
rect 24860 27338 24912 27344
rect 24768 26512 24820 26518
rect 24768 26454 24820 26460
rect 24872 26450 24900 27338
rect 25044 26512 25096 26518
rect 25044 26454 25096 26460
rect 24860 26444 24912 26450
rect 24860 26386 24912 26392
rect 24950 25936 25006 25945
rect 24950 25871 25006 25880
rect 24964 25498 24992 25871
rect 24952 25492 25004 25498
rect 24952 25434 25004 25440
rect 25056 25242 25084 26454
rect 25424 26314 25452 27662
rect 25872 27610 25924 27616
rect 25504 27600 25556 27606
rect 25504 27542 25556 27548
rect 25412 26308 25464 26314
rect 25412 26250 25464 26256
rect 25412 25968 25464 25974
rect 25412 25910 25464 25916
rect 24964 25214 25084 25242
rect 25424 25226 25452 25910
rect 25412 25220 25464 25226
rect 24676 24880 24728 24886
rect 24676 24822 24728 24828
rect 24582 24304 24638 24313
rect 24582 24239 24638 24248
rect 24584 22976 24636 22982
rect 24584 22918 24636 22924
rect 24596 22710 24624 22918
rect 24584 22704 24636 22710
rect 24584 22646 24636 22652
rect 24492 21072 24544 21078
rect 24492 21014 24544 21020
rect 24688 20874 24716 24822
rect 24964 24274 24992 25214
rect 25412 25162 25464 25168
rect 25516 24886 25544 27542
rect 25596 27328 25648 27334
rect 25648 27288 25728 27316
rect 25596 27270 25648 27276
rect 25596 26240 25648 26246
rect 25596 26182 25648 26188
rect 25504 24880 25556 24886
rect 25504 24822 25556 24828
rect 24952 24268 25004 24274
rect 24952 24210 25004 24216
rect 25044 24200 25096 24206
rect 25044 24142 25096 24148
rect 25056 23526 25084 24142
rect 25044 23520 25096 23526
rect 25044 23462 25096 23468
rect 25412 23520 25464 23526
rect 25412 23462 25464 23468
rect 24952 23112 25004 23118
rect 24952 23054 25004 23060
rect 24964 22710 24992 23054
rect 24952 22704 25004 22710
rect 24952 22646 25004 22652
rect 25056 22030 25084 23462
rect 25228 23112 25280 23118
rect 25228 23054 25280 23060
rect 25240 22778 25268 23054
rect 25424 23050 25452 23462
rect 25320 23044 25372 23050
rect 25320 22986 25372 22992
rect 25412 23044 25464 23050
rect 25412 22986 25464 22992
rect 25228 22772 25280 22778
rect 25228 22714 25280 22720
rect 25136 22704 25188 22710
rect 25136 22646 25188 22652
rect 24768 22024 24820 22030
rect 24768 21966 24820 21972
rect 25044 22024 25096 22030
rect 25148 22001 25176 22646
rect 25332 22506 25360 22986
rect 25412 22636 25464 22642
rect 25412 22578 25464 22584
rect 25320 22500 25372 22506
rect 25320 22442 25372 22448
rect 25228 22432 25280 22438
rect 25228 22374 25280 22380
rect 25044 21966 25096 21972
rect 25134 21992 25190 22001
rect 24780 21418 24808 21966
rect 25056 21622 25084 21966
rect 25134 21927 25190 21936
rect 25044 21616 25096 21622
rect 25044 21558 25096 21564
rect 24768 21412 24820 21418
rect 24768 21354 24820 21360
rect 25056 20942 25084 21558
rect 25136 21344 25188 21350
rect 25136 21286 25188 21292
rect 25148 21146 25176 21286
rect 25136 21140 25188 21146
rect 25136 21082 25188 21088
rect 25044 20936 25096 20942
rect 25044 20878 25096 20884
rect 24492 20868 24544 20874
rect 24676 20868 24728 20874
rect 24492 20810 24544 20816
rect 24596 20828 24676 20856
rect 24504 20602 24532 20810
rect 24492 20596 24544 20602
rect 24492 20538 24544 20544
rect 24492 19508 24544 19514
rect 24492 19450 24544 19456
rect 24400 16652 24452 16658
rect 24400 16594 24452 16600
rect 24308 16448 24360 16454
rect 24308 16390 24360 16396
rect 24504 16250 24532 19450
rect 24596 18698 24624 20828
rect 24676 20810 24728 20816
rect 25044 20596 25096 20602
rect 25044 20538 25096 20544
rect 24768 19712 24820 19718
rect 24768 19654 24820 19660
rect 24676 18896 24728 18902
rect 24676 18838 24728 18844
rect 24584 18692 24636 18698
rect 24584 18634 24636 18640
rect 24596 18601 24624 18634
rect 24582 18592 24638 18601
rect 24582 18527 24638 18536
rect 24584 18284 24636 18290
rect 24584 18226 24636 18232
rect 24596 16590 24624 18226
rect 24584 16584 24636 16590
rect 24584 16526 24636 16532
rect 24688 16454 24716 18838
rect 24780 16794 24808 19654
rect 25056 19446 25084 20538
rect 24952 19440 25004 19446
rect 24952 19382 25004 19388
rect 25044 19440 25096 19446
rect 25044 19382 25096 19388
rect 24860 19372 24912 19378
rect 24860 19314 24912 19320
rect 24768 16788 24820 16794
rect 24768 16730 24820 16736
rect 24768 16584 24820 16590
rect 24768 16526 24820 16532
rect 24676 16448 24728 16454
rect 24676 16390 24728 16396
rect 24492 16244 24544 16250
rect 24492 16186 24544 16192
rect 24216 15564 24268 15570
rect 24216 15506 24268 15512
rect 23848 15496 23900 15502
rect 23296 15438 23348 15444
rect 23570 15464 23626 15473
rect 23848 15438 23900 15444
rect 24032 15496 24084 15502
rect 24032 15438 24084 15444
rect 23570 15399 23626 15408
rect 22006 15056 22062 15065
rect 24780 15026 24808 16526
rect 24872 15162 24900 19314
rect 24964 18834 24992 19382
rect 24952 18828 25004 18834
rect 24952 18770 25004 18776
rect 24952 18624 25004 18630
rect 25056 18612 25084 19382
rect 25148 19174 25176 21082
rect 25240 20602 25268 22374
rect 25424 21554 25452 22578
rect 25608 22574 25636 26182
rect 25700 25770 25728 27288
rect 25780 26036 25832 26042
rect 25780 25978 25832 25984
rect 25792 25809 25820 25978
rect 25884 25906 25912 27610
rect 25976 27554 26004 28698
rect 26068 28558 26096 30126
rect 26148 29844 26200 29850
rect 26148 29786 26200 29792
rect 26056 28552 26108 28558
rect 26056 28494 26108 28500
rect 26068 28218 26096 28494
rect 26056 28212 26108 28218
rect 26056 28154 26108 28160
rect 26160 28082 26188 29786
rect 26272 29404 26580 29413
rect 26272 29402 26278 29404
rect 26334 29402 26358 29404
rect 26414 29402 26438 29404
rect 26494 29402 26518 29404
rect 26574 29402 26580 29404
rect 26334 29350 26336 29402
rect 26516 29350 26518 29402
rect 26272 29348 26278 29350
rect 26334 29348 26358 29350
rect 26414 29348 26438 29350
rect 26494 29348 26518 29350
rect 26574 29348 26580 29350
rect 26272 29339 26580 29348
rect 26424 29232 26476 29238
rect 26424 29174 26476 29180
rect 26436 29034 26464 29174
rect 26424 29028 26476 29034
rect 26424 28970 26476 28976
rect 26712 28558 26740 33254
rect 26896 32502 26924 35974
rect 26988 34678 27016 37062
rect 27172 36961 27200 37062
rect 27158 36952 27214 36961
rect 27158 36887 27214 36896
rect 27160 36576 27212 36582
rect 27160 36518 27212 36524
rect 27252 36576 27304 36582
rect 27252 36518 27304 36524
rect 27068 36372 27120 36378
rect 27068 36314 27120 36320
rect 27080 35698 27108 36314
rect 27172 36145 27200 36518
rect 27158 36136 27214 36145
rect 27158 36071 27214 36080
rect 27158 35728 27214 35737
rect 27068 35692 27120 35698
rect 27158 35663 27214 35672
rect 27068 35634 27120 35640
rect 26976 34672 27028 34678
rect 26976 34614 27028 34620
rect 27080 33862 27108 35634
rect 27172 35290 27200 35663
rect 27160 35284 27212 35290
rect 27160 35226 27212 35232
rect 27160 35080 27212 35086
rect 27160 35022 27212 35028
rect 27172 34542 27200 35022
rect 27160 34536 27212 34542
rect 27160 34478 27212 34484
rect 27068 33856 27120 33862
rect 27068 33798 27120 33804
rect 26884 32496 26936 32502
rect 26884 32438 26936 32444
rect 27264 31906 27292 36518
rect 27540 36378 27568 37742
rect 27632 36854 27660 37742
rect 28092 37641 28120 38150
rect 28078 37632 28134 37641
rect 28078 37567 28134 37576
rect 28172 37256 28224 37262
rect 28172 37198 28224 37204
rect 27988 37120 28040 37126
rect 27988 37062 28040 37068
rect 27620 36848 27672 36854
rect 27620 36790 27672 36796
rect 27896 36644 27948 36650
rect 27896 36586 27948 36592
rect 27528 36372 27580 36378
rect 27528 36314 27580 36320
rect 27344 36168 27396 36174
rect 27344 36110 27396 36116
rect 27804 36168 27856 36174
rect 27804 36110 27856 36116
rect 27356 35630 27384 36110
rect 27436 36032 27488 36038
rect 27436 35974 27488 35980
rect 27344 35624 27396 35630
rect 27344 35566 27396 35572
rect 27448 34202 27476 35974
rect 27528 35488 27580 35494
rect 27528 35430 27580 35436
rect 27620 35488 27672 35494
rect 27620 35430 27672 35436
rect 27436 34196 27488 34202
rect 27436 34138 27488 34144
rect 27344 33924 27396 33930
rect 27344 33866 27396 33872
rect 27356 33522 27384 33866
rect 27436 33856 27488 33862
rect 27436 33798 27488 33804
rect 27344 33516 27396 33522
rect 27344 33458 27396 33464
rect 27448 33402 27476 33798
rect 27356 33374 27476 33402
rect 27356 32434 27384 33374
rect 27436 32768 27488 32774
rect 27436 32710 27488 32716
rect 27344 32428 27396 32434
rect 27344 32370 27396 32376
rect 27448 32298 27476 32710
rect 27540 32434 27568 35430
rect 27632 35193 27660 35430
rect 27618 35184 27674 35193
rect 27618 35119 27674 35128
rect 27712 35012 27764 35018
rect 27712 34954 27764 34960
rect 27620 34944 27672 34950
rect 27620 34886 27672 34892
rect 27632 34513 27660 34886
rect 27618 34504 27674 34513
rect 27618 34439 27674 34448
rect 27620 34128 27672 34134
rect 27620 34070 27672 34076
rect 27632 33454 27660 34070
rect 27620 33448 27672 33454
rect 27620 33390 27672 33396
rect 27618 33280 27674 33289
rect 27724 33266 27752 34954
rect 27674 33238 27752 33266
rect 27618 33215 27674 33224
rect 27528 32428 27580 32434
rect 27528 32370 27580 32376
rect 27632 32314 27660 33215
rect 27436 32292 27488 32298
rect 27436 32234 27488 32240
rect 27540 32286 27660 32314
rect 27080 31878 27292 31906
rect 27080 31414 27108 31878
rect 27160 31816 27212 31822
rect 27212 31776 27292 31804
rect 27160 31758 27212 31764
rect 27068 31408 27120 31414
rect 27068 31350 27120 31356
rect 27264 31346 27292 31776
rect 27448 31754 27476 32234
rect 27436 31748 27488 31754
rect 27436 31690 27488 31696
rect 26976 31340 27028 31346
rect 26976 31282 27028 31288
rect 27252 31340 27304 31346
rect 27304 31300 27384 31328
rect 27252 31282 27304 31288
rect 26792 31136 26844 31142
rect 26792 31078 26844 31084
rect 26700 28552 26752 28558
rect 26700 28494 26752 28500
rect 26272 28316 26580 28325
rect 26272 28314 26278 28316
rect 26334 28314 26358 28316
rect 26414 28314 26438 28316
rect 26494 28314 26518 28316
rect 26574 28314 26580 28316
rect 26334 28262 26336 28314
rect 26516 28262 26518 28314
rect 26272 28260 26278 28262
rect 26334 28260 26358 28262
rect 26414 28260 26438 28262
rect 26494 28260 26518 28262
rect 26574 28260 26580 28262
rect 26272 28251 26580 28260
rect 26148 28076 26200 28082
rect 26148 28018 26200 28024
rect 25976 27538 26096 27554
rect 25976 27532 26108 27538
rect 25976 27526 26056 27532
rect 25976 27402 26004 27526
rect 26056 27474 26108 27480
rect 25964 27396 26016 27402
rect 25964 27338 26016 27344
rect 26148 27328 26200 27334
rect 26148 27270 26200 27276
rect 26160 26586 26188 27270
rect 26272 27228 26580 27237
rect 26272 27226 26278 27228
rect 26334 27226 26358 27228
rect 26414 27226 26438 27228
rect 26494 27226 26518 27228
rect 26574 27226 26580 27228
rect 26334 27174 26336 27226
rect 26516 27174 26518 27226
rect 26272 27172 26278 27174
rect 26334 27172 26358 27174
rect 26414 27172 26438 27174
rect 26494 27172 26518 27174
rect 26574 27172 26580 27174
rect 26272 27163 26580 27172
rect 26330 26888 26386 26897
rect 26330 26823 26332 26832
rect 26384 26823 26386 26832
rect 26332 26794 26384 26800
rect 26148 26580 26200 26586
rect 26148 26522 26200 26528
rect 26056 26308 26108 26314
rect 26056 26250 26108 26256
rect 25962 25936 26018 25945
rect 25872 25900 25924 25906
rect 25962 25871 26018 25880
rect 25872 25842 25924 25848
rect 25778 25800 25834 25809
rect 25688 25764 25740 25770
rect 25778 25735 25834 25744
rect 25688 25706 25740 25712
rect 25686 25664 25742 25673
rect 25686 25599 25742 25608
rect 25700 25294 25728 25599
rect 25688 25288 25740 25294
rect 25688 25230 25740 25236
rect 25700 23730 25728 25230
rect 25976 24290 26004 25871
rect 26068 25430 26096 26250
rect 26056 25424 26108 25430
rect 26056 25366 26108 25372
rect 26068 25294 26096 25366
rect 26160 25362 26188 26522
rect 26608 26444 26660 26450
rect 26608 26386 26660 26392
rect 26272 26140 26580 26149
rect 26272 26138 26278 26140
rect 26334 26138 26358 26140
rect 26414 26138 26438 26140
rect 26494 26138 26518 26140
rect 26574 26138 26580 26140
rect 26334 26086 26336 26138
rect 26516 26086 26518 26138
rect 26272 26084 26278 26086
rect 26334 26084 26358 26086
rect 26414 26084 26438 26086
rect 26494 26084 26518 26086
rect 26574 26084 26580 26086
rect 26272 26075 26580 26084
rect 26424 25696 26476 25702
rect 26424 25638 26476 25644
rect 26148 25356 26200 25362
rect 26332 25356 26384 25362
rect 26148 25298 26200 25304
rect 26252 25316 26332 25344
rect 26056 25288 26108 25294
rect 26252 25242 26280 25316
rect 26332 25298 26384 25304
rect 26436 25265 26464 25638
rect 26514 25392 26570 25401
rect 26514 25327 26516 25336
rect 26568 25327 26570 25336
rect 26516 25298 26568 25304
rect 26620 25294 26648 26386
rect 26804 26382 26832 31078
rect 26884 29572 26936 29578
rect 26884 29514 26936 29520
rect 26896 29170 26924 29514
rect 26884 29164 26936 29170
rect 26884 29106 26936 29112
rect 26882 29064 26938 29073
rect 26882 28999 26938 29008
rect 26896 27946 26924 28999
rect 26884 27940 26936 27946
rect 26884 27882 26936 27888
rect 26792 26376 26844 26382
rect 26792 26318 26844 26324
rect 26700 25356 26752 25362
rect 26700 25298 26752 25304
rect 26608 25288 26660 25294
rect 26056 25230 26108 25236
rect 26160 25214 26280 25242
rect 26422 25256 26478 25265
rect 26160 24936 26188 25214
rect 26608 25230 26660 25236
rect 26422 25191 26478 25200
rect 26272 25052 26580 25061
rect 26272 25050 26278 25052
rect 26334 25050 26358 25052
rect 26414 25050 26438 25052
rect 26494 25050 26518 25052
rect 26574 25050 26580 25052
rect 26334 24998 26336 25050
rect 26516 24998 26518 25050
rect 26272 24996 26278 24998
rect 26334 24996 26358 24998
rect 26414 24996 26438 24998
rect 26494 24996 26518 24998
rect 26574 24996 26580 24998
rect 26272 24987 26580 24996
rect 26620 24954 26648 25230
rect 26608 24948 26660 24954
rect 26160 24908 26280 24936
rect 25884 24262 26004 24290
rect 25688 23724 25740 23730
rect 25884 23712 25912 24262
rect 25964 24200 26016 24206
rect 26252 24188 26280 24908
rect 26608 24890 26660 24896
rect 26712 24886 26740 25298
rect 26804 25294 26832 26318
rect 26884 26240 26936 26246
rect 26884 26182 26936 26188
rect 26896 25401 26924 26182
rect 26988 25770 27016 31282
rect 27068 31272 27120 31278
rect 27068 31214 27120 31220
rect 27080 28218 27108 31214
rect 27160 30796 27212 30802
rect 27160 30738 27212 30744
rect 27068 28212 27120 28218
rect 27068 28154 27120 28160
rect 27172 28098 27200 30738
rect 27356 30598 27384 31300
rect 27344 30592 27396 30598
rect 27344 30534 27396 30540
rect 27356 30190 27384 30534
rect 27344 30184 27396 30190
rect 27344 30126 27396 30132
rect 27342 29880 27398 29889
rect 27342 29815 27398 29824
rect 27356 29646 27384 29815
rect 27448 29714 27476 31690
rect 27436 29708 27488 29714
rect 27436 29650 27488 29656
rect 27344 29640 27396 29646
rect 27344 29582 27396 29588
rect 27252 29164 27304 29170
rect 27252 29106 27304 29112
rect 27264 28422 27292 29106
rect 27356 28762 27384 29582
rect 27448 29306 27476 29650
rect 27436 29300 27488 29306
rect 27436 29242 27488 29248
rect 27344 28756 27396 28762
rect 27344 28698 27396 28704
rect 27252 28416 27304 28422
rect 27252 28358 27304 28364
rect 27080 28070 27200 28098
rect 27540 28082 27568 32286
rect 27620 32020 27672 32026
rect 27620 31962 27672 31968
rect 27632 31686 27660 31962
rect 27620 31680 27672 31686
rect 27620 31622 27672 31628
rect 27618 31376 27674 31385
rect 27816 31346 27844 36110
rect 27908 35766 27936 36586
rect 27896 35760 27948 35766
rect 27896 35702 27948 35708
rect 28000 35018 28028 37062
rect 28184 35834 28212 37198
rect 28264 36168 28316 36174
rect 28264 36110 28316 36116
rect 28276 36009 28304 36110
rect 28262 36000 28318 36009
rect 28262 35935 28318 35944
rect 28172 35828 28224 35834
rect 28172 35770 28224 35776
rect 28170 35728 28226 35737
rect 28170 35663 28226 35672
rect 28080 35624 28132 35630
rect 28080 35566 28132 35572
rect 27988 35012 28040 35018
rect 27988 34954 28040 34960
rect 28092 33998 28120 35566
rect 28080 33992 28132 33998
rect 28080 33934 28132 33940
rect 28092 32230 28120 33934
rect 27988 32224 28040 32230
rect 27988 32166 28040 32172
rect 28080 32224 28132 32230
rect 28080 32166 28132 32172
rect 27896 31680 27948 31686
rect 27894 31648 27896 31657
rect 27948 31648 27950 31657
rect 27894 31583 27950 31592
rect 27618 31311 27674 31320
rect 27804 31340 27856 31346
rect 27632 28529 27660 31311
rect 27804 31282 27856 31288
rect 27712 30048 27764 30054
rect 27712 29990 27764 29996
rect 27724 29782 27752 29990
rect 27712 29776 27764 29782
rect 27712 29718 27764 29724
rect 27816 29730 27844 31282
rect 28000 30394 28028 32166
rect 28184 31822 28212 35663
rect 28264 34944 28316 34950
rect 28264 34886 28316 34892
rect 28276 33930 28304 34886
rect 28264 33924 28316 33930
rect 28264 33866 28316 33872
rect 28276 32434 28304 33866
rect 28264 32428 28316 32434
rect 28264 32370 28316 32376
rect 28172 31816 28224 31822
rect 28172 31758 28224 31764
rect 28264 31748 28316 31754
rect 28264 31690 28316 31696
rect 28276 30666 28304 31690
rect 28172 30660 28224 30666
rect 28172 30602 28224 30608
rect 28264 30660 28316 30666
rect 28264 30602 28316 30608
rect 28080 30592 28132 30598
rect 28080 30534 28132 30540
rect 27988 30388 28040 30394
rect 27988 30330 28040 30336
rect 27816 29702 27936 29730
rect 27802 29608 27858 29617
rect 27802 29543 27858 29552
rect 27712 29300 27764 29306
rect 27712 29242 27764 29248
rect 27724 29209 27752 29242
rect 27710 29200 27766 29209
rect 27816 29170 27844 29543
rect 27908 29510 27936 29702
rect 27988 29708 28040 29714
rect 27988 29650 28040 29656
rect 27896 29504 27948 29510
rect 27896 29446 27948 29452
rect 27710 29135 27766 29144
rect 27804 29164 27856 29170
rect 27804 29106 27856 29112
rect 27896 29164 27948 29170
rect 28000 29152 28028 29650
rect 27948 29124 28028 29152
rect 27896 29106 27948 29112
rect 27908 29034 27936 29106
rect 27896 29028 27948 29034
rect 27896 28970 27948 28976
rect 27988 29028 28040 29034
rect 27988 28970 28040 28976
rect 27802 28928 27858 28937
rect 27802 28863 27858 28872
rect 27816 28762 27844 28863
rect 27804 28756 27856 28762
rect 27804 28698 27856 28704
rect 27618 28520 27674 28529
rect 27618 28455 27674 28464
rect 27528 28076 27580 28082
rect 27080 27402 27108 28070
rect 27528 28018 27580 28024
rect 27160 28008 27212 28014
rect 27160 27950 27212 27956
rect 27172 27470 27200 27950
rect 27540 27674 27568 28018
rect 27528 27668 27580 27674
rect 27528 27610 27580 27616
rect 28000 27470 28028 28970
rect 28092 28966 28120 30534
rect 28184 29238 28212 30602
rect 28276 29730 28304 30602
rect 28368 30326 28396 38150
rect 28540 36780 28592 36786
rect 28540 36722 28592 36728
rect 28552 36582 28580 36722
rect 28448 36576 28500 36582
rect 28448 36518 28500 36524
rect 28540 36576 28592 36582
rect 28540 36518 28592 36524
rect 28460 32842 28488 36518
rect 28644 35737 28672 39222
rect 29012 37806 29040 41200
rect 32496 40044 32548 40050
rect 32496 39986 32548 39992
rect 30493 39740 30801 39749
rect 30493 39738 30499 39740
rect 30555 39738 30579 39740
rect 30635 39738 30659 39740
rect 30715 39738 30739 39740
rect 30795 39738 30801 39740
rect 30555 39686 30557 39738
rect 30737 39686 30739 39738
rect 30493 39684 30499 39686
rect 30555 39684 30579 39686
rect 30635 39684 30659 39686
rect 30715 39684 30739 39686
rect 30795 39684 30801 39686
rect 30493 39675 30801 39684
rect 32404 39636 32456 39642
rect 32404 39578 32456 39584
rect 29460 39568 29512 39574
rect 29460 39510 29512 39516
rect 31300 39568 31352 39574
rect 31300 39510 31352 39516
rect 32218 39536 32274 39545
rect 29472 38962 29500 39510
rect 29828 39432 29880 39438
rect 29828 39374 29880 39380
rect 30564 39432 30616 39438
rect 30564 39374 30616 39380
rect 29644 39296 29696 39302
rect 29644 39238 29696 39244
rect 29656 39030 29684 39238
rect 29644 39024 29696 39030
rect 29644 38966 29696 38972
rect 29460 38956 29512 38962
rect 29460 38898 29512 38904
rect 29368 38548 29420 38554
rect 29368 38490 29420 38496
rect 29380 38418 29408 38490
rect 29368 38412 29420 38418
rect 29368 38354 29420 38360
rect 29000 37800 29052 37806
rect 29000 37742 29052 37748
rect 29644 37800 29696 37806
rect 29644 37742 29696 37748
rect 29090 37496 29146 37505
rect 29090 37431 29146 37440
rect 29104 36786 29132 37431
rect 29184 37256 29236 37262
rect 29184 37198 29236 37204
rect 29092 36780 29144 36786
rect 29092 36722 29144 36728
rect 29196 36553 29224 37198
rect 29368 37120 29420 37126
rect 29368 37062 29420 37068
rect 29276 36576 29328 36582
rect 29182 36544 29238 36553
rect 29276 36518 29328 36524
rect 29182 36479 29238 36488
rect 29090 36408 29146 36417
rect 29090 36343 29146 36352
rect 28724 36304 28776 36310
rect 28724 36246 28776 36252
rect 28736 36156 28764 36246
rect 28908 36168 28960 36174
rect 28736 36128 28856 36156
rect 28724 36032 28776 36038
rect 28828 36009 28856 36128
rect 28908 36110 28960 36116
rect 28724 35974 28776 35980
rect 28814 36000 28870 36009
rect 28630 35728 28686 35737
rect 28630 35663 28686 35672
rect 28540 35624 28592 35630
rect 28540 35566 28592 35572
rect 28552 34746 28580 35566
rect 28632 35556 28684 35562
rect 28632 35498 28684 35504
rect 28644 35154 28672 35498
rect 28632 35148 28684 35154
rect 28632 35090 28684 35096
rect 28540 34740 28592 34746
rect 28540 34682 28592 34688
rect 28538 34096 28594 34105
rect 28538 34031 28594 34040
rect 28552 33998 28580 34031
rect 28540 33992 28592 33998
rect 28540 33934 28592 33940
rect 28540 33856 28592 33862
rect 28540 33798 28592 33804
rect 28632 33856 28684 33862
rect 28632 33798 28684 33804
rect 28552 33153 28580 33798
rect 28538 33144 28594 33153
rect 28538 33079 28594 33088
rect 28448 32836 28500 32842
rect 28448 32778 28500 32784
rect 28446 32736 28502 32745
rect 28446 32671 28502 32680
rect 28460 32178 28488 32671
rect 28552 32366 28580 33079
rect 28644 32502 28672 33798
rect 28632 32496 28684 32502
rect 28632 32438 28684 32444
rect 28540 32360 28592 32366
rect 28540 32302 28592 32308
rect 28460 32150 28672 32178
rect 28448 31816 28500 31822
rect 28500 31776 28580 31804
rect 28448 31758 28500 31764
rect 28448 30728 28500 30734
rect 28448 30670 28500 30676
rect 28356 30320 28408 30326
rect 28356 30262 28408 30268
rect 28460 30054 28488 30670
rect 28552 30666 28580 31776
rect 28540 30660 28592 30666
rect 28540 30602 28592 30608
rect 28540 30184 28592 30190
rect 28540 30126 28592 30132
rect 28448 30048 28500 30054
rect 28448 29990 28500 29996
rect 28552 29730 28580 30126
rect 28644 30122 28672 32150
rect 28736 31464 28764 35974
rect 28814 35935 28870 35944
rect 28816 35624 28868 35630
rect 28816 35566 28868 35572
rect 28828 34950 28856 35566
rect 28816 34944 28868 34950
rect 28816 34886 28868 34892
rect 28816 34604 28868 34610
rect 28816 34546 28868 34552
rect 28828 33289 28856 34546
rect 28814 33280 28870 33289
rect 28814 33215 28870 33224
rect 28814 33144 28870 33153
rect 28814 33079 28816 33088
rect 28868 33079 28870 33088
rect 28816 33050 28868 33056
rect 28920 31929 28948 36110
rect 29104 36106 29132 36343
rect 29182 36272 29238 36281
rect 29182 36207 29184 36216
rect 29236 36207 29238 36216
rect 29184 36178 29236 36184
rect 29092 36100 29144 36106
rect 29092 36042 29144 36048
rect 29182 35864 29238 35873
rect 29182 35799 29184 35808
rect 29236 35799 29238 35808
rect 29184 35770 29236 35776
rect 29184 35624 29236 35630
rect 29184 35566 29236 35572
rect 29000 35216 29052 35222
rect 29000 35158 29052 35164
rect 28906 31920 28962 31929
rect 28906 31855 28962 31864
rect 29012 31804 29040 35158
rect 29092 34128 29144 34134
rect 29092 34070 29144 34076
rect 29104 33930 29132 34070
rect 29092 33924 29144 33930
rect 29092 33866 29144 33872
rect 29196 33862 29224 35566
rect 29288 34746 29316 36518
rect 29380 36394 29408 37062
rect 29460 36780 29512 36786
rect 29460 36722 29512 36728
rect 29552 36780 29604 36786
rect 29552 36722 29604 36728
rect 29472 36553 29500 36722
rect 29458 36544 29514 36553
rect 29458 36479 29514 36488
rect 29380 36366 29500 36394
rect 29368 36032 29420 36038
rect 29368 35974 29420 35980
rect 29380 35222 29408 35974
rect 29368 35216 29420 35222
rect 29368 35158 29420 35164
rect 29366 35048 29422 35057
rect 29366 34983 29422 34992
rect 29380 34950 29408 34983
rect 29368 34944 29420 34950
rect 29368 34886 29420 34892
rect 29276 34740 29328 34746
rect 29276 34682 29328 34688
rect 29472 34626 29500 36366
rect 29288 34598 29500 34626
rect 29184 33856 29236 33862
rect 29184 33798 29236 33804
rect 29196 33318 29224 33798
rect 29288 33522 29316 34598
rect 29368 34536 29420 34542
rect 29368 34478 29420 34484
rect 29276 33516 29328 33522
rect 29276 33458 29328 33464
rect 29276 33380 29328 33386
rect 29276 33322 29328 33328
rect 29184 33312 29236 33318
rect 29184 33254 29236 33260
rect 29288 33114 29316 33322
rect 29276 33108 29328 33114
rect 29276 33050 29328 33056
rect 29184 32904 29236 32910
rect 29182 32872 29184 32881
rect 29236 32872 29238 32881
rect 29182 32807 29238 32816
rect 29184 32496 29236 32502
rect 29184 32438 29236 32444
rect 28920 31776 29040 31804
rect 28816 31748 28868 31754
rect 28816 31690 28868 31696
rect 28828 31657 28856 31690
rect 28814 31648 28870 31657
rect 28814 31583 28870 31592
rect 28736 31436 28856 31464
rect 28724 31340 28776 31346
rect 28724 31282 28776 31288
rect 28736 31142 28764 31282
rect 28724 31136 28776 31142
rect 28724 31078 28776 31084
rect 28828 30734 28856 31436
rect 28920 31226 28948 31776
rect 28920 31198 29040 31226
rect 28908 30932 28960 30938
rect 28908 30874 28960 30880
rect 28816 30728 28868 30734
rect 28816 30670 28868 30676
rect 28724 30592 28776 30598
rect 28724 30534 28776 30540
rect 28632 30116 28684 30122
rect 28632 30058 28684 30064
rect 28632 29844 28684 29850
rect 28632 29786 28684 29792
rect 28276 29702 28580 29730
rect 28264 29504 28316 29510
rect 28264 29446 28316 29452
rect 28172 29232 28224 29238
rect 28172 29174 28224 29180
rect 28080 28960 28132 28966
rect 28080 28902 28132 28908
rect 28078 27976 28134 27985
rect 28078 27911 28134 27920
rect 28092 27878 28120 27911
rect 28080 27872 28132 27878
rect 28080 27814 28132 27820
rect 27160 27464 27212 27470
rect 27160 27406 27212 27412
rect 27988 27464 28040 27470
rect 27988 27406 28040 27412
rect 27068 27396 27120 27402
rect 27068 27338 27120 27344
rect 27080 26790 27108 27338
rect 27620 27328 27672 27334
rect 27620 27270 27672 27276
rect 27160 26988 27212 26994
rect 27160 26930 27212 26936
rect 27068 26784 27120 26790
rect 27068 26726 27120 26732
rect 26976 25764 27028 25770
rect 26976 25706 27028 25712
rect 26882 25392 26938 25401
rect 26882 25327 26938 25336
rect 26792 25288 26844 25294
rect 26792 25230 26844 25236
rect 26700 24880 26752 24886
rect 26700 24822 26752 24828
rect 26804 24818 26832 25230
rect 26976 25220 27028 25226
rect 26976 25162 27028 25168
rect 26884 25152 26936 25158
rect 26884 25094 26936 25100
rect 26792 24812 26844 24818
rect 26792 24754 26844 24760
rect 26896 24206 26924 25094
rect 26988 24954 27016 25162
rect 26976 24948 27028 24954
rect 26976 24890 27028 24896
rect 27080 24886 27108 26726
rect 27068 24880 27120 24886
rect 27068 24822 27120 24828
rect 27068 24608 27120 24614
rect 27068 24550 27120 24556
rect 26976 24404 27028 24410
rect 26976 24346 27028 24352
rect 26988 24206 27016 24346
rect 27080 24274 27108 24550
rect 27068 24268 27120 24274
rect 27068 24210 27120 24216
rect 26016 24160 26280 24188
rect 26884 24200 26936 24206
rect 25964 24142 26016 24148
rect 26884 24142 26936 24148
rect 26976 24200 27028 24206
rect 26976 24142 27028 24148
rect 26700 24132 26752 24138
rect 26700 24074 26752 24080
rect 26272 23964 26580 23973
rect 26272 23962 26278 23964
rect 26334 23962 26358 23964
rect 26414 23962 26438 23964
rect 26494 23962 26518 23964
rect 26574 23962 26580 23964
rect 26334 23910 26336 23962
rect 26516 23910 26518 23962
rect 26272 23908 26278 23910
rect 26334 23908 26358 23910
rect 26414 23908 26438 23910
rect 26494 23908 26518 23910
rect 26574 23908 26580 23910
rect 26272 23899 26580 23908
rect 25964 23724 26016 23730
rect 25884 23684 25964 23712
rect 25688 23666 25740 23672
rect 25964 23666 26016 23672
rect 26608 23656 26660 23662
rect 26608 23598 26660 23604
rect 26272 22876 26580 22885
rect 26272 22874 26278 22876
rect 26334 22874 26358 22876
rect 26414 22874 26438 22876
rect 26494 22874 26518 22876
rect 26574 22874 26580 22876
rect 26334 22822 26336 22874
rect 26516 22822 26518 22874
rect 26272 22820 26278 22822
rect 26334 22820 26358 22822
rect 26414 22820 26438 22822
rect 26494 22820 26518 22822
rect 26574 22820 26580 22822
rect 26272 22811 26580 22820
rect 26620 22778 26648 23598
rect 26608 22772 26660 22778
rect 26608 22714 26660 22720
rect 26712 22710 26740 24074
rect 26884 23792 26936 23798
rect 26884 23734 26936 23740
rect 26896 23254 26924 23734
rect 26976 23724 27028 23730
rect 26976 23666 27028 23672
rect 26884 23248 26936 23254
rect 26884 23190 26936 23196
rect 26896 22778 26924 23190
rect 26884 22772 26936 22778
rect 26884 22714 26936 22720
rect 26700 22704 26752 22710
rect 26700 22646 26752 22652
rect 25596 22568 25648 22574
rect 25596 22510 25648 22516
rect 25608 21554 25636 22510
rect 26896 21962 26924 22714
rect 25688 21956 25740 21962
rect 25688 21898 25740 21904
rect 26884 21956 26936 21962
rect 26884 21898 26936 21904
rect 25412 21548 25464 21554
rect 25412 21490 25464 21496
rect 25596 21548 25648 21554
rect 25596 21490 25648 21496
rect 25424 20806 25452 21490
rect 25412 20800 25464 20806
rect 25412 20742 25464 20748
rect 25228 20596 25280 20602
rect 25228 20538 25280 20544
rect 25136 19168 25188 19174
rect 25136 19110 25188 19116
rect 25320 19168 25372 19174
rect 25320 19110 25372 19116
rect 25148 18766 25176 19110
rect 25136 18760 25188 18766
rect 25136 18702 25188 18708
rect 25004 18584 25084 18612
rect 24952 18566 25004 18572
rect 24964 18426 24992 18566
rect 24952 18420 25004 18426
rect 24952 18362 25004 18368
rect 25332 18290 25360 19110
rect 25424 18970 25452 20742
rect 25608 19786 25636 21490
rect 25700 20777 25728 21898
rect 25780 21888 25832 21894
rect 25780 21830 25832 21836
rect 25686 20768 25742 20777
rect 25686 20703 25742 20712
rect 25792 20466 25820 21830
rect 26272 21788 26580 21797
rect 26272 21786 26278 21788
rect 26334 21786 26358 21788
rect 26414 21786 26438 21788
rect 26494 21786 26518 21788
rect 26574 21786 26580 21788
rect 26334 21734 26336 21786
rect 26516 21734 26518 21786
rect 26272 21732 26278 21734
rect 26334 21732 26358 21734
rect 26414 21732 26438 21734
rect 26494 21732 26518 21734
rect 26574 21732 26580 21734
rect 26272 21723 26580 21732
rect 26896 21622 26924 21898
rect 26884 21616 26936 21622
rect 26884 21558 26936 21564
rect 26056 21344 26108 21350
rect 26056 21286 26108 21292
rect 26516 21344 26568 21350
rect 26516 21286 26568 21292
rect 26884 21344 26936 21350
rect 26884 21286 26936 21292
rect 25964 20800 26016 20806
rect 25964 20742 26016 20748
rect 25976 20466 26004 20742
rect 26068 20602 26096 21286
rect 26528 20874 26556 21286
rect 26516 20868 26568 20874
rect 26568 20828 26648 20856
rect 26516 20810 26568 20816
rect 26272 20700 26580 20709
rect 26272 20698 26278 20700
rect 26334 20698 26358 20700
rect 26414 20698 26438 20700
rect 26494 20698 26518 20700
rect 26574 20698 26580 20700
rect 26334 20646 26336 20698
rect 26516 20646 26518 20698
rect 26272 20644 26278 20646
rect 26334 20644 26358 20646
rect 26414 20644 26438 20646
rect 26494 20644 26518 20646
rect 26574 20644 26580 20646
rect 26272 20635 26580 20644
rect 26056 20596 26108 20602
rect 26056 20538 26108 20544
rect 26332 20596 26384 20602
rect 26332 20538 26384 20544
rect 26344 20466 26372 20538
rect 26620 20534 26648 20828
rect 26896 20806 26924 21286
rect 26884 20800 26936 20806
rect 26884 20742 26936 20748
rect 26608 20528 26660 20534
rect 26608 20470 26660 20476
rect 25780 20460 25832 20466
rect 25780 20402 25832 20408
rect 25964 20460 26016 20466
rect 25964 20402 26016 20408
rect 26332 20460 26384 20466
rect 26332 20402 26384 20408
rect 26424 20460 26476 20466
rect 26424 20402 26476 20408
rect 26056 20324 26108 20330
rect 26056 20266 26108 20272
rect 25596 19780 25648 19786
rect 25596 19722 25648 19728
rect 25964 19712 26016 19718
rect 25964 19654 26016 19660
rect 25976 19514 26004 19654
rect 25964 19508 26016 19514
rect 25964 19450 26016 19456
rect 25872 19304 25924 19310
rect 25872 19246 25924 19252
rect 25780 19236 25832 19242
rect 25780 19178 25832 19184
rect 25412 18964 25464 18970
rect 25412 18906 25464 18912
rect 25320 18284 25372 18290
rect 25320 18226 25372 18232
rect 25136 18148 25188 18154
rect 25136 18090 25188 18096
rect 24952 17536 25004 17542
rect 24952 17478 25004 17484
rect 24964 16998 24992 17478
rect 25044 17264 25096 17270
rect 25044 17206 25096 17212
rect 24952 16992 25004 16998
rect 24952 16934 25004 16940
rect 24952 16516 25004 16522
rect 24952 16458 25004 16464
rect 24964 15910 24992 16458
rect 24952 15904 25004 15910
rect 24952 15846 25004 15852
rect 25056 15502 25084 17206
rect 25148 16590 25176 18090
rect 25320 17604 25372 17610
rect 25320 17546 25372 17552
rect 25228 16992 25280 16998
rect 25228 16934 25280 16940
rect 25240 16658 25268 16934
rect 25228 16652 25280 16658
rect 25228 16594 25280 16600
rect 25136 16584 25188 16590
rect 25136 16526 25188 16532
rect 25240 16114 25268 16594
rect 25332 16250 25360 17546
rect 25688 17536 25740 17542
rect 25688 17478 25740 17484
rect 25700 17338 25728 17478
rect 25688 17332 25740 17338
rect 25688 17274 25740 17280
rect 25596 17264 25648 17270
rect 25596 17206 25648 17212
rect 25504 17060 25556 17066
rect 25504 17002 25556 17008
rect 25516 16590 25544 17002
rect 25608 16590 25636 17206
rect 25504 16584 25556 16590
rect 25504 16526 25556 16532
rect 25596 16584 25648 16590
rect 25596 16526 25648 16532
rect 25412 16448 25464 16454
rect 25412 16390 25464 16396
rect 25320 16244 25372 16250
rect 25320 16186 25372 16192
rect 25424 16114 25452 16390
rect 25516 16182 25544 16526
rect 25700 16522 25728 17274
rect 25688 16516 25740 16522
rect 25688 16458 25740 16464
rect 25504 16176 25556 16182
rect 25504 16118 25556 16124
rect 25228 16108 25280 16114
rect 25228 16050 25280 16056
rect 25412 16108 25464 16114
rect 25412 16050 25464 16056
rect 25044 15496 25096 15502
rect 25044 15438 25096 15444
rect 25412 15360 25464 15366
rect 25412 15302 25464 15308
rect 24860 15156 24912 15162
rect 24860 15098 24912 15104
rect 25424 15026 25452 15302
rect 22006 14991 22008 15000
rect 22060 14991 22062 15000
rect 24768 15020 24820 15026
rect 22008 14962 22060 14968
rect 24768 14962 24820 14968
rect 25412 15020 25464 15026
rect 25412 14962 25464 14968
rect 22020 14906 22048 14962
rect 19076 6886 19196 6914
rect 21928 14878 22048 14906
rect 17831 6556 18139 6565
rect 17831 6554 17837 6556
rect 17893 6554 17917 6556
rect 17973 6554 17997 6556
rect 18053 6554 18077 6556
rect 18133 6554 18139 6556
rect 17893 6502 17895 6554
rect 18075 6502 18077 6554
rect 17831 6500 17837 6502
rect 17893 6500 17917 6502
rect 17973 6500 17997 6502
rect 18053 6500 18077 6502
rect 18133 6500 18139 6502
rect 17831 6491 18139 6500
rect 17831 5468 18139 5477
rect 17831 5466 17837 5468
rect 17893 5466 17917 5468
rect 17973 5466 17997 5468
rect 18053 5466 18077 5468
rect 18133 5466 18139 5468
rect 17893 5414 17895 5466
rect 18075 5414 18077 5466
rect 17831 5412 17837 5414
rect 17893 5412 17917 5414
rect 17973 5412 17997 5414
rect 18053 5412 18077 5414
rect 18133 5412 18139 5414
rect 17831 5403 18139 5412
rect 17831 4380 18139 4389
rect 17831 4378 17837 4380
rect 17893 4378 17917 4380
rect 17973 4378 17997 4380
rect 18053 4378 18077 4380
rect 18133 4378 18139 4380
rect 17893 4326 17895 4378
rect 18075 4326 18077 4378
rect 17831 4324 17837 4326
rect 17893 4324 17917 4326
rect 17973 4324 17997 4326
rect 18053 4324 18077 4326
rect 18133 4324 18139 4326
rect 17831 4315 18139 4324
rect 15660 4004 15712 4010
rect 15660 3946 15712 3952
rect 15568 3936 15620 3942
rect 15568 3878 15620 3884
rect 14372 3664 14424 3670
rect 14372 3606 14424 3612
rect 14384 3534 14412 3606
rect 15580 3602 15608 3878
rect 15568 3596 15620 3602
rect 15568 3538 15620 3544
rect 14280 3528 14332 3534
rect 14280 3470 14332 3476
rect 14372 3528 14424 3534
rect 14372 3470 14424 3476
rect 14292 3058 14320 3470
rect 14464 3392 14516 3398
rect 14464 3334 14516 3340
rect 14476 3126 14504 3334
rect 14464 3120 14516 3126
rect 14464 3062 14516 3068
rect 14280 3052 14332 3058
rect 14280 2994 14332 3000
rect 14832 2984 14884 2990
rect 14832 2926 14884 2932
rect 13611 2748 13919 2757
rect 13611 2746 13617 2748
rect 13673 2746 13697 2748
rect 13753 2746 13777 2748
rect 13833 2746 13857 2748
rect 13913 2746 13919 2748
rect 13673 2694 13675 2746
rect 13855 2694 13857 2746
rect 13611 2692 13617 2694
rect 13673 2692 13697 2694
rect 13753 2692 13777 2694
rect 13833 2692 13857 2694
rect 13913 2692 13919 2694
rect 13611 2683 13919 2692
rect 13464 2230 13584 2258
rect 13556 800 13584 2230
rect 14844 800 14872 2926
rect 15672 2446 15700 3946
rect 16856 3936 16908 3942
rect 16856 3878 16908 3884
rect 16120 3596 16172 3602
rect 16120 3538 16172 3544
rect 15752 3460 15804 3466
rect 15752 3402 15804 3408
rect 15764 2650 15792 3402
rect 15752 2644 15804 2650
rect 15752 2586 15804 2592
rect 15660 2440 15712 2446
rect 15660 2382 15712 2388
rect 16132 800 16160 3538
rect 16868 3058 16896 3878
rect 17831 3292 18139 3301
rect 17831 3290 17837 3292
rect 17893 3290 17917 3292
rect 17973 3290 17997 3292
rect 18053 3290 18077 3292
rect 18133 3290 18139 3292
rect 17893 3238 17895 3290
rect 18075 3238 18077 3290
rect 17831 3236 17837 3238
rect 17893 3236 17917 3238
rect 17973 3236 17997 3238
rect 18053 3236 18077 3238
rect 18133 3236 18139 3238
rect 17831 3227 18139 3236
rect 16856 3052 16908 3058
rect 16856 2994 16908 3000
rect 17040 2984 17092 2990
rect 17040 2926 17092 2932
rect 17408 2984 17460 2990
rect 17408 2926 17460 2932
rect 17052 2650 17080 2926
rect 17040 2644 17092 2650
rect 17040 2586 17092 2592
rect 17420 800 17448 2926
rect 19076 2650 19104 6886
rect 19984 6792 20036 6798
rect 19984 6734 20036 6740
rect 19996 4622 20024 6734
rect 19984 4616 20036 4622
rect 19984 4558 20036 4564
rect 19800 4480 19852 4486
rect 19800 4422 19852 4428
rect 19812 4214 19840 4422
rect 19800 4208 19852 4214
rect 19800 4150 19852 4156
rect 20260 4072 20312 4078
rect 20260 4014 20312 4020
rect 20628 4072 20680 4078
rect 20628 4014 20680 4020
rect 20076 3936 20128 3942
rect 20076 3878 20128 3884
rect 20088 3738 20116 3878
rect 20272 3738 20300 4014
rect 20076 3732 20128 3738
rect 20076 3674 20128 3680
rect 20260 3732 20312 3738
rect 20260 3674 20312 3680
rect 19432 3528 19484 3534
rect 19432 3470 19484 3476
rect 19340 3188 19392 3194
rect 19340 3130 19392 3136
rect 19064 2644 19116 2650
rect 19064 2586 19116 2592
rect 19352 2446 19380 3130
rect 19444 3058 19472 3470
rect 19432 3052 19484 3058
rect 19432 2994 19484 3000
rect 19616 2984 19668 2990
rect 19616 2926 19668 2932
rect 19984 2984 20036 2990
rect 19984 2926 20036 2932
rect 19628 2650 19656 2926
rect 19616 2644 19668 2650
rect 19616 2586 19668 2592
rect 18236 2440 18288 2446
rect 18236 2382 18288 2388
rect 19340 2440 19392 2446
rect 19340 2382 19392 2388
rect 17831 2204 18139 2213
rect 17831 2202 17837 2204
rect 17893 2202 17917 2204
rect 17973 2202 17997 2204
rect 18053 2202 18077 2204
rect 18133 2202 18139 2204
rect 17893 2150 17895 2202
rect 18075 2150 18077 2202
rect 17831 2148 17837 2150
rect 17893 2148 17917 2150
rect 17973 2148 17997 2150
rect 18053 2148 18077 2150
rect 18133 2148 18139 2150
rect 17831 2139 18139 2148
rect 18248 1442 18276 2382
rect 18064 1414 18276 1442
rect 18064 800 18092 1414
rect 19996 800 20024 2926
rect 20640 800 20668 4014
rect 21272 3596 21324 3602
rect 21272 3538 21324 3544
rect 20720 3528 20772 3534
rect 20720 3470 20772 3476
rect 20732 2650 20760 3470
rect 20720 2644 20772 2650
rect 20720 2586 20772 2592
rect 21284 800 21312 3538
rect 21928 3058 21956 14878
rect 22052 14716 22360 14725
rect 22052 14714 22058 14716
rect 22114 14714 22138 14716
rect 22194 14714 22218 14716
rect 22274 14714 22298 14716
rect 22354 14714 22360 14716
rect 22114 14662 22116 14714
rect 22296 14662 22298 14714
rect 22052 14660 22058 14662
rect 22114 14660 22138 14662
rect 22194 14660 22218 14662
rect 22274 14660 22298 14662
rect 22354 14660 22360 14662
rect 22052 14651 22360 14660
rect 25516 14414 25544 16118
rect 25596 16040 25648 16046
rect 25596 15982 25648 15988
rect 25608 15910 25636 15982
rect 25596 15904 25648 15910
rect 25596 15846 25648 15852
rect 25608 15434 25636 15846
rect 25700 15570 25728 16458
rect 25688 15564 25740 15570
rect 25688 15506 25740 15512
rect 25596 15428 25648 15434
rect 25596 15370 25648 15376
rect 25594 15328 25650 15337
rect 25594 15263 25650 15272
rect 25608 15162 25636 15263
rect 25596 15156 25648 15162
rect 25596 15098 25648 15104
rect 25594 15056 25650 15065
rect 25792 15026 25820 19178
rect 25884 17134 25912 19246
rect 25872 17128 25924 17134
rect 25872 17070 25924 17076
rect 25870 16552 25926 16561
rect 25870 16487 25926 16496
rect 25884 15502 25912 16487
rect 25872 15496 25924 15502
rect 25872 15438 25924 15444
rect 25594 14991 25596 15000
rect 25648 14991 25650 15000
rect 25780 15020 25832 15026
rect 25596 14962 25648 14968
rect 25780 14962 25832 14968
rect 25976 14414 26004 19450
rect 26068 19378 26096 20266
rect 26344 19836 26372 20402
rect 26436 20330 26464 20402
rect 26424 20324 26476 20330
rect 26424 20266 26476 20272
rect 26516 20256 26568 20262
rect 26568 20216 26648 20244
rect 26516 20198 26568 20204
rect 26160 19808 26372 19836
rect 26160 19378 26188 19808
rect 26272 19612 26580 19621
rect 26272 19610 26278 19612
rect 26334 19610 26358 19612
rect 26414 19610 26438 19612
rect 26494 19610 26518 19612
rect 26574 19610 26580 19612
rect 26334 19558 26336 19610
rect 26516 19558 26518 19610
rect 26272 19556 26278 19558
rect 26334 19556 26358 19558
rect 26414 19556 26438 19558
rect 26494 19556 26518 19558
rect 26574 19556 26580 19558
rect 26272 19547 26580 19556
rect 26332 19508 26384 19514
rect 26332 19450 26384 19456
rect 26056 19372 26108 19378
rect 26056 19314 26108 19320
rect 26148 19372 26200 19378
rect 26148 19314 26200 19320
rect 26148 19168 26200 19174
rect 26148 19110 26200 19116
rect 26160 18766 26188 19110
rect 26148 18760 26200 18766
rect 26148 18702 26200 18708
rect 26344 18698 26372 19450
rect 26620 18766 26648 20216
rect 26792 19848 26844 19854
rect 26792 19790 26844 19796
rect 26804 19378 26832 19790
rect 26792 19372 26844 19378
rect 26792 19314 26844 19320
rect 26608 18760 26660 18766
rect 26608 18702 26660 18708
rect 26332 18692 26384 18698
rect 26332 18634 26384 18640
rect 26272 18524 26580 18533
rect 26272 18522 26278 18524
rect 26334 18522 26358 18524
rect 26414 18522 26438 18524
rect 26494 18522 26518 18524
rect 26574 18522 26580 18524
rect 26334 18470 26336 18522
rect 26516 18470 26518 18522
rect 26272 18468 26278 18470
rect 26334 18468 26358 18470
rect 26414 18468 26438 18470
rect 26494 18468 26518 18470
rect 26574 18468 26580 18470
rect 26272 18459 26580 18468
rect 26608 18420 26660 18426
rect 26608 18362 26660 18368
rect 26056 18080 26108 18086
rect 26056 18022 26108 18028
rect 26068 17882 26096 18022
rect 26056 17876 26108 17882
rect 26056 17818 26108 17824
rect 26068 17270 26096 17818
rect 26148 17536 26200 17542
rect 26148 17478 26200 17484
rect 26056 17264 26108 17270
rect 26056 17206 26108 17212
rect 26056 17128 26108 17134
rect 26056 17070 26108 17076
rect 25504 14408 25556 14414
rect 25504 14350 25556 14356
rect 25964 14408 26016 14414
rect 25964 14350 26016 14356
rect 26068 14346 26096 17070
rect 26160 16590 26188 17478
rect 26272 17436 26580 17445
rect 26272 17434 26278 17436
rect 26334 17434 26358 17436
rect 26414 17434 26438 17436
rect 26494 17434 26518 17436
rect 26574 17434 26580 17436
rect 26334 17382 26336 17434
rect 26516 17382 26518 17434
rect 26272 17380 26278 17382
rect 26334 17380 26358 17382
rect 26414 17380 26438 17382
rect 26494 17380 26518 17382
rect 26574 17380 26580 17382
rect 26272 17371 26580 17380
rect 26516 16992 26568 16998
rect 26516 16934 26568 16940
rect 26148 16584 26200 16590
rect 26148 16526 26200 16532
rect 26160 16114 26188 16526
rect 26528 16454 26556 16934
rect 26516 16448 26568 16454
rect 26516 16390 26568 16396
rect 26272 16348 26580 16357
rect 26272 16346 26278 16348
rect 26334 16346 26358 16348
rect 26414 16346 26438 16348
rect 26494 16346 26518 16348
rect 26574 16346 26580 16348
rect 26334 16294 26336 16346
rect 26516 16294 26518 16346
rect 26272 16292 26278 16294
rect 26334 16292 26358 16294
rect 26414 16292 26438 16294
rect 26494 16292 26518 16294
rect 26574 16292 26580 16294
rect 26272 16283 26580 16292
rect 26148 16108 26200 16114
rect 26148 16050 26200 16056
rect 26160 15026 26188 16050
rect 26620 15994 26648 18362
rect 26700 17604 26752 17610
rect 26700 17546 26752 17552
rect 26528 15966 26648 15994
rect 26424 15632 26476 15638
rect 26424 15574 26476 15580
rect 26436 15473 26464 15574
rect 26422 15464 26478 15473
rect 26422 15399 26424 15408
rect 26476 15399 26478 15408
rect 26424 15370 26476 15376
rect 26528 15366 26556 15966
rect 26608 15904 26660 15910
rect 26608 15846 26660 15852
rect 26516 15360 26568 15366
rect 26516 15302 26568 15308
rect 26272 15260 26580 15269
rect 26272 15258 26278 15260
rect 26334 15258 26358 15260
rect 26414 15258 26438 15260
rect 26494 15258 26518 15260
rect 26574 15258 26580 15260
rect 26334 15206 26336 15258
rect 26516 15206 26518 15258
rect 26272 15204 26278 15206
rect 26334 15204 26358 15206
rect 26414 15204 26438 15206
rect 26494 15204 26518 15206
rect 26574 15204 26580 15206
rect 26272 15195 26580 15204
rect 26148 15020 26200 15026
rect 26148 14962 26200 14968
rect 26620 14414 26648 15846
rect 26712 14618 26740 17546
rect 26896 17338 26924 20742
rect 26988 20602 27016 23666
rect 27080 23662 27108 24210
rect 27068 23656 27120 23662
rect 27068 23598 27120 23604
rect 27080 23050 27108 23598
rect 27068 23044 27120 23050
rect 27068 22986 27120 22992
rect 27068 22024 27120 22030
rect 27068 21966 27120 21972
rect 27080 21486 27108 21966
rect 27172 21690 27200 26930
rect 27528 26308 27580 26314
rect 27528 26250 27580 26256
rect 27436 26036 27488 26042
rect 27436 25978 27488 25984
rect 27344 25900 27396 25906
rect 27344 25842 27396 25848
rect 27252 25764 27304 25770
rect 27252 25706 27304 25712
rect 27264 25226 27292 25706
rect 27356 25537 27384 25842
rect 27448 25809 27476 25978
rect 27540 25974 27568 26250
rect 27528 25968 27580 25974
rect 27528 25910 27580 25916
rect 27632 25906 27660 27270
rect 28000 26858 28028 27406
rect 28080 27396 28132 27402
rect 28080 27338 28132 27344
rect 27988 26852 28040 26858
rect 27988 26794 28040 26800
rect 27804 26240 27856 26246
rect 27804 26182 27856 26188
rect 27816 25906 27844 26182
rect 27620 25900 27672 25906
rect 27620 25842 27672 25848
rect 27804 25900 27856 25906
rect 27804 25842 27856 25848
rect 27988 25900 28040 25906
rect 27988 25842 28040 25848
rect 27434 25800 27490 25809
rect 27434 25735 27490 25744
rect 27434 25664 27490 25673
rect 27434 25599 27490 25608
rect 27342 25528 27398 25537
rect 27342 25463 27398 25472
rect 27448 25294 27476 25599
rect 27528 25424 27580 25430
rect 27528 25366 27580 25372
rect 27436 25288 27488 25294
rect 27436 25230 27488 25236
rect 27252 25220 27304 25226
rect 27252 25162 27304 25168
rect 27540 24857 27568 25366
rect 27632 24954 27660 25842
rect 27896 25764 27948 25770
rect 27896 25706 27948 25712
rect 27620 24948 27672 24954
rect 27620 24890 27672 24896
rect 27526 24848 27582 24857
rect 27526 24783 27582 24792
rect 27436 24404 27488 24410
rect 27436 24346 27488 24352
rect 27252 22636 27304 22642
rect 27252 22578 27304 22584
rect 27264 22166 27292 22578
rect 27252 22160 27304 22166
rect 27252 22102 27304 22108
rect 27264 21962 27292 22102
rect 27448 22030 27476 24346
rect 27632 23866 27660 24890
rect 27620 23860 27672 23866
rect 27620 23802 27672 23808
rect 27528 23588 27580 23594
rect 27528 23530 27580 23536
rect 27540 23050 27568 23530
rect 27618 23080 27674 23089
rect 27528 23044 27580 23050
rect 27618 23015 27620 23024
rect 27528 22986 27580 22992
rect 27672 23015 27674 23024
rect 27620 22986 27672 22992
rect 27540 22642 27568 22986
rect 27528 22636 27580 22642
rect 27528 22578 27580 22584
rect 27804 22432 27856 22438
rect 27804 22374 27856 22380
rect 27816 22030 27844 22374
rect 27436 22024 27488 22030
rect 27436 21966 27488 21972
rect 27804 22024 27856 22030
rect 27804 21966 27856 21972
rect 27252 21956 27304 21962
rect 27252 21898 27304 21904
rect 27160 21684 27212 21690
rect 27160 21626 27212 21632
rect 27068 21480 27120 21486
rect 27068 21422 27120 21428
rect 26976 20596 27028 20602
rect 26976 20538 27028 20544
rect 26976 19236 27028 19242
rect 26976 19178 27028 19184
rect 26988 18698 27016 19178
rect 26976 18692 27028 18698
rect 26976 18634 27028 18640
rect 26884 17332 26936 17338
rect 26884 17274 26936 17280
rect 26792 17196 26844 17202
rect 26792 17138 26844 17144
rect 26804 15706 26832 17138
rect 26884 16448 26936 16454
rect 26884 16390 26936 16396
rect 26792 15700 26844 15706
rect 26792 15642 26844 15648
rect 26896 15502 26924 16390
rect 26988 15706 27016 18634
rect 26976 15700 27028 15706
rect 26976 15642 27028 15648
rect 26884 15496 26936 15502
rect 26884 15438 26936 15444
rect 26700 14612 26752 14618
rect 26700 14554 26752 14560
rect 26896 14414 26924 15438
rect 27080 15162 27108 21422
rect 27264 20584 27292 21898
rect 27344 21888 27396 21894
rect 27344 21830 27396 21836
rect 27356 21622 27384 21830
rect 27344 21616 27396 21622
rect 27344 21558 27396 21564
rect 27448 21350 27476 21966
rect 27908 21962 27936 25706
rect 28000 25498 28028 25842
rect 27988 25492 28040 25498
rect 27988 25434 28040 25440
rect 28092 25294 28120 27338
rect 28184 27130 28212 29174
rect 28276 27470 28304 29446
rect 28368 28014 28396 29702
rect 28540 29640 28592 29646
rect 28644 29628 28672 29786
rect 28736 29714 28764 30534
rect 28724 29708 28776 29714
rect 28724 29650 28776 29656
rect 28592 29600 28672 29628
rect 28540 29582 28592 29588
rect 28736 29510 28764 29650
rect 28828 29578 28856 30670
rect 28816 29572 28868 29578
rect 28816 29514 28868 29520
rect 28724 29504 28776 29510
rect 28724 29446 28776 29452
rect 28828 29170 28856 29514
rect 28816 29164 28868 29170
rect 28816 29106 28868 29112
rect 28448 28960 28500 28966
rect 28448 28902 28500 28908
rect 28460 28422 28488 28902
rect 28448 28416 28500 28422
rect 28920 28393 28948 30874
rect 29012 30161 29040 31198
rect 29196 30870 29224 32438
rect 29380 31754 29408 34478
rect 29460 34060 29512 34066
rect 29460 34002 29512 34008
rect 29472 33522 29500 34002
rect 29460 33516 29512 33522
rect 29460 33458 29512 33464
rect 29460 32564 29512 32570
rect 29460 32506 29512 32512
rect 29472 32473 29500 32506
rect 29458 32464 29514 32473
rect 29458 32399 29514 32408
rect 29472 32366 29500 32399
rect 29460 32360 29512 32366
rect 29460 32302 29512 32308
rect 29460 32224 29512 32230
rect 29460 32166 29512 32172
rect 29368 31748 29420 31754
rect 29368 31690 29420 31696
rect 29380 31362 29408 31690
rect 29288 31334 29408 31362
rect 29184 30864 29236 30870
rect 29184 30806 29236 30812
rect 29092 30796 29144 30802
rect 29092 30738 29144 30744
rect 29104 30705 29132 30738
rect 29090 30696 29146 30705
rect 29090 30631 29146 30640
rect 28998 30152 29054 30161
rect 28998 30087 29054 30096
rect 29092 30048 29144 30054
rect 29092 29990 29144 29996
rect 29104 29646 29132 29990
rect 29288 29850 29316 31334
rect 29472 31226 29500 32166
rect 29380 31210 29500 31226
rect 29368 31204 29500 31210
rect 29420 31198 29500 31204
rect 29368 31146 29420 31152
rect 29458 31104 29514 31113
rect 29458 31039 29514 31048
rect 29368 30932 29420 30938
rect 29368 30874 29420 30880
rect 29276 29844 29328 29850
rect 29276 29786 29328 29792
rect 29092 29640 29144 29646
rect 29092 29582 29144 29588
rect 29184 29640 29236 29646
rect 29184 29582 29236 29588
rect 29092 29164 29144 29170
rect 29092 29106 29144 29112
rect 29000 28756 29052 28762
rect 29000 28698 29052 28704
rect 29012 28626 29040 28698
rect 29000 28620 29052 28626
rect 29000 28562 29052 28568
rect 29104 28558 29132 29106
rect 29196 28966 29224 29582
rect 29274 29472 29330 29481
rect 29274 29407 29330 29416
rect 29184 28960 29236 28966
rect 29184 28902 29236 28908
rect 29092 28552 29144 28558
rect 29092 28494 29144 28500
rect 28448 28358 28500 28364
rect 28906 28384 28962 28393
rect 28356 28008 28408 28014
rect 28356 27950 28408 27956
rect 28264 27464 28316 27470
rect 28264 27406 28316 27412
rect 28172 27124 28224 27130
rect 28172 27066 28224 27072
rect 28172 26852 28224 26858
rect 28172 26794 28224 26800
rect 28184 25945 28212 26794
rect 28460 26518 28488 28358
rect 28906 28319 28962 28328
rect 29104 28234 29132 28494
rect 29184 28484 29236 28490
rect 29184 28426 29236 28432
rect 28920 28206 29132 28234
rect 28816 28144 28868 28150
rect 28816 28086 28868 28092
rect 28828 27713 28856 28086
rect 28814 27704 28870 27713
rect 28814 27639 28870 27648
rect 28920 27470 28948 28206
rect 29090 28112 29146 28121
rect 29000 28076 29052 28082
rect 29090 28047 29146 28056
rect 29000 28018 29052 28024
rect 29012 27985 29040 28018
rect 29104 28014 29132 28047
rect 29092 28008 29144 28014
rect 28998 27976 29054 27985
rect 29092 27950 29144 27956
rect 28998 27911 29054 27920
rect 28908 27464 28960 27470
rect 28908 27406 28960 27412
rect 28724 27328 28776 27334
rect 28724 27270 28776 27276
rect 28540 27124 28592 27130
rect 28540 27066 28592 27072
rect 28264 26512 28316 26518
rect 28264 26454 28316 26460
rect 28448 26512 28500 26518
rect 28448 26454 28500 26460
rect 28276 26246 28304 26454
rect 28264 26240 28316 26246
rect 28264 26182 28316 26188
rect 28170 25936 28226 25945
rect 28226 25880 28304 25888
rect 28170 25871 28172 25880
rect 28224 25860 28304 25880
rect 28172 25842 28224 25848
rect 28172 25764 28224 25770
rect 28172 25706 28224 25712
rect 28080 25288 28132 25294
rect 28080 25230 28132 25236
rect 28184 24818 28212 25706
rect 28172 24812 28224 24818
rect 28172 24754 28224 24760
rect 28276 24698 28304 25860
rect 28356 25492 28408 25498
rect 28356 25434 28408 25440
rect 28368 25294 28396 25434
rect 28356 25288 28408 25294
rect 28356 25230 28408 25236
rect 28356 25152 28408 25158
rect 28356 25094 28408 25100
rect 28448 25152 28500 25158
rect 28448 25094 28500 25100
rect 28368 24954 28396 25094
rect 28356 24948 28408 24954
rect 28356 24890 28408 24896
rect 28460 24886 28488 25094
rect 28448 24880 28500 24886
rect 28448 24822 28500 24828
rect 28092 24670 28304 24698
rect 28092 22030 28120 24670
rect 28448 24268 28500 24274
rect 28448 24210 28500 24216
rect 28356 24200 28408 24206
rect 28356 24142 28408 24148
rect 28172 24064 28224 24070
rect 28172 24006 28224 24012
rect 28080 22024 28132 22030
rect 28080 21966 28132 21972
rect 27896 21956 27948 21962
rect 27896 21898 27948 21904
rect 27988 21888 28040 21894
rect 27988 21830 28040 21836
rect 27896 21616 27948 21622
rect 27896 21558 27948 21564
rect 27528 21548 27580 21554
rect 27528 21490 27580 21496
rect 27436 21344 27488 21350
rect 27436 21286 27488 21292
rect 27436 20868 27488 20874
rect 27436 20810 27488 20816
rect 27264 20556 27384 20584
rect 27252 20460 27304 20466
rect 27252 20402 27304 20408
rect 27264 20058 27292 20402
rect 27252 20052 27304 20058
rect 27252 19994 27304 20000
rect 27356 19922 27384 20556
rect 27344 19916 27396 19922
rect 27344 19858 27396 19864
rect 27344 19372 27396 19378
rect 27344 19314 27396 19320
rect 27252 19304 27304 19310
rect 27252 19246 27304 19252
rect 27264 18902 27292 19246
rect 27356 19174 27384 19314
rect 27344 19168 27396 19174
rect 27344 19110 27396 19116
rect 27252 18896 27304 18902
rect 27252 18838 27304 18844
rect 27160 18760 27212 18766
rect 27212 18720 27292 18748
rect 27160 18702 27212 18708
rect 27264 18358 27292 18720
rect 27344 18624 27396 18630
rect 27344 18566 27396 18572
rect 27252 18352 27304 18358
rect 27252 18294 27304 18300
rect 27160 17672 27212 17678
rect 27160 17614 27212 17620
rect 27172 17202 27200 17614
rect 27160 17196 27212 17202
rect 27160 17138 27212 17144
rect 27160 16720 27212 16726
rect 27160 16662 27212 16668
rect 27172 16046 27200 16662
rect 27160 16040 27212 16046
rect 27160 15982 27212 15988
rect 27264 15162 27292 18294
rect 27356 18290 27384 18566
rect 27344 18284 27396 18290
rect 27344 18226 27396 18232
rect 27068 15156 27120 15162
rect 27068 15098 27120 15104
rect 27252 15156 27304 15162
rect 27252 15098 27304 15104
rect 27448 14550 27476 20810
rect 27540 20806 27568 21490
rect 27528 20800 27580 20806
rect 27528 20742 27580 20748
rect 27540 20534 27568 20742
rect 27528 20528 27580 20534
rect 27528 20470 27580 20476
rect 27908 19854 27936 21558
rect 27896 19848 27948 19854
rect 27896 19790 27948 19796
rect 27712 19712 27764 19718
rect 27710 19680 27712 19689
rect 27804 19712 27856 19718
rect 27764 19680 27766 19689
rect 27804 19654 27856 19660
rect 27710 19615 27766 19624
rect 27816 19378 27844 19654
rect 27804 19372 27856 19378
rect 27804 19314 27856 19320
rect 27712 19304 27764 19310
rect 27712 19246 27764 19252
rect 27724 18834 27752 19246
rect 27712 18828 27764 18834
rect 27712 18770 27764 18776
rect 27620 18760 27672 18766
rect 27620 18702 27672 18708
rect 27632 18222 27660 18702
rect 27712 18284 27764 18290
rect 27712 18226 27764 18232
rect 27620 18216 27672 18222
rect 27620 18158 27672 18164
rect 27724 16794 27752 18226
rect 27908 17542 27936 19790
rect 28000 18426 28028 21830
rect 28092 21622 28120 21966
rect 28080 21616 28132 21622
rect 28080 21558 28132 21564
rect 28184 20466 28212 24006
rect 28368 23526 28396 24142
rect 28460 24070 28488 24210
rect 28448 24064 28500 24070
rect 28448 24006 28500 24012
rect 28552 23798 28580 27066
rect 28736 27062 28764 27270
rect 28724 27056 28776 27062
rect 28724 26998 28776 27004
rect 28724 26240 28776 26246
rect 29012 26234 29040 27911
rect 29104 27538 29132 27950
rect 29092 27532 29144 27538
rect 29092 27474 29144 27480
rect 29196 27470 29224 28426
rect 29184 27464 29236 27470
rect 29184 27406 29236 27412
rect 29184 26920 29236 26926
rect 29184 26862 29236 26868
rect 29196 26586 29224 26862
rect 29184 26580 29236 26586
rect 29184 26522 29236 26528
rect 28724 26182 28776 26188
rect 28828 26206 29040 26234
rect 28736 25906 28764 26182
rect 28724 25900 28776 25906
rect 28724 25842 28776 25848
rect 28724 24268 28776 24274
rect 28724 24210 28776 24216
rect 28736 24138 28764 24210
rect 28724 24132 28776 24138
rect 28724 24074 28776 24080
rect 28540 23792 28592 23798
rect 28540 23734 28592 23740
rect 28448 23656 28500 23662
rect 28448 23598 28500 23604
rect 28356 23520 28408 23526
rect 28356 23462 28408 23468
rect 28264 23316 28316 23322
rect 28264 23258 28316 23264
rect 28276 21554 28304 23258
rect 28460 23118 28488 23598
rect 28448 23112 28500 23118
rect 28448 23054 28500 23060
rect 28356 23044 28408 23050
rect 28356 22986 28408 22992
rect 28368 22166 28396 22986
rect 28356 22160 28408 22166
rect 28356 22102 28408 22108
rect 28448 22092 28500 22098
rect 28448 22034 28500 22040
rect 28264 21548 28316 21554
rect 28264 21490 28316 21496
rect 28356 21004 28408 21010
rect 28356 20946 28408 20952
rect 28172 20460 28224 20466
rect 28172 20402 28224 20408
rect 28368 19242 28396 20946
rect 28356 19236 28408 19242
rect 28356 19178 28408 19184
rect 28368 18834 28396 19178
rect 28460 18970 28488 22034
rect 28552 20942 28580 23734
rect 28828 23662 28856 26206
rect 29092 25968 29144 25974
rect 29092 25910 29144 25916
rect 29001 25424 29053 25430
rect 28998 25392 29001 25401
rect 29053 25392 29054 25401
rect 28998 25327 29054 25336
rect 29104 24614 29132 25910
rect 29288 25498 29316 29407
rect 29380 27878 29408 30874
rect 29368 27872 29420 27878
rect 29368 27814 29420 27820
rect 29380 26994 29408 27814
rect 29472 27606 29500 31039
rect 29564 29850 29592 36722
rect 29656 36156 29684 37742
rect 29734 37360 29790 37369
rect 29734 37295 29790 37304
rect 29748 37126 29776 37295
rect 29736 37120 29788 37126
rect 29736 37062 29788 37068
rect 29656 36128 29776 36156
rect 29644 35216 29696 35222
rect 29644 35158 29696 35164
rect 29656 30938 29684 35158
rect 29748 34134 29776 36128
rect 29840 35222 29868 39374
rect 30196 39364 30248 39370
rect 30196 39306 30248 39312
rect 30012 37936 30064 37942
rect 30010 37904 30012 37913
rect 30104 37936 30156 37942
rect 30064 37904 30066 37913
rect 30104 37878 30156 37884
rect 30010 37839 30066 37848
rect 29918 37768 29974 37777
rect 29918 37703 29974 37712
rect 29932 37330 29960 37703
rect 30116 37466 30144 37878
rect 30104 37460 30156 37466
rect 30104 37402 30156 37408
rect 30010 37360 30066 37369
rect 29920 37324 29972 37330
rect 30010 37295 30066 37304
rect 29920 37266 29972 37272
rect 30024 37194 30052 37295
rect 30104 37256 30156 37262
rect 30104 37198 30156 37204
rect 30012 37188 30064 37194
rect 30012 37130 30064 37136
rect 30012 36848 30064 36854
rect 30012 36790 30064 36796
rect 29920 36576 29972 36582
rect 29920 36518 29972 36524
rect 29932 36417 29960 36518
rect 29918 36408 29974 36417
rect 29918 36343 29974 36352
rect 29920 36168 29972 36174
rect 29920 36110 29972 36116
rect 29932 35873 29960 36110
rect 29918 35864 29974 35873
rect 30024 35834 30052 36790
rect 29918 35799 29974 35808
rect 30012 35828 30064 35834
rect 30012 35770 30064 35776
rect 29920 35692 29972 35698
rect 29920 35634 29972 35640
rect 29828 35216 29880 35222
rect 29828 35158 29880 35164
rect 29932 35086 29960 35634
rect 30116 35136 30144 37198
rect 30208 36378 30236 39306
rect 30380 39296 30432 39302
rect 30380 39238 30432 39244
rect 30288 38276 30340 38282
rect 30288 38218 30340 38224
rect 30300 38010 30328 38218
rect 30288 38004 30340 38010
rect 30288 37946 30340 37952
rect 30288 37256 30340 37262
rect 30288 37198 30340 37204
rect 30300 36582 30328 37198
rect 30288 36576 30340 36582
rect 30288 36518 30340 36524
rect 30196 36372 30248 36378
rect 30196 36314 30248 36320
rect 30300 36310 30328 36518
rect 30288 36304 30340 36310
rect 30288 36246 30340 36252
rect 30196 36100 30248 36106
rect 30196 36042 30248 36048
rect 30208 35698 30236 36042
rect 30196 35692 30248 35698
rect 30196 35634 30248 35640
rect 30392 35272 30420 39238
rect 30576 38894 30604 39374
rect 30932 39296 30984 39302
rect 30932 39238 30984 39244
rect 30564 38888 30616 38894
rect 30564 38830 30616 38836
rect 30493 38652 30801 38661
rect 30493 38650 30499 38652
rect 30555 38650 30579 38652
rect 30635 38650 30659 38652
rect 30715 38650 30739 38652
rect 30795 38650 30801 38652
rect 30555 38598 30557 38650
rect 30737 38598 30739 38650
rect 30493 38596 30499 38598
rect 30555 38596 30579 38598
rect 30635 38596 30659 38598
rect 30715 38596 30739 38598
rect 30795 38596 30801 38598
rect 30493 38587 30801 38596
rect 30944 37806 30972 39238
rect 31208 38208 31260 38214
rect 31208 38150 31260 38156
rect 30932 37800 30984 37806
rect 30932 37742 30984 37748
rect 30493 37564 30801 37573
rect 30493 37562 30499 37564
rect 30555 37562 30579 37564
rect 30635 37562 30659 37564
rect 30715 37562 30739 37564
rect 30795 37562 30801 37564
rect 30555 37510 30557 37562
rect 30737 37510 30739 37562
rect 30493 37508 30499 37510
rect 30555 37508 30579 37510
rect 30635 37508 30659 37510
rect 30715 37508 30739 37510
rect 30795 37508 30801 37510
rect 30493 37499 30801 37508
rect 30748 37324 30800 37330
rect 30800 37272 30880 37274
rect 30748 37266 30880 37272
rect 30760 37246 30880 37266
rect 30564 37120 30616 37126
rect 30564 37062 30616 37068
rect 30576 36854 30604 37062
rect 30564 36848 30616 36854
rect 30564 36790 30616 36796
rect 30852 36718 30880 37246
rect 31022 37224 31078 37233
rect 31022 37159 31078 37168
rect 31116 37188 31168 37194
rect 30932 37120 30984 37126
rect 30930 37088 30932 37097
rect 30984 37088 30986 37097
rect 30930 37023 30986 37032
rect 30840 36712 30892 36718
rect 30840 36654 30892 36660
rect 30493 36476 30801 36485
rect 30493 36474 30499 36476
rect 30555 36474 30579 36476
rect 30635 36474 30659 36476
rect 30715 36474 30739 36476
rect 30795 36474 30801 36476
rect 30555 36422 30557 36474
rect 30737 36422 30739 36474
rect 30493 36420 30499 36422
rect 30555 36420 30579 36422
rect 30635 36420 30659 36422
rect 30715 36420 30739 36422
rect 30795 36420 30801 36422
rect 30493 36411 30801 36420
rect 30852 36310 30880 36654
rect 30932 36644 30984 36650
rect 30932 36586 30984 36592
rect 30840 36304 30892 36310
rect 30840 36246 30892 36252
rect 30852 35562 30880 36246
rect 30944 36145 30972 36586
rect 31036 36378 31064 37159
rect 31116 37130 31168 37136
rect 31128 36417 31156 37130
rect 31220 36854 31248 38150
rect 31312 37233 31340 39510
rect 32218 39471 32274 39480
rect 31852 38888 31904 38894
rect 31852 38830 31904 38836
rect 31576 37868 31628 37874
rect 31576 37810 31628 37816
rect 31392 37800 31444 37806
rect 31392 37742 31444 37748
rect 31298 37224 31354 37233
rect 31298 37159 31354 37168
rect 31208 36848 31260 36854
rect 31208 36790 31260 36796
rect 31114 36408 31170 36417
rect 31024 36372 31076 36378
rect 31114 36343 31170 36352
rect 31024 36314 31076 36320
rect 31116 36236 31168 36242
rect 31116 36178 31168 36184
rect 30930 36136 30986 36145
rect 30930 36071 30986 36080
rect 31024 35624 31076 35630
rect 31024 35566 31076 35572
rect 30840 35556 30892 35562
rect 30840 35498 30892 35504
rect 30932 35488 30984 35494
rect 30930 35456 30932 35465
rect 30984 35456 30986 35465
rect 30493 35388 30801 35397
rect 30930 35391 30986 35400
rect 30493 35386 30499 35388
rect 30555 35386 30579 35388
rect 30635 35386 30659 35388
rect 30715 35386 30739 35388
rect 30795 35386 30801 35388
rect 30555 35334 30557 35386
rect 30737 35334 30739 35386
rect 30493 35332 30499 35334
rect 30555 35332 30579 35334
rect 30635 35332 30659 35334
rect 30715 35332 30739 35334
rect 30795 35332 30801 35334
rect 30493 35323 30801 35332
rect 30392 35244 30604 35272
rect 30116 35108 30328 35136
rect 29828 35080 29880 35086
rect 29828 35022 29880 35028
rect 29920 35080 29972 35086
rect 29920 35022 29972 35028
rect 29840 34746 29868 35022
rect 30104 35012 30156 35018
rect 30104 34954 30156 34960
rect 29828 34740 29880 34746
rect 29828 34682 29880 34688
rect 30116 34678 30144 34954
rect 29920 34672 29972 34678
rect 29920 34614 29972 34620
rect 30104 34672 30156 34678
rect 30104 34614 30156 34620
rect 29828 34400 29880 34406
rect 29828 34342 29880 34348
rect 29736 34128 29788 34134
rect 29736 34070 29788 34076
rect 29736 33992 29788 33998
rect 29736 33934 29788 33940
rect 29748 33590 29776 33934
rect 29736 33584 29788 33590
rect 29736 33526 29788 33532
rect 29748 32298 29776 33526
rect 29840 33318 29868 34342
rect 29932 33454 29960 34614
rect 30012 34604 30064 34610
rect 30012 34546 30064 34552
rect 29920 33448 29972 33454
rect 29920 33390 29972 33396
rect 29828 33312 29880 33318
rect 29828 33254 29880 33260
rect 29932 33046 29960 33390
rect 29828 33040 29880 33046
rect 29828 32982 29880 32988
rect 29920 33040 29972 33046
rect 29920 32982 29972 32988
rect 29840 32774 29868 32982
rect 29920 32904 29972 32910
rect 30024 32892 30052 34546
rect 30194 34504 30250 34513
rect 30194 34439 30250 34448
rect 30104 34400 30156 34406
rect 30104 34342 30156 34348
rect 30116 34202 30144 34342
rect 30104 34196 30156 34202
rect 30104 34138 30156 34144
rect 30104 33924 30156 33930
rect 30104 33866 30156 33872
rect 29972 32864 30052 32892
rect 29920 32846 29972 32852
rect 29828 32768 29880 32774
rect 29828 32710 29880 32716
rect 29828 32428 29880 32434
rect 29828 32370 29880 32376
rect 29736 32292 29788 32298
rect 29736 32234 29788 32240
rect 29748 31634 29776 32234
rect 29840 32026 29868 32370
rect 30116 32026 30144 33866
rect 30208 32570 30236 34439
rect 30196 32564 30248 32570
rect 30196 32506 30248 32512
rect 29828 32020 29880 32026
rect 29828 31962 29880 31968
rect 30104 32020 30156 32026
rect 30104 31962 30156 31968
rect 29748 31606 29868 31634
rect 29734 31512 29790 31521
rect 29734 31447 29790 31456
rect 29644 30932 29696 30938
rect 29644 30874 29696 30880
rect 29552 29844 29604 29850
rect 29552 29786 29604 29792
rect 29564 29034 29592 29786
rect 29644 29640 29696 29646
rect 29642 29608 29644 29617
rect 29696 29608 29698 29617
rect 29642 29543 29698 29552
rect 29748 29492 29776 31447
rect 29840 31414 29868 31606
rect 29828 31408 29880 31414
rect 29828 31350 29880 31356
rect 30300 31124 30328 35108
rect 30576 34678 30604 35244
rect 30564 34672 30616 34678
rect 30564 34614 30616 34620
rect 30493 34300 30801 34309
rect 30493 34298 30499 34300
rect 30555 34298 30579 34300
rect 30635 34298 30659 34300
rect 30715 34298 30739 34300
rect 30795 34298 30801 34300
rect 30555 34246 30557 34298
rect 30737 34246 30739 34298
rect 30493 34244 30499 34246
rect 30555 34244 30579 34246
rect 30635 34244 30659 34246
rect 30715 34244 30739 34246
rect 30795 34244 30801 34246
rect 30493 34235 30801 34244
rect 30932 33992 30984 33998
rect 30932 33934 30984 33940
rect 30840 33924 30892 33930
rect 30840 33866 30892 33872
rect 30564 33856 30616 33862
rect 30564 33798 30616 33804
rect 30576 33590 30604 33798
rect 30564 33584 30616 33590
rect 30564 33526 30616 33532
rect 30493 33212 30801 33221
rect 30493 33210 30499 33212
rect 30555 33210 30579 33212
rect 30635 33210 30659 33212
rect 30715 33210 30739 33212
rect 30795 33210 30801 33212
rect 30555 33158 30557 33210
rect 30737 33158 30739 33210
rect 30493 33156 30499 33158
rect 30555 33156 30579 33158
rect 30635 33156 30659 33158
rect 30715 33156 30739 33158
rect 30795 33156 30801 33158
rect 30493 33147 30801 33156
rect 30748 32904 30800 32910
rect 30852 32892 30880 33866
rect 30800 32864 30880 32892
rect 30748 32846 30800 32852
rect 30944 32774 30972 33934
rect 30932 32768 30984 32774
rect 30932 32710 30984 32716
rect 30840 32360 30892 32366
rect 30840 32302 30892 32308
rect 30493 32124 30801 32133
rect 30493 32122 30499 32124
rect 30555 32122 30579 32124
rect 30635 32122 30659 32124
rect 30715 32122 30739 32124
rect 30795 32122 30801 32124
rect 30555 32070 30557 32122
rect 30737 32070 30739 32122
rect 30493 32068 30499 32070
rect 30555 32068 30579 32070
rect 30635 32068 30659 32070
rect 30715 32068 30739 32070
rect 30795 32068 30801 32070
rect 30493 32059 30801 32068
rect 30656 32020 30708 32026
rect 30656 31962 30708 31968
rect 30668 31822 30696 31962
rect 30656 31816 30708 31822
rect 30656 31758 30708 31764
rect 30852 31736 30880 32302
rect 30760 31708 30880 31736
rect 30930 31784 30986 31793
rect 31036 31754 31064 35566
rect 31128 34202 31156 36178
rect 31298 35864 31354 35873
rect 31298 35799 31354 35808
rect 31312 34746 31340 35799
rect 31208 34740 31260 34746
rect 31208 34682 31260 34688
rect 31300 34740 31352 34746
rect 31300 34682 31352 34688
rect 31116 34196 31168 34202
rect 31116 34138 31168 34144
rect 31128 33998 31156 34138
rect 31116 33992 31168 33998
rect 31116 33934 31168 33940
rect 31116 32768 31168 32774
rect 31116 32710 31168 32716
rect 31128 31890 31156 32710
rect 31220 32230 31248 34682
rect 31300 34060 31352 34066
rect 31300 34002 31352 34008
rect 31312 33658 31340 34002
rect 31300 33652 31352 33658
rect 31300 33594 31352 33600
rect 31312 32910 31340 33594
rect 31300 32904 31352 32910
rect 31300 32846 31352 32852
rect 31298 32600 31354 32609
rect 31298 32535 31354 32544
rect 31312 32502 31340 32535
rect 31404 32502 31432 37742
rect 31484 37324 31536 37330
rect 31484 37266 31536 37272
rect 31496 32774 31524 37266
rect 31588 37262 31616 37810
rect 31576 37256 31628 37262
rect 31576 37198 31628 37204
rect 31588 36174 31616 37198
rect 31864 36394 31892 38830
rect 32232 38350 32260 39471
rect 32220 38344 32272 38350
rect 32220 38286 32272 38292
rect 32218 37904 32274 37913
rect 32218 37839 32274 37848
rect 32126 37768 32182 37777
rect 32126 37703 32182 37712
rect 31942 37496 31998 37505
rect 31942 37431 31998 37440
rect 31956 36718 31984 37431
rect 32036 37120 32088 37126
rect 32036 37062 32088 37068
rect 32048 36825 32076 37062
rect 32034 36816 32090 36825
rect 32034 36751 32090 36760
rect 31944 36712 31996 36718
rect 31944 36654 31996 36660
rect 31772 36378 31892 36394
rect 31760 36372 31892 36378
rect 31812 36366 31892 36372
rect 31760 36314 31812 36320
rect 31576 36168 31628 36174
rect 31576 36110 31628 36116
rect 32036 36100 32088 36106
rect 32036 36042 32088 36048
rect 31944 35760 31996 35766
rect 31758 35728 31814 35737
rect 31668 35692 31720 35698
rect 31588 35652 31668 35680
rect 31588 34406 31616 35652
rect 31944 35702 31996 35708
rect 31758 35663 31760 35672
rect 31668 35634 31720 35640
rect 31812 35663 31814 35672
rect 31760 35634 31812 35640
rect 31852 35624 31904 35630
rect 31852 35566 31904 35572
rect 31760 35488 31812 35494
rect 31758 35456 31760 35465
rect 31812 35456 31814 35465
rect 31758 35391 31814 35400
rect 31668 34944 31720 34950
rect 31668 34886 31720 34892
rect 31576 34400 31628 34406
rect 31576 34342 31628 34348
rect 31576 34128 31628 34134
rect 31680 34116 31708 34886
rect 31760 34740 31812 34746
rect 31760 34682 31812 34688
rect 31628 34088 31708 34116
rect 31576 34070 31628 34076
rect 31588 32842 31616 34070
rect 31772 34066 31800 34682
rect 31760 34060 31812 34066
rect 31760 34002 31812 34008
rect 31864 33946 31892 35566
rect 31772 33918 31892 33946
rect 31666 33688 31722 33697
rect 31666 33623 31722 33632
rect 31576 32836 31628 32842
rect 31576 32778 31628 32784
rect 31484 32768 31536 32774
rect 31484 32710 31536 32716
rect 31300 32496 31352 32502
rect 31300 32438 31352 32444
rect 31392 32496 31444 32502
rect 31392 32438 31444 32444
rect 31496 32434 31524 32710
rect 31680 32570 31708 33623
rect 31772 32570 31800 33918
rect 31956 33862 31984 35702
rect 32048 34950 32076 36042
rect 32140 35086 32168 37703
rect 32232 36378 32260 37839
rect 32310 36952 32366 36961
rect 32310 36887 32366 36896
rect 32220 36372 32272 36378
rect 32220 36314 32272 36320
rect 32218 36136 32274 36145
rect 32218 36071 32274 36080
rect 32128 35080 32180 35086
rect 32128 35022 32180 35028
rect 32036 34944 32088 34950
rect 32036 34886 32088 34892
rect 32034 34096 32090 34105
rect 32034 34031 32036 34040
rect 32088 34031 32090 34040
rect 32036 34002 32088 34008
rect 32128 33924 32180 33930
rect 32128 33866 32180 33872
rect 31944 33856 31996 33862
rect 31944 33798 31996 33804
rect 32140 33590 32168 33866
rect 32128 33584 32180 33590
rect 31850 33552 31906 33561
rect 32128 33526 32180 33532
rect 31850 33487 31906 33496
rect 31576 32564 31628 32570
rect 31576 32506 31628 32512
rect 31668 32564 31720 32570
rect 31668 32506 31720 32512
rect 31760 32564 31812 32570
rect 31760 32506 31812 32512
rect 31484 32428 31536 32434
rect 31484 32370 31536 32376
rect 31208 32224 31260 32230
rect 31208 32166 31260 32172
rect 31392 32224 31444 32230
rect 31392 32166 31444 32172
rect 31300 31952 31352 31958
rect 31300 31894 31352 31900
rect 31116 31884 31168 31890
rect 31116 31826 31168 31832
rect 31208 31794 31260 31800
rect 30930 31719 30932 31728
rect 30760 31278 30788 31708
rect 30984 31719 30986 31728
rect 31024 31748 31076 31754
rect 30932 31690 30984 31696
rect 31208 31736 31260 31742
rect 31024 31690 31076 31696
rect 31220 31482 31248 31736
rect 31208 31476 31260 31482
rect 31208 31418 31260 31424
rect 30748 31272 30800 31278
rect 30748 31214 30800 31220
rect 30380 31136 30432 31142
rect 30300 31096 30380 31124
rect 30380 31078 30432 31084
rect 30932 31136 30984 31142
rect 30932 31078 30984 31084
rect 30493 31036 30801 31045
rect 30493 31034 30499 31036
rect 30555 31034 30579 31036
rect 30635 31034 30659 31036
rect 30715 31034 30739 31036
rect 30795 31034 30801 31036
rect 30555 30982 30557 31034
rect 30737 30982 30739 31034
rect 30493 30980 30499 30982
rect 30555 30980 30579 30982
rect 30635 30980 30659 30982
rect 30715 30980 30739 30982
rect 30795 30980 30801 30982
rect 30493 30971 30801 30980
rect 30748 30796 30800 30802
rect 30748 30738 30800 30744
rect 30760 30598 30788 30738
rect 30944 30734 30972 31078
rect 31312 30818 31340 31894
rect 31404 31346 31432 32166
rect 31496 31414 31524 32370
rect 31588 31890 31616 32506
rect 31760 32020 31812 32026
rect 31760 31962 31812 31968
rect 31576 31884 31628 31890
rect 31576 31826 31628 31832
rect 31588 31482 31616 31826
rect 31668 31816 31720 31822
rect 31668 31758 31720 31764
rect 31576 31476 31628 31482
rect 31576 31418 31628 31424
rect 31484 31408 31536 31414
rect 31484 31350 31536 31356
rect 31392 31340 31444 31346
rect 31392 31282 31444 31288
rect 31220 30790 31340 30818
rect 30932 30728 30984 30734
rect 30932 30670 30984 30676
rect 31022 30696 31078 30705
rect 31022 30631 31024 30640
rect 31076 30631 31078 30640
rect 31024 30602 31076 30608
rect 30748 30592 30800 30598
rect 30748 30534 30800 30540
rect 30380 30388 30432 30394
rect 30380 30330 30432 30336
rect 30472 30388 30524 30394
rect 30472 30330 30524 30336
rect 30012 30252 30064 30258
rect 30012 30194 30064 30200
rect 29920 30184 29972 30190
rect 29920 30126 29972 30132
rect 29656 29464 29776 29492
rect 29552 29028 29604 29034
rect 29552 28970 29604 28976
rect 29656 28490 29684 29464
rect 29736 28960 29788 28966
rect 29736 28902 29788 28908
rect 29748 28558 29776 28902
rect 29736 28552 29788 28558
rect 29736 28494 29788 28500
rect 29828 28552 29880 28558
rect 29932 28540 29960 30126
rect 30024 28608 30052 30194
rect 30104 29708 30156 29714
rect 30104 29650 30156 29656
rect 30116 29102 30144 29650
rect 30392 29646 30420 30330
rect 30484 30190 30512 30330
rect 30472 30184 30524 30190
rect 30472 30126 30524 30132
rect 30932 30184 30984 30190
rect 30932 30126 30984 30132
rect 30493 29948 30801 29957
rect 30493 29946 30499 29948
rect 30555 29946 30579 29948
rect 30635 29946 30659 29948
rect 30715 29946 30739 29948
rect 30795 29946 30801 29948
rect 30555 29894 30557 29946
rect 30737 29894 30739 29946
rect 30493 29892 30499 29894
rect 30555 29892 30579 29894
rect 30635 29892 30659 29894
rect 30715 29892 30739 29894
rect 30795 29892 30801 29894
rect 30493 29883 30801 29892
rect 30380 29640 30432 29646
rect 30380 29582 30432 29588
rect 30838 29608 30894 29617
rect 30196 29572 30248 29578
rect 30838 29543 30894 29552
rect 30196 29514 30248 29520
rect 30104 29096 30156 29102
rect 30104 29038 30156 29044
rect 30208 28966 30236 29514
rect 30748 29504 30800 29510
rect 30748 29446 30800 29452
rect 30760 29306 30788 29446
rect 30748 29300 30800 29306
rect 30748 29242 30800 29248
rect 30852 29170 30880 29543
rect 30944 29209 30972 30126
rect 31220 29594 31248 30790
rect 31300 30728 31352 30734
rect 31300 30670 31352 30676
rect 31312 30002 31340 30670
rect 31404 30122 31432 31282
rect 31484 31272 31536 31278
rect 31484 31214 31536 31220
rect 31496 30938 31524 31214
rect 31484 30932 31536 30938
rect 31484 30874 31536 30880
rect 31680 30394 31708 31758
rect 31772 31482 31800 31962
rect 31760 31476 31812 31482
rect 31760 31418 31812 31424
rect 31864 31414 31892 33487
rect 32232 31890 32260 36071
rect 32324 33590 32352 36887
rect 32312 33584 32364 33590
rect 32312 33526 32364 33532
rect 32312 32292 32364 32298
rect 32312 32234 32364 32240
rect 32324 31890 32352 32234
rect 32220 31884 32272 31890
rect 32220 31826 32272 31832
rect 32312 31884 32364 31890
rect 32312 31826 32364 31832
rect 32232 31521 32260 31826
rect 32218 31512 32274 31521
rect 32218 31447 32274 31456
rect 31852 31408 31904 31414
rect 31852 31350 31904 31356
rect 32324 30938 32352 31826
rect 32416 31686 32444 39578
rect 32508 39438 32536 39986
rect 32588 39840 32640 39846
rect 32588 39782 32640 39788
rect 32496 39432 32548 39438
rect 32496 39374 32548 39380
rect 32600 39030 32628 39782
rect 32588 39024 32640 39030
rect 32588 38966 32640 38972
rect 32876 38894 32904 41200
rect 33046 40896 33102 40905
rect 33046 40831 33102 40840
rect 32864 38888 32916 38894
rect 32864 38830 32916 38836
rect 32772 38752 32824 38758
rect 32772 38694 32824 38700
rect 32784 38654 32812 38694
rect 32784 38626 32904 38654
rect 32496 37800 32548 37806
rect 32496 37742 32548 37748
rect 32508 37398 32536 37742
rect 32588 37732 32640 37738
rect 32588 37674 32640 37680
rect 32496 37392 32548 37398
rect 32496 37334 32548 37340
rect 32496 37256 32548 37262
rect 32496 37198 32548 37204
rect 32508 36689 32536 37198
rect 32494 36680 32550 36689
rect 32494 36615 32550 36624
rect 32494 35184 32550 35193
rect 32494 35119 32550 35128
rect 32508 34610 32536 35119
rect 32496 34604 32548 34610
rect 32496 34546 32548 34552
rect 32600 34490 32628 37674
rect 32680 37188 32732 37194
rect 32680 37130 32732 37136
rect 32692 36922 32720 37130
rect 32680 36916 32732 36922
rect 32680 36858 32732 36864
rect 32876 35630 32904 38626
rect 33060 37330 33088 40831
rect 33048 37324 33100 37330
rect 33048 37266 33100 37272
rect 33520 36718 33548 41200
rect 34164 38418 34192 41200
rect 34336 39364 34388 39370
rect 34336 39306 34388 39312
rect 34348 38865 34376 39306
rect 34713 39196 35021 39205
rect 34713 39194 34719 39196
rect 34775 39194 34799 39196
rect 34855 39194 34879 39196
rect 34935 39194 34959 39196
rect 35015 39194 35021 39196
rect 34775 39142 34777 39194
rect 34957 39142 34959 39194
rect 34713 39140 34719 39142
rect 34775 39140 34799 39142
rect 34855 39140 34879 39142
rect 34935 39140 34959 39142
rect 35015 39140 35021 39142
rect 34713 39131 35021 39140
rect 34334 38856 34390 38865
rect 34334 38791 34390 38800
rect 34152 38412 34204 38418
rect 34152 38354 34204 38360
rect 34713 38108 35021 38117
rect 34713 38106 34719 38108
rect 34775 38106 34799 38108
rect 34855 38106 34879 38108
rect 34935 38106 34959 38108
rect 35015 38106 35021 38108
rect 34775 38054 34777 38106
rect 34957 38054 34959 38106
rect 34713 38052 34719 38054
rect 34775 38052 34799 38054
rect 34855 38052 34879 38054
rect 34935 38052 34959 38054
rect 35015 38052 35021 38054
rect 34713 38043 35021 38052
rect 34336 37936 34388 37942
rect 34334 37904 34336 37913
rect 34388 37904 34390 37913
rect 34334 37839 34390 37848
rect 34060 37460 34112 37466
rect 34060 37402 34112 37408
rect 33508 36712 33560 36718
rect 33508 36654 33560 36660
rect 32956 36576 33008 36582
rect 32956 36518 33008 36524
rect 32968 35698 32996 36518
rect 34072 35766 34100 37402
rect 34713 37020 35021 37029
rect 34713 37018 34719 37020
rect 34775 37018 34799 37020
rect 34855 37018 34879 37020
rect 34935 37018 34959 37020
rect 35015 37018 35021 37020
rect 34775 36966 34777 37018
rect 34957 36966 34959 37018
rect 34713 36964 34719 36966
rect 34775 36964 34799 36966
rect 34855 36964 34879 36966
rect 34935 36964 34959 36966
rect 35015 36964 35021 36966
rect 34713 36955 35021 36964
rect 34334 36816 34390 36825
rect 34334 36751 34390 36760
rect 34348 36242 34376 36751
rect 34336 36236 34388 36242
rect 34336 36178 34388 36184
rect 34713 35932 35021 35941
rect 34713 35930 34719 35932
rect 34775 35930 34799 35932
rect 34855 35930 34879 35932
rect 34935 35930 34959 35932
rect 35015 35930 35021 35932
rect 34775 35878 34777 35930
rect 34957 35878 34959 35930
rect 34713 35876 34719 35878
rect 34775 35876 34799 35878
rect 34855 35876 34879 35878
rect 34935 35876 34959 35878
rect 35015 35876 35021 35878
rect 34713 35867 35021 35876
rect 34060 35760 34112 35766
rect 34060 35702 34112 35708
rect 32956 35692 33008 35698
rect 32956 35634 33008 35640
rect 32864 35624 32916 35630
rect 32864 35566 32916 35572
rect 32772 35488 32824 35494
rect 32770 35456 32772 35465
rect 32824 35456 32826 35465
rect 32770 35391 32826 35400
rect 32508 34462 32628 34490
rect 32404 31680 32456 31686
rect 32404 31622 32456 31628
rect 32312 30932 32364 30938
rect 32312 30874 32364 30880
rect 31760 30796 31812 30802
rect 31760 30738 31812 30744
rect 32036 30796 32088 30802
rect 32036 30738 32088 30744
rect 31668 30388 31720 30394
rect 31668 30330 31720 30336
rect 31576 30320 31628 30326
rect 31576 30262 31628 30268
rect 31392 30116 31444 30122
rect 31392 30058 31444 30064
rect 31484 30048 31536 30054
rect 31312 29974 31432 30002
rect 31484 29990 31536 29996
rect 31036 29566 31248 29594
rect 30930 29200 30986 29209
rect 30840 29164 30892 29170
rect 30930 29135 30986 29144
rect 30840 29106 30892 29112
rect 30288 29028 30340 29034
rect 30288 28970 30340 28976
rect 30196 28960 30248 28966
rect 30196 28902 30248 28908
rect 30024 28580 30144 28608
rect 29880 28512 29960 28540
rect 29828 28494 29880 28500
rect 29644 28484 29696 28490
rect 29644 28426 29696 28432
rect 29552 28416 29604 28422
rect 29552 28358 29604 28364
rect 29564 27878 29592 28358
rect 29642 28248 29698 28257
rect 29642 28183 29698 28192
rect 29656 28150 29684 28183
rect 29644 28144 29696 28150
rect 29644 28086 29696 28092
rect 29644 28008 29696 28014
rect 29644 27950 29696 27956
rect 29552 27872 29604 27878
rect 29552 27814 29604 27820
rect 29656 27713 29684 27950
rect 29642 27704 29698 27713
rect 29642 27639 29698 27648
rect 29460 27600 29512 27606
rect 29460 27542 29512 27548
rect 29460 27328 29512 27334
rect 29656 27316 29684 27639
rect 29748 27606 29776 28494
rect 29828 28416 29880 28422
rect 29828 28358 29880 28364
rect 29840 28082 29868 28358
rect 29828 28076 29880 28082
rect 29828 28018 29880 28024
rect 29736 27600 29788 27606
rect 29736 27542 29788 27548
rect 29460 27270 29512 27276
rect 29564 27288 29684 27316
rect 29368 26988 29420 26994
rect 29368 26930 29420 26936
rect 29368 26784 29420 26790
rect 29368 26726 29420 26732
rect 29380 25906 29408 26726
rect 29368 25900 29420 25906
rect 29368 25842 29420 25848
rect 29276 25492 29328 25498
rect 29276 25434 29328 25440
rect 29092 24608 29144 24614
rect 29092 24550 29144 24556
rect 29000 23724 29052 23730
rect 29000 23666 29052 23672
rect 28816 23656 28868 23662
rect 28816 23598 28868 23604
rect 28632 23588 28684 23594
rect 28632 23530 28684 23536
rect 28644 22982 28672 23530
rect 28908 23520 28960 23526
rect 28908 23462 28960 23468
rect 28816 23180 28868 23186
rect 28816 23122 28868 23128
rect 28828 23089 28856 23122
rect 28814 23080 28870 23089
rect 28814 23015 28870 23024
rect 28632 22976 28684 22982
rect 28632 22918 28684 22924
rect 28644 22012 28672 22918
rect 28920 22642 28948 23462
rect 29012 23118 29040 23666
rect 29104 23662 29132 24550
rect 29092 23656 29144 23662
rect 29092 23598 29144 23604
rect 29104 23322 29132 23598
rect 29092 23316 29144 23322
rect 29092 23258 29144 23264
rect 29368 23248 29420 23254
rect 29368 23190 29420 23196
rect 29000 23112 29052 23118
rect 29000 23054 29052 23060
rect 29184 22976 29236 22982
rect 29184 22918 29236 22924
rect 28998 22808 29054 22817
rect 28998 22743 29054 22752
rect 29012 22710 29040 22743
rect 29000 22704 29052 22710
rect 29000 22646 29052 22652
rect 28908 22636 28960 22642
rect 28908 22578 28960 22584
rect 28724 22432 28776 22438
rect 28724 22374 28776 22380
rect 28736 22273 28764 22374
rect 28722 22264 28778 22273
rect 28722 22199 28778 22208
rect 28816 22228 28868 22234
rect 28816 22170 28868 22176
rect 28644 21984 28764 22012
rect 28736 21010 28764 21984
rect 28724 21004 28776 21010
rect 28724 20946 28776 20952
rect 28540 20936 28592 20942
rect 28540 20878 28592 20884
rect 28828 20482 28856 22170
rect 28920 21554 28948 22578
rect 29196 22030 29224 22918
rect 29276 22704 29328 22710
rect 29276 22646 29328 22652
rect 29184 22024 29236 22030
rect 29184 21966 29236 21972
rect 29000 21888 29052 21894
rect 28998 21856 29000 21865
rect 29052 21856 29054 21865
rect 28998 21791 29054 21800
rect 29288 21622 29316 22646
rect 29276 21616 29328 21622
rect 29276 21558 29328 21564
rect 28908 21548 28960 21554
rect 28908 21490 28960 21496
rect 29288 21078 29316 21558
rect 29276 21072 29328 21078
rect 29276 21014 29328 21020
rect 29000 21004 29052 21010
rect 29000 20946 29052 20952
rect 28736 20454 28856 20482
rect 29012 20466 29040 20946
rect 29092 20936 29144 20942
rect 29092 20878 29144 20884
rect 28908 20460 28960 20466
rect 28736 20448 28764 20454
rect 28552 20420 28764 20448
rect 28448 18964 28500 18970
rect 28448 18906 28500 18912
rect 28356 18828 28408 18834
rect 28356 18770 28408 18776
rect 28264 18760 28316 18766
rect 28262 18728 28264 18737
rect 28316 18728 28318 18737
rect 28262 18663 28318 18672
rect 28368 18630 28396 18770
rect 28552 18698 28580 20420
rect 28908 20402 28960 20408
rect 29000 20460 29052 20466
rect 29000 20402 29052 20408
rect 28816 20392 28868 20398
rect 28816 20334 28868 20340
rect 28724 20324 28776 20330
rect 28724 20266 28776 20272
rect 28632 20256 28684 20262
rect 28632 20198 28684 20204
rect 28540 18692 28592 18698
rect 28540 18634 28592 18640
rect 28356 18624 28408 18630
rect 28184 18584 28356 18612
rect 27988 18420 28040 18426
rect 27988 18362 28040 18368
rect 28080 18284 28132 18290
rect 28080 18226 28132 18232
rect 27896 17536 27948 17542
rect 27896 17478 27948 17484
rect 27804 16992 27856 16998
rect 27804 16934 27856 16940
rect 27712 16788 27764 16794
rect 27712 16730 27764 16736
rect 27816 16590 27844 16934
rect 27804 16584 27856 16590
rect 27804 16526 27856 16532
rect 27816 15434 27844 16526
rect 27804 15428 27856 15434
rect 27804 15370 27856 15376
rect 27816 15026 27844 15370
rect 28092 15162 28120 18226
rect 28184 16658 28212 18584
rect 28356 18566 28408 18572
rect 28356 18284 28408 18290
rect 28356 18226 28408 18232
rect 28264 18216 28316 18222
rect 28264 18158 28316 18164
rect 28276 18086 28304 18158
rect 28264 18080 28316 18086
rect 28264 18022 28316 18028
rect 28276 17610 28304 18022
rect 28368 17882 28396 18226
rect 28448 18216 28500 18222
rect 28448 18158 28500 18164
rect 28460 17882 28488 18158
rect 28356 17876 28408 17882
rect 28356 17818 28408 17824
rect 28448 17876 28500 17882
rect 28448 17818 28500 17824
rect 28460 17678 28488 17818
rect 28448 17672 28500 17678
rect 28448 17614 28500 17620
rect 28264 17604 28316 17610
rect 28264 17546 28316 17552
rect 28172 16652 28224 16658
rect 28172 16594 28224 16600
rect 28184 16114 28212 16594
rect 28276 16182 28304 17546
rect 28448 17264 28500 17270
rect 28448 17206 28500 17212
rect 28460 16794 28488 17206
rect 28448 16788 28500 16794
rect 28448 16730 28500 16736
rect 28460 16590 28488 16730
rect 28448 16584 28500 16590
rect 28448 16526 28500 16532
rect 28552 16454 28580 18634
rect 28540 16448 28592 16454
rect 28540 16390 28592 16396
rect 28264 16176 28316 16182
rect 28264 16118 28316 16124
rect 28172 16108 28224 16114
rect 28172 16050 28224 16056
rect 28356 16108 28408 16114
rect 28356 16050 28408 16056
rect 28080 15156 28132 15162
rect 28080 15098 28132 15104
rect 28184 15026 28212 16050
rect 28368 15366 28396 16050
rect 28644 16046 28672 20198
rect 28736 19310 28764 20266
rect 28828 19786 28856 20334
rect 28920 20330 28948 20402
rect 28908 20324 28960 20330
rect 28908 20266 28960 20272
rect 28920 19786 28948 20266
rect 28816 19780 28868 19786
rect 28816 19722 28868 19728
rect 28908 19780 28960 19786
rect 28908 19722 28960 19728
rect 28724 19304 28776 19310
rect 28724 19246 28776 19252
rect 28736 18902 28764 19246
rect 28724 18896 28776 18902
rect 28724 18838 28776 18844
rect 28828 18834 28856 19722
rect 28816 18828 28868 18834
rect 28816 18770 28868 18776
rect 28920 18714 28948 19722
rect 29104 19718 29132 20878
rect 29380 20516 29408 23190
rect 29472 21146 29500 27270
rect 29564 26926 29592 27288
rect 29644 26988 29696 26994
rect 29644 26930 29696 26936
rect 29552 26920 29604 26926
rect 29552 26862 29604 26868
rect 29564 26246 29592 26862
rect 29656 26790 29684 26930
rect 29644 26784 29696 26790
rect 29644 26726 29696 26732
rect 29644 26512 29696 26518
rect 29644 26454 29696 26460
rect 29552 26240 29604 26246
rect 29552 26182 29604 26188
rect 29656 25158 29684 26454
rect 29748 26450 29776 27542
rect 29932 27538 29960 28512
rect 30012 28484 30064 28490
rect 30012 28426 30064 28432
rect 30024 28150 30052 28426
rect 30116 28422 30144 28580
rect 30300 28558 30328 28970
rect 30493 28860 30801 28869
rect 30493 28858 30499 28860
rect 30555 28858 30579 28860
rect 30635 28858 30659 28860
rect 30715 28858 30739 28860
rect 30795 28858 30801 28860
rect 30555 28806 30557 28858
rect 30737 28806 30739 28858
rect 30493 28804 30499 28806
rect 30555 28804 30579 28806
rect 30635 28804 30659 28806
rect 30715 28804 30739 28806
rect 30795 28804 30801 28806
rect 30493 28795 30801 28804
rect 30288 28552 30340 28558
rect 30288 28494 30340 28500
rect 30104 28416 30156 28422
rect 30104 28358 30156 28364
rect 30840 28416 30892 28422
rect 30840 28358 30892 28364
rect 30012 28144 30064 28150
rect 30012 28086 30064 28092
rect 30380 27872 30432 27878
rect 30380 27814 30432 27820
rect 30012 27668 30064 27674
rect 30012 27610 30064 27616
rect 29920 27532 29972 27538
rect 29920 27474 29972 27480
rect 29828 27464 29880 27470
rect 29828 27406 29880 27412
rect 30024 27452 30052 27610
rect 30196 27532 30248 27538
rect 30196 27474 30248 27480
rect 30288 27532 30340 27538
rect 30288 27474 30340 27480
rect 30104 27464 30156 27470
rect 30024 27424 30104 27452
rect 29736 26444 29788 26450
rect 29736 26386 29788 26392
rect 29736 26240 29788 26246
rect 29736 26182 29788 26188
rect 29644 25152 29696 25158
rect 29644 25094 29696 25100
rect 29748 24886 29776 26182
rect 29736 24880 29788 24886
rect 29736 24822 29788 24828
rect 29552 24744 29604 24750
rect 29552 24686 29604 24692
rect 29564 24274 29592 24686
rect 29736 24608 29788 24614
rect 29736 24550 29788 24556
rect 29552 24268 29604 24274
rect 29552 24210 29604 24216
rect 29748 23866 29776 24550
rect 29736 23860 29788 23866
rect 29736 23802 29788 23808
rect 29736 22568 29788 22574
rect 29736 22510 29788 22516
rect 29644 22160 29696 22166
rect 29644 22102 29696 22108
rect 29656 21418 29684 22102
rect 29644 21412 29696 21418
rect 29644 21354 29696 21360
rect 29748 21350 29776 22510
rect 29736 21344 29788 21350
rect 29736 21286 29788 21292
rect 29460 21140 29512 21146
rect 29460 21082 29512 21088
rect 29748 20641 29776 21286
rect 29840 20942 29868 27406
rect 29920 26784 29972 26790
rect 29920 26726 29972 26732
rect 29932 26518 29960 26726
rect 29920 26512 29972 26518
rect 29920 26454 29972 26460
rect 29932 25702 29960 26454
rect 29920 25696 29972 25702
rect 29920 25638 29972 25644
rect 30024 25106 30052 27424
rect 30104 27406 30156 27412
rect 30104 27328 30156 27334
rect 30104 27270 30156 27276
rect 30116 25294 30144 27270
rect 30208 26586 30236 27474
rect 30196 26580 30248 26586
rect 30196 26522 30248 26528
rect 30300 26382 30328 27474
rect 30288 26376 30340 26382
rect 30288 26318 30340 26324
rect 30392 25344 30420 27814
rect 30493 27772 30801 27781
rect 30493 27770 30499 27772
rect 30555 27770 30579 27772
rect 30635 27770 30659 27772
rect 30715 27770 30739 27772
rect 30795 27770 30801 27772
rect 30555 27718 30557 27770
rect 30737 27718 30739 27770
rect 30493 27716 30499 27718
rect 30555 27716 30579 27718
rect 30635 27716 30659 27718
rect 30715 27716 30739 27718
rect 30795 27716 30801 27718
rect 30493 27707 30801 27716
rect 30493 26684 30801 26693
rect 30493 26682 30499 26684
rect 30555 26682 30579 26684
rect 30635 26682 30659 26684
rect 30715 26682 30739 26684
rect 30795 26682 30801 26684
rect 30555 26630 30557 26682
rect 30737 26630 30739 26682
rect 30493 26628 30499 26630
rect 30555 26628 30579 26630
rect 30635 26628 30659 26630
rect 30715 26628 30739 26630
rect 30795 26628 30801 26630
rect 30493 26619 30801 26628
rect 30852 26450 30880 28358
rect 30944 28218 30972 29135
rect 31036 28257 31064 29566
rect 31116 29504 31168 29510
rect 31116 29446 31168 29452
rect 31128 29306 31156 29446
rect 31116 29300 31168 29306
rect 31300 29300 31352 29306
rect 31116 29242 31168 29248
rect 31220 29260 31300 29288
rect 31116 29164 31168 29170
rect 31116 29106 31168 29112
rect 31128 28694 31156 29106
rect 31116 28688 31168 28694
rect 31116 28630 31168 28636
rect 31022 28248 31078 28257
rect 30932 28212 30984 28218
rect 31022 28183 31078 28192
rect 30932 28154 30984 28160
rect 31024 28144 31076 28150
rect 31024 28086 31076 28092
rect 30932 28008 30984 28014
rect 30932 27950 30984 27956
rect 30944 27577 30972 27950
rect 30930 27568 30986 27577
rect 30930 27503 30986 27512
rect 30932 26852 30984 26858
rect 30932 26794 30984 26800
rect 30840 26444 30892 26450
rect 30840 26386 30892 26392
rect 30944 26314 30972 26794
rect 30932 26308 30984 26314
rect 30932 26250 30984 26256
rect 31036 26246 31064 28086
rect 31128 28082 31156 28630
rect 31116 28076 31168 28082
rect 31116 28018 31168 28024
rect 31116 27464 31168 27470
rect 31116 27406 31168 27412
rect 31128 26994 31156 27406
rect 31116 26988 31168 26994
rect 31116 26930 31168 26936
rect 31220 26330 31248 29260
rect 31300 29242 31352 29248
rect 31300 27872 31352 27878
rect 31300 27814 31352 27820
rect 31312 27538 31340 27814
rect 31300 27532 31352 27538
rect 31300 27474 31352 27480
rect 31298 26344 31354 26353
rect 31220 26302 31298 26330
rect 31298 26279 31354 26288
rect 31024 26240 31076 26246
rect 31024 26182 31076 26188
rect 31024 25900 31076 25906
rect 31024 25842 31076 25848
rect 30493 25596 30801 25605
rect 30493 25594 30499 25596
rect 30555 25594 30579 25596
rect 30635 25594 30659 25596
rect 30715 25594 30739 25596
rect 30795 25594 30801 25596
rect 30555 25542 30557 25594
rect 30737 25542 30739 25594
rect 30493 25540 30499 25542
rect 30555 25540 30579 25542
rect 30635 25540 30659 25542
rect 30715 25540 30739 25542
rect 30795 25540 30801 25542
rect 30493 25531 30801 25540
rect 31036 25498 31064 25842
rect 31208 25696 31260 25702
rect 31208 25638 31260 25644
rect 31024 25492 31076 25498
rect 31024 25434 31076 25440
rect 31114 25392 31170 25401
rect 30392 25316 30512 25344
rect 31114 25327 31170 25336
rect 30104 25288 30156 25294
rect 30104 25230 30156 25236
rect 30380 25220 30432 25226
rect 30380 25162 30432 25168
rect 30024 25078 30144 25106
rect 29920 24608 29972 24614
rect 29920 24550 29972 24556
rect 29932 22506 29960 24550
rect 30116 24188 30144 25078
rect 30196 24812 30248 24818
rect 30196 24754 30248 24760
rect 30024 24160 30144 24188
rect 29920 22500 29972 22506
rect 29920 22442 29972 22448
rect 30024 22094 30052 24160
rect 30208 24070 30236 24754
rect 30288 24200 30340 24206
rect 30288 24142 30340 24148
rect 30196 24064 30248 24070
rect 30196 24006 30248 24012
rect 30104 23656 30156 23662
rect 30104 23598 30156 23604
rect 30116 22982 30144 23598
rect 30104 22976 30156 22982
rect 30104 22918 30156 22924
rect 30116 22642 30144 22918
rect 30104 22636 30156 22642
rect 30104 22578 30156 22584
rect 30116 22234 30144 22578
rect 30104 22228 30156 22234
rect 30104 22170 30156 22176
rect 30024 22066 30144 22094
rect 29920 21072 29972 21078
rect 29920 21014 29972 21020
rect 29828 20936 29880 20942
rect 29828 20878 29880 20884
rect 29734 20632 29790 20641
rect 29734 20567 29790 20576
rect 29828 20528 29880 20534
rect 29380 20488 29592 20516
rect 29460 20392 29512 20398
rect 29460 20334 29512 20340
rect 29276 19848 29328 19854
rect 29276 19790 29328 19796
rect 29092 19712 29144 19718
rect 29092 19654 29144 19660
rect 29288 19378 29316 19790
rect 29366 19680 29422 19689
rect 29366 19615 29422 19624
rect 29380 19378 29408 19615
rect 29276 19372 29328 19378
rect 29276 19314 29328 19320
rect 29368 19372 29420 19378
rect 29368 19314 29420 19320
rect 29092 18828 29144 18834
rect 29092 18770 29144 18776
rect 28736 18686 28948 18714
rect 29000 18760 29052 18766
rect 29000 18702 29052 18708
rect 28736 16114 28764 18686
rect 29012 18358 29040 18702
rect 29000 18352 29052 18358
rect 29000 18294 29052 18300
rect 28908 17672 28960 17678
rect 28908 17614 28960 17620
rect 28816 17128 28868 17134
rect 28816 17070 28868 17076
rect 28828 16794 28856 17070
rect 28816 16788 28868 16794
rect 28816 16730 28868 16736
rect 28920 16250 28948 17614
rect 29104 16522 29132 18770
rect 29184 17196 29236 17202
rect 29184 17138 29236 17144
rect 29092 16516 29144 16522
rect 29092 16458 29144 16464
rect 28908 16244 28960 16250
rect 28908 16186 28960 16192
rect 28816 16176 28868 16182
rect 28816 16118 28868 16124
rect 29090 16144 29146 16153
rect 28724 16108 28776 16114
rect 28724 16050 28776 16056
rect 28632 16040 28684 16046
rect 28632 15982 28684 15988
rect 28448 15904 28500 15910
rect 28448 15846 28500 15852
rect 28460 15502 28488 15846
rect 28644 15502 28672 15982
rect 28448 15496 28500 15502
rect 28448 15438 28500 15444
rect 28632 15496 28684 15502
rect 28632 15438 28684 15444
rect 28356 15360 28408 15366
rect 28356 15302 28408 15308
rect 28828 15026 28856 16118
rect 29090 16079 29092 16088
rect 29144 16079 29146 16088
rect 29092 16050 29144 16056
rect 29090 16008 29146 16017
rect 29090 15943 29092 15952
rect 29144 15943 29146 15952
rect 29092 15914 29144 15920
rect 29000 15904 29052 15910
rect 29000 15846 29052 15852
rect 29012 15609 29040 15846
rect 29196 15706 29224 17138
rect 29288 16182 29316 19314
rect 29380 17134 29408 19314
rect 29472 18970 29500 20334
rect 29460 18964 29512 18970
rect 29460 18906 29512 18912
rect 29460 17808 29512 17814
rect 29460 17750 29512 17756
rect 29368 17128 29420 17134
rect 29368 17070 29420 17076
rect 29368 16992 29420 16998
rect 29368 16934 29420 16940
rect 29380 16726 29408 16934
rect 29368 16720 29420 16726
rect 29368 16662 29420 16668
rect 29472 16454 29500 17750
rect 29564 16697 29592 20488
rect 29828 20470 29880 20476
rect 29736 19984 29788 19990
rect 29736 19926 29788 19932
rect 29748 19174 29776 19926
rect 29840 19854 29868 20470
rect 29828 19848 29880 19854
rect 29828 19790 29880 19796
rect 29840 19310 29868 19790
rect 29828 19304 29880 19310
rect 29828 19246 29880 19252
rect 29736 19168 29788 19174
rect 29736 19110 29788 19116
rect 29748 18873 29776 19110
rect 29734 18864 29790 18873
rect 29644 18828 29696 18834
rect 29734 18799 29790 18808
rect 29644 18770 29696 18776
rect 29656 17202 29684 18770
rect 29748 17814 29776 18799
rect 29840 17882 29868 19246
rect 29828 17876 29880 17882
rect 29828 17818 29880 17824
rect 29736 17808 29788 17814
rect 29736 17750 29788 17756
rect 29736 17604 29788 17610
rect 29736 17546 29788 17552
rect 29644 17196 29696 17202
rect 29644 17138 29696 17144
rect 29748 16794 29776 17546
rect 29828 17332 29880 17338
rect 29828 17274 29880 17280
rect 29840 16794 29868 17274
rect 29736 16788 29788 16794
rect 29736 16730 29788 16736
rect 29828 16788 29880 16794
rect 29828 16730 29880 16736
rect 29550 16688 29606 16697
rect 29550 16623 29606 16632
rect 29552 16516 29604 16522
rect 29552 16458 29604 16464
rect 29460 16448 29512 16454
rect 29460 16390 29512 16396
rect 29472 16182 29500 16390
rect 29276 16176 29328 16182
rect 29460 16176 29512 16182
rect 29276 16118 29328 16124
rect 29366 16144 29422 16153
rect 29460 16118 29512 16124
rect 29366 16079 29368 16088
rect 29420 16079 29422 16088
rect 29368 16050 29420 16056
rect 29564 16046 29592 16458
rect 29932 16436 29960 21014
rect 30116 20942 30144 22066
rect 30104 20936 30156 20942
rect 30104 20878 30156 20884
rect 30012 20868 30064 20874
rect 30012 20810 30064 20816
rect 30024 17184 30052 20810
rect 30208 20602 30236 24006
rect 30300 23594 30328 24142
rect 30288 23588 30340 23594
rect 30288 23530 30340 23536
rect 30300 22982 30328 23530
rect 30288 22976 30340 22982
rect 30288 22918 30340 22924
rect 30288 21888 30340 21894
rect 30288 21830 30340 21836
rect 30300 21622 30328 21830
rect 30288 21616 30340 21622
rect 30288 21558 30340 21564
rect 30392 20777 30420 25162
rect 30484 24868 30512 25316
rect 31128 25294 31156 25327
rect 30656 25288 30708 25294
rect 30656 25230 30708 25236
rect 31116 25288 31168 25294
rect 31116 25230 31168 25236
rect 30668 24886 30696 25230
rect 30748 25220 30800 25226
rect 30748 25162 30800 25168
rect 30564 24880 30616 24886
rect 30484 24840 30564 24868
rect 30564 24822 30616 24828
rect 30656 24880 30708 24886
rect 30656 24822 30708 24828
rect 30760 24682 30788 25162
rect 31024 24812 31076 24818
rect 31024 24754 31076 24760
rect 30748 24676 30800 24682
rect 30748 24618 30800 24624
rect 30493 24508 30801 24517
rect 30493 24506 30499 24508
rect 30555 24506 30579 24508
rect 30635 24506 30659 24508
rect 30715 24506 30739 24508
rect 30795 24506 30801 24508
rect 30555 24454 30557 24506
rect 30737 24454 30739 24506
rect 30493 24452 30499 24454
rect 30555 24452 30579 24454
rect 30635 24452 30659 24454
rect 30715 24452 30739 24454
rect 30795 24452 30801 24454
rect 30493 24443 30801 24452
rect 31036 24274 31064 24754
rect 31220 24750 31248 25638
rect 31208 24744 31260 24750
rect 31208 24686 31260 24692
rect 31116 24608 31168 24614
rect 31116 24550 31168 24556
rect 30932 24268 30984 24274
rect 30932 24210 30984 24216
rect 31024 24268 31076 24274
rect 31024 24210 31076 24216
rect 30656 24200 30708 24206
rect 30656 24142 30708 24148
rect 30944 24154 30972 24210
rect 31128 24206 31156 24550
rect 31116 24200 31168 24206
rect 30668 23662 30696 24142
rect 30944 24126 31064 24154
rect 31116 24142 31168 24148
rect 30656 23656 30708 23662
rect 30656 23598 30708 23604
rect 30840 23520 30892 23526
rect 30840 23462 30892 23468
rect 30932 23520 30984 23526
rect 30932 23462 30984 23468
rect 30493 23420 30801 23429
rect 30493 23418 30499 23420
rect 30555 23418 30579 23420
rect 30635 23418 30659 23420
rect 30715 23418 30739 23420
rect 30795 23418 30801 23420
rect 30555 23366 30557 23418
rect 30737 23366 30739 23418
rect 30493 23364 30499 23366
rect 30555 23364 30579 23366
rect 30635 23364 30659 23366
rect 30715 23364 30739 23366
rect 30795 23364 30801 23366
rect 30493 23355 30801 23364
rect 30472 22976 30524 22982
rect 30472 22918 30524 22924
rect 30484 22778 30512 22918
rect 30472 22772 30524 22778
rect 30472 22714 30524 22720
rect 30852 22710 30880 23462
rect 30840 22704 30892 22710
rect 30840 22646 30892 22652
rect 30493 22332 30801 22341
rect 30493 22330 30499 22332
rect 30555 22330 30579 22332
rect 30635 22330 30659 22332
rect 30715 22330 30739 22332
rect 30795 22330 30801 22332
rect 30555 22278 30557 22330
rect 30737 22278 30739 22330
rect 30493 22276 30499 22278
rect 30555 22276 30579 22278
rect 30635 22276 30659 22278
rect 30715 22276 30739 22278
rect 30795 22276 30801 22278
rect 30493 22267 30801 22276
rect 30944 22094 30972 23462
rect 31036 23118 31064 24126
rect 31312 23254 31340 26279
rect 31404 25906 31432 29974
rect 31496 29173 31524 29990
rect 31588 29481 31616 30262
rect 31668 30252 31720 30258
rect 31668 30194 31720 30200
rect 31574 29472 31630 29481
rect 31574 29407 31630 29416
rect 31576 29300 31628 29306
rect 31680 29288 31708 30194
rect 31772 29617 31800 30738
rect 31942 29880 31998 29889
rect 31942 29815 31998 29824
rect 31758 29608 31814 29617
rect 31758 29543 31814 29552
rect 31628 29260 31708 29288
rect 31576 29242 31628 29248
rect 31481 29167 31533 29173
rect 31481 29109 31533 29115
rect 31772 29050 31800 29543
rect 31852 29232 31904 29238
rect 31850 29200 31852 29209
rect 31904 29200 31906 29209
rect 31956 29170 31984 29815
rect 32048 29646 32076 30738
rect 32128 30592 32180 30598
rect 32128 30534 32180 30540
rect 32036 29640 32088 29646
rect 32036 29582 32088 29588
rect 32036 29504 32088 29510
rect 32036 29446 32088 29452
rect 31850 29135 31906 29144
rect 31944 29164 31996 29170
rect 31944 29106 31996 29112
rect 32048 29050 32076 29446
rect 32140 29170 32168 30534
rect 32416 29714 32444 31622
rect 32508 31346 32536 34462
rect 32680 33312 32732 33318
rect 32680 33254 32732 33260
rect 32588 33108 32640 33114
rect 32588 33050 32640 33056
rect 32600 32314 32628 33050
rect 32692 32502 32720 33254
rect 32680 32496 32732 32502
rect 32680 32438 32732 32444
rect 32600 32286 32720 32314
rect 32586 31920 32642 31929
rect 32586 31855 32642 31864
rect 32496 31340 32548 31346
rect 32496 31282 32548 31288
rect 32496 30252 32548 30258
rect 32496 30194 32548 30200
rect 32404 29708 32456 29714
rect 32404 29650 32456 29656
rect 32220 29572 32272 29578
rect 32220 29514 32272 29520
rect 32128 29164 32180 29170
rect 32128 29106 32180 29112
rect 31668 29028 31720 29034
rect 31772 29022 31892 29050
rect 31668 28970 31720 28976
rect 31576 28960 31628 28966
rect 31576 28902 31628 28908
rect 31484 28484 31536 28490
rect 31484 28426 31536 28432
rect 31496 27470 31524 28426
rect 31588 28014 31616 28902
rect 31680 28370 31708 28970
rect 31864 28626 31892 29022
rect 31956 29022 32076 29050
rect 31956 28762 31984 29022
rect 32232 28994 32260 29514
rect 32402 29200 32458 29209
rect 32402 29135 32404 29144
rect 32456 29135 32458 29144
rect 32404 29106 32456 29112
rect 32048 28966 32260 28994
rect 32404 29028 32456 29034
rect 32404 28970 32456 28976
rect 31944 28756 31996 28762
rect 31944 28698 31996 28704
rect 31852 28620 31904 28626
rect 31852 28562 31904 28568
rect 31680 28342 31800 28370
rect 31668 28212 31720 28218
rect 31668 28154 31720 28160
rect 31576 28008 31628 28014
rect 31576 27950 31628 27956
rect 31484 27464 31536 27470
rect 31484 27406 31536 27412
rect 31496 26246 31524 27406
rect 31588 27402 31616 27950
rect 31680 27538 31708 28154
rect 31772 27985 31800 28342
rect 31758 27976 31814 27985
rect 31758 27911 31814 27920
rect 31668 27532 31720 27538
rect 31668 27474 31720 27480
rect 31576 27396 31628 27402
rect 31576 27338 31628 27344
rect 31668 27396 31720 27402
rect 31668 27338 31720 27344
rect 31576 26376 31628 26382
rect 31680 26364 31708 27338
rect 31772 26994 31800 27911
rect 31864 27878 31892 28562
rect 31852 27872 31904 27878
rect 31852 27814 31904 27820
rect 32048 27690 32076 28966
rect 32128 28756 32180 28762
rect 32128 28698 32180 28704
rect 32140 28422 32168 28698
rect 32128 28416 32180 28422
rect 32128 28358 32180 28364
rect 31956 27662 32076 27690
rect 31760 26988 31812 26994
rect 31760 26930 31812 26936
rect 31628 26336 31708 26364
rect 31760 26376 31812 26382
rect 31576 26318 31628 26324
rect 31812 26336 31892 26364
rect 31760 26318 31812 26324
rect 31484 26240 31536 26246
rect 31484 26182 31536 26188
rect 31760 25968 31812 25974
rect 31760 25910 31812 25916
rect 31392 25900 31444 25906
rect 31392 25842 31444 25848
rect 31484 25900 31536 25906
rect 31484 25842 31536 25848
rect 31404 24410 31432 25842
rect 31496 24993 31524 25842
rect 31668 25696 31720 25702
rect 31668 25638 31720 25644
rect 31576 25356 31628 25362
rect 31576 25298 31628 25304
rect 31588 25265 31616 25298
rect 31574 25256 31630 25265
rect 31574 25191 31630 25200
rect 31576 25152 31628 25158
rect 31574 25120 31576 25129
rect 31628 25120 31630 25129
rect 31574 25055 31630 25064
rect 31482 24984 31538 24993
rect 31482 24919 31538 24928
rect 31576 24880 31628 24886
rect 31576 24822 31628 24828
rect 31484 24812 31536 24818
rect 31484 24754 31536 24760
rect 31496 24682 31524 24754
rect 31484 24676 31536 24682
rect 31484 24618 31536 24624
rect 31392 24404 31444 24410
rect 31392 24346 31444 24352
rect 31484 23724 31536 23730
rect 31484 23666 31536 23672
rect 31392 23656 31444 23662
rect 31392 23598 31444 23604
rect 31300 23248 31352 23254
rect 31300 23190 31352 23196
rect 31024 23112 31076 23118
rect 31024 23054 31076 23060
rect 31036 22234 31064 23054
rect 31116 22976 31168 22982
rect 31116 22918 31168 22924
rect 31024 22228 31076 22234
rect 31024 22170 31076 22176
rect 30852 22066 30972 22094
rect 30852 21350 30880 22066
rect 31128 21486 31156 22918
rect 31404 22778 31432 23598
rect 31392 22772 31444 22778
rect 31392 22714 31444 22720
rect 31300 22500 31352 22506
rect 31300 22442 31352 22448
rect 30932 21480 30984 21486
rect 30932 21422 30984 21428
rect 31116 21480 31168 21486
rect 31116 21422 31168 21428
rect 30840 21344 30892 21350
rect 30840 21286 30892 21292
rect 30493 21244 30801 21253
rect 30493 21242 30499 21244
rect 30555 21242 30579 21244
rect 30635 21242 30659 21244
rect 30715 21242 30739 21244
rect 30795 21242 30801 21244
rect 30555 21190 30557 21242
rect 30737 21190 30739 21242
rect 30493 21188 30499 21190
rect 30555 21188 30579 21190
rect 30635 21188 30659 21190
rect 30715 21188 30739 21190
rect 30795 21188 30801 21190
rect 30493 21179 30801 21188
rect 30470 21040 30526 21049
rect 30470 20975 30472 20984
rect 30524 20975 30526 20984
rect 30840 21004 30892 21010
rect 30472 20946 30524 20952
rect 30840 20946 30892 20952
rect 30378 20768 30434 20777
rect 30378 20703 30434 20712
rect 30196 20596 30248 20602
rect 30196 20538 30248 20544
rect 30104 20392 30156 20398
rect 30104 20334 30156 20340
rect 30116 19514 30144 20334
rect 30493 20156 30801 20165
rect 30493 20154 30499 20156
rect 30555 20154 30579 20156
rect 30635 20154 30659 20156
rect 30715 20154 30739 20156
rect 30795 20154 30801 20156
rect 30555 20102 30557 20154
rect 30737 20102 30739 20154
rect 30493 20100 30499 20102
rect 30555 20100 30579 20102
rect 30635 20100 30659 20102
rect 30715 20100 30739 20102
rect 30795 20100 30801 20102
rect 30493 20091 30801 20100
rect 30852 19904 30880 20946
rect 30760 19876 30880 19904
rect 30196 19712 30248 19718
rect 30196 19654 30248 19660
rect 30104 19508 30156 19514
rect 30104 19450 30156 19456
rect 30208 18834 30236 19654
rect 30760 19174 30788 19876
rect 30840 19780 30892 19786
rect 30840 19722 30892 19728
rect 30748 19168 30800 19174
rect 30748 19110 30800 19116
rect 30493 19068 30801 19077
rect 30493 19066 30499 19068
rect 30555 19066 30579 19068
rect 30635 19066 30659 19068
rect 30715 19066 30739 19068
rect 30795 19066 30801 19068
rect 30555 19014 30557 19066
rect 30737 19014 30739 19066
rect 30493 19012 30499 19014
rect 30555 19012 30579 19014
rect 30635 19012 30659 19014
rect 30715 19012 30739 19014
rect 30795 19012 30801 19014
rect 30493 19003 30801 19012
rect 30852 18970 30880 19722
rect 30840 18964 30892 18970
rect 30840 18906 30892 18912
rect 30196 18828 30248 18834
rect 30196 18770 30248 18776
rect 30840 18692 30892 18698
rect 30840 18634 30892 18640
rect 30288 18624 30340 18630
rect 30288 18566 30340 18572
rect 30196 18284 30248 18290
rect 30196 18226 30248 18232
rect 30024 17156 30144 17184
rect 30012 17060 30064 17066
rect 30012 17002 30064 17008
rect 30024 16590 30052 17002
rect 30012 16584 30064 16590
rect 30012 16526 30064 16532
rect 30012 16448 30064 16454
rect 29932 16408 30012 16436
rect 30012 16390 30064 16396
rect 29828 16108 29880 16114
rect 29828 16050 29880 16056
rect 29552 16040 29604 16046
rect 29840 16017 29868 16050
rect 29552 15982 29604 15988
rect 29826 16008 29882 16017
rect 29826 15943 29882 15952
rect 29184 15700 29236 15706
rect 29184 15642 29236 15648
rect 28998 15600 29054 15609
rect 28998 15535 29054 15544
rect 29828 15496 29880 15502
rect 29828 15438 29880 15444
rect 29366 15192 29422 15201
rect 29366 15127 29368 15136
rect 29420 15127 29422 15136
rect 29368 15098 29420 15104
rect 29840 15094 29868 15438
rect 30116 15094 30144 17156
rect 30208 16182 30236 18226
rect 30300 17338 30328 18566
rect 30493 17980 30801 17989
rect 30493 17978 30499 17980
rect 30555 17978 30579 17980
rect 30635 17978 30659 17980
rect 30715 17978 30739 17980
rect 30795 17978 30801 17980
rect 30555 17926 30557 17978
rect 30737 17926 30739 17978
rect 30493 17924 30499 17926
rect 30555 17924 30579 17926
rect 30635 17924 30659 17926
rect 30715 17924 30739 17926
rect 30795 17924 30801 17926
rect 30493 17915 30801 17924
rect 30656 17536 30708 17542
rect 30656 17478 30708 17484
rect 30288 17332 30340 17338
rect 30288 17274 30340 17280
rect 30380 17332 30432 17338
rect 30380 17274 30432 17280
rect 30392 17218 30420 17274
rect 30668 17270 30696 17478
rect 30300 17190 30420 17218
rect 30656 17264 30708 17270
rect 30656 17206 30708 17212
rect 30472 17196 30524 17202
rect 30196 16176 30248 16182
rect 30196 16118 30248 16124
rect 30300 15162 30328 17190
rect 30472 17138 30524 17144
rect 30484 17105 30512 17138
rect 30470 17096 30526 17105
rect 30380 17060 30432 17066
rect 30470 17031 30526 17040
rect 30380 17002 30432 17008
rect 30392 16522 30420 17002
rect 30484 16998 30512 17031
rect 30472 16992 30524 16998
rect 30472 16934 30524 16940
rect 30493 16892 30801 16901
rect 30493 16890 30499 16892
rect 30555 16890 30579 16892
rect 30635 16890 30659 16892
rect 30715 16890 30739 16892
rect 30795 16890 30801 16892
rect 30555 16838 30557 16890
rect 30737 16838 30739 16890
rect 30493 16836 30499 16838
rect 30555 16836 30579 16838
rect 30635 16836 30659 16838
rect 30715 16836 30739 16838
rect 30795 16836 30801 16838
rect 30493 16827 30801 16836
rect 30472 16720 30524 16726
rect 30470 16688 30472 16697
rect 30524 16688 30526 16697
rect 30470 16623 30526 16632
rect 30654 16688 30710 16697
rect 30654 16623 30710 16632
rect 30380 16516 30432 16522
rect 30380 16458 30432 16464
rect 30472 16516 30524 16522
rect 30472 16458 30524 16464
rect 30484 16114 30512 16458
rect 30668 16114 30696 16623
rect 30746 16280 30802 16289
rect 30746 16215 30748 16224
rect 30800 16215 30802 16224
rect 30748 16186 30800 16192
rect 30472 16108 30524 16114
rect 30392 16068 30472 16096
rect 30392 15502 30420 16068
rect 30472 16050 30524 16056
rect 30656 16108 30708 16114
rect 30656 16050 30708 16056
rect 30493 15804 30801 15813
rect 30493 15802 30499 15804
rect 30555 15802 30579 15804
rect 30635 15802 30659 15804
rect 30715 15802 30739 15804
rect 30795 15802 30801 15804
rect 30555 15750 30557 15802
rect 30737 15750 30739 15802
rect 30493 15748 30499 15750
rect 30555 15748 30579 15750
rect 30635 15748 30659 15750
rect 30715 15748 30739 15750
rect 30795 15748 30801 15750
rect 30493 15739 30801 15748
rect 30852 15706 30880 18634
rect 30944 18358 30972 21422
rect 31116 21344 31168 21350
rect 31116 21286 31168 21292
rect 31024 20256 31076 20262
rect 31024 20198 31076 20204
rect 31036 19378 31064 20198
rect 31024 19372 31076 19378
rect 31024 19314 31076 19320
rect 31128 19174 31156 21286
rect 31312 20942 31340 22442
rect 31404 21010 31432 22714
rect 31392 21004 31444 21010
rect 31392 20946 31444 20952
rect 31300 20936 31352 20942
rect 31300 20878 31352 20884
rect 31208 20460 31260 20466
rect 31208 20402 31260 20408
rect 31024 19168 31076 19174
rect 31024 19110 31076 19116
rect 31116 19168 31168 19174
rect 31116 19110 31168 19116
rect 30932 18352 30984 18358
rect 31036 18340 31064 19110
rect 31116 18352 31168 18358
rect 31036 18312 31116 18340
rect 30932 18294 30984 18300
rect 31116 18294 31168 18300
rect 30932 18216 30984 18222
rect 30932 18158 30984 18164
rect 30944 17814 30972 18158
rect 30932 17808 30984 17814
rect 30932 17750 30984 17756
rect 30944 17202 30972 17750
rect 31024 17740 31076 17746
rect 31024 17682 31076 17688
rect 30932 17196 30984 17202
rect 30932 17138 30984 17144
rect 30930 16824 30986 16833
rect 30930 16759 30986 16768
rect 30840 15700 30892 15706
rect 30840 15642 30892 15648
rect 30838 15600 30894 15609
rect 30838 15535 30894 15544
rect 30852 15502 30880 15535
rect 30380 15496 30432 15502
rect 30380 15438 30432 15444
rect 30840 15496 30892 15502
rect 30840 15438 30892 15444
rect 30944 15178 30972 16759
rect 30288 15156 30340 15162
rect 30288 15098 30340 15104
rect 30852 15150 30972 15178
rect 29828 15088 29880 15094
rect 29828 15030 29880 15036
rect 30104 15088 30156 15094
rect 30104 15030 30156 15036
rect 27804 15020 27856 15026
rect 27804 14962 27856 14968
rect 28172 15020 28224 15026
rect 28172 14962 28224 14968
rect 28816 15020 28868 15026
rect 28816 14962 28868 14968
rect 29000 14952 29052 14958
rect 29000 14894 29052 14900
rect 27436 14544 27488 14550
rect 27436 14486 27488 14492
rect 26608 14408 26660 14414
rect 26608 14350 26660 14356
rect 26884 14408 26936 14414
rect 26884 14350 26936 14356
rect 26056 14340 26108 14346
rect 26056 14282 26108 14288
rect 26272 14172 26580 14181
rect 26272 14170 26278 14172
rect 26334 14170 26358 14172
rect 26414 14170 26438 14172
rect 26494 14170 26518 14172
rect 26574 14170 26580 14172
rect 26334 14118 26336 14170
rect 26516 14118 26518 14170
rect 26272 14116 26278 14118
rect 26334 14116 26358 14118
rect 26414 14116 26438 14118
rect 26494 14116 26518 14118
rect 26574 14116 26580 14118
rect 26272 14107 26580 14116
rect 22052 13628 22360 13637
rect 22052 13626 22058 13628
rect 22114 13626 22138 13628
rect 22194 13626 22218 13628
rect 22274 13626 22298 13628
rect 22354 13626 22360 13628
rect 22114 13574 22116 13626
rect 22296 13574 22298 13626
rect 22052 13572 22058 13574
rect 22114 13572 22138 13574
rect 22194 13572 22218 13574
rect 22274 13572 22298 13574
rect 22354 13572 22360 13574
rect 22052 13563 22360 13572
rect 26272 13084 26580 13093
rect 26272 13082 26278 13084
rect 26334 13082 26358 13084
rect 26414 13082 26438 13084
rect 26494 13082 26518 13084
rect 26574 13082 26580 13084
rect 26334 13030 26336 13082
rect 26516 13030 26518 13082
rect 26272 13028 26278 13030
rect 26334 13028 26358 13030
rect 26414 13028 26438 13030
rect 26494 13028 26518 13030
rect 26574 13028 26580 13030
rect 26272 13019 26580 13028
rect 22052 12540 22360 12549
rect 22052 12538 22058 12540
rect 22114 12538 22138 12540
rect 22194 12538 22218 12540
rect 22274 12538 22298 12540
rect 22354 12538 22360 12540
rect 22114 12486 22116 12538
rect 22296 12486 22298 12538
rect 22052 12484 22058 12486
rect 22114 12484 22138 12486
rect 22194 12484 22218 12486
rect 22274 12484 22298 12486
rect 22354 12484 22360 12486
rect 22052 12475 22360 12484
rect 26272 11996 26580 12005
rect 26272 11994 26278 11996
rect 26334 11994 26358 11996
rect 26414 11994 26438 11996
rect 26494 11994 26518 11996
rect 26574 11994 26580 11996
rect 26334 11942 26336 11994
rect 26516 11942 26518 11994
rect 26272 11940 26278 11942
rect 26334 11940 26358 11942
rect 26414 11940 26438 11942
rect 26494 11940 26518 11942
rect 26574 11940 26580 11942
rect 26272 11931 26580 11940
rect 22052 11452 22360 11461
rect 22052 11450 22058 11452
rect 22114 11450 22138 11452
rect 22194 11450 22218 11452
rect 22274 11450 22298 11452
rect 22354 11450 22360 11452
rect 22114 11398 22116 11450
rect 22296 11398 22298 11450
rect 22052 11396 22058 11398
rect 22114 11396 22138 11398
rect 22194 11396 22218 11398
rect 22274 11396 22298 11398
rect 22354 11396 22360 11398
rect 22052 11387 22360 11396
rect 26272 10908 26580 10917
rect 26272 10906 26278 10908
rect 26334 10906 26358 10908
rect 26414 10906 26438 10908
rect 26494 10906 26518 10908
rect 26574 10906 26580 10908
rect 26334 10854 26336 10906
rect 26516 10854 26518 10906
rect 26272 10852 26278 10854
rect 26334 10852 26358 10854
rect 26414 10852 26438 10854
rect 26494 10852 26518 10854
rect 26574 10852 26580 10854
rect 26272 10843 26580 10852
rect 22052 10364 22360 10373
rect 22052 10362 22058 10364
rect 22114 10362 22138 10364
rect 22194 10362 22218 10364
rect 22274 10362 22298 10364
rect 22354 10362 22360 10364
rect 22114 10310 22116 10362
rect 22296 10310 22298 10362
rect 22052 10308 22058 10310
rect 22114 10308 22138 10310
rect 22194 10308 22218 10310
rect 22274 10308 22298 10310
rect 22354 10308 22360 10310
rect 22052 10299 22360 10308
rect 26272 9820 26580 9829
rect 26272 9818 26278 9820
rect 26334 9818 26358 9820
rect 26414 9818 26438 9820
rect 26494 9818 26518 9820
rect 26574 9818 26580 9820
rect 26334 9766 26336 9818
rect 26516 9766 26518 9818
rect 26272 9764 26278 9766
rect 26334 9764 26358 9766
rect 26414 9764 26438 9766
rect 26494 9764 26518 9766
rect 26574 9764 26580 9766
rect 26272 9755 26580 9764
rect 22052 9276 22360 9285
rect 22052 9274 22058 9276
rect 22114 9274 22138 9276
rect 22194 9274 22218 9276
rect 22274 9274 22298 9276
rect 22354 9274 22360 9276
rect 22114 9222 22116 9274
rect 22296 9222 22298 9274
rect 22052 9220 22058 9222
rect 22114 9220 22138 9222
rect 22194 9220 22218 9222
rect 22274 9220 22298 9222
rect 22354 9220 22360 9222
rect 22052 9211 22360 9220
rect 26272 8732 26580 8741
rect 26272 8730 26278 8732
rect 26334 8730 26358 8732
rect 26414 8730 26438 8732
rect 26494 8730 26518 8732
rect 26574 8730 26580 8732
rect 26334 8678 26336 8730
rect 26516 8678 26518 8730
rect 26272 8676 26278 8678
rect 26334 8676 26358 8678
rect 26414 8676 26438 8678
rect 26494 8676 26518 8678
rect 26574 8676 26580 8678
rect 26272 8667 26580 8676
rect 22052 8188 22360 8197
rect 22052 8186 22058 8188
rect 22114 8186 22138 8188
rect 22194 8186 22218 8188
rect 22274 8186 22298 8188
rect 22354 8186 22360 8188
rect 22114 8134 22116 8186
rect 22296 8134 22298 8186
rect 22052 8132 22058 8134
rect 22114 8132 22138 8134
rect 22194 8132 22218 8134
rect 22274 8132 22298 8134
rect 22354 8132 22360 8134
rect 22052 8123 22360 8132
rect 26272 7644 26580 7653
rect 26272 7642 26278 7644
rect 26334 7642 26358 7644
rect 26414 7642 26438 7644
rect 26494 7642 26518 7644
rect 26574 7642 26580 7644
rect 26334 7590 26336 7642
rect 26516 7590 26518 7642
rect 26272 7588 26278 7590
rect 26334 7588 26358 7590
rect 26414 7588 26438 7590
rect 26494 7588 26518 7590
rect 26574 7588 26580 7590
rect 26272 7579 26580 7588
rect 22052 7100 22360 7109
rect 22052 7098 22058 7100
rect 22114 7098 22138 7100
rect 22194 7098 22218 7100
rect 22274 7098 22298 7100
rect 22354 7098 22360 7100
rect 22114 7046 22116 7098
rect 22296 7046 22298 7098
rect 22052 7044 22058 7046
rect 22114 7044 22138 7046
rect 22194 7044 22218 7046
rect 22274 7044 22298 7046
rect 22354 7044 22360 7046
rect 22052 7035 22360 7044
rect 26272 6556 26580 6565
rect 26272 6554 26278 6556
rect 26334 6554 26358 6556
rect 26414 6554 26438 6556
rect 26494 6554 26518 6556
rect 26574 6554 26580 6556
rect 26334 6502 26336 6554
rect 26516 6502 26518 6554
rect 26272 6500 26278 6502
rect 26334 6500 26358 6502
rect 26414 6500 26438 6502
rect 26494 6500 26518 6502
rect 26574 6500 26580 6502
rect 26272 6491 26580 6500
rect 22052 6012 22360 6021
rect 22052 6010 22058 6012
rect 22114 6010 22138 6012
rect 22194 6010 22218 6012
rect 22274 6010 22298 6012
rect 22354 6010 22360 6012
rect 22114 5958 22116 6010
rect 22296 5958 22298 6010
rect 22052 5956 22058 5958
rect 22114 5956 22138 5958
rect 22194 5956 22218 5958
rect 22274 5956 22298 5958
rect 22354 5956 22360 5958
rect 22052 5947 22360 5956
rect 28816 5772 28868 5778
rect 28816 5714 28868 5720
rect 26272 5468 26580 5477
rect 26272 5466 26278 5468
rect 26334 5466 26358 5468
rect 26414 5466 26438 5468
rect 26494 5466 26518 5468
rect 26574 5466 26580 5468
rect 26334 5414 26336 5466
rect 26516 5414 26518 5466
rect 26272 5412 26278 5414
rect 26334 5412 26358 5414
rect 26414 5412 26438 5414
rect 26494 5412 26518 5414
rect 26574 5412 26580 5414
rect 26272 5403 26580 5412
rect 28080 5228 28132 5234
rect 28080 5170 28132 5176
rect 22052 4924 22360 4933
rect 22052 4922 22058 4924
rect 22114 4922 22138 4924
rect 22194 4922 22218 4924
rect 22274 4922 22298 4924
rect 22354 4922 22360 4924
rect 22114 4870 22116 4922
rect 22296 4870 22298 4922
rect 22052 4868 22058 4870
rect 22114 4868 22138 4870
rect 22194 4868 22218 4870
rect 22274 4868 22298 4870
rect 22354 4868 22360 4870
rect 22052 4859 22360 4868
rect 28092 4622 28120 5170
rect 28080 4616 28132 4622
rect 28080 4558 28132 4564
rect 26272 4380 26580 4389
rect 26272 4378 26278 4380
rect 26334 4378 26358 4380
rect 26414 4378 26438 4380
rect 26494 4378 26518 4380
rect 26574 4378 26580 4380
rect 26334 4326 26336 4378
rect 26516 4326 26518 4378
rect 26272 4324 26278 4326
rect 26334 4324 26358 4326
rect 26414 4324 26438 4326
rect 26494 4324 26518 4326
rect 26574 4324 26580 4326
rect 26272 4315 26580 4324
rect 28828 4146 28856 5714
rect 28816 4140 28868 4146
rect 28816 4082 28868 4088
rect 27896 4072 27948 4078
rect 27896 4014 27948 4020
rect 27712 4004 27764 4010
rect 27712 3946 27764 3952
rect 27620 3936 27672 3942
rect 27620 3878 27672 3884
rect 22052 3836 22360 3845
rect 22052 3834 22058 3836
rect 22114 3834 22138 3836
rect 22194 3834 22218 3836
rect 22274 3834 22298 3836
rect 22354 3834 22360 3836
rect 22114 3782 22116 3834
rect 22296 3782 22298 3834
rect 22052 3780 22058 3782
rect 22114 3780 22138 3782
rect 22194 3780 22218 3782
rect 22274 3780 22298 3782
rect 22354 3780 22360 3782
rect 22052 3771 22360 3780
rect 23756 3732 23808 3738
rect 23756 3674 23808 3680
rect 23768 3534 23796 3674
rect 23756 3528 23808 3534
rect 23756 3470 23808 3476
rect 24768 3528 24820 3534
rect 24768 3470 24820 3476
rect 22100 3460 22152 3466
rect 22100 3402 22152 3408
rect 22112 3194 22140 3402
rect 22100 3188 22152 3194
rect 22100 3130 22152 3136
rect 23768 3126 23796 3470
rect 24032 3392 24084 3398
rect 24032 3334 24084 3340
rect 24044 3126 24072 3334
rect 24780 3194 24808 3470
rect 26272 3292 26580 3301
rect 26272 3290 26278 3292
rect 26334 3290 26358 3292
rect 26414 3290 26438 3292
rect 26494 3290 26518 3292
rect 26574 3290 26580 3292
rect 26334 3238 26336 3290
rect 26516 3238 26518 3290
rect 26272 3236 26278 3238
rect 26334 3236 26358 3238
rect 26414 3236 26438 3238
rect 26494 3236 26518 3238
rect 26574 3236 26580 3238
rect 26272 3227 26580 3236
rect 24768 3188 24820 3194
rect 24768 3130 24820 3136
rect 27632 3126 27660 3878
rect 27724 3738 27752 3946
rect 27908 3738 27936 4014
rect 27712 3732 27764 3738
rect 27712 3674 27764 3680
rect 27896 3732 27948 3738
rect 27896 3674 27948 3680
rect 28448 3528 28500 3534
rect 28448 3470 28500 3476
rect 27712 3460 27764 3466
rect 27712 3402 27764 3408
rect 23756 3120 23808 3126
rect 23756 3062 23808 3068
rect 24032 3120 24084 3126
rect 24032 3062 24084 3068
rect 27620 3120 27672 3126
rect 27620 3062 27672 3068
rect 21916 3052 21968 3058
rect 21916 2994 21968 3000
rect 24492 2984 24544 2990
rect 24492 2926 24544 2932
rect 22052 2748 22360 2757
rect 22052 2746 22058 2748
rect 22114 2746 22138 2748
rect 22194 2746 22218 2748
rect 22274 2746 22298 2748
rect 22354 2746 22360 2748
rect 22114 2694 22116 2746
rect 22296 2694 22298 2746
rect 22052 2692 22058 2694
rect 22114 2692 22138 2694
rect 22194 2692 22218 2694
rect 22274 2692 22298 2694
rect 22354 2692 22360 2694
rect 22052 2683 22360 2692
rect 24504 800 24532 2926
rect 27724 2446 27752 3402
rect 28460 3058 28488 3470
rect 28540 3120 28592 3126
rect 28540 3062 28592 3068
rect 28448 3052 28500 3058
rect 28448 2994 28500 3000
rect 28552 2922 28580 3062
rect 28540 2916 28592 2922
rect 28540 2858 28592 2864
rect 28552 2446 28580 2858
rect 29012 2446 29040 14894
rect 30493 14716 30801 14725
rect 30493 14714 30499 14716
rect 30555 14714 30579 14716
rect 30635 14714 30659 14716
rect 30715 14714 30739 14716
rect 30795 14714 30801 14716
rect 30555 14662 30557 14714
rect 30737 14662 30739 14714
rect 30493 14660 30499 14662
rect 30555 14660 30579 14662
rect 30635 14660 30659 14662
rect 30715 14660 30739 14662
rect 30795 14660 30801 14662
rect 30493 14651 30801 14660
rect 30852 14074 30880 15150
rect 30932 15020 30984 15026
rect 30932 14962 30984 14968
rect 30840 14068 30892 14074
rect 30840 14010 30892 14016
rect 30944 13938 30972 14962
rect 31036 14618 31064 17682
rect 31128 16046 31156 18294
rect 31220 17882 31248 20402
rect 31312 18465 31340 20878
rect 31392 20800 31444 20806
rect 31392 20742 31444 20748
rect 31404 20466 31432 20742
rect 31392 20460 31444 20466
rect 31392 20402 31444 20408
rect 31404 19718 31432 20402
rect 31392 19712 31444 19718
rect 31392 19654 31444 19660
rect 31392 19508 31444 19514
rect 31392 19450 31444 19456
rect 31298 18456 31354 18465
rect 31298 18391 31300 18400
rect 31352 18391 31354 18400
rect 31300 18362 31352 18368
rect 31300 18284 31352 18290
rect 31300 18226 31352 18232
rect 31208 17876 31260 17882
rect 31208 17818 31260 17824
rect 31208 17672 31260 17678
rect 31312 17660 31340 18226
rect 31260 17632 31340 17660
rect 31208 17614 31260 17620
rect 31220 16980 31248 17614
rect 31220 16952 31340 16980
rect 31208 16584 31260 16590
rect 31206 16552 31208 16561
rect 31260 16552 31262 16561
rect 31206 16487 31262 16496
rect 31116 16040 31168 16046
rect 31116 15982 31168 15988
rect 31208 15972 31260 15978
rect 31208 15914 31260 15920
rect 31024 14612 31076 14618
rect 31024 14554 31076 14560
rect 30288 13932 30340 13938
rect 30288 13874 30340 13880
rect 30932 13932 30984 13938
rect 30932 13874 30984 13880
rect 30300 13308 30328 13874
rect 30493 13628 30801 13637
rect 30493 13626 30499 13628
rect 30555 13626 30579 13628
rect 30635 13626 30659 13628
rect 30715 13626 30739 13628
rect 30795 13626 30801 13628
rect 30555 13574 30557 13626
rect 30737 13574 30739 13626
rect 30493 13572 30499 13574
rect 30555 13572 30579 13574
rect 30635 13572 30659 13574
rect 30715 13572 30739 13574
rect 30795 13572 30801 13574
rect 30493 13563 30801 13572
rect 30380 13320 30432 13326
rect 30300 13280 30380 13308
rect 30300 6730 30328 13280
rect 30380 13262 30432 13268
rect 30944 12850 30972 13874
rect 31220 13530 31248 15914
rect 31312 15638 31340 16952
rect 31300 15632 31352 15638
rect 31300 15574 31352 15580
rect 31404 14074 31432 19450
rect 31496 18086 31524 23666
rect 31588 21434 31616 24822
rect 31680 21622 31708 25638
rect 31772 25362 31800 25910
rect 31760 25356 31812 25362
rect 31760 25298 31812 25304
rect 31772 24721 31800 25298
rect 31864 24886 31892 26336
rect 31956 25838 31984 27662
rect 32034 27568 32090 27577
rect 32034 27503 32090 27512
rect 32048 27470 32076 27503
rect 32036 27464 32088 27470
rect 32036 27406 32088 27412
rect 32140 26926 32168 28358
rect 32416 28014 32444 28970
rect 32508 28914 32536 30194
rect 32600 29714 32628 31855
rect 32692 31822 32720 32286
rect 32680 31816 32732 31822
rect 32680 31758 32732 31764
rect 32876 31498 32904 35566
rect 32784 31470 32904 31498
rect 32588 29708 32640 29714
rect 32588 29650 32640 29656
rect 32784 29510 32812 31470
rect 32968 31396 32996 35634
rect 33508 35624 33560 35630
rect 33508 35566 33560 35572
rect 33140 35488 33192 35494
rect 33140 35430 33192 35436
rect 32876 31368 32996 31396
rect 32772 29504 32824 29510
rect 32772 29446 32824 29452
rect 32508 28886 32628 28914
rect 32494 28384 32550 28393
rect 32494 28319 32550 28328
rect 32508 28082 32536 28319
rect 32496 28076 32548 28082
rect 32496 28018 32548 28024
rect 32404 28008 32456 28014
rect 32404 27950 32456 27956
rect 32404 27872 32456 27878
rect 32404 27814 32456 27820
rect 32220 27532 32272 27538
rect 32220 27474 32272 27480
rect 32128 26920 32180 26926
rect 32128 26862 32180 26868
rect 32128 26376 32180 26382
rect 32128 26318 32180 26324
rect 32140 26246 32168 26318
rect 32128 26240 32180 26246
rect 32128 26182 32180 26188
rect 31944 25832 31996 25838
rect 31944 25774 31996 25780
rect 31956 25294 31984 25774
rect 32034 25528 32090 25537
rect 32034 25463 32090 25472
rect 32048 25362 32076 25463
rect 32036 25356 32088 25362
rect 32036 25298 32088 25304
rect 31944 25288 31996 25294
rect 31944 25230 31996 25236
rect 32034 25120 32090 25129
rect 32034 25055 32090 25064
rect 31944 24948 31996 24954
rect 31944 24890 31996 24896
rect 31852 24880 31904 24886
rect 31852 24822 31904 24828
rect 31758 24712 31814 24721
rect 31758 24647 31814 24656
rect 31852 24608 31904 24614
rect 31852 24550 31904 24556
rect 31864 24206 31892 24550
rect 31852 24200 31904 24206
rect 31852 24142 31904 24148
rect 31852 24064 31904 24070
rect 31852 24006 31904 24012
rect 31760 23860 31812 23866
rect 31760 23802 31812 23808
rect 31772 22030 31800 23802
rect 31760 22024 31812 22030
rect 31760 21966 31812 21972
rect 31668 21616 31720 21622
rect 31668 21558 31720 21564
rect 31760 21548 31812 21554
rect 31760 21490 31812 21496
rect 31588 21406 31708 21434
rect 31576 21344 31628 21350
rect 31576 21286 31628 21292
rect 31588 21146 31616 21286
rect 31576 21140 31628 21146
rect 31576 21082 31628 21088
rect 31574 21040 31630 21049
rect 31574 20975 31576 20984
rect 31628 20975 31630 20984
rect 31576 20946 31628 20952
rect 31680 19530 31708 21406
rect 31772 19854 31800 21490
rect 31864 21418 31892 24006
rect 31956 23322 31984 24890
rect 32048 24206 32076 25055
rect 32128 24676 32180 24682
rect 32128 24618 32180 24624
rect 32036 24200 32088 24206
rect 32036 24142 32088 24148
rect 32036 23588 32088 23594
rect 32036 23530 32088 23536
rect 31944 23316 31996 23322
rect 31944 23258 31996 23264
rect 32048 23118 32076 23530
rect 32036 23112 32088 23118
rect 32036 23054 32088 23060
rect 32140 22094 32168 24618
rect 32232 24070 32260 27474
rect 32416 26926 32444 27814
rect 32496 27464 32548 27470
rect 32496 27406 32548 27412
rect 32600 27418 32628 28886
rect 32876 28762 32904 31368
rect 32956 30932 33008 30938
rect 32956 30874 33008 30880
rect 32968 30258 32996 30874
rect 32956 30252 33008 30258
rect 32956 30194 33008 30200
rect 33048 30252 33100 30258
rect 33048 30194 33100 30200
rect 33060 29170 33088 30194
rect 33152 29306 33180 35430
rect 33230 33824 33286 33833
rect 33230 33759 33286 33768
rect 33244 30326 33272 33759
rect 33416 32360 33468 32366
rect 33416 32302 33468 32308
rect 33428 30938 33456 32302
rect 33520 31278 33548 35566
rect 33692 35488 33744 35494
rect 33692 35430 33744 35436
rect 33508 31272 33560 31278
rect 33508 31214 33560 31220
rect 33704 31210 33732 35430
rect 34612 35012 34664 35018
rect 34612 34954 34664 34960
rect 34336 34672 34388 34678
rect 34334 34640 34336 34649
rect 34388 34640 34390 34649
rect 34334 34575 34390 34584
rect 34426 34096 34482 34105
rect 34426 34031 34482 34040
rect 34336 33924 34388 33930
rect 34336 33866 34388 33872
rect 34348 33425 34376 33866
rect 34440 33590 34468 34031
rect 34428 33584 34480 33590
rect 34428 33526 34480 33532
rect 34334 33416 34390 33425
rect 34334 33351 34390 33360
rect 34624 32881 34652 34954
rect 34713 34844 35021 34853
rect 34713 34842 34719 34844
rect 34775 34842 34799 34844
rect 34855 34842 34879 34844
rect 34935 34842 34959 34844
rect 35015 34842 35021 34844
rect 34775 34790 34777 34842
rect 34957 34790 34959 34842
rect 34713 34788 34719 34790
rect 34775 34788 34799 34790
rect 34855 34788 34879 34790
rect 34935 34788 34959 34790
rect 35015 34788 35021 34790
rect 34713 34779 35021 34788
rect 34713 33756 35021 33765
rect 34713 33754 34719 33756
rect 34775 33754 34799 33756
rect 34855 33754 34879 33756
rect 34935 33754 34959 33756
rect 35015 33754 35021 33756
rect 34775 33702 34777 33754
rect 34957 33702 34959 33754
rect 34713 33700 34719 33702
rect 34775 33700 34799 33702
rect 34855 33700 34879 33702
rect 34935 33700 34959 33702
rect 35015 33700 35021 33702
rect 34713 33691 35021 33700
rect 34610 32872 34666 32881
rect 33784 32836 33836 32842
rect 33784 32778 33836 32784
rect 34244 32836 34296 32842
rect 34610 32807 34666 32816
rect 34244 32778 34296 32784
rect 33692 31204 33744 31210
rect 33692 31146 33744 31152
rect 33416 30932 33468 30938
rect 33416 30874 33468 30880
rect 33416 30728 33468 30734
rect 33416 30670 33468 30676
rect 33232 30320 33284 30326
rect 33232 30262 33284 30268
rect 33230 29880 33286 29889
rect 33230 29815 33286 29824
rect 33244 29782 33272 29815
rect 33232 29776 33284 29782
rect 33232 29718 33284 29724
rect 33324 29640 33376 29646
rect 33322 29608 33324 29617
rect 33376 29608 33378 29617
rect 33322 29543 33378 29552
rect 33140 29300 33192 29306
rect 33140 29242 33192 29248
rect 33048 29164 33100 29170
rect 33048 29106 33100 29112
rect 33324 29164 33376 29170
rect 33324 29106 33376 29112
rect 32968 29034 33272 29050
rect 32968 29028 33284 29034
rect 32968 29022 33232 29028
rect 32864 28756 32916 28762
rect 32864 28698 32916 28704
rect 32770 28656 32826 28665
rect 32770 28591 32826 28600
rect 32678 28520 32734 28529
rect 32678 28455 32734 28464
rect 32692 28150 32720 28455
rect 32680 28144 32732 28150
rect 32680 28086 32732 28092
rect 32404 26920 32456 26926
rect 32404 26862 32456 26868
rect 32404 26784 32456 26790
rect 32404 26726 32456 26732
rect 32416 26450 32444 26726
rect 32404 26444 32456 26450
rect 32404 26386 32456 26392
rect 32312 26376 32364 26382
rect 32312 26318 32364 26324
rect 32220 24064 32272 24070
rect 32220 24006 32272 24012
rect 32324 23526 32352 26318
rect 32404 26308 32456 26314
rect 32404 26250 32456 26256
rect 32416 24682 32444 26250
rect 32508 24698 32536 27406
rect 32600 27390 32720 27418
rect 32588 27328 32640 27334
rect 32588 27270 32640 27276
rect 32600 27130 32628 27270
rect 32588 27124 32640 27130
rect 32588 27066 32640 27072
rect 32692 26602 32720 27390
rect 32784 26738 32812 28591
rect 32864 28552 32916 28558
rect 32864 28494 32916 28500
rect 32876 27946 32904 28494
rect 32864 27940 32916 27946
rect 32864 27882 32916 27888
rect 32876 26926 32904 27882
rect 32968 27062 32996 29022
rect 33232 28970 33284 28976
rect 33336 28694 33364 29106
rect 33428 29073 33456 30670
rect 33796 29646 33824 32778
rect 34060 32768 34112 32774
rect 34060 32710 34112 32716
rect 34072 31226 34100 32710
rect 33980 31198 34100 31226
rect 33874 29744 33930 29753
rect 33874 29679 33930 29688
rect 33600 29640 33652 29646
rect 33600 29582 33652 29588
rect 33784 29640 33836 29646
rect 33784 29582 33836 29588
rect 33414 29064 33470 29073
rect 33414 28999 33470 29008
rect 33324 28688 33376 28694
rect 33324 28630 33376 28636
rect 33612 28422 33640 29582
rect 33784 29504 33836 29510
rect 33784 29446 33836 29452
rect 33796 29170 33824 29446
rect 33784 29164 33836 29170
rect 33784 29106 33836 29112
rect 33796 28490 33824 29106
rect 33888 28762 33916 29679
rect 33980 29306 34008 31198
rect 34060 31136 34112 31142
rect 34060 31078 34112 31084
rect 34072 30734 34100 31078
rect 34060 30728 34112 30734
rect 34060 30670 34112 30676
rect 34256 30682 34284 32778
rect 34713 32668 35021 32677
rect 34713 32666 34719 32668
rect 34775 32666 34799 32668
rect 34855 32666 34879 32668
rect 34935 32666 34959 32668
rect 35015 32666 35021 32668
rect 34775 32614 34777 32666
rect 34957 32614 34959 32666
rect 34713 32612 34719 32614
rect 34775 32612 34799 32614
rect 34855 32612 34879 32614
rect 34935 32612 34959 32614
rect 35015 32612 35021 32614
rect 34713 32603 35021 32612
rect 34336 32360 34388 32366
rect 34336 32302 34388 32308
rect 34348 32065 34376 32302
rect 34334 32056 34390 32065
rect 34334 31991 34390 32000
rect 34713 31580 35021 31589
rect 34713 31578 34719 31580
rect 34775 31578 34799 31580
rect 34855 31578 34879 31580
rect 34935 31578 34959 31580
rect 35015 31578 35021 31580
rect 34775 31526 34777 31578
rect 34957 31526 34959 31578
rect 34713 31524 34719 31526
rect 34775 31524 34799 31526
rect 34855 31524 34879 31526
rect 34935 31524 34959 31526
rect 35015 31524 35021 31526
rect 34713 31515 35021 31524
rect 34334 31376 34390 31385
rect 34334 31311 34336 31320
rect 34388 31311 34390 31320
rect 34336 31282 34388 31288
rect 34256 30654 34376 30682
rect 34244 30592 34296 30598
rect 34244 30534 34296 30540
rect 34256 29850 34284 30534
rect 34244 29844 34296 29850
rect 34244 29786 34296 29792
rect 34244 29708 34296 29714
rect 34244 29650 34296 29656
rect 34060 29640 34112 29646
rect 34060 29582 34112 29588
rect 33968 29300 34020 29306
rect 33968 29242 34020 29248
rect 33876 28756 33928 28762
rect 33876 28698 33928 28704
rect 33784 28484 33836 28490
rect 33784 28426 33836 28432
rect 33600 28416 33652 28422
rect 33600 28358 33652 28364
rect 34072 28218 34100 29582
rect 34060 28212 34112 28218
rect 34060 28154 34112 28160
rect 34256 27674 34284 29650
rect 34348 29646 34376 30654
rect 34713 30492 35021 30501
rect 34713 30490 34719 30492
rect 34775 30490 34799 30492
rect 34855 30490 34879 30492
rect 34935 30490 34959 30492
rect 35015 30490 35021 30492
rect 34775 30438 34777 30490
rect 34957 30438 34959 30490
rect 34713 30436 34719 30438
rect 34775 30436 34799 30438
rect 34855 30436 34879 30438
rect 34935 30436 34959 30438
rect 35015 30436 35021 30438
rect 34713 30427 35021 30436
rect 34336 29640 34388 29646
rect 34336 29582 34388 29588
rect 34348 29034 34376 29582
rect 34713 29404 35021 29413
rect 34713 29402 34719 29404
rect 34775 29402 34799 29404
rect 34855 29402 34879 29404
rect 34935 29402 34959 29404
rect 35015 29402 35021 29404
rect 34775 29350 34777 29402
rect 34957 29350 34959 29402
rect 34713 29348 34719 29350
rect 34775 29348 34799 29350
rect 34855 29348 34879 29350
rect 34935 29348 34959 29350
rect 35015 29348 35021 29350
rect 34713 29339 35021 29348
rect 34336 29028 34388 29034
rect 34336 28970 34388 28976
rect 34713 28316 35021 28325
rect 34713 28314 34719 28316
rect 34775 28314 34799 28316
rect 34855 28314 34879 28316
rect 34935 28314 34959 28316
rect 35015 28314 35021 28316
rect 34775 28262 34777 28314
rect 34957 28262 34959 28314
rect 34713 28260 34719 28262
rect 34775 28260 34799 28262
rect 34855 28260 34879 28262
rect 34935 28260 34959 28262
rect 35015 28260 35021 28262
rect 34713 28251 35021 28260
rect 34336 28008 34388 28014
rect 34334 27976 34336 27985
rect 34388 27976 34390 27985
rect 34334 27911 34390 27920
rect 34244 27668 34296 27674
rect 34244 27610 34296 27616
rect 34256 27062 34284 27610
rect 34713 27228 35021 27237
rect 34713 27226 34719 27228
rect 34775 27226 34799 27228
rect 34855 27226 34879 27228
rect 34935 27226 34959 27228
rect 35015 27226 35021 27228
rect 34775 27174 34777 27226
rect 34957 27174 34959 27226
rect 34713 27172 34719 27174
rect 34775 27172 34799 27174
rect 34855 27172 34879 27174
rect 34935 27172 34959 27174
rect 35015 27172 35021 27174
rect 34713 27163 35021 27172
rect 32956 27056 33008 27062
rect 32956 26998 33008 27004
rect 33600 27056 33652 27062
rect 33600 26998 33652 27004
rect 34244 27056 34296 27062
rect 34244 26998 34296 27004
rect 33508 26988 33560 26994
rect 33508 26930 33560 26936
rect 32864 26920 32916 26926
rect 32864 26862 32916 26868
rect 33048 26920 33100 26926
rect 33048 26862 33100 26868
rect 32784 26710 32904 26738
rect 32600 26574 32720 26602
rect 32600 24970 32628 26574
rect 32680 26512 32732 26518
rect 32680 26454 32732 26460
rect 32692 26314 32720 26454
rect 32680 26308 32732 26314
rect 32680 26250 32732 26256
rect 32876 25362 32904 26710
rect 32864 25356 32916 25362
rect 32864 25298 32916 25304
rect 32600 24942 32904 24970
rect 32680 24812 32732 24818
rect 32680 24754 32732 24760
rect 32692 24721 32720 24754
rect 32678 24712 32734 24721
rect 32404 24676 32456 24682
rect 32508 24670 32628 24698
rect 32404 24618 32456 24624
rect 32404 24336 32456 24342
rect 32404 24278 32456 24284
rect 32416 23866 32444 24278
rect 32496 24200 32548 24206
rect 32496 24142 32548 24148
rect 32508 23905 32536 24142
rect 32494 23896 32550 23905
rect 32404 23860 32456 23866
rect 32494 23831 32550 23840
rect 32404 23802 32456 23808
rect 32496 23656 32548 23662
rect 32496 23598 32548 23604
rect 32312 23520 32364 23526
rect 32508 23497 32536 23598
rect 32312 23462 32364 23468
rect 32494 23488 32550 23497
rect 32324 22642 32352 23462
rect 32494 23423 32550 23432
rect 32496 23112 32548 23118
rect 32496 23054 32548 23060
rect 32508 22681 32536 23054
rect 32494 22672 32550 22681
rect 32312 22636 32364 22642
rect 32494 22607 32550 22616
rect 32312 22578 32364 22584
rect 32600 22098 32628 24670
rect 32678 24647 32734 24656
rect 32680 24132 32732 24138
rect 32680 24074 32732 24080
rect 32692 23769 32720 24074
rect 32678 23760 32734 23769
rect 32678 23695 32734 23704
rect 32680 23656 32732 23662
rect 32678 23624 32680 23633
rect 32732 23624 32734 23633
rect 32876 23594 32904 24942
rect 33060 24410 33088 26862
rect 33324 26784 33376 26790
rect 33324 26726 33376 26732
rect 33232 26240 33284 26246
rect 33232 26182 33284 26188
rect 33244 24818 33272 26182
rect 33336 25401 33364 26726
rect 33416 26308 33468 26314
rect 33416 26250 33468 26256
rect 33322 25392 33378 25401
rect 33322 25327 33378 25336
rect 33428 24818 33456 26250
rect 33232 24812 33284 24818
rect 33232 24754 33284 24760
rect 33416 24812 33468 24818
rect 33416 24754 33468 24760
rect 33048 24404 33100 24410
rect 33048 24346 33100 24352
rect 32678 23559 32734 23568
rect 32864 23588 32916 23594
rect 32864 23530 32916 23536
rect 32680 23044 32732 23050
rect 32680 22986 32732 22992
rect 32048 22066 32168 22094
rect 32588 22092 32640 22098
rect 31944 22024 31996 22030
rect 31944 21966 31996 21972
rect 31852 21412 31904 21418
rect 31852 21354 31904 21360
rect 31850 20904 31906 20913
rect 31956 20890 31984 21966
rect 31906 20862 31984 20890
rect 31850 20839 31906 20848
rect 31864 20806 31892 20839
rect 31852 20800 31904 20806
rect 31852 20742 31904 20748
rect 31852 20392 31904 20398
rect 31852 20334 31904 20340
rect 31864 20058 31892 20334
rect 31944 20324 31996 20330
rect 31944 20266 31996 20272
rect 31956 20058 31984 20266
rect 31852 20052 31904 20058
rect 31852 19994 31904 20000
rect 31944 20052 31996 20058
rect 31944 19994 31996 20000
rect 31864 19938 31892 19994
rect 31864 19910 31984 19938
rect 31760 19848 31812 19854
rect 31760 19790 31812 19796
rect 31588 19502 31708 19530
rect 31772 19530 31800 19790
rect 31772 19502 31892 19530
rect 31484 18080 31536 18086
rect 31484 18022 31536 18028
rect 31482 16824 31538 16833
rect 31482 16759 31538 16768
rect 31496 16250 31524 16759
rect 31484 16244 31536 16250
rect 31484 16186 31536 16192
rect 31588 15706 31616 19502
rect 31760 19372 31812 19378
rect 31680 19332 31760 19360
rect 31680 18766 31708 19332
rect 31760 19314 31812 19320
rect 31758 18864 31814 18873
rect 31758 18799 31814 18808
rect 31772 18766 31800 18799
rect 31668 18760 31720 18766
rect 31668 18702 31720 18708
rect 31760 18760 31812 18766
rect 31760 18702 31812 18708
rect 31666 18456 31722 18465
rect 31666 18391 31722 18400
rect 31576 15700 31628 15706
rect 31576 15642 31628 15648
rect 31680 15502 31708 18391
rect 31864 18222 31892 19502
rect 31956 19310 31984 19910
rect 31944 19304 31996 19310
rect 31944 19246 31996 19252
rect 31944 19168 31996 19174
rect 31944 19110 31996 19116
rect 31956 18290 31984 19110
rect 31944 18284 31996 18290
rect 31944 18226 31996 18232
rect 31852 18216 31904 18222
rect 31852 18158 31904 18164
rect 31852 18080 31904 18086
rect 31852 18022 31904 18028
rect 31864 17814 31892 18022
rect 31852 17808 31904 17814
rect 31852 17750 31904 17756
rect 31852 17672 31904 17678
rect 31852 17614 31904 17620
rect 31864 17202 31892 17614
rect 31852 17196 31904 17202
rect 31852 17138 31904 17144
rect 31758 17096 31814 17105
rect 31758 17031 31814 17040
rect 31772 16590 31800 17031
rect 31760 16584 31812 16590
rect 31760 16526 31812 16532
rect 31864 15638 31892 17138
rect 31956 16182 31984 18226
rect 31944 16176 31996 16182
rect 31944 16118 31996 16124
rect 32048 15706 32076 22066
rect 32588 22034 32640 22040
rect 32404 22024 32456 22030
rect 32404 21966 32456 21972
rect 32416 21894 32444 21966
rect 32404 21888 32456 21894
rect 32404 21830 32456 21836
rect 32128 21072 32180 21078
rect 32128 21014 32180 21020
rect 32140 20806 32168 21014
rect 32416 21010 32444 21830
rect 32404 21004 32456 21010
rect 32404 20946 32456 20952
rect 32128 20800 32180 20806
rect 32416 20788 32444 20946
rect 32496 20936 32548 20942
rect 32548 20896 32628 20924
rect 32496 20878 32548 20884
rect 32416 20760 32536 20788
rect 32128 20742 32180 20748
rect 32312 20460 32364 20466
rect 32312 20402 32364 20408
rect 32220 19780 32272 19786
rect 32220 19722 32272 19728
rect 32128 19372 32180 19378
rect 32128 19314 32180 19320
rect 32036 15700 32088 15706
rect 32036 15642 32088 15648
rect 31852 15632 31904 15638
rect 31852 15574 31904 15580
rect 31668 15496 31720 15502
rect 31668 15438 31720 15444
rect 31668 15020 31720 15026
rect 31668 14962 31720 14968
rect 31392 14068 31444 14074
rect 31392 14010 31444 14016
rect 31574 13968 31630 13977
rect 31574 13903 31576 13912
rect 31628 13903 31630 13912
rect 31576 13874 31628 13880
rect 31208 13524 31260 13530
rect 31208 13466 31260 13472
rect 30932 12844 30984 12850
rect 30932 12786 30984 12792
rect 31484 12844 31536 12850
rect 31484 12786 31536 12792
rect 30493 12540 30801 12549
rect 30493 12538 30499 12540
rect 30555 12538 30579 12540
rect 30635 12538 30659 12540
rect 30715 12538 30739 12540
rect 30795 12538 30801 12540
rect 30555 12486 30557 12538
rect 30737 12486 30739 12538
rect 30493 12484 30499 12486
rect 30555 12484 30579 12486
rect 30635 12484 30659 12486
rect 30715 12484 30739 12486
rect 30795 12484 30801 12486
rect 30493 12475 30801 12484
rect 30493 11452 30801 11461
rect 30493 11450 30499 11452
rect 30555 11450 30579 11452
rect 30635 11450 30659 11452
rect 30715 11450 30739 11452
rect 30795 11450 30801 11452
rect 30555 11398 30557 11450
rect 30737 11398 30739 11450
rect 30493 11396 30499 11398
rect 30555 11396 30579 11398
rect 30635 11396 30659 11398
rect 30715 11396 30739 11398
rect 30795 11396 30801 11398
rect 30493 11387 30801 11396
rect 31496 10606 31524 12786
rect 31588 12238 31616 13874
rect 31576 12232 31628 12238
rect 31576 12174 31628 12180
rect 31484 10600 31536 10606
rect 31484 10542 31536 10548
rect 30493 10364 30801 10373
rect 30493 10362 30499 10364
rect 30555 10362 30579 10364
rect 30635 10362 30659 10364
rect 30715 10362 30739 10364
rect 30795 10362 30801 10364
rect 30555 10310 30557 10362
rect 30737 10310 30739 10362
rect 30493 10308 30499 10310
rect 30555 10308 30579 10310
rect 30635 10308 30659 10310
rect 30715 10308 30739 10310
rect 30795 10308 30801 10310
rect 30493 10299 30801 10308
rect 30493 9276 30801 9285
rect 30493 9274 30499 9276
rect 30555 9274 30579 9276
rect 30635 9274 30659 9276
rect 30715 9274 30739 9276
rect 30795 9274 30801 9276
rect 30555 9222 30557 9274
rect 30737 9222 30739 9274
rect 30493 9220 30499 9222
rect 30555 9220 30579 9222
rect 30635 9220 30659 9222
rect 30715 9220 30739 9222
rect 30795 9220 30801 9222
rect 30493 9211 30801 9220
rect 30493 8188 30801 8197
rect 30493 8186 30499 8188
rect 30555 8186 30579 8188
rect 30635 8186 30659 8188
rect 30715 8186 30739 8188
rect 30795 8186 30801 8188
rect 30555 8134 30557 8186
rect 30737 8134 30739 8186
rect 30493 8132 30499 8134
rect 30555 8132 30579 8134
rect 30635 8132 30659 8134
rect 30715 8132 30739 8134
rect 30795 8132 30801 8134
rect 30493 8123 30801 8132
rect 30493 7100 30801 7109
rect 30493 7098 30499 7100
rect 30555 7098 30579 7100
rect 30635 7098 30659 7100
rect 30715 7098 30739 7100
rect 30795 7098 30801 7100
rect 30555 7046 30557 7098
rect 30737 7046 30739 7098
rect 30493 7044 30499 7046
rect 30555 7044 30579 7046
rect 30635 7044 30659 7046
rect 30715 7044 30739 7046
rect 30795 7044 30801 7046
rect 30493 7035 30801 7044
rect 30288 6724 30340 6730
rect 30288 6666 30340 6672
rect 31496 6322 31524 10542
rect 31680 8090 31708 14962
rect 32140 14958 32168 19314
rect 32232 17678 32260 19722
rect 32324 19446 32352 20402
rect 32312 19440 32364 19446
rect 32312 19382 32364 19388
rect 32312 19304 32364 19310
rect 32312 19246 32364 19252
rect 32220 17672 32272 17678
rect 32220 17614 32272 17620
rect 32220 17536 32272 17542
rect 32324 17490 32352 19246
rect 32402 19000 32458 19009
rect 32402 18935 32458 18944
rect 32416 18902 32444 18935
rect 32404 18896 32456 18902
rect 32404 18838 32456 18844
rect 32416 18426 32444 18838
rect 32404 18420 32456 18426
rect 32404 18362 32456 18368
rect 32272 17484 32352 17490
rect 32220 17478 32352 17484
rect 32232 17462 32352 17478
rect 32232 17270 32260 17462
rect 32416 17320 32444 18362
rect 32508 18358 32536 20760
rect 32496 18352 32548 18358
rect 32496 18294 32548 18300
rect 32324 17292 32444 17320
rect 32220 17264 32272 17270
rect 32220 17206 32272 17212
rect 32324 17116 32352 17292
rect 32508 17252 32536 18294
rect 32232 17088 32352 17116
rect 32416 17224 32536 17252
rect 32232 16522 32260 17088
rect 32416 16980 32444 17224
rect 32496 17128 32548 17134
rect 32496 17070 32548 17076
rect 32324 16952 32444 16980
rect 32220 16516 32272 16522
rect 32220 16458 32272 16464
rect 32324 15570 32352 16952
rect 32402 16280 32458 16289
rect 32402 16215 32404 16224
rect 32456 16215 32458 16224
rect 32404 16186 32456 16192
rect 32312 15564 32364 15570
rect 32312 15506 32364 15512
rect 32128 14952 32180 14958
rect 32128 14894 32180 14900
rect 32508 14618 32536 17070
rect 32496 14612 32548 14618
rect 32496 14554 32548 14560
rect 32496 13864 32548 13870
rect 32496 13806 32548 13812
rect 31850 13560 31906 13569
rect 31850 13495 31852 13504
rect 31904 13495 31906 13504
rect 31852 13466 31904 13472
rect 31760 13320 31812 13326
rect 31760 13262 31812 13268
rect 31668 8084 31720 8090
rect 31668 8026 31720 8032
rect 31484 6316 31536 6322
rect 31484 6258 31536 6264
rect 30493 6012 30801 6021
rect 30493 6010 30499 6012
rect 30555 6010 30579 6012
rect 30635 6010 30659 6012
rect 30715 6010 30739 6012
rect 30795 6010 30801 6012
rect 30555 5958 30557 6010
rect 30737 5958 30739 6010
rect 30493 5956 30499 5958
rect 30555 5956 30579 5958
rect 30635 5956 30659 5958
rect 30715 5956 30739 5958
rect 30795 5956 30801 5958
rect 30493 5947 30801 5956
rect 31300 5704 31352 5710
rect 31300 5646 31352 5652
rect 31024 5024 31076 5030
rect 31024 4966 31076 4972
rect 31208 5024 31260 5030
rect 31208 4966 31260 4972
rect 30493 4924 30801 4933
rect 30493 4922 30499 4924
rect 30555 4922 30579 4924
rect 30635 4922 30659 4924
rect 30715 4922 30739 4924
rect 30795 4922 30801 4924
rect 30555 4870 30557 4922
rect 30737 4870 30739 4922
rect 30493 4868 30499 4870
rect 30555 4868 30579 4870
rect 30635 4868 30659 4870
rect 30715 4868 30739 4870
rect 30795 4868 30801 4870
rect 30493 4859 30801 4868
rect 30840 4548 30892 4554
rect 30840 4490 30892 4496
rect 30104 4072 30156 4078
rect 30104 4014 30156 4020
rect 30116 3738 30144 4014
rect 30493 3836 30801 3845
rect 30493 3834 30499 3836
rect 30555 3834 30579 3836
rect 30635 3834 30659 3836
rect 30715 3834 30739 3836
rect 30795 3834 30801 3836
rect 30555 3782 30557 3834
rect 30737 3782 30739 3834
rect 30493 3780 30499 3782
rect 30555 3780 30579 3782
rect 30635 3780 30659 3782
rect 30715 3780 30739 3782
rect 30795 3780 30801 3782
rect 30493 3771 30801 3780
rect 30104 3732 30156 3738
rect 30104 3674 30156 3680
rect 29644 3528 29696 3534
rect 29644 3470 29696 3476
rect 30380 3528 30432 3534
rect 30380 3470 30432 3476
rect 29656 3058 29684 3470
rect 29920 3120 29972 3126
rect 29920 3062 29972 3068
rect 29644 3052 29696 3058
rect 29644 2994 29696 3000
rect 29932 2990 29960 3062
rect 29092 2984 29144 2990
rect 29092 2926 29144 2932
rect 29920 2984 29972 2990
rect 29920 2926 29972 2932
rect 30288 2984 30340 2990
rect 30288 2926 30340 2932
rect 29104 2514 29132 2926
rect 30196 2848 30248 2854
rect 30196 2790 30248 2796
rect 29092 2508 29144 2514
rect 29092 2450 29144 2456
rect 27712 2440 27764 2446
rect 27712 2382 27764 2388
rect 28540 2440 28592 2446
rect 28540 2382 28592 2388
rect 29000 2440 29052 2446
rect 29000 2382 29052 2388
rect 30208 2378 30236 2790
rect 30196 2372 30248 2378
rect 30196 2314 30248 2320
rect 26272 2204 26580 2213
rect 26272 2202 26278 2204
rect 26334 2202 26358 2204
rect 26414 2202 26438 2204
rect 26494 2202 26518 2204
rect 26574 2202 26580 2204
rect 26334 2150 26336 2202
rect 26516 2150 26518 2202
rect 26272 2148 26278 2150
rect 26334 2148 26358 2150
rect 26414 2148 26438 2150
rect 26494 2148 26518 2150
rect 26574 2148 26580 2150
rect 26272 2139 26580 2148
rect 30300 800 30328 2926
rect 30392 2514 30420 3470
rect 30493 2748 30801 2757
rect 30493 2746 30499 2748
rect 30555 2746 30579 2748
rect 30635 2746 30659 2748
rect 30715 2746 30739 2748
rect 30795 2746 30801 2748
rect 30555 2694 30557 2746
rect 30737 2694 30739 2746
rect 30493 2692 30499 2694
rect 30555 2692 30579 2694
rect 30635 2692 30659 2694
rect 30715 2692 30739 2694
rect 30795 2692 30801 2694
rect 30493 2683 30801 2692
rect 30852 2650 30880 4490
rect 31036 3466 31064 4966
rect 31220 3602 31248 4966
rect 31312 4146 31340 5646
rect 31300 4140 31352 4146
rect 31300 4082 31352 4088
rect 31668 3936 31720 3942
rect 31668 3878 31720 3884
rect 31208 3596 31260 3602
rect 31208 3538 31260 3544
rect 31300 3596 31352 3602
rect 31300 3538 31352 3544
rect 31024 3460 31076 3466
rect 31024 3402 31076 3408
rect 31312 3126 31340 3538
rect 31300 3120 31352 3126
rect 31300 3062 31352 3068
rect 30840 2644 30892 2650
rect 30840 2586 30892 2592
rect 31680 2514 31708 3878
rect 31772 3670 31800 13262
rect 32508 12442 32536 13806
rect 32600 13530 32628 20896
rect 32692 20777 32720 22986
rect 33140 22636 33192 22642
rect 33192 22596 33364 22624
rect 33140 22578 33192 22584
rect 32772 22024 32824 22030
rect 32772 21966 32824 21972
rect 32784 21554 32812 21966
rect 33048 21684 33100 21690
rect 33048 21626 33100 21632
rect 32772 21548 32824 21554
rect 32772 21490 32824 21496
rect 32678 20768 32734 20777
rect 32678 20703 32734 20712
rect 32784 20534 32812 21490
rect 33060 21185 33088 21626
rect 33140 21548 33192 21554
rect 33140 21490 33192 21496
rect 33046 21176 33102 21185
rect 33046 21111 33102 21120
rect 32956 20800 33008 20806
rect 32956 20742 33008 20748
rect 32772 20528 32824 20534
rect 32772 20470 32824 20476
rect 32968 20380 32996 20742
rect 32876 20352 32996 20380
rect 32772 19780 32824 19786
rect 32772 19722 32824 19728
rect 32680 18828 32732 18834
rect 32680 18770 32732 18776
rect 32692 17066 32720 18770
rect 32680 17060 32732 17066
rect 32680 17002 32732 17008
rect 32680 16516 32732 16522
rect 32680 16458 32732 16464
rect 32692 15978 32720 16458
rect 32680 15972 32732 15978
rect 32680 15914 32732 15920
rect 32680 15632 32732 15638
rect 32680 15574 32732 15580
rect 32692 15502 32720 15574
rect 32680 15496 32732 15502
rect 32680 15438 32732 15444
rect 32784 15162 32812 19722
rect 32876 18290 32904 20352
rect 32956 19780 33008 19786
rect 32956 19722 33008 19728
rect 32968 18426 32996 19722
rect 33048 19712 33100 19718
rect 33048 19654 33100 19660
rect 33060 18698 33088 19654
rect 33048 18692 33100 18698
rect 33048 18634 33100 18640
rect 32956 18420 33008 18426
rect 32956 18362 33008 18368
rect 32864 18284 32916 18290
rect 32864 18226 32916 18232
rect 33046 18048 33102 18057
rect 33046 17983 33102 17992
rect 32956 17536 33008 17542
rect 32956 17478 33008 17484
rect 32864 16652 32916 16658
rect 32864 16594 32916 16600
rect 32772 15156 32824 15162
rect 32772 15098 32824 15104
rect 32772 15020 32824 15026
rect 32772 14962 32824 14968
rect 32680 14340 32732 14346
rect 32680 14282 32732 14288
rect 32588 13524 32640 13530
rect 32588 13466 32640 13472
rect 32496 12436 32548 12442
rect 32496 12378 32548 12384
rect 32692 10810 32720 14282
rect 32680 10804 32732 10810
rect 32680 10746 32732 10752
rect 32496 8968 32548 8974
rect 32496 8910 32548 8916
rect 32508 8498 32536 8910
rect 32496 8492 32548 8498
rect 32496 8434 32548 8440
rect 31944 6792 31996 6798
rect 31944 6734 31996 6740
rect 31852 5704 31904 5710
rect 31852 5646 31904 5652
rect 31864 4690 31892 5646
rect 31852 4684 31904 4690
rect 31852 4626 31904 4632
rect 31852 4072 31904 4078
rect 31852 4014 31904 4020
rect 31760 3664 31812 3670
rect 31760 3606 31812 3612
rect 30380 2508 30432 2514
rect 30380 2450 30432 2456
rect 30932 2508 30984 2514
rect 30932 2450 30984 2456
rect 31668 2508 31720 2514
rect 31668 2450 31720 2456
rect 30944 800 30972 2450
rect -10 200 102 800
rect 634 200 746 800
rect 1278 200 1390 800
rect 1922 200 2034 800
rect 2566 200 2678 800
rect 3210 200 3322 800
rect 3854 200 3966 800
rect 4498 200 4610 800
rect 5142 200 5254 800
rect 6430 200 6542 800
rect 7074 200 7186 800
rect 7718 200 7830 800
rect 8362 200 8474 800
rect 9006 200 9118 800
rect 9650 200 9762 800
rect 10294 200 10406 800
rect 10938 200 11050 800
rect 11582 200 11694 800
rect 12870 200 12982 800
rect 13514 200 13626 800
rect 14158 200 14270 800
rect 14802 200 14914 800
rect 15446 200 15558 800
rect 16090 200 16202 800
rect 16734 200 16846 800
rect 17378 200 17490 800
rect 18022 200 18134 800
rect 19310 200 19422 800
rect 19954 200 20066 800
rect 20598 200 20710 800
rect 21242 200 21354 800
rect 21886 200 21998 800
rect 22530 200 22642 800
rect 23174 200 23286 800
rect 23818 200 23930 800
rect 24462 200 24574 800
rect 25750 200 25862 800
rect 26394 200 26506 800
rect 27038 200 27150 800
rect 27682 200 27794 800
rect 28326 200 28438 800
rect 28970 200 29082 800
rect 29614 200 29726 800
rect 30258 200 30370 800
rect 30902 200 31014 800
rect 31864 105 31892 4014
rect 31956 3738 31984 6734
rect 32680 6656 32732 6662
rect 32680 6598 32732 6604
rect 32036 5704 32088 5710
rect 32036 5646 32088 5652
rect 32048 5234 32076 5646
rect 32128 5636 32180 5642
rect 32128 5578 32180 5584
rect 32036 5228 32088 5234
rect 32036 5170 32088 5176
rect 31944 3732 31996 3738
rect 31944 3674 31996 3680
rect 32140 2582 32168 5578
rect 32692 4690 32720 6598
rect 32680 4684 32732 4690
rect 32680 4626 32732 4632
rect 32680 4072 32732 4078
rect 32680 4014 32732 4020
rect 32496 3392 32548 3398
rect 32496 3334 32548 3340
rect 32508 3126 32536 3334
rect 32692 3194 32720 4014
rect 32680 3188 32732 3194
rect 32680 3130 32732 3136
rect 32496 3120 32548 3126
rect 32496 3062 32548 3068
rect 32220 2916 32272 2922
rect 32220 2858 32272 2864
rect 32128 2576 32180 2582
rect 32128 2518 32180 2524
rect 32232 800 32260 2858
rect 32784 2854 32812 14962
rect 32876 11762 32904 16594
rect 32968 16114 32996 17478
rect 32956 16108 33008 16114
rect 32956 16050 33008 16056
rect 33060 15162 33088 17983
rect 33152 15706 33180 21490
rect 33232 20052 33284 20058
rect 33232 19994 33284 20000
rect 33244 18766 33272 19994
rect 33336 19786 33364 22596
rect 33428 22094 33456 24754
rect 33520 24682 33548 26930
rect 33612 25265 33640 26998
rect 33692 26988 33744 26994
rect 33692 26930 33744 26936
rect 33704 26586 33732 26930
rect 34244 26852 34296 26858
rect 34244 26794 34296 26800
rect 33692 26580 33744 26586
rect 33692 26522 33744 26528
rect 33598 25256 33654 25265
rect 33598 25191 33654 25200
rect 34060 25220 34112 25226
rect 33612 24886 33640 25191
rect 34060 25162 34112 25168
rect 33600 24880 33652 24886
rect 33600 24822 33652 24828
rect 34072 24818 34100 25162
rect 34060 24812 34112 24818
rect 34060 24754 34112 24760
rect 33508 24676 33560 24682
rect 33508 24618 33560 24624
rect 33428 22066 33548 22094
rect 33416 19916 33468 19922
rect 33416 19858 33468 19864
rect 33324 19780 33376 19786
rect 33324 19722 33376 19728
rect 33232 18760 33284 18766
rect 33232 18702 33284 18708
rect 33232 18216 33284 18222
rect 33284 18164 33364 18170
rect 33232 18158 33364 18164
rect 33244 18142 33364 18158
rect 33232 17604 33284 17610
rect 33232 17546 33284 17552
rect 33140 15700 33192 15706
rect 33140 15642 33192 15648
rect 33048 15156 33100 15162
rect 33048 15098 33100 15104
rect 33140 12776 33192 12782
rect 33140 12718 33192 12724
rect 32864 11756 32916 11762
rect 32864 11698 32916 11704
rect 33152 11354 33180 12718
rect 33244 11762 33272 17546
rect 33336 16114 33364 18142
rect 33324 16108 33376 16114
rect 33324 16050 33376 16056
rect 33324 12300 33376 12306
rect 33324 12242 33376 12248
rect 33232 11756 33284 11762
rect 33232 11698 33284 11704
rect 33140 11348 33192 11354
rect 33140 11290 33192 11296
rect 33336 10674 33364 12242
rect 33428 11354 33456 19858
rect 33520 16250 33548 22066
rect 33600 21344 33652 21350
rect 33600 21286 33652 21292
rect 33612 18290 33640 21286
rect 33692 20460 33744 20466
rect 33692 20402 33744 20408
rect 33704 18970 33732 20402
rect 33784 20256 33836 20262
rect 33784 20198 33836 20204
rect 33796 19990 33824 20198
rect 33784 19984 33836 19990
rect 33784 19926 33836 19932
rect 33692 18964 33744 18970
rect 33692 18906 33744 18912
rect 33692 18624 33744 18630
rect 33692 18566 33744 18572
rect 33704 18358 33732 18566
rect 33692 18352 33744 18358
rect 33692 18294 33744 18300
rect 33600 18284 33652 18290
rect 33600 18226 33652 18232
rect 33508 16244 33560 16250
rect 33508 16186 33560 16192
rect 33612 15026 33640 18226
rect 33704 15609 33732 18294
rect 33796 16998 33824 19926
rect 33968 18080 34020 18086
rect 33968 18022 34020 18028
rect 33784 16992 33836 16998
rect 33784 16934 33836 16940
rect 33690 15600 33746 15609
rect 33690 15535 33746 15544
rect 33796 15502 33824 16934
rect 33980 15570 34008 18022
rect 34072 15706 34100 24754
rect 34152 24268 34204 24274
rect 34152 24210 34204 24216
rect 34164 20448 34192 24210
rect 34256 22778 34284 26794
rect 34713 26140 35021 26149
rect 34713 26138 34719 26140
rect 34775 26138 34799 26140
rect 34855 26138 34879 26140
rect 34935 26138 34959 26140
rect 35015 26138 35021 26140
rect 34775 26086 34777 26138
rect 34957 26086 34959 26138
rect 34713 26084 34719 26086
rect 34775 26084 34799 26086
rect 34855 26084 34879 26086
rect 34935 26084 34959 26086
rect 35015 26084 35021 26086
rect 34713 26075 35021 26084
rect 34334 25936 34390 25945
rect 34334 25871 34336 25880
rect 34388 25871 34390 25880
rect 34336 25842 34388 25848
rect 34334 25256 34390 25265
rect 34334 25191 34336 25200
rect 34388 25191 34390 25200
rect 34336 25162 34388 25168
rect 34713 25052 35021 25061
rect 34713 25050 34719 25052
rect 34775 25050 34799 25052
rect 34855 25050 34879 25052
rect 34935 25050 34959 25052
rect 35015 25050 35021 25052
rect 34775 24998 34777 25050
rect 34957 24998 34959 25050
rect 34713 24996 34719 24998
rect 34775 24996 34799 24998
rect 34855 24996 34879 24998
rect 34935 24996 34959 24998
rect 35015 24996 35021 24998
rect 34713 24987 35021 24996
rect 34426 24576 34482 24585
rect 34426 24511 34482 24520
rect 34336 24132 34388 24138
rect 34336 24074 34388 24080
rect 34348 23769 34376 24074
rect 34440 23798 34468 24511
rect 34713 23964 35021 23973
rect 34713 23962 34719 23964
rect 34775 23962 34799 23964
rect 34855 23962 34879 23964
rect 34935 23962 34959 23964
rect 35015 23962 35021 23964
rect 34775 23910 34777 23962
rect 34957 23910 34959 23962
rect 34713 23908 34719 23910
rect 34775 23908 34799 23910
rect 34855 23908 34879 23910
rect 34935 23908 34959 23910
rect 35015 23908 35021 23910
rect 34713 23899 35021 23908
rect 34428 23792 34480 23798
rect 34334 23760 34390 23769
rect 34428 23734 34480 23740
rect 34334 23695 34390 23704
rect 34334 23216 34390 23225
rect 34334 23151 34336 23160
rect 34388 23151 34390 23160
rect 34336 23122 34388 23128
rect 34520 22976 34572 22982
rect 34520 22918 34572 22924
rect 34334 22808 34390 22817
rect 34244 22772 34296 22778
rect 34334 22743 34390 22752
rect 34244 22714 34296 22720
rect 34348 22642 34376 22743
rect 34336 22636 34388 22642
rect 34336 22578 34388 22584
rect 34336 20868 34388 20874
rect 34336 20810 34388 20816
rect 34242 20632 34298 20641
rect 34242 20567 34244 20576
rect 34296 20567 34298 20576
rect 34244 20538 34296 20544
rect 34348 20505 34376 20810
rect 34334 20496 34390 20505
rect 34244 20460 34296 20466
rect 34164 20420 34244 20448
rect 34334 20431 34390 20440
rect 34244 20402 34296 20408
rect 34336 19848 34388 19854
rect 34334 19816 34336 19825
rect 34388 19816 34390 19825
rect 34334 19751 34390 19760
rect 34336 19304 34388 19310
rect 34336 19246 34388 19252
rect 34348 19145 34376 19246
rect 34334 19136 34390 19145
rect 34334 19071 34390 19080
rect 34334 17776 34390 17785
rect 34334 17711 34336 17720
rect 34388 17711 34390 17720
rect 34336 17682 34388 17688
rect 34336 17128 34388 17134
rect 34334 17096 34336 17105
rect 34388 17096 34390 17105
rect 34334 17031 34390 17040
rect 34532 16250 34560 22918
rect 34713 22876 35021 22885
rect 34713 22874 34719 22876
rect 34775 22874 34799 22876
rect 34855 22874 34879 22876
rect 34935 22874 34959 22876
rect 35015 22874 35021 22876
rect 34775 22822 34777 22874
rect 34957 22822 34959 22874
rect 34713 22820 34719 22822
rect 34775 22820 34799 22822
rect 34855 22820 34879 22822
rect 34935 22820 34959 22822
rect 35015 22820 35021 22822
rect 34713 22811 35021 22820
rect 34713 21788 35021 21797
rect 34713 21786 34719 21788
rect 34775 21786 34799 21788
rect 34855 21786 34879 21788
rect 34935 21786 34959 21788
rect 35015 21786 35021 21788
rect 34775 21734 34777 21786
rect 34957 21734 34959 21786
rect 34713 21732 34719 21734
rect 34775 21732 34799 21734
rect 34855 21732 34879 21734
rect 34935 21732 34959 21734
rect 35015 21732 35021 21734
rect 34713 21723 35021 21732
rect 34713 20700 35021 20709
rect 34713 20698 34719 20700
rect 34775 20698 34799 20700
rect 34855 20698 34879 20700
rect 34935 20698 34959 20700
rect 35015 20698 35021 20700
rect 34775 20646 34777 20698
rect 34957 20646 34959 20698
rect 34713 20644 34719 20646
rect 34775 20644 34799 20646
rect 34855 20644 34879 20646
rect 34935 20644 34959 20646
rect 35015 20644 35021 20646
rect 34713 20635 35021 20644
rect 34713 19612 35021 19621
rect 34713 19610 34719 19612
rect 34775 19610 34799 19612
rect 34855 19610 34879 19612
rect 34935 19610 34959 19612
rect 35015 19610 35021 19612
rect 34775 19558 34777 19610
rect 34957 19558 34959 19610
rect 34713 19556 34719 19558
rect 34775 19556 34799 19558
rect 34855 19556 34879 19558
rect 34935 19556 34959 19558
rect 35015 19556 35021 19558
rect 34713 19547 35021 19556
rect 34713 18524 35021 18533
rect 34713 18522 34719 18524
rect 34775 18522 34799 18524
rect 34855 18522 34879 18524
rect 34935 18522 34959 18524
rect 35015 18522 35021 18524
rect 34775 18470 34777 18522
rect 34957 18470 34959 18522
rect 34713 18468 34719 18470
rect 34775 18468 34799 18470
rect 34855 18468 34879 18470
rect 34935 18468 34959 18470
rect 35015 18468 35021 18470
rect 34713 18459 35021 18468
rect 34713 17436 35021 17445
rect 34713 17434 34719 17436
rect 34775 17434 34799 17436
rect 34855 17434 34879 17436
rect 34935 17434 34959 17436
rect 35015 17434 35021 17436
rect 34775 17382 34777 17434
rect 34957 17382 34959 17434
rect 34713 17380 34719 17382
rect 34775 17380 34799 17382
rect 34855 17380 34879 17382
rect 34935 17380 34959 17382
rect 35015 17380 35021 17382
rect 34713 17371 35021 17380
rect 35164 16516 35216 16522
rect 35164 16458 35216 16464
rect 35176 16425 35204 16458
rect 35162 16416 35218 16425
rect 34713 16348 35021 16357
rect 35162 16351 35218 16360
rect 34713 16346 34719 16348
rect 34775 16346 34799 16348
rect 34855 16346 34879 16348
rect 34935 16346 34959 16348
rect 35015 16346 35021 16348
rect 34775 16294 34777 16346
rect 34957 16294 34959 16346
rect 34713 16292 34719 16294
rect 34775 16292 34799 16294
rect 34855 16292 34879 16294
rect 34935 16292 34959 16294
rect 35015 16292 35021 16294
rect 34713 16283 35021 16292
rect 34520 16244 34572 16250
rect 34520 16186 34572 16192
rect 34060 15700 34112 15706
rect 34060 15642 34112 15648
rect 33968 15564 34020 15570
rect 33968 15506 34020 15512
rect 33784 15496 33836 15502
rect 33784 15438 33836 15444
rect 34244 15428 34296 15434
rect 34244 15370 34296 15376
rect 33782 15056 33838 15065
rect 33600 15020 33652 15026
rect 33782 14991 33784 15000
rect 33600 14962 33652 14968
rect 33836 14991 33838 15000
rect 33784 14962 33836 14968
rect 33508 14272 33560 14278
rect 33508 14214 33560 14220
rect 33416 11348 33468 11354
rect 33416 11290 33468 11296
rect 33520 11150 33548 14214
rect 33598 13560 33654 13569
rect 33598 13495 33600 13504
rect 33652 13495 33654 13504
rect 33600 13466 33652 13472
rect 33782 13424 33838 13433
rect 33782 13359 33838 13368
rect 33796 13326 33824 13359
rect 33784 13320 33836 13326
rect 33784 13262 33836 13268
rect 33966 11792 34022 11801
rect 33966 11727 33968 11736
rect 34020 11727 34022 11736
rect 33968 11698 34020 11704
rect 33508 11144 33560 11150
rect 33508 11086 33560 11092
rect 33324 10668 33376 10674
rect 33324 10610 33376 10616
rect 33140 8084 33192 8090
rect 33140 8026 33192 8032
rect 33048 5160 33100 5166
rect 33048 5102 33100 5108
rect 33060 4185 33088 5102
rect 33046 4176 33102 4185
rect 33046 4111 33102 4120
rect 33152 4010 33180 8026
rect 33324 7880 33376 7886
rect 33324 7822 33376 7828
rect 33232 7200 33284 7206
rect 33232 7142 33284 7148
rect 33244 6866 33272 7142
rect 33232 6860 33284 6866
rect 33232 6802 33284 6808
rect 33336 6254 33364 7822
rect 33520 7410 33548 11086
rect 34256 10266 34284 15370
rect 34713 15260 35021 15269
rect 34713 15258 34719 15260
rect 34775 15258 34799 15260
rect 34855 15258 34879 15260
rect 34935 15258 34959 15260
rect 35015 15258 35021 15260
rect 34775 15206 34777 15258
rect 34957 15206 34959 15258
rect 34713 15204 34719 15206
rect 34775 15204 34799 15206
rect 34855 15204 34879 15206
rect 34935 15204 34959 15206
rect 35015 15204 35021 15206
rect 34713 15195 35021 15204
rect 34336 14408 34388 14414
rect 34334 14376 34336 14385
rect 34388 14376 34390 14385
rect 34334 14311 34390 14320
rect 34713 14172 35021 14181
rect 34713 14170 34719 14172
rect 34775 14170 34799 14172
rect 34855 14170 34879 14172
rect 34935 14170 34959 14172
rect 35015 14170 35021 14172
rect 34775 14118 34777 14170
rect 34957 14118 34959 14170
rect 34713 14116 34719 14118
rect 34775 14116 34799 14118
rect 34855 14116 34879 14118
rect 34935 14116 34959 14118
rect 35015 14116 35021 14118
rect 34713 14107 35021 14116
rect 34336 13864 34388 13870
rect 34336 13806 34388 13812
rect 34348 13705 34376 13806
rect 34334 13696 34390 13705
rect 34334 13631 34390 13640
rect 34713 13084 35021 13093
rect 34713 13082 34719 13084
rect 34775 13082 34799 13084
rect 34855 13082 34879 13084
rect 34935 13082 34959 13084
rect 35015 13082 35021 13084
rect 34775 13030 34777 13082
rect 34957 13030 34959 13082
rect 34713 13028 34719 13030
rect 34775 13028 34799 13030
rect 34855 13028 34879 13030
rect 34935 13028 34959 13030
rect 35015 13028 35021 13030
rect 34713 13019 35021 13028
rect 34336 12912 34388 12918
rect 34334 12880 34336 12889
rect 34388 12880 34390 12889
rect 34334 12815 34390 12824
rect 34334 12336 34390 12345
rect 34334 12271 34336 12280
rect 34388 12271 34390 12280
rect 34336 12242 34388 12248
rect 34713 11996 35021 12005
rect 34713 11994 34719 11996
rect 34775 11994 34799 11996
rect 34855 11994 34879 11996
rect 34935 11994 34959 11996
rect 35015 11994 35021 11996
rect 34775 11942 34777 11994
rect 34957 11942 34959 11994
rect 34713 11940 34719 11942
rect 34775 11940 34799 11942
rect 34855 11940 34879 11942
rect 34935 11940 34959 11942
rect 35015 11940 35021 11942
rect 34713 11931 35021 11940
rect 34713 10908 35021 10917
rect 34713 10906 34719 10908
rect 34775 10906 34799 10908
rect 34855 10906 34879 10908
rect 34935 10906 34959 10908
rect 35015 10906 35021 10908
rect 34775 10854 34777 10906
rect 34957 10854 34959 10906
rect 34713 10852 34719 10854
rect 34775 10852 34799 10854
rect 34855 10852 34879 10854
rect 34935 10852 34959 10854
rect 35015 10852 35021 10854
rect 34713 10843 35021 10852
rect 34244 10260 34296 10266
rect 34244 10202 34296 10208
rect 34060 10056 34112 10062
rect 34060 9998 34112 10004
rect 34072 9625 34100 9998
rect 34713 9820 35021 9829
rect 34713 9818 34719 9820
rect 34775 9818 34799 9820
rect 34855 9818 34879 9820
rect 34935 9818 34959 9820
rect 35015 9818 35021 9820
rect 34775 9766 34777 9818
rect 34957 9766 34959 9818
rect 34713 9764 34719 9766
rect 34775 9764 34799 9766
rect 34855 9764 34879 9766
rect 34935 9764 34959 9766
rect 35015 9764 35021 9766
rect 34713 9755 35021 9764
rect 34058 9616 34114 9625
rect 34058 9551 34114 9560
rect 34334 8936 34390 8945
rect 34334 8871 34390 8880
rect 34348 8566 34376 8871
rect 34713 8732 35021 8741
rect 34713 8730 34719 8732
rect 34775 8730 34799 8732
rect 34855 8730 34879 8732
rect 34935 8730 34959 8732
rect 35015 8730 35021 8732
rect 34775 8678 34777 8730
rect 34957 8678 34959 8730
rect 34713 8676 34719 8678
rect 34775 8676 34799 8678
rect 34855 8676 34879 8678
rect 34935 8676 34959 8678
rect 35015 8676 35021 8678
rect 34713 8667 35021 8676
rect 34336 8560 34388 8566
rect 34336 8502 34388 8508
rect 33876 8424 33928 8430
rect 33876 8366 33928 8372
rect 33888 8090 33916 8366
rect 33876 8084 33928 8090
rect 33876 8026 33928 8032
rect 33784 7880 33836 7886
rect 33784 7822 33836 7828
rect 33508 7404 33560 7410
rect 33508 7346 33560 7352
rect 33520 6914 33548 7346
rect 33428 6886 33548 6914
rect 33324 6248 33376 6254
rect 33324 6190 33376 6196
rect 33140 4004 33192 4010
rect 33140 3946 33192 3952
rect 33152 3670 33180 3946
rect 33140 3664 33192 3670
rect 33140 3606 33192 3612
rect 32772 2848 32824 2854
rect 32772 2790 32824 2796
rect 32864 2508 32916 2514
rect 32864 2450 32916 2456
rect 32876 800 32904 2450
rect 33428 2310 33456 6886
rect 33796 3602 33824 7822
rect 34713 7644 35021 7653
rect 34713 7642 34719 7644
rect 34775 7642 34799 7644
rect 34855 7642 34879 7644
rect 34935 7642 34959 7644
rect 35015 7642 35021 7644
rect 34775 7590 34777 7642
rect 34957 7590 34959 7642
rect 34713 7588 34719 7590
rect 34775 7588 34799 7590
rect 34855 7588 34879 7590
rect 34935 7588 34959 7590
rect 35015 7588 35021 7590
rect 34713 7579 35021 7588
rect 33968 7200 34020 7206
rect 33968 7142 34020 7148
rect 33980 6730 34008 7142
rect 34334 6896 34390 6905
rect 34334 6831 34336 6840
rect 34388 6831 34390 6840
rect 34336 6802 34388 6808
rect 33968 6724 34020 6730
rect 33968 6666 34020 6672
rect 34713 6556 35021 6565
rect 34713 6554 34719 6556
rect 34775 6554 34799 6556
rect 34855 6554 34879 6556
rect 34935 6554 34959 6556
rect 35015 6554 35021 6556
rect 34775 6502 34777 6554
rect 34957 6502 34959 6554
rect 34713 6500 34719 6502
rect 34775 6500 34799 6502
rect 34855 6500 34879 6502
rect 34935 6500 34959 6502
rect 35015 6500 35021 6502
rect 34713 6491 35021 6500
rect 34336 6248 34388 6254
rect 34336 6190 34388 6196
rect 34060 5296 34112 5302
rect 34060 5238 34112 5244
rect 34072 3738 34100 5238
rect 34348 4865 34376 6190
rect 34612 5636 34664 5642
rect 34612 5578 34664 5584
rect 34334 4856 34390 4865
rect 34334 4791 34390 4800
rect 34336 4548 34388 4554
rect 34336 4490 34388 4496
rect 34060 3732 34112 3738
rect 34060 3674 34112 3680
rect 33784 3596 33836 3602
rect 33784 3538 33836 3544
rect 33508 3528 33560 3534
rect 34348 3505 34376 4490
rect 34520 4480 34572 4486
rect 34520 4422 34572 4428
rect 33508 3470 33560 3476
rect 34334 3496 34390 3505
rect 33520 2990 33548 3470
rect 34334 3431 34390 3440
rect 33508 2984 33560 2990
rect 33508 2926 33560 2932
rect 33416 2304 33468 2310
rect 33416 2246 33468 2252
rect 34532 1154 34560 4422
rect 34520 1148 34572 1154
rect 34520 1090 34572 1096
rect 34624 921 34652 5578
rect 34713 5468 35021 5477
rect 34713 5466 34719 5468
rect 34775 5466 34799 5468
rect 34855 5466 34879 5468
rect 34935 5466 34959 5468
rect 35015 5466 35021 5468
rect 34775 5414 34777 5466
rect 34957 5414 34959 5466
rect 34713 5412 34719 5414
rect 34775 5412 34799 5414
rect 34855 5412 34879 5414
rect 34935 5412 34959 5414
rect 35015 5412 35021 5414
rect 34713 5403 35021 5412
rect 34713 4380 35021 4389
rect 34713 4378 34719 4380
rect 34775 4378 34799 4380
rect 34855 4378 34879 4380
rect 34935 4378 34959 4380
rect 35015 4378 35021 4380
rect 34775 4326 34777 4378
rect 34957 4326 34959 4378
rect 34713 4324 34719 4326
rect 34775 4324 34799 4326
rect 34855 4324 34879 4326
rect 34935 4324 34959 4326
rect 35015 4324 35021 4326
rect 34713 4315 35021 4324
rect 35440 4072 35492 4078
rect 35440 4014 35492 4020
rect 34713 3292 35021 3301
rect 34713 3290 34719 3292
rect 34775 3290 34799 3292
rect 34855 3290 34879 3292
rect 34935 3290 34959 3292
rect 35015 3290 35021 3292
rect 34775 3238 34777 3290
rect 34957 3238 34959 3290
rect 34713 3236 34719 3238
rect 34775 3236 34799 3238
rect 34855 3236 34879 3238
rect 34935 3236 34959 3238
rect 35015 3236 35021 3238
rect 34713 3227 35021 3236
rect 34713 2204 35021 2213
rect 34713 2202 34719 2204
rect 34775 2202 34799 2204
rect 34855 2202 34879 2204
rect 34935 2202 34959 2204
rect 35015 2202 35021 2204
rect 34775 2150 34777 2202
rect 34957 2150 34959 2202
rect 34713 2148 34719 2150
rect 34775 2148 34799 2150
rect 34855 2148 34879 2150
rect 34935 2148 34959 2150
rect 35015 2148 35021 2150
rect 34713 2139 35021 2148
rect 34796 1148 34848 1154
rect 34796 1090 34848 1096
rect 34610 912 34666 921
rect 34610 847 34666 856
rect 34808 800 34836 1090
rect 35452 800 35480 4014
rect 35900 3460 35952 3466
rect 35900 3402 35952 3408
rect 35912 2145 35940 3402
rect 35898 2136 35954 2145
rect 35898 2071 35954 2080
rect 32190 200 32302 800
rect 32834 200 32946 800
rect 33478 200 33590 800
rect 34122 200 34234 800
rect 34766 200 34878 800
rect 35410 200 35522 800
rect 31850 96 31906 105
rect 31850 31 31906 40
<< via2 >>
rect 2778 41520 2834 41576
rect 3422 40840 3478 40896
rect 2042 37440 2098 37496
rect 5176 39738 5232 39740
rect 5256 39738 5312 39740
rect 5336 39738 5392 39740
rect 5416 39738 5472 39740
rect 5176 39686 5222 39738
rect 5222 39686 5232 39738
rect 5256 39686 5286 39738
rect 5286 39686 5298 39738
rect 5298 39686 5312 39738
rect 5336 39686 5350 39738
rect 5350 39686 5362 39738
rect 5362 39686 5392 39738
rect 5416 39686 5426 39738
rect 5426 39686 5472 39738
rect 5176 39684 5232 39686
rect 5256 39684 5312 39686
rect 5336 39684 5392 39686
rect 5416 39684 5472 39686
rect 3514 38800 3570 38856
rect 2778 36760 2834 36816
rect 2870 36080 2926 36136
rect 2778 35400 2834 35456
rect 2778 34040 2834 34096
rect 2226 19080 2282 19136
rect 2778 31320 2834 31376
rect 2778 25200 2834 25256
rect 3514 32000 3570 32056
rect 2778 18400 2834 18456
rect 2778 17076 2780 17096
rect 2780 17076 2832 17096
rect 2832 17076 2834 17096
rect 2778 17040 2834 17076
rect 2778 15680 2834 15736
rect 2778 14320 2834 14376
rect 2778 13640 2834 13696
rect 2778 11636 2780 11656
rect 2780 11636 2832 11656
rect 2832 11636 2834 11656
rect 2778 11600 2834 11636
rect 2778 10920 2834 10976
rect 2778 8880 2834 8936
rect 2778 8200 2834 8256
rect 2778 7520 2834 7576
rect 2778 4800 2834 4856
rect 2778 4120 2834 4176
rect 2870 3440 2926 3496
rect 3422 5480 3478 5536
rect 2778 2080 2834 2136
rect 3974 2760 4030 2816
rect 5176 38650 5232 38652
rect 5256 38650 5312 38652
rect 5336 38650 5392 38652
rect 5416 38650 5472 38652
rect 5176 38598 5222 38650
rect 5222 38598 5232 38650
rect 5256 38598 5286 38650
rect 5286 38598 5298 38650
rect 5298 38598 5312 38650
rect 5336 38598 5350 38650
rect 5350 38598 5362 38650
rect 5362 38598 5392 38650
rect 5416 38598 5426 38650
rect 5426 38598 5472 38650
rect 5176 38596 5232 38598
rect 5256 38596 5312 38598
rect 5336 38596 5392 38598
rect 5416 38596 5472 38598
rect 5176 37562 5232 37564
rect 5256 37562 5312 37564
rect 5336 37562 5392 37564
rect 5416 37562 5472 37564
rect 5176 37510 5222 37562
rect 5222 37510 5232 37562
rect 5256 37510 5286 37562
rect 5286 37510 5298 37562
rect 5298 37510 5312 37562
rect 5336 37510 5350 37562
rect 5350 37510 5362 37562
rect 5362 37510 5392 37562
rect 5416 37510 5426 37562
rect 5426 37510 5472 37562
rect 5176 37508 5232 37510
rect 5256 37508 5312 37510
rect 5336 37508 5392 37510
rect 5416 37508 5472 37510
rect 13617 39738 13673 39740
rect 13697 39738 13753 39740
rect 13777 39738 13833 39740
rect 13857 39738 13913 39740
rect 13617 39686 13663 39738
rect 13663 39686 13673 39738
rect 13697 39686 13727 39738
rect 13727 39686 13739 39738
rect 13739 39686 13753 39738
rect 13777 39686 13791 39738
rect 13791 39686 13803 39738
rect 13803 39686 13833 39738
rect 13857 39686 13867 39738
rect 13867 39686 13913 39738
rect 13617 39684 13673 39686
rect 13697 39684 13753 39686
rect 13777 39684 13833 39686
rect 13857 39684 13913 39686
rect 13726 39380 13728 39400
rect 13728 39380 13780 39400
rect 13780 39380 13782 39400
rect 5176 36474 5232 36476
rect 5256 36474 5312 36476
rect 5336 36474 5392 36476
rect 5416 36474 5472 36476
rect 5176 36422 5222 36474
rect 5222 36422 5232 36474
rect 5256 36422 5286 36474
rect 5286 36422 5298 36474
rect 5298 36422 5312 36474
rect 5336 36422 5350 36474
rect 5350 36422 5362 36474
rect 5362 36422 5392 36474
rect 5416 36422 5426 36474
rect 5426 36422 5472 36474
rect 5176 36420 5232 36422
rect 5256 36420 5312 36422
rect 5336 36420 5392 36422
rect 5416 36420 5472 36422
rect 4066 1400 4122 1456
rect 5176 35386 5232 35388
rect 5256 35386 5312 35388
rect 5336 35386 5392 35388
rect 5416 35386 5472 35388
rect 5176 35334 5222 35386
rect 5222 35334 5232 35386
rect 5256 35334 5286 35386
rect 5286 35334 5298 35386
rect 5298 35334 5312 35386
rect 5336 35334 5350 35386
rect 5350 35334 5362 35386
rect 5362 35334 5392 35386
rect 5416 35334 5426 35386
rect 5426 35334 5472 35386
rect 5176 35332 5232 35334
rect 5256 35332 5312 35334
rect 5336 35332 5392 35334
rect 5416 35332 5472 35334
rect 5176 34298 5232 34300
rect 5256 34298 5312 34300
rect 5336 34298 5392 34300
rect 5416 34298 5472 34300
rect 5176 34246 5222 34298
rect 5222 34246 5232 34298
rect 5256 34246 5286 34298
rect 5286 34246 5298 34298
rect 5298 34246 5312 34298
rect 5336 34246 5350 34298
rect 5350 34246 5362 34298
rect 5362 34246 5392 34298
rect 5416 34246 5426 34298
rect 5426 34246 5472 34298
rect 5176 34244 5232 34246
rect 5256 34244 5312 34246
rect 5336 34244 5392 34246
rect 5416 34244 5472 34246
rect 5176 33210 5232 33212
rect 5256 33210 5312 33212
rect 5336 33210 5392 33212
rect 5416 33210 5472 33212
rect 5176 33158 5222 33210
rect 5222 33158 5232 33210
rect 5256 33158 5286 33210
rect 5286 33158 5298 33210
rect 5298 33158 5312 33210
rect 5336 33158 5350 33210
rect 5350 33158 5362 33210
rect 5362 33158 5392 33210
rect 5416 33158 5426 33210
rect 5426 33158 5472 33210
rect 5176 33156 5232 33158
rect 5256 33156 5312 33158
rect 5336 33156 5392 33158
rect 5416 33156 5472 33158
rect 5176 32122 5232 32124
rect 5256 32122 5312 32124
rect 5336 32122 5392 32124
rect 5416 32122 5472 32124
rect 5176 32070 5222 32122
rect 5222 32070 5232 32122
rect 5256 32070 5286 32122
rect 5286 32070 5298 32122
rect 5298 32070 5312 32122
rect 5336 32070 5350 32122
rect 5350 32070 5362 32122
rect 5362 32070 5392 32122
rect 5416 32070 5426 32122
rect 5426 32070 5472 32122
rect 5176 32068 5232 32070
rect 5256 32068 5312 32070
rect 5336 32068 5392 32070
rect 5416 32068 5472 32070
rect 5176 31034 5232 31036
rect 5256 31034 5312 31036
rect 5336 31034 5392 31036
rect 5416 31034 5472 31036
rect 5176 30982 5222 31034
rect 5222 30982 5232 31034
rect 5256 30982 5286 31034
rect 5286 30982 5298 31034
rect 5298 30982 5312 31034
rect 5336 30982 5350 31034
rect 5350 30982 5362 31034
rect 5362 30982 5392 31034
rect 5416 30982 5426 31034
rect 5426 30982 5472 31034
rect 5176 30980 5232 30982
rect 5256 30980 5312 30982
rect 5336 30980 5392 30982
rect 5416 30980 5472 30982
rect 5176 29946 5232 29948
rect 5256 29946 5312 29948
rect 5336 29946 5392 29948
rect 5416 29946 5472 29948
rect 5176 29894 5222 29946
rect 5222 29894 5232 29946
rect 5256 29894 5286 29946
rect 5286 29894 5298 29946
rect 5298 29894 5312 29946
rect 5336 29894 5350 29946
rect 5350 29894 5362 29946
rect 5362 29894 5392 29946
rect 5416 29894 5426 29946
rect 5426 29894 5472 29946
rect 5176 29892 5232 29894
rect 5256 29892 5312 29894
rect 5336 29892 5392 29894
rect 5416 29892 5472 29894
rect 5176 28858 5232 28860
rect 5256 28858 5312 28860
rect 5336 28858 5392 28860
rect 5416 28858 5472 28860
rect 5176 28806 5222 28858
rect 5222 28806 5232 28858
rect 5256 28806 5286 28858
rect 5286 28806 5298 28858
rect 5298 28806 5312 28858
rect 5336 28806 5350 28858
rect 5350 28806 5362 28858
rect 5362 28806 5392 28858
rect 5416 28806 5426 28858
rect 5426 28806 5472 28858
rect 5176 28804 5232 28806
rect 5256 28804 5312 28806
rect 5336 28804 5392 28806
rect 5416 28804 5472 28806
rect 5176 27770 5232 27772
rect 5256 27770 5312 27772
rect 5336 27770 5392 27772
rect 5416 27770 5472 27772
rect 5176 27718 5222 27770
rect 5222 27718 5232 27770
rect 5256 27718 5286 27770
rect 5286 27718 5298 27770
rect 5298 27718 5312 27770
rect 5336 27718 5350 27770
rect 5350 27718 5362 27770
rect 5362 27718 5392 27770
rect 5416 27718 5426 27770
rect 5426 27718 5472 27770
rect 5176 27716 5232 27718
rect 5256 27716 5312 27718
rect 5336 27716 5392 27718
rect 5416 27716 5472 27718
rect 5176 26682 5232 26684
rect 5256 26682 5312 26684
rect 5336 26682 5392 26684
rect 5416 26682 5472 26684
rect 5176 26630 5222 26682
rect 5222 26630 5232 26682
rect 5256 26630 5286 26682
rect 5286 26630 5298 26682
rect 5298 26630 5312 26682
rect 5336 26630 5350 26682
rect 5350 26630 5362 26682
rect 5362 26630 5392 26682
rect 5416 26630 5426 26682
rect 5426 26630 5472 26682
rect 5176 26628 5232 26630
rect 5256 26628 5312 26630
rect 5336 26628 5392 26630
rect 5416 26628 5472 26630
rect 5176 25594 5232 25596
rect 5256 25594 5312 25596
rect 5336 25594 5392 25596
rect 5416 25594 5472 25596
rect 5176 25542 5222 25594
rect 5222 25542 5232 25594
rect 5256 25542 5286 25594
rect 5286 25542 5298 25594
rect 5298 25542 5312 25594
rect 5336 25542 5350 25594
rect 5350 25542 5362 25594
rect 5362 25542 5392 25594
rect 5416 25542 5426 25594
rect 5426 25542 5472 25594
rect 5176 25540 5232 25542
rect 5256 25540 5312 25542
rect 5336 25540 5392 25542
rect 5416 25540 5472 25542
rect 5176 24506 5232 24508
rect 5256 24506 5312 24508
rect 5336 24506 5392 24508
rect 5416 24506 5472 24508
rect 5176 24454 5222 24506
rect 5222 24454 5232 24506
rect 5256 24454 5286 24506
rect 5286 24454 5298 24506
rect 5298 24454 5312 24506
rect 5336 24454 5350 24506
rect 5350 24454 5362 24506
rect 5362 24454 5392 24506
rect 5416 24454 5426 24506
rect 5426 24454 5472 24506
rect 5176 24452 5232 24454
rect 5256 24452 5312 24454
rect 5336 24452 5392 24454
rect 5416 24452 5472 24454
rect 5176 23418 5232 23420
rect 5256 23418 5312 23420
rect 5336 23418 5392 23420
rect 5416 23418 5472 23420
rect 5176 23366 5222 23418
rect 5222 23366 5232 23418
rect 5256 23366 5286 23418
rect 5286 23366 5298 23418
rect 5298 23366 5312 23418
rect 5336 23366 5350 23418
rect 5350 23366 5362 23418
rect 5362 23366 5392 23418
rect 5416 23366 5426 23418
rect 5426 23366 5472 23418
rect 5176 23364 5232 23366
rect 5256 23364 5312 23366
rect 5336 23364 5392 23366
rect 5416 23364 5472 23366
rect 5176 22330 5232 22332
rect 5256 22330 5312 22332
rect 5336 22330 5392 22332
rect 5416 22330 5472 22332
rect 5176 22278 5222 22330
rect 5222 22278 5232 22330
rect 5256 22278 5286 22330
rect 5286 22278 5298 22330
rect 5298 22278 5312 22330
rect 5336 22278 5350 22330
rect 5350 22278 5362 22330
rect 5362 22278 5392 22330
rect 5416 22278 5426 22330
rect 5426 22278 5472 22330
rect 5176 22276 5232 22278
rect 5256 22276 5312 22278
rect 5336 22276 5392 22278
rect 5416 22276 5472 22278
rect 5176 21242 5232 21244
rect 5256 21242 5312 21244
rect 5336 21242 5392 21244
rect 5416 21242 5472 21244
rect 5176 21190 5222 21242
rect 5222 21190 5232 21242
rect 5256 21190 5286 21242
rect 5286 21190 5298 21242
rect 5298 21190 5312 21242
rect 5336 21190 5350 21242
rect 5350 21190 5362 21242
rect 5362 21190 5392 21242
rect 5416 21190 5426 21242
rect 5426 21190 5472 21242
rect 5176 21188 5232 21190
rect 5256 21188 5312 21190
rect 5336 21188 5392 21190
rect 5416 21188 5472 21190
rect 5176 20154 5232 20156
rect 5256 20154 5312 20156
rect 5336 20154 5392 20156
rect 5416 20154 5472 20156
rect 5176 20102 5222 20154
rect 5222 20102 5232 20154
rect 5256 20102 5286 20154
rect 5286 20102 5298 20154
rect 5298 20102 5312 20154
rect 5336 20102 5350 20154
rect 5350 20102 5362 20154
rect 5362 20102 5392 20154
rect 5416 20102 5426 20154
rect 5426 20102 5472 20154
rect 5176 20100 5232 20102
rect 5256 20100 5312 20102
rect 5336 20100 5392 20102
rect 5416 20100 5472 20102
rect 5176 19066 5232 19068
rect 5256 19066 5312 19068
rect 5336 19066 5392 19068
rect 5416 19066 5472 19068
rect 5176 19014 5222 19066
rect 5222 19014 5232 19066
rect 5256 19014 5286 19066
rect 5286 19014 5298 19066
rect 5298 19014 5312 19066
rect 5336 19014 5350 19066
rect 5350 19014 5362 19066
rect 5362 19014 5392 19066
rect 5416 19014 5426 19066
rect 5426 19014 5472 19066
rect 5176 19012 5232 19014
rect 5256 19012 5312 19014
rect 5336 19012 5392 19014
rect 5416 19012 5472 19014
rect 5176 17978 5232 17980
rect 5256 17978 5312 17980
rect 5336 17978 5392 17980
rect 5416 17978 5472 17980
rect 5176 17926 5222 17978
rect 5222 17926 5232 17978
rect 5256 17926 5286 17978
rect 5286 17926 5298 17978
rect 5298 17926 5312 17978
rect 5336 17926 5350 17978
rect 5350 17926 5362 17978
rect 5362 17926 5392 17978
rect 5416 17926 5426 17978
rect 5426 17926 5472 17978
rect 5176 17924 5232 17926
rect 5256 17924 5312 17926
rect 5336 17924 5392 17926
rect 5416 17924 5472 17926
rect 5176 16890 5232 16892
rect 5256 16890 5312 16892
rect 5336 16890 5392 16892
rect 5416 16890 5472 16892
rect 5176 16838 5222 16890
rect 5222 16838 5232 16890
rect 5256 16838 5286 16890
rect 5286 16838 5298 16890
rect 5298 16838 5312 16890
rect 5336 16838 5350 16890
rect 5350 16838 5362 16890
rect 5362 16838 5392 16890
rect 5416 16838 5426 16890
rect 5426 16838 5472 16890
rect 5176 16836 5232 16838
rect 5256 16836 5312 16838
rect 5336 16836 5392 16838
rect 5416 16836 5472 16838
rect 5176 15802 5232 15804
rect 5256 15802 5312 15804
rect 5336 15802 5392 15804
rect 5416 15802 5472 15804
rect 5176 15750 5222 15802
rect 5222 15750 5232 15802
rect 5256 15750 5286 15802
rect 5286 15750 5298 15802
rect 5298 15750 5312 15802
rect 5336 15750 5350 15802
rect 5350 15750 5362 15802
rect 5362 15750 5392 15802
rect 5416 15750 5426 15802
rect 5426 15750 5472 15802
rect 5176 15748 5232 15750
rect 5256 15748 5312 15750
rect 5336 15748 5392 15750
rect 5416 15748 5472 15750
rect 5176 14714 5232 14716
rect 5256 14714 5312 14716
rect 5336 14714 5392 14716
rect 5416 14714 5472 14716
rect 5176 14662 5222 14714
rect 5222 14662 5232 14714
rect 5256 14662 5286 14714
rect 5286 14662 5298 14714
rect 5298 14662 5312 14714
rect 5336 14662 5350 14714
rect 5350 14662 5362 14714
rect 5362 14662 5392 14714
rect 5416 14662 5426 14714
rect 5426 14662 5472 14714
rect 5176 14660 5232 14662
rect 5256 14660 5312 14662
rect 5336 14660 5392 14662
rect 5416 14660 5472 14662
rect 5176 13626 5232 13628
rect 5256 13626 5312 13628
rect 5336 13626 5392 13628
rect 5416 13626 5472 13628
rect 5176 13574 5222 13626
rect 5222 13574 5232 13626
rect 5256 13574 5286 13626
rect 5286 13574 5298 13626
rect 5298 13574 5312 13626
rect 5336 13574 5350 13626
rect 5350 13574 5362 13626
rect 5362 13574 5392 13626
rect 5416 13574 5426 13626
rect 5426 13574 5472 13626
rect 5176 13572 5232 13574
rect 5256 13572 5312 13574
rect 5336 13572 5392 13574
rect 5416 13572 5472 13574
rect 5176 12538 5232 12540
rect 5256 12538 5312 12540
rect 5336 12538 5392 12540
rect 5416 12538 5472 12540
rect 5176 12486 5222 12538
rect 5222 12486 5232 12538
rect 5256 12486 5286 12538
rect 5286 12486 5298 12538
rect 5298 12486 5312 12538
rect 5336 12486 5350 12538
rect 5350 12486 5362 12538
rect 5362 12486 5392 12538
rect 5416 12486 5426 12538
rect 5426 12486 5472 12538
rect 5176 12484 5232 12486
rect 5256 12484 5312 12486
rect 5336 12484 5392 12486
rect 5416 12484 5472 12486
rect 5176 11450 5232 11452
rect 5256 11450 5312 11452
rect 5336 11450 5392 11452
rect 5416 11450 5472 11452
rect 5176 11398 5222 11450
rect 5222 11398 5232 11450
rect 5256 11398 5286 11450
rect 5286 11398 5298 11450
rect 5298 11398 5312 11450
rect 5336 11398 5350 11450
rect 5350 11398 5362 11450
rect 5362 11398 5392 11450
rect 5416 11398 5426 11450
rect 5426 11398 5472 11450
rect 5176 11396 5232 11398
rect 5256 11396 5312 11398
rect 5336 11396 5392 11398
rect 5416 11396 5472 11398
rect 5176 10362 5232 10364
rect 5256 10362 5312 10364
rect 5336 10362 5392 10364
rect 5416 10362 5472 10364
rect 5176 10310 5222 10362
rect 5222 10310 5232 10362
rect 5256 10310 5286 10362
rect 5286 10310 5298 10362
rect 5298 10310 5312 10362
rect 5336 10310 5350 10362
rect 5350 10310 5362 10362
rect 5362 10310 5392 10362
rect 5416 10310 5426 10362
rect 5426 10310 5472 10362
rect 5176 10308 5232 10310
rect 5256 10308 5312 10310
rect 5336 10308 5392 10310
rect 5416 10308 5472 10310
rect 5176 9274 5232 9276
rect 5256 9274 5312 9276
rect 5336 9274 5392 9276
rect 5416 9274 5472 9276
rect 5176 9222 5222 9274
rect 5222 9222 5232 9274
rect 5256 9222 5286 9274
rect 5286 9222 5298 9274
rect 5298 9222 5312 9274
rect 5336 9222 5350 9274
rect 5350 9222 5362 9274
rect 5362 9222 5392 9274
rect 5416 9222 5426 9274
rect 5426 9222 5472 9274
rect 5176 9220 5232 9222
rect 5256 9220 5312 9222
rect 5336 9220 5392 9222
rect 5416 9220 5472 9222
rect 5176 8186 5232 8188
rect 5256 8186 5312 8188
rect 5336 8186 5392 8188
rect 5416 8186 5472 8188
rect 5176 8134 5222 8186
rect 5222 8134 5232 8186
rect 5256 8134 5286 8186
rect 5286 8134 5298 8186
rect 5298 8134 5312 8186
rect 5336 8134 5350 8186
rect 5350 8134 5362 8186
rect 5362 8134 5392 8186
rect 5416 8134 5426 8186
rect 5426 8134 5472 8186
rect 5176 8132 5232 8134
rect 5256 8132 5312 8134
rect 5336 8132 5392 8134
rect 5416 8132 5472 8134
rect 13726 39344 13782 39380
rect 9396 39194 9452 39196
rect 9476 39194 9532 39196
rect 9556 39194 9612 39196
rect 9636 39194 9692 39196
rect 9396 39142 9442 39194
rect 9442 39142 9452 39194
rect 9476 39142 9506 39194
rect 9506 39142 9518 39194
rect 9518 39142 9532 39194
rect 9556 39142 9570 39194
rect 9570 39142 9582 39194
rect 9582 39142 9612 39194
rect 9636 39142 9646 39194
rect 9646 39142 9692 39194
rect 9396 39140 9452 39142
rect 9476 39140 9532 39142
rect 9556 39140 9612 39142
rect 9636 39140 9692 39142
rect 9396 38106 9452 38108
rect 9476 38106 9532 38108
rect 9556 38106 9612 38108
rect 9636 38106 9692 38108
rect 9396 38054 9442 38106
rect 9442 38054 9452 38106
rect 9476 38054 9506 38106
rect 9506 38054 9518 38106
rect 9518 38054 9532 38106
rect 9556 38054 9570 38106
rect 9570 38054 9582 38106
rect 9582 38054 9612 38106
rect 9636 38054 9646 38106
rect 9646 38054 9692 38106
rect 9396 38052 9452 38054
rect 9476 38052 9532 38054
rect 9556 38052 9612 38054
rect 9636 38052 9692 38054
rect 9396 37018 9452 37020
rect 9476 37018 9532 37020
rect 9556 37018 9612 37020
rect 9636 37018 9692 37020
rect 9396 36966 9442 37018
rect 9442 36966 9452 37018
rect 9476 36966 9506 37018
rect 9506 36966 9518 37018
rect 9518 36966 9532 37018
rect 9556 36966 9570 37018
rect 9570 36966 9582 37018
rect 9582 36966 9612 37018
rect 9636 36966 9646 37018
rect 9646 36966 9692 37018
rect 9396 36964 9452 36966
rect 9476 36964 9532 36966
rect 9556 36964 9612 36966
rect 9636 36964 9692 36966
rect 9396 35930 9452 35932
rect 9476 35930 9532 35932
rect 9556 35930 9612 35932
rect 9636 35930 9692 35932
rect 9396 35878 9442 35930
rect 9442 35878 9452 35930
rect 9476 35878 9506 35930
rect 9506 35878 9518 35930
rect 9518 35878 9532 35930
rect 9556 35878 9570 35930
rect 9570 35878 9582 35930
rect 9582 35878 9612 35930
rect 9636 35878 9646 35930
rect 9646 35878 9692 35930
rect 9396 35876 9452 35878
rect 9476 35876 9532 35878
rect 9556 35876 9612 35878
rect 9636 35876 9692 35878
rect 9396 34842 9452 34844
rect 9476 34842 9532 34844
rect 9556 34842 9612 34844
rect 9636 34842 9692 34844
rect 9396 34790 9442 34842
rect 9442 34790 9452 34842
rect 9476 34790 9506 34842
rect 9506 34790 9518 34842
rect 9518 34790 9532 34842
rect 9556 34790 9570 34842
rect 9570 34790 9582 34842
rect 9582 34790 9612 34842
rect 9636 34790 9646 34842
rect 9646 34790 9692 34842
rect 9396 34788 9452 34790
rect 9476 34788 9532 34790
rect 9556 34788 9612 34790
rect 9636 34788 9692 34790
rect 9396 33754 9452 33756
rect 9476 33754 9532 33756
rect 9556 33754 9612 33756
rect 9636 33754 9692 33756
rect 9396 33702 9442 33754
rect 9442 33702 9452 33754
rect 9476 33702 9506 33754
rect 9506 33702 9518 33754
rect 9518 33702 9532 33754
rect 9556 33702 9570 33754
rect 9570 33702 9582 33754
rect 9582 33702 9612 33754
rect 9636 33702 9646 33754
rect 9646 33702 9692 33754
rect 9396 33700 9452 33702
rect 9476 33700 9532 33702
rect 9556 33700 9612 33702
rect 9636 33700 9692 33702
rect 13617 38650 13673 38652
rect 13697 38650 13753 38652
rect 13777 38650 13833 38652
rect 13857 38650 13913 38652
rect 13617 38598 13663 38650
rect 13663 38598 13673 38650
rect 13697 38598 13727 38650
rect 13727 38598 13739 38650
rect 13739 38598 13753 38650
rect 13777 38598 13791 38650
rect 13791 38598 13803 38650
rect 13803 38598 13833 38650
rect 13857 38598 13867 38650
rect 13867 38598 13913 38650
rect 13617 38596 13673 38598
rect 13697 38596 13753 38598
rect 13777 38596 13833 38598
rect 13857 38596 13913 38598
rect 13617 37562 13673 37564
rect 13697 37562 13753 37564
rect 13777 37562 13833 37564
rect 13857 37562 13913 37564
rect 13617 37510 13663 37562
rect 13663 37510 13673 37562
rect 13697 37510 13727 37562
rect 13727 37510 13739 37562
rect 13739 37510 13753 37562
rect 13777 37510 13791 37562
rect 13791 37510 13803 37562
rect 13803 37510 13833 37562
rect 13857 37510 13867 37562
rect 13867 37510 13913 37562
rect 13617 37508 13673 37510
rect 13697 37508 13753 37510
rect 13777 37508 13833 37510
rect 13857 37508 13913 37510
rect 13617 36474 13673 36476
rect 13697 36474 13753 36476
rect 13777 36474 13833 36476
rect 13857 36474 13913 36476
rect 13617 36422 13663 36474
rect 13663 36422 13673 36474
rect 13697 36422 13727 36474
rect 13727 36422 13739 36474
rect 13739 36422 13753 36474
rect 13777 36422 13791 36474
rect 13791 36422 13803 36474
rect 13803 36422 13833 36474
rect 13857 36422 13867 36474
rect 13867 36422 13913 36474
rect 13617 36420 13673 36422
rect 13697 36420 13753 36422
rect 13777 36420 13833 36422
rect 13857 36420 13913 36422
rect 13617 35386 13673 35388
rect 13697 35386 13753 35388
rect 13777 35386 13833 35388
rect 13857 35386 13913 35388
rect 13617 35334 13663 35386
rect 13663 35334 13673 35386
rect 13697 35334 13727 35386
rect 13727 35334 13739 35386
rect 13739 35334 13753 35386
rect 13777 35334 13791 35386
rect 13791 35334 13803 35386
rect 13803 35334 13833 35386
rect 13857 35334 13867 35386
rect 13867 35334 13913 35386
rect 13617 35332 13673 35334
rect 13697 35332 13753 35334
rect 13777 35332 13833 35334
rect 13857 35332 13913 35334
rect 13617 34298 13673 34300
rect 13697 34298 13753 34300
rect 13777 34298 13833 34300
rect 13857 34298 13913 34300
rect 13617 34246 13663 34298
rect 13663 34246 13673 34298
rect 13697 34246 13727 34298
rect 13727 34246 13739 34298
rect 13739 34246 13753 34298
rect 13777 34246 13791 34298
rect 13791 34246 13803 34298
rect 13803 34246 13833 34298
rect 13857 34246 13867 34298
rect 13867 34246 13913 34298
rect 13617 34244 13673 34246
rect 13697 34244 13753 34246
rect 13777 34244 13833 34246
rect 13857 34244 13913 34246
rect 13617 33210 13673 33212
rect 13697 33210 13753 33212
rect 13777 33210 13833 33212
rect 13857 33210 13913 33212
rect 13617 33158 13663 33210
rect 13663 33158 13673 33210
rect 13697 33158 13727 33210
rect 13727 33158 13739 33210
rect 13739 33158 13753 33210
rect 13777 33158 13791 33210
rect 13791 33158 13803 33210
rect 13803 33158 13833 33210
rect 13857 33158 13867 33210
rect 13867 33158 13913 33210
rect 13617 33156 13673 33158
rect 13697 33156 13753 33158
rect 13777 33156 13833 33158
rect 13857 33156 13913 33158
rect 9396 32666 9452 32668
rect 9476 32666 9532 32668
rect 9556 32666 9612 32668
rect 9636 32666 9692 32668
rect 9396 32614 9442 32666
rect 9442 32614 9452 32666
rect 9476 32614 9506 32666
rect 9506 32614 9518 32666
rect 9518 32614 9532 32666
rect 9556 32614 9570 32666
rect 9570 32614 9582 32666
rect 9582 32614 9612 32666
rect 9636 32614 9646 32666
rect 9646 32614 9692 32666
rect 9396 32612 9452 32614
rect 9476 32612 9532 32614
rect 9556 32612 9612 32614
rect 9636 32612 9692 32614
rect 13617 32122 13673 32124
rect 13697 32122 13753 32124
rect 13777 32122 13833 32124
rect 13857 32122 13913 32124
rect 13617 32070 13663 32122
rect 13663 32070 13673 32122
rect 13697 32070 13727 32122
rect 13727 32070 13739 32122
rect 13739 32070 13753 32122
rect 13777 32070 13791 32122
rect 13791 32070 13803 32122
rect 13803 32070 13833 32122
rect 13857 32070 13867 32122
rect 13867 32070 13913 32122
rect 13617 32068 13673 32070
rect 13697 32068 13753 32070
rect 13777 32068 13833 32070
rect 13857 32068 13913 32070
rect 9396 31578 9452 31580
rect 9476 31578 9532 31580
rect 9556 31578 9612 31580
rect 9636 31578 9692 31580
rect 9396 31526 9442 31578
rect 9442 31526 9452 31578
rect 9476 31526 9506 31578
rect 9506 31526 9518 31578
rect 9518 31526 9532 31578
rect 9556 31526 9570 31578
rect 9570 31526 9582 31578
rect 9582 31526 9612 31578
rect 9636 31526 9646 31578
rect 9646 31526 9692 31578
rect 9396 31524 9452 31526
rect 9476 31524 9532 31526
rect 9556 31524 9612 31526
rect 9636 31524 9692 31526
rect 13617 31034 13673 31036
rect 13697 31034 13753 31036
rect 13777 31034 13833 31036
rect 13857 31034 13913 31036
rect 13617 30982 13663 31034
rect 13663 30982 13673 31034
rect 13697 30982 13727 31034
rect 13727 30982 13739 31034
rect 13739 30982 13753 31034
rect 13777 30982 13791 31034
rect 13791 30982 13803 31034
rect 13803 30982 13833 31034
rect 13857 30982 13867 31034
rect 13867 30982 13913 31034
rect 13617 30980 13673 30982
rect 13697 30980 13753 30982
rect 13777 30980 13833 30982
rect 13857 30980 13913 30982
rect 9396 30490 9452 30492
rect 9476 30490 9532 30492
rect 9556 30490 9612 30492
rect 9636 30490 9692 30492
rect 9396 30438 9442 30490
rect 9442 30438 9452 30490
rect 9476 30438 9506 30490
rect 9506 30438 9518 30490
rect 9518 30438 9532 30490
rect 9556 30438 9570 30490
rect 9570 30438 9582 30490
rect 9582 30438 9612 30490
rect 9636 30438 9646 30490
rect 9646 30438 9692 30490
rect 9396 30436 9452 30438
rect 9476 30436 9532 30438
rect 9556 30436 9612 30438
rect 9636 30436 9692 30438
rect 13617 29946 13673 29948
rect 13697 29946 13753 29948
rect 13777 29946 13833 29948
rect 13857 29946 13913 29948
rect 13617 29894 13663 29946
rect 13663 29894 13673 29946
rect 13697 29894 13727 29946
rect 13727 29894 13739 29946
rect 13739 29894 13753 29946
rect 13777 29894 13791 29946
rect 13791 29894 13803 29946
rect 13803 29894 13833 29946
rect 13857 29894 13867 29946
rect 13867 29894 13913 29946
rect 13617 29892 13673 29894
rect 13697 29892 13753 29894
rect 13777 29892 13833 29894
rect 13857 29892 13913 29894
rect 9396 29402 9452 29404
rect 9476 29402 9532 29404
rect 9556 29402 9612 29404
rect 9636 29402 9692 29404
rect 9396 29350 9442 29402
rect 9442 29350 9452 29402
rect 9476 29350 9506 29402
rect 9506 29350 9518 29402
rect 9518 29350 9532 29402
rect 9556 29350 9570 29402
rect 9570 29350 9582 29402
rect 9582 29350 9612 29402
rect 9636 29350 9646 29402
rect 9646 29350 9692 29402
rect 9396 29348 9452 29350
rect 9476 29348 9532 29350
rect 9556 29348 9612 29350
rect 9636 29348 9692 29350
rect 13617 28858 13673 28860
rect 13697 28858 13753 28860
rect 13777 28858 13833 28860
rect 13857 28858 13913 28860
rect 13617 28806 13663 28858
rect 13663 28806 13673 28858
rect 13697 28806 13727 28858
rect 13727 28806 13739 28858
rect 13739 28806 13753 28858
rect 13777 28806 13791 28858
rect 13791 28806 13803 28858
rect 13803 28806 13833 28858
rect 13857 28806 13867 28858
rect 13867 28806 13913 28858
rect 13617 28804 13673 28806
rect 13697 28804 13753 28806
rect 13777 28804 13833 28806
rect 13857 28804 13913 28806
rect 9396 28314 9452 28316
rect 9476 28314 9532 28316
rect 9556 28314 9612 28316
rect 9636 28314 9692 28316
rect 9396 28262 9442 28314
rect 9442 28262 9452 28314
rect 9476 28262 9506 28314
rect 9506 28262 9518 28314
rect 9518 28262 9532 28314
rect 9556 28262 9570 28314
rect 9570 28262 9582 28314
rect 9582 28262 9612 28314
rect 9636 28262 9646 28314
rect 9646 28262 9692 28314
rect 9396 28260 9452 28262
rect 9476 28260 9532 28262
rect 9556 28260 9612 28262
rect 9636 28260 9692 28262
rect 13617 27770 13673 27772
rect 13697 27770 13753 27772
rect 13777 27770 13833 27772
rect 13857 27770 13913 27772
rect 13617 27718 13663 27770
rect 13663 27718 13673 27770
rect 13697 27718 13727 27770
rect 13727 27718 13739 27770
rect 13739 27718 13753 27770
rect 13777 27718 13791 27770
rect 13791 27718 13803 27770
rect 13803 27718 13833 27770
rect 13857 27718 13867 27770
rect 13867 27718 13913 27770
rect 13617 27716 13673 27718
rect 13697 27716 13753 27718
rect 13777 27716 13833 27718
rect 13857 27716 13913 27718
rect 9396 27226 9452 27228
rect 9476 27226 9532 27228
rect 9556 27226 9612 27228
rect 9636 27226 9692 27228
rect 9396 27174 9442 27226
rect 9442 27174 9452 27226
rect 9476 27174 9506 27226
rect 9506 27174 9518 27226
rect 9518 27174 9532 27226
rect 9556 27174 9570 27226
rect 9570 27174 9582 27226
rect 9582 27174 9612 27226
rect 9636 27174 9646 27226
rect 9646 27174 9692 27226
rect 9396 27172 9452 27174
rect 9476 27172 9532 27174
rect 9556 27172 9612 27174
rect 9636 27172 9692 27174
rect 13617 26682 13673 26684
rect 13697 26682 13753 26684
rect 13777 26682 13833 26684
rect 13857 26682 13913 26684
rect 13617 26630 13663 26682
rect 13663 26630 13673 26682
rect 13697 26630 13727 26682
rect 13727 26630 13739 26682
rect 13739 26630 13753 26682
rect 13777 26630 13791 26682
rect 13791 26630 13803 26682
rect 13803 26630 13833 26682
rect 13857 26630 13867 26682
rect 13867 26630 13913 26682
rect 13617 26628 13673 26630
rect 13697 26628 13753 26630
rect 13777 26628 13833 26630
rect 13857 26628 13913 26630
rect 9396 26138 9452 26140
rect 9476 26138 9532 26140
rect 9556 26138 9612 26140
rect 9636 26138 9692 26140
rect 9396 26086 9442 26138
rect 9442 26086 9452 26138
rect 9476 26086 9506 26138
rect 9506 26086 9518 26138
rect 9518 26086 9532 26138
rect 9556 26086 9570 26138
rect 9570 26086 9582 26138
rect 9582 26086 9612 26138
rect 9636 26086 9646 26138
rect 9646 26086 9692 26138
rect 9396 26084 9452 26086
rect 9476 26084 9532 26086
rect 9556 26084 9612 26086
rect 9636 26084 9692 26086
rect 13617 25594 13673 25596
rect 13697 25594 13753 25596
rect 13777 25594 13833 25596
rect 13857 25594 13913 25596
rect 13617 25542 13663 25594
rect 13663 25542 13673 25594
rect 13697 25542 13727 25594
rect 13727 25542 13739 25594
rect 13739 25542 13753 25594
rect 13777 25542 13791 25594
rect 13791 25542 13803 25594
rect 13803 25542 13833 25594
rect 13857 25542 13867 25594
rect 13867 25542 13913 25594
rect 13617 25540 13673 25542
rect 13697 25540 13753 25542
rect 13777 25540 13833 25542
rect 13857 25540 13913 25542
rect 16118 28464 16174 28520
rect 9396 25050 9452 25052
rect 9476 25050 9532 25052
rect 9556 25050 9612 25052
rect 9636 25050 9692 25052
rect 9396 24998 9442 25050
rect 9442 24998 9452 25050
rect 9476 24998 9506 25050
rect 9506 24998 9518 25050
rect 9518 24998 9532 25050
rect 9556 24998 9570 25050
rect 9570 24998 9582 25050
rect 9582 24998 9612 25050
rect 9636 24998 9646 25050
rect 9646 24998 9692 25050
rect 9396 24996 9452 24998
rect 9476 24996 9532 24998
rect 9556 24996 9612 24998
rect 9636 24996 9692 24998
rect 13617 24506 13673 24508
rect 13697 24506 13753 24508
rect 13777 24506 13833 24508
rect 13857 24506 13913 24508
rect 13617 24454 13663 24506
rect 13663 24454 13673 24506
rect 13697 24454 13727 24506
rect 13727 24454 13739 24506
rect 13739 24454 13753 24506
rect 13777 24454 13791 24506
rect 13791 24454 13803 24506
rect 13803 24454 13833 24506
rect 13857 24454 13867 24506
rect 13867 24454 13913 24506
rect 13617 24452 13673 24454
rect 13697 24452 13753 24454
rect 13777 24452 13833 24454
rect 13857 24452 13913 24454
rect 9396 23962 9452 23964
rect 9476 23962 9532 23964
rect 9556 23962 9612 23964
rect 9636 23962 9692 23964
rect 9396 23910 9442 23962
rect 9442 23910 9452 23962
rect 9476 23910 9506 23962
rect 9506 23910 9518 23962
rect 9518 23910 9532 23962
rect 9556 23910 9570 23962
rect 9570 23910 9582 23962
rect 9582 23910 9612 23962
rect 9636 23910 9646 23962
rect 9646 23910 9692 23962
rect 9396 23908 9452 23910
rect 9476 23908 9532 23910
rect 9556 23908 9612 23910
rect 9636 23908 9692 23910
rect 13617 23418 13673 23420
rect 13697 23418 13753 23420
rect 13777 23418 13833 23420
rect 13857 23418 13913 23420
rect 13617 23366 13663 23418
rect 13663 23366 13673 23418
rect 13697 23366 13727 23418
rect 13727 23366 13739 23418
rect 13739 23366 13753 23418
rect 13777 23366 13791 23418
rect 13791 23366 13803 23418
rect 13803 23366 13833 23418
rect 13857 23366 13867 23418
rect 13867 23366 13913 23418
rect 13617 23364 13673 23366
rect 13697 23364 13753 23366
rect 13777 23364 13833 23366
rect 13857 23364 13913 23366
rect 9396 22874 9452 22876
rect 9476 22874 9532 22876
rect 9556 22874 9612 22876
rect 9636 22874 9692 22876
rect 9396 22822 9442 22874
rect 9442 22822 9452 22874
rect 9476 22822 9506 22874
rect 9506 22822 9518 22874
rect 9518 22822 9532 22874
rect 9556 22822 9570 22874
rect 9570 22822 9582 22874
rect 9582 22822 9612 22874
rect 9636 22822 9646 22874
rect 9646 22822 9692 22874
rect 9396 22820 9452 22822
rect 9476 22820 9532 22822
rect 9556 22820 9612 22822
rect 9636 22820 9692 22822
rect 13617 22330 13673 22332
rect 13697 22330 13753 22332
rect 13777 22330 13833 22332
rect 13857 22330 13913 22332
rect 13617 22278 13663 22330
rect 13663 22278 13673 22330
rect 13697 22278 13727 22330
rect 13727 22278 13739 22330
rect 13739 22278 13753 22330
rect 13777 22278 13791 22330
rect 13791 22278 13803 22330
rect 13803 22278 13833 22330
rect 13857 22278 13867 22330
rect 13867 22278 13913 22330
rect 13617 22276 13673 22278
rect 13697 22276 13753 22278
rect 13777 22276 13833 22278
rect 13857 22276 13913 22278
rect 9396 21786 9452 21788
rect 9476 21786 9532 21788
rect 9556 21786 9612 21788
rect 9636 21786 9692 21788
rect 9396 21734 9442 21786
rect 9442 21734 9452 21786
rect 9476 21734 9506 21786
rect 9506 21734 9518 21786
rect 9518 21734 9532 21786
rect 9556 21734 9570 21786
rect 9570 21734 9582 21786
rect 9582 21734 9612 21786
rect 9636 21734 9646 21786
rect 9646 21734 9692 21786
rect 9396 21732 9452 21734
rect 9476 21732 9532 21734
rect 9556 21732 9612 21734
rect 9636 21732 9692 21734
rect 13617 21242 13673 21244
rect 13697 21242 13753 21244
rect 13777 21242 13833 21244
rect 13857 21242 13913 21244
rect 13617 21190 13663 21242
rect 13663 21190 13673 21242
rect 13697 21190 13727 21242
rect 13727 21190 13739 21242
rect 13739 21190 13753 21242
rect 13777 21190 13791 21242
rect 13791 21190 13803 21242
rect 13803 21190 13833 21242
rect 13857 21190 13867 21242
rect 13867 21190 13913 21242
rect 13617 21188 13673 21190
rect 13697 21188 13753 21190
rect 13777 21188 13833 21190
rect 13857 21188 13913 21190
rect 9396 20698 9452 20700
rect 9476 20698 9532 20700
rect 9556 20698 9612 20700
rect 9636 20698 9692 20700
rect 9396 20646 9442 20698
rect 9442 20646 9452 20698
rect 9476 20646 9506 20698
rect 9506 20646 9518 20698
rect 9518 20646 9532 20698
rect 9556 20646 9570 20698
rect 9570 20646 9582 20698
rect 9582 20646 9612 20698
rect 9636 20646 9646 20698
rect 9646 20646 9692 20698
rect 9396 20644 9452 20646
rect 9476 20644 9532 20646
rect 9556 20644 9612 20646
rect 9636 20644 9692 20646
rect 13617 20154 13673 20156
rect 13697 20154 13753 20156
rect 13777 20154 13833 20156
rect 13857 20154 13913 20156
rect 13617 20102 13663 20154
rect 13663 20102 13673 20154
rect 13697 20102 13727 20154
rect 13727 20102 13739 20154
rect 13739 20102 13753 20154
rect 13777 20102 13791 20154
rect 13791 20102 13803 20154
rect 13803 20102 13833 20154
rect 13857 20102 13867 20154
rect 13867 20102 13913 20154
rect 13617 20100 13673 20102
rect 13697 20100 13753 20102
rect 13777 20100 13833 20102
rect 13857 20100 13913 20102
rect 9396 19610 9452 19612
rect 9476 19610 9532 19612
rect 9556 19610 9612 19612
rect 9636 19610 9692 19612
rect 9396 19558 9442 19610
rect 9442 19558 9452 19610
rect 9476 19558 9506 19610
rect 9506 19558 9518 19610
rect 9518 19558 9532 19610
rect 9556 19558 9570 19610
rect 9570 19558 9582 19610
rect 9582 19558 9612 19610
rect 9636 19558 9646 19610
rect 9646 19558 9692 19610
rect 9396 19556 9452 19558
rect 9476 19556 9532 19558
rect 9556 19556 9612 19558
rect 9636 19556 9692 19558
rect 13617 19066 13673 19068
rect 13697 19066 13753 19068
rect 13777 19066 13833 19068
rect 13857 19066 13913 19068
rect 13617 19014 13663 19066
rect 13663 19014 13673 19066
rect 13697 19014 13727 19066
rect 13727 19014 13739 19066
rect 13739 19014 13753 19066
rect 13777 19014 13791 19066
rect 13791 19014 13803 19066
rect 13803 19014 13833 19066
rect 13857 19014 13867 19066
rect 13867 19014 13913 19066
rect 13617 19012 13673 19014
rect 13697 19012 13753 19014
rect 13777 19012 13833 19014
rect 13857 19012 13913 19014
rect 9396 18522 9452 18524
rect 9476 18522 9532 18524
rect 9556 18522 9612 18524
rect 9636 18522 9692 18524
rect 9396 18470 9442 18522
rect 9442 18470 9452 18522
rect 9476 18470 9506 18522
rect 9506 18470 9518 18522
rect 9518 18470 9532 18522
rect 9556 18470 9570 18522
rect 9570 18470 9582 18522
rect 9582 18470 9612 18522
rect 9636 18470 9646 18522
rect 9646 18470 9692 18522
rect 9396 18468 9452 18470
rect 9476 18468 9532 18470
rect 9556 18468 9612 18470
rect 9636 18468 9692 18470
rect 13617 17978 13673 17980
rect 13697 17978 13753 17980
rect 13777 17978 13833 17980
rect 13857 17978 13913 17980
rect 13617 17926 13663 17978
rect 13663 17926 13673 17978
rect 13697 17926 13727 17978
rect 13727 17926 13739 17978
rect 13739 17926 13753 17978
rect 13777 17926 13791 17978
rect 13791 17926 13803 17978
rect 13803 17926 13833 17978
rect 13857 17926 13867 17978
rect 13867 17926 13913 17978
rect 13617 17924 13673 17926
rect 13697 17924 13753 17926
rect 13777 17924 13833 17926
rect 13857 17924 13913 17926
rect 9396 17434 9452 17436
rect 9476 17434 9532 17436
rect 9556 17434 9612 17436
rect 9636 17434 9692 17436
rect 9396 17382 9442 17434
rect 9442 17382 9452 17434
rect 9476 17382 9506 17434
rect 9506 17382 9518 17434
rect 9518 17382 9532 17434
rect 9556 17382 9570 17434
rect 9570 17382 9582 17434
rect 9582 17382 9612 17434
rect 9636 17382 9646 17434
rect 9646 17382 9692 17434
rect 9396 17380 9452 17382
rect 9476 17380 9532 17382
rect 9556 17380 9612 17382
rect 9636 17380 9692 17382
rect 13617 16890 13673 16892
rect 13697 16890 13753 16892
rect 13777 16890 13833 16892
rect 13857 16890 13913 16892
rect 13617 16838 13663 16890
rect 13663 16838 13673 16890
rect 13697 16838 13727 16890
rect 13727 16838 13739 16890
rect 13739 16838 13753 16890
rect 13777 16838 13791 16890
rect 13791 16838 13803 16890
rect 13803 16838 13833 16890
rect 13857 16838 13867 16890
rect 13867 16838 13913 16890
rect 13617 16836 13673 16838
rect 13697 16836 13753 16838
rect 13777 16836 13833 16838
rect 13857 16836 13913 16838
rect 9396 16346 9452 16348
rect 9476 16346 9532 16348
rect 9556 16346 9612 16348
rect 9636 16346 9692 16348
rect 9396 16294 9442 16346
rect 9442 16294 9452 16346
rect 9476 16294 9506 16346
rect 9506 16294 9518 16346
rect 9518 16294 9532 16346
rect 9556 16294 9570 16346
rect 9570 16294 9582 16346
rect 9582 16294 9612 16346
rect 9636 16294 9646 16346
rect 9646 16294 9692 16346
rect 9396 16292 9452 16294
rect 9476 16292 9532 16294
rect 9556 16292 9612 16294
rect 9636 16292 9692 16294
rect 13617 15802 13673 15804
rect 13697 15802 13753 15804
rect 13777 15802 13833 15804
rect 13857 15802 13913 15804
rect 13617 15750 13663 15802
rect 13663 15750 13673 15802
rect 13697 15750 13727 15802
rect 13727 15750 13739 15802
rect 13739 15750 13753 15802
rect 13777 15750 13791 15802
rect 13791 15750 13803 15802
rect 13803 15750 13833 15802
rect 13857 15750 13867 15802
rect 13867 15750 13913 15802
rect 13617 15748 13673 15750
rect 13697 15748 13753 15750
rect 13777 15748 13833 15750
rect 13857 15748 13913 15750
rect 9396 15258 9452 15260
rect 9476 15258 9532 15260
rect 9556 15258 9612 15260
rect 9636 15258 9692 15260
rect 9396 15206 9442 15258
rect 9442 15206 9452 15258
rect 9476 15206 9506 15258
rect 9506 15206 9518 15258
rect 9518 15206 9532 15258
rect 9556 15206 9570 15258
rect 9570 15206 9582 15258
rect 9582 15206 9612 15258
rect 9636 15206 9646 15258
rect 9646 15206 9692 15258
rect 9396 15204 9452 15206
rect 9476 15204 9532 15206
rect 9556 15204 9612 15206
rect 9636 15204 9692 15206
rect 15750 24148 15752 24168
rect 15752 24148 15804 24168
rect 15804 24148 15806 24168
rect 15750 24112 15806 24148
rect 17837 39194 17893 39196
rect 17917 39194 17973 39196
rect 17997 39194 18053 39196
rect 18077 39194 18133 39196
rect 17837 39142 17883 39194
rect 17883 39142 17893 39194
rect 17917 39142 17947 39194
rect 17947 39142 17959 39194
rect 17959 39142 17973 39194
rect 17997 39142 18011 39194
rect 18011 39142 18023 39194
rect 18023 39142 18053 39194
rect 18077 39142 18087 39194
rect 18087 39142 18133 39194
rect 17837 39140 17893 39142
rect 17917 39140 17973 39142
rect 17997 39140 18053 39142
rect 18077 39140 18133 39142
rect 17837 38106 17893 38108
rect 17917 38106 17973 38108
rect 17997 38106 18053 38108
rect 18077 38106 18133 38108
rect 17837 38054 17883 38106
rect 17883 38054 17893 38106
rect 17917 38054 17947 38106
rect 17947 38054 17959 38106
rect 17959 38054 17973 38106
rect 17997 38054 18011 38106
rect 18011 38054 18023 38106
rect 18023 38054 18053 38106
rect 18077 38054 18087 38106
rect 18087 38054 18133 38106
rect 17837 38052 17893 38054
rect 17917 38052 17973 38054
rect 17997 38052 18053 38054
rect 18077 38052 18133 38054
rect 17837 37018 17893 37020
rect 17917 37018 17973 37020
rect 17997 37018 18053 37020
rect 18077 37018 18133 37020
rect 17837 36966 17883 37018
rect 17883 36966 17893 37018
rect 17917 36966 17947 37018
rect 17947 36966 17959 37018
rect 17959 36966 17973 37018
rect 17997 36966 18011 37018
rect 18011 36966 18023 37018
rect 18023 36966 18053 37018
rect 18077 36966 18087 37018
rect 18087 36966 18133 37018
rect 17837 36964 17893 36966
rect 17917 36964 17973 36966
rect 17997 36964 18053 36966
rect 18077 36964 18133 36966
rect 17590 36780 17646 36816
rect 17590 36760 17592 36780
rect 17592 36760 17644 36780
rect 17644 36760 17646 36780
rect 17837 35930 17893 35932
rect 17917 35930 17973 35932
rect 17997 35930 18053 35932
rect 18077 35930 18133 35932
rect 17837 35878 17883 35930
rect 17883 35878 17893 35930
rect 17917 35878 17947 35930
rect 17947 35878 17959 35930
rect 17959 35878 17973 35930
rect 17997 35878 18011 35930
rect 18011 35878 18023 35930
rect 18023 35878 18053 35930
rect 18077 35878 18087 35930
rect 18087 35878 18133 35930
rect 17837 35876 17893 35878
rect 17917 35876 17973 35878
rect 17997 35876 18053 35878
rect 18077 35876 18133 35878
rect 18878 37204 18880 37224
rect 18880 37204 18932 37224
rect 18932 37204 18934 37224
rect 18878 37168 18934 37204
rect 17837 34842 17893 34844
rect 17917 34842 17973 34844
rect 17997 34842 18053 34844
rect 18077 34842 18133 34844
rect 17837 34790 17883 34842
rect 17883 34790 17893 34842
rect 17917 34790 17947 34842
rect 17947 34790 17959 34842
rect 17959 34790 17973 34842
rect 17997 34790 18011 34842
rect 18011 34790 18023 34842
rect 18023 34790 18053 34842
rect 18077 34790 18087 34842
rect 18087 34790 18133 34842
rect 17837 34788 17893 34790
rect 17917 34788 17973 34790
rect 17997 34788 18053 34790
rect 18077 34788 18133 34790
rect 17590 34584 17646 34640
rect 17837 33754 17893 33756
rect 17917 33754 17973 33756
rect 17997 33754 18053 33756
rect 18077 33754 18133 33756
rect 17837 33702 17883 33754
rect 17883 33702 17893 33754
rect 17917 33702 17947 33754
rect 17947 33702 17959 33754
rect 17959 33702 17973 33754
rect 17997 33702 18011 33754
rect 18011 33702 18023 33754
rect 18023 33702 18053 33754
rect 18077 33702 18087 33754
rect 18087 33702 18133 33754
rect 17837 33700 17893 33702
rect 17917 33700 17973 33702
rect 17997 33700 18053 33702
rect 18077 33700 18133 33702
rect 17837 32666 17893 32668
rect 17917 32666 17973 32668
rect 17997 32666 18053 32668
rect 18077 32666 18133 32668
rect 17837 32614 17883 32666
rect 17883 32614 17893 32666
rect 17917 32614 17947 32666
rect 17947 32614 17959 32666
rect 17959 32614 17973 32666
rect 17997 32614 18011 32666
rect 18011 32614 18023 32666
rect 18023 32614 18053 32666
rect 18077 32614 18087 32666
rect 18087 32614 18133 32666
rect 17837 32612 17893 32614
rect 17917 32612 17973 32614
rect 17997 32612 18053 32614
rect 18077 32612 18133 32614
rect 16854 29144 16910 29200
rect 17590 28872 17646 28928
rect 17837 31578 17893 31580
rect 17917 31578 17973 31580
rect 17997 31578 18053 31580
rect 18077 31578 18133 31580
rect 17837 31526 17883 31578
rect 17883 31526 17893 31578
rect 17917 31526 17947 31578
rect 17947 31526 17959 31578
rect 17959 31526 17973 31578
rect 17997 31526 18011 31578
rect 18011 31526 18023 31578
rect 18023 31526 18053 31578
rect 18077 31526 18087 31578
rect 18087 31526 18133 31578
rect 17837 31524 17893 31526
rect 17917 31524 17973 31526
rect 17997 31524 18053 31526
rect 18077 31524 18133 31526
rect 17837 30490 17893 30492
rect 17917 30490 17973 30492
rect 17997 30490 18053 30492
rect 18077 30490 18133 30492
rect 17837 30438 17883 30490
rect 17883 30438 17893 30490
rect 17917 30438 17947 30490
rect 17947 30438 17959 30490
rect 17959 30438 17973 30490
rect 17997 30438 18011 30490
rect 18011 30438 18023 30490
rect 18023 30438 18053 30490
rect 18077 30438 18087 30490
rect 18087 30438 18133 30490
rect 17837 30436 17893 30438
rect 17917 30436 17973 30438
rect 17997 30436 18053 30438
rect 18077 30436 18133 30438
rect 17866 29688 17922 29744
rect 17837 29402 17893 29404
rect 17917 29402 17973 29404
rect 17997 29402 18053 29404
rect 18077 29402 18133 29404
rect 17837 29350 17883 29402
rect 17883 29350 17893 29402
rect 17917 29350 17947 29402
rect 17947 29350 17959 29402
rect 17959 29350 17973 29402
rect 17997 29350 18011 29402
rect 18011 29350 18023 29402
rect 18023 29350 18053 29402
rect 18077 29350 18087 29402
rect 18087 29350 18133 29402
rect 17837 29348 17893 29350
rect 17917 29348 17973 29350
rect 17997 29348 18053 29350
rect 18077 29348 18133 29350
rect 18326 29144 18382 29200
rect 18326 28600 18382 28656
rect 17837 28314 17893 28316
rect 17917 28314 17973 28316
rect 17997 28314 18053 28316
rect 18077 28314 18133 28316
rect 17837 28262 17883 28314
rect 17883 28262 17893 28314
rect 17917 28262 17947 28314
rect 17947 28262 17959 28314
rect 17959 28262 17973 28314
rect 17997 28262 18011 28314
rect 18011 28262 18023 28314
rect 18023 28262 18053 28314
rect 18077 28262 18087 28314
rect 18087 28262 18133 28314
rect 17837 28260 17893 28262
rect 17917 28260 17973 28262
rect 17997 28260 18053 28262
rect 18077 28260 18133 28262
rect 22058 39738 22114 39740
rect 22138 39738 22194 39740
rect 22218 39738 22274 39740
rect 22298 39738 22354 39740
rect 22058 39686 22104 39738
rect 22104 39686 22114 39738
rect 22138 39686 22168 39738
rect 22168 39686 22180 39738
rect 22180 39686 22194 39738
rect 22218 39686 22232 39738
rect 22232 39686 22244 39738
rect 22244 39686 22274 39738
rect 22298 39686 22308 39738
rect 22308 39686 22354 39738
rect 22058 39684 22114 39686
rect 22138 39684 22194 39686
rect 22218 39684 22274 39686
rect 22298 39684 22354 39686
rect 21454 38936 21510 38992
rect 21362 38256 21418 38312
rect 20626 36660 20628 36680
rect 20628 36660 20680 36680
rect 20680 36660 20682 36680
rect 20626 36624 20682 36660
rect 19798 35536 19854 35592
rect 19338 35128 19394 35184
rect 19430 32988 19432 33008
rect 19432 32988 19484 33008
rect 19484 32988 19486 33008
rect 19430 32952 19486 32988
rect 18694 29572 18750 29608
rect 18694 29552 18696 29572
rect 18696 29552 18748 29572
rect 18748 29552 18750 29572
rect 18602 29452 18604 29472
rect 18604 29452 18656 29472
rect 18656 29452 18658 29472
rect 18602 29416 18658 29452
rect 18970 28908 18972 28928
rect 18972 28908 19024 28928
rect 19024 28908 19026 28928
rect 18970 28872 19026 28908
rect 18970 28600 19026 28656
rect 17837 27226 17893 27228
rect 17917 27226 17973 27228
rect 17997 27226 18053 27228
rect 18077 27226 18133 27228
rect 17837 27174 17883 27226
rect 17883 27174 17893 27226
rect 17917 27174 17947 27226
rect 17947 27174 17959 27226
rect 17959 27174 17973 27226
rect 17997 27174 18011 27226
rect 18011 27174 18023 27226
rect 18023 27174 18053 27226
rect 18077 27174 18087 27226
rect 18087 27174 18133 27226
rect 17837 27172 17893 27174
rect 17917 27172 17973 27174
rect 17997 27172 18053 27174
rect 18077 27172 18133 27174
rect 18694 27512 18750 27568
rect 17837 26138 17893 26140
rect 17917 26138 17973 26140
rect 17997 26138 18053 26140
rect 18077 26138 18133 26140
rect 17837 26086 17883 26138
rect 17883 26086 17893 26138
rect 17917 26086 17947 26138
rect 17947 26086 17959 26138
rect 17959 26086 17973 26138
rect 17997 26086 18011 26138
rect 18011 26086 18023 26138
rect 18023 26086 18053 26138
rect 18077 26086 18087 26138
rect 18087 26086 18133 26138
rect 17837 26084 17893 26086
rect 17917 26084 17973 26086
rect 17997 26084 18053 26086
rect 18077 26084 18133 26086
rect 18050 25220 18106 25256
rect 18050 25200 18052 25220
rect 18052 25200 18104 25220
rect 18104 25200 18106 25220
rect 17130 24112 17186 24168
rect 17837 25050 17893 25052
rect 17917 25050 17973 25052
rect 17997 25050 18053 25052
rect 18077 25050 18133 25052
rect 17837 24998 17883 25050
rect 17883 24998 17893 25050
rect 17917 24998 17947 25050
rect 17947 24998 17959 25050
rect 17959 24998 17973 25050
rect 17997 24998 18011 25050
rect 18011 24998 18023 25050
rect 18023 24998 18053 25050
rect 18077 24998 18087 25050
rect 18087 24998 18133 25050
rect 17837 24996 17893 24998
rect 17917 24996 17973 24998
rect 17997 24996 18053 24998
rect 18077 24996 18133 24998
rect 19614 30268 19616 30288
rect 19616 30268 19668 30288
rect 19668 30268 19670 30288
rect 19614 30232 19670 30268
rect 19614 30096 19670 30152
rect 19246 29572 19302 29608
rect 19246 29552 19248 29572
rect 19248 29552 19300 29572
rect 19300 29552 19302 29572
rect 19062 26832 19118 26888
rect 18970 26460 18972 26480
rect 18972 26460 19024 26480
rect 19024 26460 19026 26480
rect 18970 26424 19026 26460
rect 17837 23962 17893 23964
rect 17917 23962 17973 23964
rect 17997 23962 18053 23964
rect 18077 23962 18133 23964
rect 17837 23910 17883 23962
rect 17883 23910 17893 23962
rect 17917 23910 17947 23962
rect 17947 23910 17959 23962
rect 17959 23910 17973 23962
rect 17997 23910 18011 23962
rect 18011 23910 18023 23962
rect 18023 23910 18053 23962
rect 18077 23910 18087 23962
rect 18087 23910 18133 23962
rect 17837 23908 17893 23910
rect 17917 23908 17973 23910
rect 17997 23908 18053 23910
rect 18077 23908 18133 23910
rect 17958 23724 18014 23760
rect 17958 23704 17960 23724
rect 17960 23704 18012 23724
rect 18012 23704 18014 23724
rect 17837 22874 17893 22876
rect 17917 22874 17973 22876
rect 17997 22874 18053 22876
rect 18077 22874 18133 22876
rect 17837 22822 17883 22874
rect 17883 22822 17893 22874
rect 17917 22822 17947 22874
rect 17947 22822 17959 22874
rect 17959 22822 17973 22874
rect 17997 22822 18011 22874
rect 18011 22822 18023 22874
rect 18023 22822 18053 22874
rect 18077 22822 18087 22874
rect 18087 22822 18133 22874
rect 17837 22820 17893 22822
rect 17917 22820 17973 22822
rect 17997 22820 18053 22822
rect 18077 22820 18133 22822
rect 17837 21786 17893 21788
rect 17917 21786 17973 21788
rect 17997 21786 18053 21788
rect 18077 21786 18133 21788
rect 17837 21734 17883 21786
rect 17883 21734 17893 21786
rect 17917 21734 17947 21786
rect 17947 21734 17959 21786
rect 17959 21734 17973 21786
rect 17997 21734 18011 21786
rect 18011 21734 18023 21786
rect 18023 21734 18053 21786
rect 18077 21734 18087 21786
rect 18087 21734 18133 21786
rect 17837 21732 17893 21734
rect 17917 21732 17973 21734
rect 17997 21732 18053 21734
rect 18077 21732 18133 21734
rect 17837 20698 17893 20700
rect 17917 20698 17973 20700
rect 17997 20698 18053 20700
rect 18077 20698 18133 20700
rect 17837 20646 17883 20698
rect 17883 20646 17893 20698
rect 17917 20646 17947 20698
rect 17947 20646 17959 20698
rect 17959 20646 17973 20698
rect 17997 20646 18011 20698
rect 18011 20646 18023 20698
rect 18023 20646 18053 20698
rect 18077 20646 18087 20698
rect 18087 20646 18133 20698
rect 17837 20644 17893 20646
rect 17917 20644 17973 20646
rect 17997 20644 18053 20646
rect 18077 20644 18133 20646
rect 17837 19610 17893 19612
rect 17917 19610 17973 19612
rect 17997 19610 18053 19612
rect 18077 19610 18133 19612
rect 17837 19558 17883 19610
rect 17883 19558 17893 19610
rect 17917 19558 17947 19610
rect 17947 19558 17959 19610
rect 17959 19558 17973 19610
rect 17997 19558 18011 19610
rect 18011 19558 18023 19610
rect 18023 19558 18053 19610
rect 18077 19558 18087 19610
rect 18087 19558 18133 19610
rect 17837 19556 17893 19558
rect 17917 19556 17973 19558
rect 17997 19556 18053 19558
rect 18077 19556 18133 19558
rect 17837 18522 17893 18524
rect 17917 18522 17973 18524
rect 17997 18522 18053 18524
rect 18077 18522 18133 18524
rect 17837 18470 17883 18522
rect 17883 18470 17893 18522
rect 17917 18470 17947 18522
rect 17947 18470 17959 18522
rect 17959 18470 17973 18522
rect 17997 18470 18011 18522
rect 18011 18470 18023 18522
rect 18023 18470 18053 18522
rect 18077 18470 18087 18522
rect 18087 18470 18133 18522
rect 17837 18468 17893 18470
rect 17917 18468 17973 18470
rect 17997 18468 18053 18470
rect 18077 18468 18133 18470
rect 17837 17434 17893 17436
rect 17917 17434 17973 17436
rect 17997 17434 18053 17436
rect 18077 17434 18133 17436
rect 17837 17382 17883 17434
rect 17883 17382 17893 17434
rect 17917 17382 17947 17434
rect 17947 17382 17959 17434
rect 17959 17382 17973 17434
rect 17997 17382 18011 17434
rect 18011 17382 18023 17434
rect 18023 17382 18053 17434
rect 18077 17382 18087 17434
rect 18087 17382 18133 17434
rect 17837 17380 17893 17382
rect 17917 17380 17973 17382
rect 17997 17380 18053 17382
rect 18077 17380 18133 17382
rect 17837 16346 17893 16348
rect 17917 16346 17973 16348
rect 17997 16346 18053 16348
rect 18077 16346 18133 16348
rect 17837 16294 17883 16346
rect 17883 16294 17893 16346
rect 17917 16294 17947 16346
rect 17947 16294 17959 16346
rect 17959 16294 17973 16346
rect 17997 16294 18011 16346
rect 18011 16294 18023 16346
rect 18023 16294 18053 16346
rect 18077 16294 18087 16346
rect 18087 16294 18133 16346
rect 17837 16292 17893 16294
rect 17917 16292 17973 16294
rect 17997 16292 18053 16294
rect 18077 16292 18133 16294
rect 17837 15258 17893 15260
rect 17917 15258 17973 15260
rect 17997 15258 18053 15260
rect 18077 15258 18133 15260
rect 17837 15206 17883 15258
rect 17883 15206 17893 15258
rect 17917 15206 17947 15258
rect 17947 15206 17959 15258
rect 17959 15206 17973 15258
rect 17997 15206 18011 15258
rect 18011 15206 18023 15258
rect 18023 15206 18053 15258
rect 18077 15206 18087 15258
rect 18087 15206 18133 15258
rect 17837 15204 17893 15206
rect 17917 15204 17973 15206
rect 17997 15204 18053 15206
rect 18077 15204 18133 15206
rect 13617 14714 13673 14716
rect 13697 14714 13753 14716
rect 13777 14714 13833 14716
rect 13857 14714 13913 14716
rect 13617 14662 13663 14714
rect 13663 14662 13673 14714
rect 13697 14662 13727 14714
rect 13727 14662 13739 14714
rect 13739 14662 13753 14714
rect 13777 14662 13791 14714
rect 13791 14662 13803 14714
rect 13803 14662 13833 14714
rect 13857 14662 13867 14714
rect 13867 14662 13913 14714
rect 13617 14660 13673 14662
rect 13697 14660 13753 14662
rect 13777 14660 13833 14662
rect 13857 14660 13913 14662
rect 9396 14170 9452 14172
rect 9476 14170 9532 14172
rect 9556 14170 9612 14172
rect 9636 14170 9692 14172
rect 9396 14118 9442 14170
rect 9442 14118 9452 14170
rect 9476 14118 9506 14170
rect 9506 14118 9518 14170
rect 9518 14118 9532 14170
rect 9556 14118 9570 14170
rect 9570 14118 9582 14170
rect 9582 14118 9612 14170
rect 9636 14118 9646 14170
rect 9646 14118 9692 14170
rect 9396 14116 9452 14118
rect 9476 14116 9532 14118
rect 9556 14116 9612 14118
rect 9636 14116 9692 14118
rect 17837 14170 17893 14172
rect 17917 14170 17973 14172
rect 17997 14170 18053 14172
rect 18077 14170 18133 14172
rect 17837 14118 17883 14170
rect 17883 14118 17893 14170
rect 17917 14118 17947 14170
rect 17947 14118 17959 14170
rect 17959 14118 17973 14170
rect 17997 14118 18011 14170
rect 18011 14118 18023 14170
rect 18023 14118 18053 14170
rect 18077 14118 18087 14170
rect 18087 14118 18133 14170
rect 17837 14116 17893 14118
rect 17917 14116 17973 14118
rect 17997 14116 18053 14118
rect 18077 14116 18133 14118
rect 13617 13626 13673 13628
rect 13697 13626 13753 13628
rect 13777 13626 13833 13628
rect 13857 13626 13913 13628
rect 13617 13574 13663 13626
rect 13663 13574 13673 13626
rect 13697 13574 13727 13626
rect 13727 13574 13739 13626
rect 13739 13574 13753 13626
rect 13777 13574 13791 13626
rect 13791 13574 13803 13626
rect 13803 13574 13833 13626
rect 13857 13574 13867 13626
rect 13867 13574 13913 13626
rect 13617 13572 13673 13574
rect 13697 13572 13753 13574
rect 13777 13572 13833 13574
rect 13857 13572 13913 13574
rect 9396 13082 9452 13084
rect 9476 13082 9532 13084
rect 9556 13082 9612 13084
rect 9636 13082 9692 13084
rect 9396 13030 9442 13082
rect 9442 13030 9452 13082
rect 9476 13030 9506 13082
rect 9506 13030 9518 13082
rect 9518 13030 9532 13082
rect 9556 13030 9570 13082
rect 9570 13030 9582 13082
rect 9582 13030 9612 13082
rect 9636 13030 9646 13082
rect 9646 13030 9692 13082
rect 9396 13028 9452 13030
rect 9476 13028 9532 13030
rect 9556 13028 9612 13030
rect 9636 13028 9692 13030
rect 17837 13082 17893 13084
rect 17917 13082 17973 13084
rect 17997 13082 18053 13084
rect 18077 13082 18133 13084
rect 17837 13030 17883 13082
rect 17883 13030 17893 13082
rect 17917 13030 17947 13082
rect 17947 13030 17959 13082
rect 17959 13030 17973 13082
rect 17997 13030 18011 13082
rect 18011 13030 18023 13082
rect 18023 13030 18053 13082
rect 18077 13030 18087 13082
rect 18087 13030 18133 13082
rect 17837 13028 17893 13030
rect 17917 13028 17973 13030
rect 17997 13028 18053 13030
rect 18077 13028 18133 13030
rect 13617 12538 13673 12540
rect 13697 12538 13753 12540
rect 13777 12538 13833 12540
rect 13857 12538 13913 12540
rect 13617 12486 13663 12538
rect 13663 12486 13673 12538
rect 13697 12486 13727 12538
rect 13727 12486 13739 12538
rect 13739 12486 13753 12538
rect 13777 12486 13791 12538
rect 13791 12486 13803 12538
rect 13803 12486 13833 12538
rect 13857 12486 13867 12538
rect 13867 12486 13913 12538
rect 13617 12484 13673 12486
rect 13697 12484 13753 12486
rect 13777 12484 13833 12486
rect 13857 12484 13913 12486
rect 9396 11994 9452 11996
rect 9476 11994 9532 11996
rect 9556 11994 9612 11996
rect 9636 11994 9692 11996
rect 9396 11942 9442 11994
rect 9442 11942 9452 11994
rect 9476 11942 9506 11994
rect 9506 11942 9518 11994
rect 9518 11942 9532 11994
rect 9556 11942 9570 11994
rect 9570 11942 9582 11994
rect 9582 11942 9612 11994
rect 9636 11942 9646 11994
rect 9646 11942 9692 11994
rect 9396 11940 9452 11942
rect 9476 11940 9532 11942
rect 9556 11940 9612 11942
rect 9636 11940 9692 11942
rect 13617 11450 13673 11452
rect 13697 11450 13753 11452
rect 13777 11450 13833 11452
rect 13857 11450 13913 11452
rect 13617 11398 13663 11450
rect 13663 11398 13673 11450
rect 13697 11398 13727 11450
rect 13727 11398 13739 11450
rect 13739 11398 13753 11450
rect 13777 11398 13791 11450
rect 13791 11398 13803 11450
rect 13803 11398 13833 11450
rect 13857 11398 13867 11450
rect 13867 11398 13913 11450
rect 13617 11396 13673 11398
rect 13697 11396 13753 11398
rect 13777 11396 13833 11398
rect 13857 11396 13913 11398
rect 9396 10906 9452 10908
rect 9476 10906 9532 10908
rect 9556 10906 9612 10908
rect 9636 10906 9692 10908
rect 9396 10854 9442 10906
rect 9442 10854 9452 10906
rect 9476 10854 9506 10906
rect 9506 10854 9518 10906
rect 9518 10854 9532 10906
rect 9556 10854 9570 10906
rect 9570 10854 9582 10906
rect 9582 10854 9612 10906
rect 9636 10854 9646 10906
rect 9646 10854 9692 10906
rect 9396 10852 9452 10854
rect 9476 10852 9532 10854
rect 9556 10852 9612 10854
rect 9636 10852 9692 10854
rect 13617 10362 13673 10364
rect 13697 10362 13753 10364
rect 13777 10362 13833 10364
rect 13857 10362 13913 10364
rect 13617 10310 13663 10362
rect 13663 10310 13673 10362
rect 13697 10310 13727 10362
rect 13727 10310 13739 10362
rect 13739 10310 13753 10362
rect 13777 10310 13791 10362
rect 13791 10310 13803 10362
rect 13803 10310 13833 10362
rect 13857 10310 13867 10362
rect 13867 10310 13913 10362
rect 13617 10308 13673 10310
rect 13697 10308 13753 10310
rect 13777 10308 13833 10310
rect 13857 10308 13913 10310
rect 9396 9818 9452 9820
rect 9476 9818 9532 9820
rect 9556 9818 9612 9820
rect 9636 9818 9692 9820
rect 9396 9766 9442 9818
rect 9442 9766 9452 9818
rect 9476 9766 9506 9818
rect 9506 9766 9518 9818
rect 9518 9766 9532 9818
rect 9556 9766 9570 9818
rect 9570 9766 9582 9818
rect 9582 9766 9612 9818
rect 9636 9766 9646 9818
rect 9646 9766 9692 9818
rect 9396 9764 9452 9766
rect 9476 9764 9532 9766
rect 9556 9764 9612 9766
rect 9636 9764 9692 9766
rect 5176 7098 5232 7100
rect 5256 7098 5312 7100
rect 5336 7098 5392 7100
rect 5416 7098 5472 7100
rect 5176 7046 5222 7098
rect 5222 7046 5232 7098
rect 5256 7046 5286 7098
rect 5286 7046 5298 7098
rect 5298 7046 5312 7098
rect 5336 7046 5350 7098
rect 5350 7046 5362 7098
rect 5362 7046 5392 7098
rect 5416 7046 5426 7098
rect 5426 7046 5472 7098
rect 5176 7044 5232 7046
rect 5256 7044 5312 7046
rect 5336 7044 5392 7046
rect 5416 7044 5472 7046
rect 13617 9274 13673 9276
rect 13697 9274 13753 9276
rect 13777 9274 13833 9276
rect 13857 9274 13913 9276
rect 13617 9222 13663 9274
rect 13663 9222 13673 9274
rect 13697 9222 13727 9274
rect 13727 9222 13739 9274
rect 13739 9222 13753 9274
rect 13777 9222 13791 9274
rect 13791 9222 13803 9274
rect 13803 9222 13833 9274
rect 13857 9222 13867 9274
rect 13867 9222 13913 9274
rect 13617 9220 13673 9222
rect 13697 9220 13753 9222
rect 13777 9220 13833 9222
rect 13857 9220 13913 9222
rect 9396 8730 9452 8732
rect 9476 8730 9532 8732
rect 9556 8730 9612 8732
rect 9636 8730 9692 8732
rect 9396 8678 9442 8730
rect 9442 8678 9452 8730
rect 9476 8678 9506 8730
rect 9506 8678 9518 8730
rect 9518 8678 9532 8730
rect 9556 8678 9570 8730
rect 9570 8678 9582 8730
rect 9582 8678 9612 8730
rect 9636 8678 9646 8730
rect 9646 8678 9692 8730
rect 9396 8676 9452 8678
rect 9476 8676 9532 8678
rect 9556 8676 9612 8678
rect 9636 8676 9692 8678
rect 13617 8186 13673 8188
rect 13697 8186 13753 8188
rect 13777 8186 13833 8188
rect 13857 8186 13913 8188
rect 13617 8134 13663 8186
rect 13663 8134 13673 8186
rect 13697 8134 13727 8186
rect 13727 8134 13739 8186
rect 13739 8134 13753 8186
rect 13777 8134 13791 8186
rect 13791 8134 13803 8186
rect 13803 8134 13833 8186
rect 13857 8134 13867 8186
rect 13867 8134 13913 8186
rect 13617 8132 13673 8134
rect 13697 8132 13753 8134
rect 13777 8132 13833 8134
rect 13857 8132 13913 8134
rect 9396 7642 9452 7644
rect 9476 7642 9532 7644
rect 9556 7642 9612 7644
rect 9636 7642 9692 7644
rect 9396 7590 9442 7642
rect 9442 7590 9452 7642
rect 9476 7590 9506 7642
rect 9506 7590 9518 7642
rect 9518 7590 9532 7642
rect 9556 7590 9570 7642
rect 9570 7590 9582 7642
rect 9582 7590 9612 7642
rect 9636 7590 9646 7642
rect 9646 7590 9692 7642
rect 9396 7588 9452 7590
rect 9476 7588 9532 7590
rect 9556 7588 9612 7590
rect 9636 7588 9692 7590
rect 13617 7098 13673 7100
rect 13697 7098 13753 7100
rect 13777 7098 13833 7100
rect 13857 7098 13913 7100
rect 13617 7046 13663 7098
rect 13663 7046 13673 7098
rect 13697 7046 13727 7098
rect 13727 7046 13739 7098
rect 13739 7046 13753 7098
rect 13777 7046 13791 7098
rect 13791 7046 13803 7098
rect 13803 7046 13833 7098
rect 13857 7046 13867 7098
rect 13867 7046 13913 7098
rect 13617 7044 13673 7046
rect 13697 7044 13753 7046
rect 13777 7044 13833 7046
rect 13857 7044 13913 7046
rect 5176 6010 5232 6012
rect 5256 6010 5312 6012
rect 5336 6010 5392 6012
rect 5416 6010 5472 6012
rect 5176 5958 5222 6010
rect 5222 5958 5232 6010
rect 5256 5958 5286 6010
rect 5286 5958 5298 6010
rect 5298 5958 5312 6010
rect 5336 5958 5350 6010
rect 5350 5958 5362 6010
rect 5362 5958 5392 6010
rect 5416 5958 5426 6010
rect 5426 5958 5472 6010
rect 5176 5956 5232 5958
rect 5256 5956 5312 5958
rect 5336 5956 5392 5958
rect 5416 5956 5472 5958
rect 5176 4922 5232 4924
rect 5256 4922 5312 4924
rect 5336 4922 5392 4924
rect 5416 4922 5472 4924
rect 5176 4870 5222 4922
rect 5222 4870 5232 4922
rect 5256 4870 5286 4922
rect 5286 4870 5298 4922
rect 5298 4870 5312 4922
rect 5336 4870 5350 4922
rect 5350 4870 5362 4922
rect 5362 4870 5392 4922
rect 5416 4870 5426 4922
rect 5426 4870 5472 4922
rect 5176 4868 5232 4870
rect 5256 4868 5312 4870
rect 5336 4868 5392 4870
rect 5416 4868 5472 4870
rect 5176 3834 5232 3836
rect 5256 3834 5312 3836
rect 5336 3834 5392 3836
rect 5416 3834 5472 3836
rect 5176 3782 5222 3834
rect 5222 3782 5232 3834
rect 5256 3782 5286 3834
rect 5286 3782 5298 3834
rect 5298 3782 5312 3834
rect 5336 3782 5350 3834
rect 5350 3782 5362 3834
rect 5362 3782 5392 3834
rect 5416 3782 5426 3834
rect 5426 3782 5472 3834
rect 5176 3780 5232 3782
rect 5256 3780 5312 3782
rect 5336 3780 5392 3782
rect 5416 3780 5472 3782
rect 5176 2746 5232 2748
rect 5256 2746 5312 2748
rect 5336 2746 5392 2748
rect 5416 2746 5472 2748
rect 5176 2694 5222 2746
rect 5222 2694 5232 2746
rect 5256 2694 5286 2746
rect 5286 2694 5298 2746
rect 5298 2694 5312 2746
rect 5336 2694 5350 2746
rect 5350 2694 5362 2746
rect 5362 2694 5392 2746
rect 5416 2694 5426 2746
rect 5426 2694 5472 2746
rect 5176 2692 5232 2694
rect 5256 2692 5312 2694
rect 5336 2692 5392 2694
rect 5416 2692 5472 2694
rect 9396 6554 9452 6556
rect 9476 6554 9532 6556
rect 9556 6554 9612 6556
rect 9636 6554 9692 6556
rect 9396 6502 9442 6554
rect 9442 6502 9452 6554
rect 9476 6502 9506 6554
rect 9506 6502 9518 6554
rect 9518 6502 9532 6554
rect 9556 6502 9570 6554
rect 9570 6502 9582 6554
rect 9582 6502 9612 6554
rect 9636 6502 9646 6554
rect 9646 6502 9692 6554
rect 9396 6500 9452 6502
rect 9476 6500 9532 6502
rect 9556 6500 9612 6502
rect 9636 6500 9692 6502
rect 9396 5466 9452 5468
rect 9476 5466 9532 5468
rect 9556 5466 9612 5468
rect 9636 5466 9692 5468
rect 9396 5414 9442 5466
rect 9442 5414 9452 5466
rect 9476 5414 9506 5466
rect 9506 5414 9518 5466
rect 9518 5414 9532 5466
rect 9556 5414 9570 5466
rect 9570 5414 9582 5466
rect 9582 5414 9612 5466
rect 9636 5414 9646 5466
rect 9646 5414 9692 5466
rect 9396 5412 9452 5414
rect 9476 5412 9532 5414
rect 9556 5412 9612 5414
rect 9636 5412 9692 5414
rect 9396 4378 9452 4380
rect 9476 4378 9532 4380
rect 9556 4378 9612 4380
rect 9636 4378 9692 4380
rect 9396 4326 9442 4378
rect 9442 4326 9452 4378
rect 9476 4326 9506 4378
rect 9506 4326 9518 4378
rect 9518 4326 9532 4378
rect 9556 4326 9570 4378
rect 9570 4326 9582 4378
rect 9582 4326 9612 4378
rect 9636 4326 9646 4378
rect 9646 4326 9692 4378
rect 9396 4324 9452 4326
rect 9476 4324 9532 4326
rect 9556 4324 9612 4326
rect 9636 4324 9692 4326
rect 13617 6010 13673 6012
rect 13697 6010 13753 6012
rect 13777 6010 13833 6012
rect 13857 6010 13913 6012
rect 13617 5958 13663 6010
rect 13663 5958 13673 6010
rect 13697 5958 13727 6010
rect 13727 5958 13739 6010
rect 13739 5958 13753 6010
rect 13777 5958 13791 6010
rect 13791 5958 13803 6010
rect 13803 5958 13833 6010
rect 13857 5958 13867 6010
rect 13867 5958 13913 6010
rect 13617 5956 13673 5958
rect 13697 5956 13753 5958
rect 13777 5956 13833 5958
rect 13857 5956 13913 5958
rect 9396 3290 9452 3292
rect 9476 3290 9532 3292
rect 9556 3290 9612 3292
rect 9636 3290 9692 3292
rect 9396 3238 9442 3290
rect 9442 3238 9452 3290
rect 9476 3238 9506 3290
rect 9506 3238 9518 3290
rect 9518 3238 9532 3290
rect 9556 3238 9570 3290
rect 9570 3238 9582 3290
rect 9582 3238 9612 3290
rect 9636 3238 9646 3290
rect 9646 3238 9692 3290
rect 9396 3236 9452 3238
rect 9476 3236 9532 3238
rect 9556 3236 9612 3238
rect 9636 3236 9692 3238
rect 13617 4922 13673 4924
rect 13697 4922 13753 4924
rect 13777 4922 13833 4924
rect 13857 4922 13913 4924
rect 13617 4870 13663 4922
rect 13663 4870 13673 4922
rect 13697 4870 13727 4922
rect 13727 4870 13739 4922
rect 13739 4870 13753 4922
rect 13777 4870 13791 4922
rect 13791 4870 13803 4922
rect 13803 4870 13833 4922
rect 13857 4870 13867 4922
rect 13867 4870 13913 4922
rect 13617 4868 13673 4870
rect 13697 4868 13753 4870
rect 13777 4868 13833 4870
rect 13857 4868 13913 4870
rect 9396 2202 9452 2204
rect 9476 2202 9532 2204
rect 9556 2202 9612 2204
rect 9636 2202 9692 2204
rect 9396 2150 9442 2202
rect 9442 2150 9452 2202
rect 9476 2150 9506 2202
rect 9506 2150 9518 2202
rect 9518 2150 9532 2202
rect 9556 2150 9570 2202
rect 9570 2150 9582 2202
rect 9582 2150 9612 2202
rect 9636 2150 9646 2202
rect 9646 2150 9692 2202
rect 9396 2148 9452 2150
rect 9476 2148 9532 2150
rect 9556 2148 9612 2150
rect 9636 2148 9692 2150
rect 13617 3834 13673 3836
rect 13697 3834 13753 3836
rect 13777 3834 13833 3836
rect 13857 3834 13913 3836
rect 13617 3782 13663 3834
rect 13663 3782 13673 3834
rect 13697 3782 13727 3834
rect 13727 3782 13739 3834
rect 13739 3782 13753 3834
rect 13777 3782 13791 3834
rect 13791 3782 13803 3834
rect 13803 3782 13833 3834
rect 13857 3782 13867 3834
rect 13867 3782 13913 3834
rect 13617 3780 13673 3782
rect 13697 3780 13753 3782
rect 13777 3780 13833 3782
rect 13857 3780 13913 3782
rect 17837 11994 17893 11996
rect 17917 11994 17973 11996
rect 17997 11994 18053 11996
rect 18077 11994 18133 11996
rect 17837 11942 17883 11994
rect 17883 11942 17893 11994
rect 17917 11942 17947 11994
rect 17947 11942 17959 11994
rect 17959 11942 17973 11994
rect 17997 11942 18011 11994
rect 18011 11942 18023 11994
rect 18023 11942 18053 11994
rect 18077 11942 18087 11994
rect 18087 11942 18133 11994
rect 17837 11940 17893 11942
rect 17917 11940 17973 11942
rect 17997 11940 18053 11942
rect 18077 11940 18133 11942
rect 17837 10906 17893 10908
rect 17917 10906 17973 10908
rect 17997 10906 18053 10908
rect 18077 10906 18133 10908
rect 17837 10854 17883 10906
rect 17883 10854 17893 10906
rect 17917 10854 17947 10906
rect 17947 10854 17959 10906
rect 17959 10854 17973 10906
rect 17997 10854 18011 10906
rect 18011 10854 18023 10906
rect 18023 10854 18053 10906
rect 18077 10854 18087 10906
rect 18087 10854 18133 10906
rect 17837 10852 17893 10854
rect 17917 10852 17973 10854
rect 17997 10852 18053 10854
rect 18077 10852 18133 10854
rect 17837 9818 17893 9820
rect 17917 9818 17973 9820
rect 17997 9818 18053 9820
rect 18077 9818 18133 9820
rect 17837 9766 17883 9818
rect 17883 9766 17893 9818
rect 17917 9766 17947 9818
rect 17947 9766 17959 9818
rect 17959 9766 17973 9818
rect 17997 9766 18011 9818
rect 18011 9766 18023 9818
rect 18023 9766 18053 9818
rect 18077 9766 18087 9818
rect 18087 9766 18133 9818
rect 17837 9764 17893 9766
rect 17917 9764 17973 9766
rect 17997 9764 18053 9766
rect 18077 9764 18133 9766
rect 17837 8730 17893 8732
rect 17917 8730 17973 8732
rect 17997 8730 18053 8732
rect 18077 8730 18133 8732
rect 17837 8678 17883 8730
rect 17883 8678 17893 8730
rect 17917 8678 17947 8730
rect 17947 8678 17959 8730
rect 17959 8678 17973 8730
rect 17997 8678 18011 8730
rect 18011 8678 18023 8730
rect 18023 8678 18053 8730
rect 18077 8678 18087 8730
rect 18087 8678 18133 8730
rect 17837 8676 17893 8678
rect 17917 8676 17973 8678
rect 17997 8676 18053 8678
rect 18077 8676 18133 8678
rect 17837 7642 17893 7644
rect 17917 7642 17973 7644
rect 17997 7642 18053 7644
rect 18077 7642 18133 7644
rect 17837 7590 17883 7642
rect 17883 7590 17893 7642
rect 17917 7590 17947 7642
rect 17947 7590 17959 7642
rect 17959 7590 17973 7642
rect 17997 7590 18011 7642
rect 18011 7590 18023 7642
rect 18023 7590 18053 7642
rect 18077 7590 18087 7642
rect 18087 7590 18133 7642
rect 17837 7588 17893 7590
rect 17917 7588 17973 7590
rect 17997 7588 18053 7590
rect 18077 7588 18133 7590
rect 19982 33652 20038 33688
rect 19982 33632 19984 33652
rect 19984 33632 20036 33652
rect 20036 33632 20038 33652
rect 20626 35672 20682 35728
rect 22058 38650 22114 38652
rect 22138 38650 22194 38652
rect 22218 38650 22274 38652
rect 22298 38650 22354 38652
rect 22058 38598 22104 38650
rect 22104 38598 22114 38650
rect 22138 38598 22168 38650
rect 22168 38598 22180 38650
rect 22180 38598 22194 38650
rect 22218 38598 22232 38650
rect 22232 38598 22244 38650
rect 22244 38598 22274 38650
rect 22298 38598 22308 38650
rect 22308 38598 22354 38650
rect 22058 38596 22114 38598
rect 22138 38596 22194 38598
rect 22218 38596 22274 38598
rect 22298 38596 22354 38598
rect 23754 37848 23810 37904
rect 22058 37562 22114 37564
rect 22138 37562 22194 37564
rect 22218 37562 22274 37564
rect 22298 37562 22354 37564
rect 22058 37510 22104 37562
rect 22104 37510 22114 37562
rect 22138 37510 22168 37562
rect 22168 37510 22180 37562
rect 22180 37510 22194 37562
rect 22218 37510 22232 37562
rect 22232 37510 22244 37562
rect 22244 37510 22274 37562
rect 22298 37510 22308 37562
rect 22308 37510 22354 37562
rect 22058 37508 22114 37510
rect 22138 37508 22194 37510
rect 22218 37508 22274 37510
rect 22298 37508 22354 37510
rect 22058 36474 22114 36476
rect 22138 36474 22194 36476
rect 22218 36474 22274 36476
rect 22298 36474 22354 36476
rect 22058 36422 22104 36474
rect 22104 36422 22114 36474
rect 22138 36422 22168 36474
rect 22168 36422 22180 36474
rect 22180 36422 22194 36474
rect 22218 36422 22232 36474
rect 22232 36422 22244 36474
rect 22244 36422 22274 36474
rect 22298 36422 22308 36474
rect 22308 36422 22354 36474
rect 22058 36420 22114 36422
rect 22138 36420 22194 36422
rect 22218 36420 22274 36422
rect 22298 36420 22354 36422
rect 21178 33904 21234 33960
rect 21270 33516 21326 33552
rect 21270 33496 21272 33516
rect 21272 33496 21324 33516
rect 21324 33496 21326 33516
rect 20626 32972 20682 33008
rect 20626 32952 20628 32972
rect 20628 32952 20680 32972
rect 20680 32952 20682 32972
rect 21454 34992 21510 35048
rect 21730 33652 21786 33688
rect 21730 33632 21732 33652
rect 21732 33632 21784 33652
rect 21784 33632 21786 33652
rect 22282 35808 22338 35864
rect 22466 36352 22522 36408
rect 22058 35386 22114 35388
rect 22138 35386 22194 35388
rect 22218 35386 22274 35388
rect 22298 35386 22354 35388
rect 22058 35334 22104 35386
rect 22104 35334 22114 35386
rect 22138 35334 22168 35386
rect 22168 35334 22180 35386
rect 22180 35334 22194 35386
rect 22218 35334 22232 35386
rect 22232 35334 22244 35386
rect 22244 35334 22274 35386
rect 22298 35334 22308 35386
rect 22308 35334 22354 35386
rect 22058 35332 22114 35334
rect 22138 35332 22194 35334
rect 22218 35332 22274 35334
rect 22298 35332 22354 35334
rect 22058 34298 22114 34300
rect 22138 34298 22194 34300
rect 22218 34298 22274 34300
rect 22298 34298 22354 34300
rect 22058 34246 22104 34298
rect 22104 34246 22114 34298
rect 22138 34246 22168 34298
rect 22168 34246 22180 34298
rect 22180 34246 22194 34298
rect 22218 34246 22232 34298
rect 22232 34246 22244 34298
rect 22244 34246 22274 34298
rect 22298 34246 22308 34298
rect 22308 34246 22354 34298
rect 22058 34244 22114 34246
rect 22138 34244 22194 34246
rect 22218 34244 22274 34246
rect 22298 34244 22354 34246
rect 22058 33210 22114 33212
rect 22138 33210 22194 33212
rect 22218 33210 22274 33212
rect 22298 33210 22354 33212
rect 22058 33158 22104 33210
rect 22104 33158 22114 33210
rect 22138 33158 22168 33210
rect 22168 33158 22180 33210
rect 22180 33158 22194 33210
rect 22218 33158 22232 33210
rect 22232 33158 22244 33210
rect 22244 33158 22274 33210
rect 22298 33158 22308 33210
rect 22308 33158 22354 33210
rect 22058 33156 22114 33158
rect 22138 33156 22194 33158
rect 22218 33156 22274 33158
rect 22298 33156 22354 33158
rect 23478 37032 23534 37088
rect 22742 34992 22798 35048
rect 23294 36216 23350 36272
rect 23478 34176 23534 34232
rect 24030 37440 24086 37496
rect 25042 37712 25098 37768
rect 24674 37032 24730 37088
rect 24490 35808 24546 35864
rect 24122 34992 24178 35048
rect 23662 33496 23718 33552
rect 22650 32308 22652 32328
rect 22652 32308 22704 32328
rect 22704 32308 22706 32328
rect 22650 32272 22706 32308
rect 20626 31320 20682 31376
rect 22058 32122 22114 32124
rect 22138 32122 22194 32124
rect 22218 32122 22274 32124
rect 22298 32122 22354 32124
rect 22058 32070 22104 32122
rect 22104 32070 22114 32122
rect 22138 32070 22168 32122
rect 22168 32070 22180 32122
rect 22180 32070 22194 32122
rect 22218 32070 22232 32122
rect 22232 32070 22244 32122
rect 22244 32070 22274 32122
rect 22298 32070 22308 32122
rect 22308 32070 22354 32122
rect 22058 32068 22114 32070
rect 22138 32068 22194 32070
rect 22218 32068 22274 32070
rect 22298 32068 22354 32070
rect 22742 31864 22798 31920
rect 22926 31864 22982 31920
rect 22058 31034 22114 31036
rect 22138 31034 22194 31036
rect 22218 31034 22274 31036
rect 22298 31034 22354 31036
rect 22058 30982 22104 31034
rect 22104 30982 22114 31034
rect 22138 30982 22168 31034
rect 22168 30982 22180 31034
rect 22180 30982 22194 31034
rect 22218 30982 22232 31034
rect 22232 30982 22244 31034
rect 22244 30982 22274 31034
rect 22298 30982 22308 31034
rect 22308 30982 22354 31034
rect 22058 30980 22114 30982
rect 22138 30980 22194 30982
rect 22218 30980 22274 30982
rect 22298 30980 22354 30982
rect 21914 30268 21916 30288
rect 21916 30268 21968 30288
rect 21968 30268 21970 30288
rect 21914 30232 21970 30268
rect 22058 29946 22114 29948
rect 22138 29946 22194 29948
rect 22218 29946 22274 29948
rect 22298 29946 22354 29948
rect 22058 29894 22104 29946
rect 22104 29894 22114 29946
rect 22138 29894 22168 29946
rect 22168 29894 22180 29946
rect 22180 29894 22194 29946
rect 22218 29894 22232 29946
rect 22232 29894 22244 29946
rect 22244 29894 22274 29946
rect 22298 29894 22308 29946
rect 22308 29894 22354 29946
rect 22058 29892 22114 29894
rect 22138 29892 22194 29894
rect 22218 29892 22274 29894
rect 22298 29892 22354 29894
rect 20442 28092 20444 28112
rect 20444 28092 20496 28112
rect 20496 28092 20498 28112
rect 20442 28056 20498 28092
rect 22006 29164 22062 29200
rect 22006 29144 22008 29164
rect 22008 29144 22060 29164
rect 22060 29144 22062 29164
rect 22282 29008 22338 29064
rect 22058 28858 22114 28860
rect 22138 28858 22194 28860
rect 22218 28858 22274 28860
rect 22298 28858 22354 28860
rect 22058 28806 22104 28858
rect 22104 28806 22114 28858
rect 22138 28806 22168 28858
rect 22168 28806 22180 28858
rect 22180 28806 22194 28858
rect 22218 28806 22232 28858
rect 22232 28806 22244 28858
rect 22244 28806 22274 28858
rect 22298 28806 22308 28858
rect 22308 28806 22354 28858
rect 22058 28804 22114 28806
rect 22138 28804 22194 28806
rect 22218 28804 22274 28806
rect 22298 28804 22354 28806
rect 22466 29144 22522 29200
rect 22058 27770 22114 27772
rect 22138 27770 22194 27772
rect 22218 27770 22274 27772
rect 22298 27770 22354 27772
rect 22058 27718 22104 27770
rect 22104 27718 22114 27770
rect 22138 27718 22168 27770
rect 22168 27718 22180 27770
rect 22180 27718 22194 27770
rect 22218 27718 22232 27770
rect 22232 27718 22244 27770
rect 22244 27718 22274 27770
rect 22298 27718 22308 27770
rect 22308 27718 22354 27770
rect 22058 27716 22114 27718
rect 22138 27716 22194 27718
rect 22218 27716 22274 27718
rect 22298 27716 22354 27718
rect 19246 26288 19302 26344
rect 20074 25880 20130 25936
rect 19338 24792 19394 24848
rect 19246 23704 19302 23760
rect 19522 18672 19578 18728
rect 20626 25372 20628 25392
rect 20628 25372 20680 25392
rect 20680 25372 20682 25392
rect 20626 25336 20682 25372
rect 21178 24928 21234 24984
rect 22058 26682 22114 26684
rect 22138 26682 22194 26684
rect 22218 26682 22274 26684
rect 22298 26682 22354 26684
rect 22058 26630 22104 26682
rect 22104 26630 22114 26682
rect 22138 26630 22168 26682
rect 22168 26630 22180 26682
rect 22180 26630 22194 26682
rect 22218 26630 22232 26682
rect 22232 26630 22244 26682
rect 22244 26630 22274 26682
rect 22298 26630 22308 26682
rect 22308 26630 22354 26682
rect 22058 26628 22114 26630
rect 22138 26628 22194 26630
rect 22218 26628 22274 26630
rect 22298 26628 22354 26630
rect 22926 29552 22982 29608
rect 23478 29164 23534 29200
rect 23478 29144 23480 29164
rect 23480 29144 23532 29164
rect 23532 29144 23534 29164
rect 22058 25594 22114 25596
rect 22138 25594 22194 25596
rect 22218 25594 22274 25596
rect 22298 25594 22354 25596
rect 22058 25542 22104 25594
rect 22104 25542 22114 25594
rect 22138 25542 22168 25594
rect 22168 25542 22180 25594
rect 22180 25542 22194 25594
rect 22218 25542 22232 25594
rect 22232 25542 22244 25594
rect 22244 25542 22274 25594
rect 22298 25542 22308 25594
rect 22308 25542 22354 25594
rect 22058 25540 22114 25542
rect 22138 25540 22194 25542
rect 22218 25540 22274 25542
rect 22298 25540 22354 25542
rect 20534 21936 20590 21992
rect 20994 21548 21050 21584
rect 20994 21528 20996 21548
rect 20996 21528 21048 21548
rect 21048 21528 21050 21548
rect 22058 24506 22114 24508
rect 22138 24506 22194 24508
rect 22218 24506 22274 24508
rect 22298 24506 22354 24508
rect 22058 24454 22104 24506
rect 22104 24454 22114 24506
rect 22138 24454 22168 24506
rect 22168 24454 22180 24506
rect 22180 24454 22194 24506
rect 22218 24454 22232 24506
rect 22232 24454 22244 24506
rect 22244 24454 22274 24506
rect 22298 24454 22308 24506
rect 22308 24454 22354 24506
rect 22058 24452 22114 24454
rect 22138 24452 22194 24454
rect 22218 24452 22274 24454
rect 22298 24452 22354 24454
rect 22282 24248 22338 24304
rect 22058 23418 22114 23420
rect 22138 23418 22194 23420
rect 22218 23418 22274 23420
rect 22298 23418 22354 23420
rect 22058 23366 22104 23418
rect 22104 23366 22114 23418
rect 22138 23366 22168 23418
rect 22168 23366 22180 23418
rect 22180 23366 22194 23418
rect 22218 23366 22232 23418
rect 22232 23366 22244 23418
rect 22244 23366 22274 23418
rect 22298 23366 22308 23418
rect 22308 23366 22354 23418
rect 22058 23364 22114 23366
rect 22138 23364 22194 23366
rect 22218 23364 22274 23366
rect 22298 23364 22354 23366
rect 21362 21392 21418 21448
rect 22058 22330 22114 22332
rect 22138 22330 22194 22332
rect 22218 22330 22274 22332
rect 22298 22330 22354 22332
rect 22058 22278 22104 22330
rect 22104 22278 22114 22330
rect 22138 22278 22168 22330
rect 22168 22278 22180 22330
rect 22180 22278 22194 22330
rect 22218 22278 22232 22330
rect 22232 22278 22244 22330
rect 22244 22278 22274 22330
rect 22298 22278 22308 22330
rect 22308 22278 22354 22330
rect 22058 22276 22114 22278
rect 22138 22276 22194 22278
rect 22218 22276 22274 22278
rect 22298 22276 22354 22278
rect 23478 28464 23534 28520
rect 24122 31728 24178 31784
rect 23386 26308 23442 26344
rect 23386 26288 23388 26308
rect 23388 26288 23440 26308
rect 23440 26288 23442 26308
rect 22834 23432 22890 23488
rect 22006 21392 22062 21448
rect 22058 21242 22114 21244
rect 22138 21242 22194 21244
rect 22218 21242 22274 21244
rect 22298 21242 22354 21244
rect 22058 21190 22104 21242
rect 22104 21190 22114 21242
rect 22138 21190 22168 21242
rect 22168 21190 22180 21242
rect 22180 21190 22194 21242
rect 22218 21190 22232 21242
rect 22232 21190 22244 21242
rect 22244 21190 22274 21242
rect 22298 21190 22308 21242
rect 22308 21190 22354 21242
rect 22058 21188 22114 21190
rect 22138 21188 22194 21190
rect 22218 21188 22274 21190
rect 22298 21188 22354 21190
rect 22098 20868 22154 20904
rect 22098 20848 22100 20868
rect 22100 20848 22152 20868
rect 22152 20848 22154 20868
rect 22058 20154 22114 20156
rect 22138 20154 22194 20156
rect 22218 20154 22274 20156
rect 22298 20154 22354 20156
rect 22058 20102 22104 20154
rect 22104 20102 22114 20154
rect 22138 20102 22168 20154
rect 22168 20102 22180 20154
rect 22180 20102 22194 20154
rect 22218 20102 22232 20154
rect 22232 20102 22244 20154
rect 22244 20102 22274 20154
rect 22298 20102 22308 20154
rect 22308 20102 22354 20154
rect 22058 20100 22114 20102
rect 22138 20100 22194 20102
rect 22218 20100 22274 20102
rect 22298 20100 22354 20102
rect 22058 19066 22114 19068
rect 22138 19066 22194 19068
rect 22218 19066 22274 19068
rect 22298 19066 22354 19068
rect 22058 19014 22104 19066
rect 22104 19014 22114 19066
rect 22138 19014 22168 19066
rect 22168 19014 22180 19066
rect 22180 19014 22194 19066
rect 22218 19014 22232 19066
rect 22232 19014 22244 19066
rect 22244 19014 22274 19066
rect 22298 19014 22308 19066
rect 22308 19014 22354 19066
rect 22058 19012 22114 19014
rect 22138 19012 22194 19014
rect 22218 19012 22274 19014
rect 22298 19012 22354 19014
rect 22058 17978 22114 17980
rect 22138 17978 22194 17980
rect 22218 17978 22274 17980
rect 22298 17978 22354 17980
rect 22058 17926 22104 17978
rect 22104 17926 22114 17978
rect 22138 17926 22168 17978
rect 22168 17926 22180 17978
rect 22180 17926 22194 17978
rect 22218 17926 22232 17978
rect 22232 17926 22244 17978
rect 22244 17926 22274 17978
rect 22298 17926 22308 17978
rect 22308 17926 22354 17978
rect 22058 17924 22114 17926
rect 22138 17924 22194 17926
rect 22218 17924 22274 17926
rect 22298 17924 22354 17926
rect 22058 16890 22114 16892
rect 22138 16890 22194 16892
rect 22218 16890 22274 16892
rect 22298 16890 22354 16892
rect 22058 16838 22104 16890
rect 22104 16838 22114 16890
rect 22138 16838 22168 16890
rect 22168 16838 22180 16890
rect 22180 16838 22194 16890
rect 22218 16838 22232 16890
rect 22232 16838 22244 16890
rect 22244 16838 22274 16890
rect 22298 16838 22308 16890
rect 22308 16838 22354 16890
rect 22058 16836 22114 16838
rect 22138 16836 22194 16838
rect 22218 16836 22274 16838
rect 22298 16836 22354 16838
rect 23294 21528 23350 21584
rect 24950 36216 25006 36272
rect 24766 34040 24822 34096
rect 24582 32272 24638 32328
rect 26278 39194 26334 39196
rect 26358 39194 26414 39196
rect 26438 39194 26494 39196
rect 26518 39194 26574 39196
rect 26278 39142 26324 39194
rect 26324 39142 26334 39194
rect 26358 39142 26388 39194
rect 26388 39142 26400 39194
rect 26400 39142 26414 39194
rect 26438 39142 26452 39194
rect 26452 39142 26464 39194
rect 26464 39142 26494 39194
rect 26518 39142 26528 39194
rect 26528 39142 26574 39194
rect 26278 39140 26334 39142
rect 26358 39140 26414 39142
rect 26438 39140 26494 39142
rect 26518 39140 26574 39142
rect 27618 38936 27674 38992
rect 26422 38256 26478 38312
rect 26278 38106 26334 38108
rect 26358 38106 26414 38108
rect 26438 38106 26494 38108
rect 26518 38106 26574 38108
rect 26278 38054 26324 38106
rect 26324 38054 26334 38106
rect 26358 38054 26388 38106
rect 26388 38054 26400 38106
rect 26400 38054 26414 38106
rect 26438 38054 26452 38106
rect 26452 38054 26464 38106
rect 26464 38054 26494 38106
rect 26518 38054 26528 38106
rect 26528 38054 26574 38106
rect 26278 38052 26334 38054
rect 26358 38052 26414 38054
rect 26438 38052 26494 38054
rect 26518 38052 26574 38054
rect 25318 37884 25320 37904
rect 25320 37884 25372 37904
rect 25372 37884 25374 37904
rect 25318 37848 25374 37884
rect 25686 37304 25742 37360
rect 25318 36080 25374 36136
rect 25134 32408 25190 32464
rect 25134 31864 25190 31920
rect 25502 32816 25558 32872
rect 24214 28056 24270 28112
rect 27158 37712 27214 37768
rect 26278 37018 26334 37020
rect 26358 37018 26414 37020
rect 26438 37018 26494 37020
rect 26518 37018 26574 37020
rect 26278 36966 26324 37018
rect 26324 36966 26334 37018
rect 26358 36966 26388 37018
rect 26388 36966 26400 37018
rect 26400 36966 26414 37018
rect 26438 36966 26452 37018
rect 26452 36966 26464 37018
rect 26464 36966 26494 37018
rect 26518 36966 26528 37018
rect 26528 36966 26574 37018
rect 26278 36964 26334 36966
rect 26358 36964 26414 36966
rect 26438 36964 26494 36966
rect 26518 36964 26574 36966
rect 25778 31864 25834 31920
rect 26278 35930 26334 35932
rect 26358 35930 26414 35932
rect 26438 35930 26494 35932
rect 26518 35930 26574 35932
rect 26278 35878 26324 35930
rect 26324 35878 26334 35930
rect 26358 35878 26388 35930
rect 26388 35878 26400 35930
rect 26400 35878 26414 35930
rect 26438 35878 26452 35930
rect 26452 35878 26464 35930
rect 26464 35878 26494 35930
rect 26518 35878 26528 35930
rect 26528 35878 26574 35930
rect 26278 35876 26334 35878
rect 26358 35876 26414 35878
rect 26438 35876 26494 35878
rect 26518 35876 26574 35878
rect 26278 34842 26334 34844
rect 26358 34842 26414 34844
rect 26438 34842 26494 34844
rect 26518 34842 26574 34844
rect 26278 34790 26324 34842
rect 26324 34790 26334 34842
rect 26358 34790 26388 34842
rect 26388 34790 26400 34842
rect 26400 34790 26414 34842
rect 26438 34790 26452 34842
rect 26452 34790 26464 34842
rect 26464 34790 26494 34842
rect 26518 34790 26528 34842
rect 26528 34790 26574 34842
rect 26278 34788 26334 34790
rect 26358 34788 26414 34790
rect 26438 34788 26494 34790
rect 26518 34788 26574 34790
rect 26278 33754 26334 33756
rect 26358 33754 26414 33756
rect 26438 33754 26494 33756
rect 26518 33754 26574 33756
rect 26278 33702 26324 33754
rect 26324 33702 26334 33754
rect 26358 33702 26388 33754
rect 26388 33702 26400 33754
rect 26400 33702 26414 33754
rect 26438 33702 26452 33754
rect 26452 33702 26464 33754
rect 26464 33702 26494 33754
rect 26518 33702 26528 33754
rect 26528 33702 26574 33754
rect 26278 33700 26334 33702
rect 26358 33700 26414 33702
rect 26438 33700 26494 33702
rect 26518 33700 26574 33702
rect 26698 33516 26754 33552
rect 26698 33496 26700 33516
rect 26700 33496 26752 33516
rect 26752 33496 26754 33516
rect 26278 32666 26334 32668
rect 26358 32666 26414 32668
rect 26438 32666 26494 32668
rect 26518 32666 26574 32668
rect 26278 32614 26324 32666
rect 26324 32614 26334 32666
rect 26358 32614 26388 32666
rect 26388 32614 26400 32666
rect 26400 32614 26414 32666
rect 26438 32614 26452 32666
rect 26452 32614 26464 32666
rect 26464 32614 26494 32666
rect 26518 32614 26528 32666
rect 26528 32614 26574 32666
rect 26278 32612 26334 32614
rect 26358 32612 26414 32614
rect 26438 32612 26494 32614
rect 26518 32612 26574 32614
rect 26278 31578 26334 31580
rect 26358 31578 26414 31580
rect 26438 31578 26494 31580
rect 26518 31578 26574 31580
rect 26278 31526 26324 31578
rect 26324 31526 26334 31578
rect 26358 31526 26388 31578
rect 26388 31526 26400 31578
rect 26400 31526 26414 31578
rect 26438 31526 26452 31578
rect 26452 31526 26464 31578
rect 26464 31526 26494 31578
rect 26518 31526 26528 31578
rect 26528 31526 26574 31578
rect 26278 31524 26334 31526
rect 26358 31524 26414 31526
rect 26438 31524 26494 31526
rect 26518 31524 26574 31526
rect 26278 30490 26334 30492
rect 26358 30490 26414 30492
rect 26438 30490 26494 30492
rect 26518 30490 26574 30492
rect 26278 30438 26324 30490
rect 26324 30438 26334 30490
rect 26358 30438 26388 30490
rect 26388 30438 26400 30490
rect 26400 30438 26414 30490
rect 26438 30438 26452 30490
rect 26452 30438 26464 30490
rect 26464 30438 26494 30490
rect 26518 30438 26528 30490
rect 26528 30438 26574 30490
rect 26278 30436 26334 30438
rect 26358 30436 26414 30438
rect 26438 30436 26494 30438
rect 26518 30436 26574 30438
rect 25042 29416 25098 29472
rect 24398 24928 24454 24984
rect 22058 15802 22114 15804
rect 22138 15802 22194 15804
rect 22218 15802 22274 15804
rect 22298 15802 22354 15804
rect 22058 15750 22104 15802
rect 22104 15750 22114 15802
rect 22138 15750 22168 15802
rect 22168 15750 22180 15802
rect 22180 15750 22194 15802
rect 22218 15750 22232 15802
rect 22232 15750 22244 15802
rect 22244 15750 22274 15802
rect 22298 15750 22308 15802
rect 22308 15750 22354 15802
rect 22058 15748 22114 15750
rect 22138 15748 22194 15750
rect 22218 15748 22274 15750
rect 22298 15748 22354 15750
rect 24214 20848 24270 20904
rect 24950 25880 25006 25936
rect 24582 24248 24638 24304
rect 25134 21936 25190 21992
rect 24582 18536 24638 18592
rect 23570 15408 23626 15464
rect 22006 15020 22062 15056
rect 26278 29402 26334 29404
rect 26358 29402 26414 29404
rect 26438 29402 26494 29404
rect 26518 29402 26574 29404
rect 26278 29350 26324 29402
rect 26324 29350 26334 29402
rect 26358 29350 26388 29402
rect 26388 29350 26400 29402
rect 26400 29350 26414 29402
rect 26438 29350 26452 29402
rect 26452 29350 26464 29402
rect 26464 29350 26494 29402
rect 26518 29350 26528 29402
rect 26528 29350 26574 29402
rect 26278 29348 26334 29350
rect 26358 29348 26414 29350
rect 26438 29348 26494 29350
rect 26518 29348 26574 29350
rect 27158 36896 27214 36952
rect 27158 36080 27214 36136
rect 27158 35672 27214 35728
rect 28078 37576 28134 37632
rect 27618 35128 27674 35184
rect 27618 34448 27674 34504
rect 27618 33224 27674 33280
rect 26278 28314 26334 28316
rect 26358 28314 26414 28316
rect 26438 28314 26494 28316
rect 26518 28314 26574 28316
rect 26278 28262 26324 28314
rect 26324 28262 26334 28314
rect 26358 28262 26388 28314
rect 26388 28262 26400 28314
rect 26400 28262 26414 28314
rect 26438 28262 26452 28314
rect 26452 28262 26464 28314
rect 26464 28262 26494 28314
rect 26518 28262 26528 28314
rect 26528 28262 26574 28314
rect 26278 28260 26334 28262
rect 26358 28260 26414 28262
rect 26438 28260 26494 28262
rect 26518 28260 26574 28262
rect 26278 27226 26334 27228
rect 26358 27226 26414 27228
rect 26438 27226 26494 27228
rect 26518 27226 26574 27228
rect 26278 27174 26324 27226
rect 26324 27174 26334 27226
rect 26358 27174 26388 27226
rect 26388 27174 26400 27226
rect 26400 27174 26414 27226
rect 26438 27174 26452 27226
rect 26452 27174 26464 27226
rect 26464 27174 26494 27226
rect 26518 27174 26528 27226
rect 26528 27174 26574 27226
rect 26278 27172 26334 27174
rect 26358 27172 26414 27174
rect 26438 27172 26494 27174
rect 26518 27172 26574 27174
rect 26330 26852 26386 26888
rect 26330 26832 26332 26852
rect 26332 26832 26384 26852
rect 26384 26832 26386 26852
rect 25962 25880 26018 25936
rect 25778 25744 25834 25800
rect 25686 25608 25742 25664
rect 26278 26138 26334 26140
rect 26358 26138 26414 26140
rect 26438 26138 26494 26140
rect 26518 26138 26574 26140
rect 26278 26086 26324 26138
rect 26324 26086 26334 26138
rect 26358 26086 26388 26138
rect 26388 26086 26400 26138
rect 26400 26086 26414 26138
rect 26438 26086 26452 26138
rect 26452 26086 26464 26138
rect 26464 26086 26494 26138
rect 26518 26086 26528 26138
rect 26528 26086 26574 26138
rect 26278 26084 26334 26086
rect 26358 26084 26414 26086
rect 26438 26084 26494 26086
rect 26518 26084 26574 26086
rect 26514 25356 26570 25392
rect 26514 25336 26516 25356
rect 26516 25336 26568 25356
rect 26568 25336 26570 25356
rect 26882 29008 26938 29064
rect 26422 25200 26478 25256
rect 26278 25050 26334 25052
rect 26358 25050 26414 25052
rect 26438 25050 26494 25052
rect 26518 25050 26574 25052
rect 26278 24998 26324 25050
rect 26324 24998 26334 25050
rect 26358 24998 26388 25050
rect 26388 24998 26400 25050
rect 26400 24998 26414 25050
rect 26438 24998 26452 25050
rect 26452 24998 26464 25050
rect 26464 24998 26494 25050
rect 26518 24998 26528 25050
rect 26528 24998 26574 25050
rect 26278 24996 26334 24998
rect 26358 24996 26414 24998
rect 26438 24996 26494 24998
rect 26518 24996 26574 24998
rect 27342 29824 27398 29880
rect 27618 31320 27674 31376
rect 28262 35944 28318 36000
rect 28170 35672 28226 35728
rect 27894 31628 27896 31648
rect 27896 31628 27948 31648
rect 27948 31628 27950 31648
rect 27894 31592 27950 31628
rect 27802 29552 27858 29608
rect 27710 29144 27766 29200
rect 27802 28872 27858 28928
rect 27618 28464 27674 28520
rect 30499 39738 30555 39740
rect 30579 39738 30635 39740
rect 30659 39738 30715 39740
rect 30739 39738 30795 39740
rect 30499 39686 30545 39738
rect 30545 39686 30555 39738
rect 30579 39686 30609 39738
rect 30609 39686 30621 39738
rect 30621 39686 30635 39738
rect 30659 39686 30673 39738
rect 30673 39686 30685 39738
rect 30685 39686 30715 39738
rect 30739 39686 30749 39738
rect 30749 39686 30795 39738
rect 30499 39684 30555 39686
rect 30579 39684 30635 39686
rect 30659 39684 30715 39686
rect 30739 39684 30795 39686
rect 29090 37440 29146 37496
rect 29182 36488 29238 36544
rect 29090 36352 29146 36408
rect 28630 35672 28686 35728
rect 28538 34040 28594 34096
rect 28538 33088 28594 33144
rect 28446 32680 28502 32736
rect 28814 35944 28870 36000
rect 28814 33224 28870 33280
rect 28814 33108 28870 33144
rect 28814 33088 28816 33108
rect 28816 33088 28868 33108
rect 28868 33088 28870 33108
rect 29182 36236 29238 36272
rect 29182 36216 29184 36236
rect 29184 36216 29236 36236
rect 29236 36216 29238 36236
rect 29182 35828 29238 35864
rect 29182 35808 29184 35828
rect 29184 35808 29236 35828
rect 29236 35808 29238 35828
rect 28906 31864 28962 31920
rect 29458 36488 29514 36544
rect 29366 34992 29422 35048
rect 29182 32852 29184 32872
rect 29184 32852 29236 32872
rect 29236 32852 29238 32872
rect 29182 32816 29238 32852
rect 28814 31592 28870 31648
rect 28078 27920 28134 27976
rect 26882 25336 26938 25392
rect 26278 23962 26334 23964
rect 26358 23962 26414 23964
rect 26438 23962 26494 23964
rect 26518 23962 26574 23964
rect 26278 23910 26324 23962
rect 26324 23910 26334 23962
rect 26358 23910 26388 23962
rect 26388 23910 26400 23962
rect 26400 23910 26414 23962
rect 26438 23910 26452 23962
rect 26452 23910 26464 23962
rect 26464 23910 26494 23962
rect 26518 23910 26528 23962
rect 26528 23910 26574 23962
rect 26278 23908 26334 23910
rect 26358 23908 26414 23910
rect 26438 23908 26494 23910
rect 26518 23908 26574 23910
rect 26278 22874 26334 22876
rect 26358 22874 26414 22876
rect 26438 22874 26494 22876
rect 26518 22874 26574 22876
rect 26278 22822 26324 22874
rect 26324 22822 26334 22874
rect 26358 22822 26388 22874
rect 26388 22822 26400 22874
rect 26400 22822 26414 22874
rect 26438 22822 26452 22874
rect 26452 22822 26464 22874
rect 26464 22822 26494 22874
rect 26518 22822 26528 22874
rect 26528 22822 26574 22874
rect 26278 22820 26334 22822
rect 26358 22820 26414 22822
rect 26438 22820 26494 22822
rect 26518 22820 26574 22822
rect 25686 20712 25742 20768
rect 26278 21786 26334 21788
rect 26358 21786 26414 21788
rect 26438 21786 26494 21788
rect 26518 21786 26574 21788
rect 26278 21734 26324 21786
rect 26324 21734 26334 21786
rect 26358 21734 26388 21786
rect 26388 21734 26400 21786
rect 26400 21734 26414 21786
rect 26438 21734 26452 21786
rect 26452 21734 26464 21786
rect 26464 21734 26494 21786
rect 26518 21734 26528 21786
rect 26528 21734 26574 21786
rect 26278 21732 26334 21734
rect 26358 21732 26414 21734
rect 26438 21732 26494 21734
rect 26518 21732 26574 21734
rect 26278 20698 26334 20700
rect 26358 20698 26414 20700
rect 26438 20698 26494 20700
rect 26518 20698 26574 20700
rect 26278 20646 26324 20698
rect 26324 20646 26334 20698
rect 26358 20646 26388 20698
rect 26388 20646 26400 20698
rect 26400 20646 26414 20698
rect 26438 20646 26452 20698
rect 26452 20646 26464 20698
rect 26464 20646 26494 20698
rect 26518 20646 26528 20698
rect 26528 20646 26574 20698
rect 26278 20644 26334 20646
rect 26358 20644 26414 20646
rect 26438 20644 26494 20646
rect 26518 20644 26574 20646
rect 22006 15000 22008 15020
rect 22008 15000 22060 15020
rect 22060 15000 22062 15020
rect 17837 6554 17893 6556
rect 17917 6554 17973 6556
rect 17997 6554 18053 6556
rect 18077 6554 18133 6556
rect 17837 6502 17883 6554
rect 17883 6502 17893 6554
rect 17917 6502 17947 6554
rect 17947 6502 17959 6554
rect 17959 6502 17973 6554
rect 17997 6502 18011 6554
rect 18011 6502 18023 6554
rect 18023 6502 18053 6554
rect 18077 6502 18087 6554
rect 18087 6502 18133 6554
rect 17837 6500 17893 6502
rect 17917 6500 17973 6502
rect 17997 6500 18053 6502
rect 18077 6500 18133 6502
rect 17837 5466 17893 5468
rect 17917 5466 17973 5468
rect 17997 5466 18053 5468
rect 18077 5466 18133 5468
rect 17837 5414 17883 5466
rect 17883 5414 17893 5466
rect 17917 5414 17947 5466
rect 17947 5414 17959 5466
rect 17959 5414 17973 5466
rect 17997 5414 18011 5466
rect 18011 5414 18023 5466
rect 18023 5414 18053 5466
rect 18077 5414 18087 5466
rect 18087 5414 18133 5466
rect 17837 5412 17893 5414
rect 17917 5412 17973 5414
rect 17997 5412 18053 5414
rect 18077 5412 18133 5414
rect 17837 4378 17893 4380
rect 17917 4378 17973 4380
rect 17997 4378 18053 4380
rect 18077 4378 18133 4380
rect 17837 4326 17883 4378
rect 17883 4326 17893 4378
rect 17917 4326 17947 4378
rect 17947 4326 17959 4378
rect 17959 4326 17973 4378
rect 17997 4326 18011 4378
rect 18011 4326 18023 4378
rect 18023 4326 18053 4378
rect 18077 4326 18087 4378
rect 18087 4326 18133 4378
rect 17837 4324 17893 4326
rect 17917 4324 17973 4326
rect 17997 4324 18053 4326
rect 18077 4324 18133 4326
rect 13617 2746 13673 2748
rect 13697 2746 13753 2748
rect 13777 2746 13833 2748
rect 13857 2746 13913 2748
rect 13617 2694 13663 2746
rect 13663 2694 13673 2746
rect 13697 2694 13727 2746
rect 13727 2694 13739 2746
rect 13739 2694 13753 2746
rect 13777 2694 13791 2746
rect 13791 2694 13803 2746
rect 13803 2694 13833 2746
rect 13857 2694 13867 2746
rect 13867 2694 13913 2746
rect 13617 2692 13673 2694
rect 13697 2692 13753 2694
rect 13777 2692 13833 2694
rect 13857 2692 13913 2694
rect 17837 3290 17893 3292
rect 17917 3290 17973 3292
rect 17997 3290 18053 3292
rect 18077 3290 18133 3292
rect 17837 3238 17883 3290
rect 17883 3238 17893 3290
rect 17917 3238 17947 3290
rect 17947 3238 17959 3290
rect 17959 3238 17973 3290
rect 17997 3238 18011 3290
rect 18011 3238 18023 3290
rect 18023 3238 18053 3290
rect 18077 3238 18087 3290
rect 18087 3238 18133 3290
rect 17837 3236 17893 3238
rect 17917 3236 17973 3238
rect 17997 3236 18053 3238
rect 18077 3236 18133 3238
rect 17837 2202 17893 2204
rect 17917 2202 17973 2204
rect 17997 2202 18053 2204
rect 18077 2202 18133 2204
rect 17837 2150 17883 2202
rect 17883 2150 17893 2202
rect 17917 2150 17947 2202
rect 17947 2150 17959 2202
rect 17959 2150 17973 2202
rect 17997 2150 18011 2202
rect 18011 2150 18023 2202
rect 18023 2150 18053 2202
rect 18077 2150 18087 2202
rect 18087 2150 18133 2202
rect 17837 2148 17893 2150
rect 17917 2148 17973 2150
rect 17997 2148 18053 2150
rect 18077 2148 18133 2150
rect 22058 14714 22114 14716
rect 22138 14714 22194 14716
rect 22218 14714 22274 14716
rect 22298 14714 22354 14716
rect 22058 14662 22104 14714
rect 22104 14662 22114 14714
rect 22138 14662 22168 14714
rect 22168 14662 22180 14714
rect 22180 14662 22194 14714
rect 22218 14662 22232 14714
rect 22232 14662 22244 14714
rect 22244 14662 22274 14714
rect 22298 14662 22308 14714
rect 22308 14662 22354 14714
rect 22058 14660 22114 14662
rect 22138 14660 22194 14662
rect 22218 14660 22274 14662
rect 22298 14660 22354 14662
rect 25594 15272 25650 15328
rect 25594 15020 25650 15056
rect 25870 16496 25926 16552
rect 25594 15000 25596 15020
rect 25596 15000 25648 15020
rect 25648 15000 25650 15020
rect 26278 19610 26334 19612
rect 26358 19610 26414 19612
rect 26438 19610 26494 19612
rect 26518 19610 26574 19612
rect 26278 19558 26324 19610
rect 26324 19558 26334 19610
rect 26358 19558 26388 19610
rect 26388 19558 26400 19610
rect 26400 19558 26414 19610
rect 26438 19558 26452 19610
rect 26452 19558 26464 19610
rect 26464 19558 26494 19610
rect 26518 19558 26528 19610
rect 26528 19558 26574 19610
rect 26278 19556 26334 19558
rect 26358 19556 26414 19558
rect 26438 19556 26494 19558
rect 26518 19556 26574 19558
rect 26278 18522 26334 18524
rect 26358 18522 26414 18524
rect 26438 18522 26494 18524
rect 26518 18522 26574 18524
rect 26278 18470 26324 18522
rect 26324 18470 26334 18522
rect 26358 18470 26388 18522
rect 26388 18470 26400 18522
rect 26400 18470 26414 18522
rect 26438 18470 26452 18522
rect 26452 18470 26464 18522
rect 26464 18470 26494 18522
rect 26518 18470 26528 18522
rect 26528 18470 26574 18522
rect 26278 18468 26334 18470
rect 26358 18468 26414 18470
rect 26438 18468 26494 18470
rect 26518 18468 26574 18470
rect 26278 17434 26334 17436
rect 26358 17434 26414 17436
rect 26438 17434 26494 17436
rect 26518 17434 26574 17436
rect 26278 17382 26324 17434
rect 26324 17382 26334 17434
rect 26358 17382 26388 17434
rect 26388 17382 26400 17434
rect 26400 17382 26414 17434
rect 26438 17382 26452 17434
rect 26452 17382 26464 17434
rect 26464 17382 26494 17434
rect 26518 17382 26528 17434
rect 26528 17382 26574 17434
rect 26278 17380 26334 17382
rect 26358 17380 26414 17382
rect 26438 17380 26494 17382
rect 26518 17380 26574 17382
rect 26278 16346 26334 16348
rect 26358 16346 26414 16348
rect 26438 16346 26494 16348
rect 26518 16346 26574 16348
rect 26278 16294 26324 16346
rect 26324 16294 26334 16346
rect 26358 16294 26388 16346
rect 26388 16294 26400 16346
rect 26400 16294 26414 16346
rect 26438 16294 26452 16346
rect 26452 16294 26464 16346
rect 26464 16294 26494 16346
rect 26518 16294 26528 16346
rect 26528 16294 26574 16346
rect 26278 16292 26334 16294
rect 26358 16292 26414 16294
rect 26438 16292 26494 16294
rect 26518 16292 26574 16294
rect 26422 15428 26478 15464
rect 26422 15408 26424 15428
rect 26424 15408 26476 15428
rect 26476 15408 26478 15428
rect 26278 15258 26334 15260
rect 26358 15258 26414 15260
rect 26438 15258 26494 15260
rect 26518 15258 26574 15260
rect 26278 15206 26324 15258
rect 26324 15206 26334 15258
rect 26358 15206 26388 15258
rect 26388 15206 26400 15258
rect 26400 15206 26414 15258
rect 26438 15206 26452 15258
rect 26452 15206 26464 15258
rect 26464 15206 26494 15258
rect 26518 15206 26528 15258
rect 26528 15206 26574 15258
rect 26278 15204 26334 15206
rect 26358 15204 26414 15206
rect 26438 15204 26494 15206
rect 26518 15204 26574 15206
rect 27434 25744 27490 25800
rect 27434 25608 27490 25664
rect 27342 25472 27398 25528
rect 27526 24792 27582 24848
rect 27618 23044 27674 23080
rect 27618 23024 27620 23044
rect 27620 23024 27672 23044
rect 27672 23024 27674 23044
rect 29458 32408 29514 32464
rect 29090 30640 29146 30696
rect 28998 30096 29054 30152
rect 29458 31048 29514 31104
rect 29274 29416 29330 29472
rect 28906 28328 28962 28384
rect 28814 27648 28870 27704
rect 29090 28056 29146 28112
rect 28998 27920 29054 27976
rect 28170 25900 28226 25936
rect 28170 25880 28172 25900
rect 28172 25880 28224 25900
rect 28224 25880 28226 25900
rect 27710 19660 27712 19680
rect 27712 19660 27764 19680
rect 27764 19660 27766 19680
rect 27710 19624 27766 19660
rect 28998 25372 29001 25392
rect 29001 25372 29053 25392
rect 29053 25372 29054 25392
rect 28998 25336 29054 25372
rect 29734 37304 29790 37360
rect 30010 37884 30012 37904
rect 30012 37884 30064 37904
rect 30064 37884 30066 37904
rect 30010 37848 30066 37884
rect 29918 37712 29974 37768
rect 30010 37304 30066 37360
rect 29918 36352 29974 36408
rect 29918 35808 29974 35864
rect 30499 38650 30555 38652
rect 30579 38650 30635 38652
rect 30659 38650 30715 38652
rect 30739 38650 30795 38652
rect 30499 38598 30545 38650
rect 30545 38598 30555 38650
rect 30579 38598 30609 38650
rect 30609 38598 30621 38650
rect 30621 38598 30635 38650
rect 30659 38598 30673 38650
rect 30673 38598 30685 38650
rect 30685 38598 30715 38650
rect 30739 38598 30749 38650
rect 30749 38598 30795 38650
rect 30499 38596 30555 38598
rect 30579 38596 30635 38598
rect 30659 38596 30715 38598
rect 30739 38596 30795 38598
rect 30499 37562 30555 37564
rect 30579 37562 30635 37564
rect 30659 37562 30715 37564
rect 30739 37562 30795 37564
rect 30499 37510 30545 37562
rect 30545 37510 30555 37562
rect 30579 37510 30609 37562
rect 30609 37510 30621 37562
rect 30621 37510 30635 37562
rect 30659 37510 30673 37562
rect 30673 37510 30685 37562
rect 30685 37510 30715 37562
rect 30739 37510 30749 37562
rect 30749 37510 30795 37562
rect 30499 37508 30555 37510
rect 30579 37508 30635 37510
rect 30659 37508 30715 37510
rect 30739 37508 30795 37510
rect 31022 37168 31078 37224
rect 30930 37068 30932 37088
rect 30932 37068 30984 37088
rect 30984 37068 30986 37088
rect 30930 37032 30986 37068
rect 30499 36474 30555 36476
rect 30579 36474 30635 36476
rect 30659 36474 30715 36476
rect 30739 36474 30795 36476
rect 30499 36422 30545 36474
rect 30545 36422 30555 36474
rect 30579 36422 30609 36474
rect 30609 36422 30621 36474
rect 30621 36422 30635 36474
rect 30659 36422 30673 36474
rect 30673 36422 30685 36474
rect 30685 36422 30715 36474
rect 30739 36422 30749 36474
rect 30749 36422 30795 36474
rect 30499 36420 30555 36422
rect 30579 36420 30635 36422
rect 30659 36420 30715 36422
rect 30739 36420 30795 36422
rect 32218 39480 32274 39536
rect 31298 37168 31354 37224
rect 31114 36352 31170 36408
rect 30930 36080 30986 36136
rect 30930 35436 30932 35456
rect 30932 35436 30984 35456
rect 30984 35436 30986 35456
rect 30930 35400 30986 35436
rect 30499 35386 30555 35388
rect 30579 35386 30635 35388
rect 30659 35386 30715 35388
rect 30739 35386 30795 35388
rect 30499 35334 30545 35386
rect 30545 35334 30555 35386
rect 30579 35334 30609 35386
rect 30609 35334 30621 35386
rect 30621 35334 30635 35386
rect 30659 35334 30673 35386
rect 30673 35334 30685 35386
rect 30685 35334 30715 35386
rect 30739 35334 30749 35386
rect 30749 35334 30795 35386
rect 30499 35332 30555 35334
rect 30579 35332 30635 35334
rect 30659 35332 30715 35334
rect 30739 35332 30795 35334
rect 30194 34448 30250 34504
rect 29734 31456 29790 31512
rect 29642 29588 29644 29608
rect 29644 29588 29696 29608
rect 29696 29588 29698 29608
rect 29642 29552 29698 29588
rect 30499 34298 30555 34300
rect 30579 34298 30635 34300
rect 30659 34298 30715 34300
rect 30739 34298 30795 34300
rect 30499 34246 30545 34298
rect 30545 34246 30555 34298
rect 30579 34246 30609 34298
rect 30609 34246 30621 34298
rect 30621 34246 30635 34298
rect 30659 34246 30673 34298
rect 30673 34246 30685 34298
rect 30685 34246 30715 34298
rect 30739 34246 30749 34298
rect 30749 34246 30795 34298
rect 30499 34244 30555 34246
rect 30579 34244 30635 34246
rect 30659 34244 30715 34246
rect 30739 34244 30795 34246
rect 30499 33210 30555 33212
rect 30579 33210 30635 33212
rect 30659 33210 30715 33212
rect 30739 33210 30795 33212
rect 30499 33158 30545 33210
rect 30545 33158 30555 33210
rect 30579 33158 30609 33210
rect 30609 33158 30621 33210
rect 30621 33158 30635 33210
rect 30659 33158 30673 33210
rect 30673 33158 30685 33210
rect 30685 33158 30715 33210
rect 30739 33158 30749 33210
rect 30749 33158 30795 33210
rect 30499 33156 30555 33158
rect 30579 33156 30635 33158
rect 30659 33156 30715 33158
rect 30739 33156 30795 33158
rect 30499 32122 30555 32124
rect 30579 32122 30635 32124
rect 30659 32122 30715 32124
rect 30739 32122 30795 32124
rect 30499 32070 30545 32122
rect 30545 32070 30555 32122
rect 30579 32070 30609 32122
rect 30609 32070 30621 32122
rect 30621 32070 30635 32122
rect 30659 32070 30673 32122
rect 30673 32070 30685 32122
rect 30685 32070 30715 32122
rect 30739 32070 30749 32122
rect 30749 32070 30795 32122
rect 30499 32068 30555 32070
rect 30579 32068 30635 32070
rect 30659 32068 30715 32070
rect 30739 32068 30795 32070
rect 30930 31748 30986 31784
rect 31298 35808 31354 35864
rect 31298 32544 31354 32600
rect 32218 37848 32274 37904
rect 32126 37712 32182 37768
rect 31942 37440 31998 37496
rect 32034 36760 32090 36816
rect 31758 35692 31814 35728
rect 31758 35672 31760 35692
rect 31760 35672 31812 35692
rect 31812 35672 31814 35692
rect 31758 35436 31760 35456
rect 31760 35436 31812 35456
rect 31812 35436 31814 35456
rect 31758 35400 31814 35436
rect 31666 33632 31722 33688
rect 32310 36896 32366 36952
rect 32218 36080 32274 36136
rect 32034 34060 32090 34096
rect 32034 34040 32036 34060
rect 32036 34040 32088 34060
rect 32088 34040 32090 34060
rect 31850 33496 31906 33552
rect 30930 31728 30932 31748
rect 30932 31728 30984 31748
rect 30984 31728 30986 31748
rect 30499 31034 30555 31036
rect 30579 31034 30635 31036
rect 30659 31034 30715 31036
rect 30739 31034 30795 31036
rect 30499 30982 30545 31034
rect 30545 30982 30555 31034
rect 30579 30982 30609 31034
rect 30609 30982 30621 31034
rect 30621 30982 30635 31034
rect 30659 30982 30673 31034
rect 30673 30982 30685 31034
rect 30685 30982 30715 31034
rect 30739 30982 30749 31034
rect 30749 30982 30795 31034
rect 30499 30980 30555 30982
rect 30579 30980 30635 30982
rect 30659 30980 30715 30982
rect 30739 30980 30795 30982
rect 31022 30660 31078 30696
rect 31022 30640 31024 30660
rect 31024 30640 31076 30660
rect 31076 30640 31078 30660
rect 30499 29946 30555 29948
rect 30579 29946 30635 29948
rect 30659 29946 30715 29948
rect 30739 29946 30795 29948
rect 30499 29894 30545 29946
rect 30545 29894 30555 29946
rect 30579 29894 30609 29946
rect 30609 29894 30621 29946
rect 30621 29894 30635 29946
rect 30659 29894 30673 29946
rect 30673 29894 30685 29946
rect 30685 29894 30715 29946
rect 30739 29894 30749 29946
rect 30749 29894 30795 29946
rect 30499 29892 30555 29894
rect 30579 29892 30635 29894
rect 30659 29892 30715 29894
rect 30739 29892 30795 29894
rect 30838 29552 30894 29608
rect 32218 31456 32274 31512
rect 33046 40840 33102 40896
rect 32494 36624 32550 36680
rect 32494 35128 32550 35184
rect 34719 39194 34775 39196
rect 34799 39194 34855 39196
rect 34879 39194 34935 39196
rect 34959 39194 35015 39196
rect 34719 39142 34765 39194
rect 34765 39142 34775 39194
rect 34799 39142 34829 39194
rect 34829 39142 34841 39194
rect 34841 39142 34855 39194
rect 34879 39142 34893 39194
rect 34893 39142 34905 39194
rect 34905 39142 34935 39194
rect 34959 39142 34969 39194
rect 34969 39142 35015 39194
rect 34719 39140 34775 39142
rect 34799 39140 34855 39142
rect 34879 39140 34935 39142
rect 34959 39140 35015 39142
rect 34334 38800 34390 38856
rect 34719 38106 34775 38108
rect 34799 38106 34855 38108
rect 34879 38106 34935 38108
rect 34959 38106 35015 38108
rect 34719 38054 34765 38106
rect 34765 38054 34775 38106
rect 34799 38054 34829 38106
rect 34829 38054 34841 38106
rect 34841 38054 34855 38106
rect 34879 38054 34893 38106
rect 34893 38054 34905 38106
rect 34905 38054 34935 38106
rect 34959 38054 34969 38106
rect 34969 38054 35015 38106
rect 34719 38052 34775 38054
rect 34799 38052 34855 38054
rect 34879 38052 34935 38054
rect 34959 38052 35015 38054
rect 34334 37884 34336 37904
rect 34336 37884 34388 37904
rect 34388 37884 34390 37904
rect 34334 37848 34390 37884
rect 34719 37018 34775 37020
rect 34799 37018 34855 37020
rect 34879 37018 34935 37020
rect 34959 37018 35015 37020
rect 34719 36966 34765 37018
rect 34765 36966 34775 37018
rect 34799 36966 34829 37018
rect 34829 36966 34841 37018
rect 34841 36966 34855 37018
rect 34879 36966 34893 37018
rect 34893 36966 34905 37018
rect 34905 36966 34935 37018
rect 34959 36966 34969 37018
rect 34969 36966 35015 37018
rect 34719 36964 34775 36966
rect 34799 36964 34855 36966
rect 34879 36964 34935 36966
rect 34959 36964 35015 36966
rect 34334 36760 34390 36816
rect 34719 35930 34775 35932
rect 34799 35930 34855 35932
rect 34879 35930 34935 35932
rect 34959 35930 35015 35932
rect 34719 35878 34765 35930
rect 34765 35878 34775 35930
rect 34799 35878 34829 35930
rect 34829 35878 34841 35930
rect 34841 35878 34855 35930
rect 34879 35878 34893 35930
rect 34893 35878 34905 35930
rect 34905 35878 34935 35930
rect 34959 35878 34969 35930
rect 34969 35878 35015 35930
rect 34719 35876 34775 35878
rect 34799 35876 34855 35878
rect 34879 35876 34935 35878
rect 34959 35876 35015 35878
rect 32770 35436 32772 35456
rect 32772 35436 32824 35456
rect 32824 35436 32826 35456
rect 32770 35400 32826 35436
rect 30930 29144 30986 29200
rect 29642 28192 29698 28248
rect 29642 27648 29698 27704
rect 28814 23024 28870 23080
rect 28998 22752 29054 22808
rect 28722 22208 28778 22264
rect 28998 21836 29000 21856
rect 29000 21836 29052 21856
rect 29052 21836 29054 21856
rect 28998 21800 29054 21836
rect 28262 18708 28264 18728
rect 28264 18708 28316 18728
rect 28316 18708 28318 18728
rect 28262 18672 28318 18708
rect 30499 28858 30555 28860
rect 30579 28858 30635 28860
rect 30659 28858 30715 28860
rect 30739 28858 30795 28860
rect 30499 28806 30545 28858
rect 30545 28806 30555 28858
rect 30579 28806 30609 28858
rect 30609 28806 30621 28858
rect 30621 28806 30635 28858
rect 30659 28806 30673 28858
rect 30673 28806 30685 28858
rect 30685 28806 30715 28858
rect 30739 28806 30749 28858
rect 30749 28806 30795 28858
rect 30499 28804 30555 28806
rect 30579 28804 30635 28806
rect 30659 28804 30715 28806
rect 30739 28804 30795 28806
rect 30499 27770 30555 27772
rect 30579 27770 30635 27772
rect 30659 27770 30715 27772
rect 30739 27770 30795 27772
rect 30499 27718 30545 27770
rect 30545 27718 30555 27770
rect 30579 27718 30609 27770
rect 30609 27718 30621 27770
rect 30621 27718 30635 27770
rect 30659 27718 30673 27770
rect 30673 27718 30685 27770
rect 30685 27718 30715 27770
rect 30739 27718 30749 27770
rect 30749 27718 30795 27770
rect 30499 27716 30555 27718
rect 30579 27716 30635 27718
rect 30659 27716 30715 27718
rect 30739 27716 30795 27718
rect 30499 26682 30555 26684
rect 30579 26682 30635 26684
rect 30659 26682 30715 26684
rect 30739 26682 30795 26684
rect 30499 26630 30545 26682
rect 30545 26630 30555 26682
rect 30579 26630 30609 26682
rect 30609 26630 30621 26682
rect 30621 26630 30635 26682
rect 30659 26630 30673 26682
rect 30673 26630 30685 26682
rect 30685 26630 30715 26682
rect 30739 26630 30749 26682
rect 30749 26630 30795 26682
rect 30499 26628 30555 26630
rect 30579 26628 30635 26630
rect 30659 26628 30715 26630
rect 30739 26628 30795 26630
rect 31022 28192 31078 28248
rect 30930 27512 30986 27568
rect 31298 26288 31354 26344
rect 30499 25594 30555 25596
rect 30579 25594 30635 25596
rect 30659 25594 30715 25596
rect 30739 25594 30795 25596
rect 30499 25542 30545 25594
rect 30545 25542 30555 25594
rect 30579 25542 30609 25594
rect 30609 25542 30621 25594
rect 30621 25542 30635 25594
rect 30659 25542 30673 25594
rect 30673 25542 30685 25594
rect 30685 25542 30715 25594
rect 30739 25542 30749 25594
rect 30749 25542 30795 25594
rect 30499 25540 30555 25542
rect 30579 25540 30635 25542
rect 30659 25540 30715 25542
rect 30739 25540 30795 25542
rect 31114 25336 31170 25392
rect 29734 20576 29790 20632
rect 29366 19624 29422 19680
rect 29090 16108 29146 16144
rect 29090 16088 29092 16108
rect 29092 16088 29144 16108
rect 29144 16088 29146 16108
rect 29090 15972 29146 16008
rect 29090 15952 29092 15972
rect 29092 15952 29144 15972
rect 29144 15952 29146 15972
rect 29734 18808 29790 18864
rect 29550 16632 29606 16688
rect 29366 16108 29422 16144
rect 29366 16088 29368 16108
rect 29368 16088 29420 16108
rect 29420 16088 29422 16108
rect 30499 24506 30555 24508
rect 30579 24506 30635 24508
rect 30659 24506 30715 24508
rect 30739 24506 30795 24508
rect 30499 24454 30545 24506
rect 30545 24454 30555 24506
rect 30579 24454 30609 24506
rect 30609 24454 30621 24506
rect 30621 24454 30635 24506
rect 30659 24454 30673 24506
rect 30673 24454 30685 24506
rect 30685 24454 30715 24506
rect 30739 24454 30749 24506
rect 30749 24454 30795 24506
rect 30499 24452 30555 24454
rect 30579 24452 30635 24454
rect 30659 24452 30715 24454
rect 30739 24452 30795 24454
rect 30499 23418 30555 23420
rect 30579 23418 30635 23420
rect 30659 23418 30715 23420
rect 30739 23418 30795 23420
rect 30499 23366 30545 23418
rect 30545 23366 30555 23418
rect 30579 23366 30609 23418
rect 30609 23366 30621 23418
rect 30621 23366 30635 23418
rect 30659 23366 30673 23418
rect 30673 23366 30685 23418
rect 30685 23366 30715 23418
rect 30739 23366 30749 23418
rect 30749 23366 30795 23418
rect 30499 23364 30555 23366
rect 30579 23364 30635 23366
rect 30659 23364 30715 23366
rect 30739 23364 30795 23366
rect 30499 22330 30555 22332
rect 30579 22330 30635 22332
rect 30659 22330 30715 22332
rect 30739 22330 30795 22332
rect 30499 22278 30545 22330
rect 30545 22278 30555 22330
rect 30579 22278 30609 22330
rect 30609 22278 30621 22330
rect 30621 22278 30635 22330
rect 30659 22278 30673 22330
rect 30673 22278 30685 22330
rect 30685 22278 30715 22330
rect 30739 22278 30749 22330
rect 30749 22278 30795 22330
rect 30499 22276 30555 22278
rect 30579 22276 30635 22278
rect 30659 22276 30715 22278
rect 30739 22276 30795 22278
rect 31574 29416 31630 29472
rect 31942 29824 31998 29880
rect 31758 29552 31814 29608
rect 31850 29180 31852 29200
rect 31852 29180 31904 29200
rect 31904 29180 31906 29200
rect 31850 29144 31906 29180
rect 32586 31864 32642 31920
rect 32402 29164 32458 29200
rect 32402 29144 32404 29164
rect 32404 29144 32456 29164
rect 32456 29144 32458 29164
rect 31758 27920 31814 27976
rect 31574 25200 31630 25256
rect 31574 25100 31576 25120
rect 31576 25100 31628 25120
rect 31628 25100 31630 25120
rect 31574 25064 31630 25100
rect 31482 24928 31538 24984
rect 30499 21242 30555 21244
rect 30579 21242 30635 21244
rect 30659 21242 30715 21244
rect 30739 21242 30795 21244
rect 30499 21190 30545 21242
rect 30545 21190 30555 21242
rect 30579 21190 30609 21242
rect 30609 21190 30621 21242
rect 30621 21190 30635 21242
rect 30659 21190 30673 21242
rect 30673 21190 30685 21242
rect 30685 21190 30715 21242
rect 30739 21190 30749 21242
rect 30749 21190 30795 21242
rect 30499 21188 30555 21190
rect 30579 21188 30635 21190
rect 30659 21188 30715 21190
rect 30739 21188 30795 21190
rect 30470 21004 30526 21040
rect 30470 20984 30472 21004
rect 30472 20984 30524 21004
rect 30524 20984 30526 21004
rect 30378 20712 30434 20768
rect 30499 20154 30555 20156
rect 30579 20154 30635 20156
rect 30659 20154 30715 20156
rect 30739 20154 30795 20156
rect 30499 20102 30545 20154
rect 30545 20102 30555 20154
rect 30579 20102 30609 20154
rect 30609 20102 30621 20154
rect 30621 20102 30635 20154
rect 30659 20102 30673 20154
rect 30673 20102 30685 20154
rect 30685 20102 30715 20154
rect 30739 20102 30749 20154
rect 30749 20102 30795 20154
rect 30499 20100 30555 20102
rect 30579 20100 30635 20102
rect 30659 20100 30715 20102
rect 30739 20100 30795 20102
rect 30499 19066 30555 19068
rect 30579 19066 30635 19068
rect 30659 19066 30715 19068
rect 30739 19066 30795 19068
rect 30499 19014 30545 19066
rect 30545 19014 30555 19066
rect 30579 19014 30609 19066
rect 30609 19014 30621 19066
rect 30621 19014 30635 19066
rect 30659 19014 30673 19066
rect 30673 19014 30685 19066
rect 30685 19014 30715 19066
rect 30739 19014 30749 19066
rect 30749 19014 30795 19066
rect 30499 19012 30555 19014
rect 30579 19012 30635 19014
rect 30659 19012 30715 19014
rect 30739 19012 30795 19014
rect 29826 15952 29882 16008
rect 28998 15544 29054 15600
rect 29366 15156 29422 15192
rect 29366 15136 29368 15156
rect 29368 15136 29420 15156
rect 29420 15136 29422 15156
rect 30499 17978 30555 17980
rect 30579 17978 30635 17980
rect 30659 17978 30715 17980
rect 30739 17978 30795 17980
rect 30499 17926 30545 17978
rect 30545 17926 30555 17978
rect 30579 17926 30609 17978
rect 30609 17926 30621 17978
rect 30621 17926 30635 17978
rect 30659 17926 30673 17978
rect 30673 17926 30685 17978
rect 30685 17926 30715 17978
rect 30739 17926 30749 17978
rect 30749 17926 30795 17978
rect 30499 17924 30555 17926
rect 30579 17924 30635 17926
rect 30659 17924 30715 17926
rect 30739 17924 30795 17926
rect 30470 17040 30526 17096
rect 30499 16890 30555 16892
rect 30579 16890 30635 16892
rect 30659 16890 30715 16892
rect 30739 16890 30795 16892
rect 30499 16838 30545 16890
rect 30545 16838 30555 16890
rect 30579 16838 30609 16890
rect 30609 16838 30621 16890
rect 30621 16838 30635 16890
rect 30659 16838 30673 16890
rect 30673 16838 30685 16890
rect 30685 16838 30715 16890
rect 30739 16838 30749 16890
rect 30749 16838 30795 16890
rect 30499 16836 30555 16838
rect 30579 16836 30635 16838
rect 30659 16836 30715 16838
rect 30739 16836 30795 16838
rect 30470 16668 30472 16688
rect 30472 16668 30524 16688
rect 30524 16668 30526 16688
rect 30470 16632 30526 16668
rect 30654 16632 30710 16688
rect 30746 16244 30802 16280
rect 30746 16224 30748 16244
rect 30748 16224 30800 16244
rect 30800 16224 30802 16244
rect 30499 15802 30555 15804
rect 30579 15802 30635 15804
rect 30659 15802 30715 15804
rect 30739 15802 30795 15804
rect 30499 15750 30545 15802
rect 30545 15750 30555 15802
rect 30579 15750 30609 15802
rect 30609 15750 30621 15802
rect 30621 15750 30635 15802
rect 30659 15750 30673 15802
rect 30673 15750 30685 15802
rect 30685 15750 30715 15802
rect 30739 15750 30749 15802
rect 30749 15750 30795 15802
rect 30499 15748 30555 15750
rect 30579 15748 30635 15750
rect 30659 15748 30715 15750
rect 30739 15748 30795 15750
rect 30930 16768 30986 16824
rect 30838 15544 30894 15600
rect 26278 14170 26334 14172
rect 26358 14170 26414 14172
rect 26438 14170 26494 14172
rect 26518 14170 26574 14172
rect 26278 14118 26324 14170
rect 26324 14118 26334 14170
rect 26358 14118 26388 14170
rect 26388 14118 26400 14170
rect 26400 14118 26414 14170
rect 26438 14118 26452 14170
rect 26452 14118 26464 14170
rect 26464 14118 26494 14170
rect 26518 14118 26528 14170
rect 26528 14118 26574 14170
rect 26278 14116 26334 14118
rect 26358 14116 26414 14118
rect 26438 14116 26494 14118
rect 26518 14116 26574 14118
rect 22058 13626 22114 13628
rect 22138 13626 22194 13628
rect 22218 13626 22274 13628
rect 22298 13626 22354 13628
rect 22058 13574 22104 13626
rect 22104 13574 22114 13626
rect 22138 13574 22168 13626
rect 22168 13574 22180 13626
rect 22180 13574 22194 13626
rect 22218 13574 22232 13626
rect 22232 13574 22244 13626
rect 22244 13574 22274 13626
rect 22298 13574 22308 13626
rect 22308 13574 22354 13626
rect 22058 13572 22114 13574
rect 22138 13572 22194 13574
rect 22218 13572 22274 13574
rect 22298 13572 22354 13574
rect 26278 13082 26334 13084
rect 26358 13082 26414 13084
rect 26438 13082 26494 13084
rect 26518 13082 26574 13084
rect 26278 13030 26324 13082
rect 26324 13030 26334 13082
rect 26358 13030 26388 13082
rect 26388 13030 26400 13082
rect 26400 13030 26414 13082
rect 26438 13030 26452 13082
rect 26452 13030 26464 13082
rect 26464 13030 26494 13082
rect 26518 13030 26528 13082
rect 26528 13030 26574 13082
rect 26278 13028 26334 13030
rect 26358 13028 26414 13030
rect 26438 13028 26494 13030
rect 26518 13028 26574 13030
rect 22058 12538 22114 12540
rect 22138 12538 22194 12540
rect 22218 12538 22274 12540
rect 22298 12538 22354 12540
rect 22058 12486 22104 12538
rect 22104 12486 22114 12538
rect 22138 12486 22168 12538
rect 22168 12486 22180 12538
rect 22180 12486 22194 12538
rect 22218 12486 22232 12538
rect 22232 12486 22244 12538
rect 22244 12486 22274 12538
rect 22298 12486 22308 12538
rect 22308 12486 22354 12538
rect 22058 12484 22114 12486
rect 22138 12484 22194 12486
rect 22218 12484 22274 12486
rect 22298 12484 22354 12486
rect 26278 11994 26334 11996
rect 26358 11994 26414 11996
rect 26438 11994 26494 11996
rect 26518 11994 26574 11996
rect 26278 11942 26324 11994
rect 26324 11942 26334 11994
rect 26358 11942 26388 11994
rect 26388 11942 26400 11994
rect 26400 11942 26414 11994
rect 26438 11942 26452 11994
rect 26452 11942 26464 11994
rect 26464 11942 26494 11994
rect 26518 11942 26528 11994
rect 26528 11942 26574 11994
rect 26278 11940 26334 11942
rect 26358 11940 26414 11942
rect 26438 11940 26494 11942
rect 26518 11940 26574 11942
rect 22058 11450 22114 11452
rect 22138 11450 22194 11452
rect 22218 11450 22274 11452
rect 22298 11450 22354 11452
rect 22058 11398 22104 11450
rect 22104 11398 22114 11450
rect 22138 11398 22168 11450
rect 22168 11398 22180 11450
rect 22180 11398 22194 11450
rect 22218 11398 22232 11450
rect 22232 11398 22244 11450
rect 22244 11398 22274 11450
rect 22298 11398 22308 11450
rect 22308 11398 22354 11450
rect 22058 11396 22114 11398
rect 22138 11396 22194 11398
rect 22218 11396 22274 11398
rect 22298 11396 22354 11398
rect 26278 10906 26334 10908
rect 26358 10906 26414 10908
rect 26438 10906 26494 10908
rect 26518 10906 26574 10908
rect 26278 10854 26324 10906
rect 26324 10854 26334 10906
rect 26358 10854 26388 10906
rect 26388 10854 26400 10906
rect 26400 10854 26414 10906
rect 26438 10854 26452 10906
rect 26452 10854 26464 10906
rect 26464 10854 26494 10906
rect 26518 10854 26528 10906
rect 26528 10854 26574 10906
rect 26278 10852 26334 10854
rect 26358 10852 26414 10854
rect 26438 10852 26494 10854
rect 26518 10852 26574 10854
rect 22058 10362 22114 10364
rect 22138 10362 22194 10364
rect 22218 10362 22274 10364
rect 22298 10362 22354 10364
rect 22058 10310 22104 10362
rect 22104 10310 22114 10362
rect 22138 10310 22168 10362
rect 22168 10310 22180 10362
rect 22180 10310 22194 10362
rect 22218 10310 22232 10362
rect 22232 10310 22244 10362
rect 22244 10310 22274 10362
rect 22298 10310 22308 10362
rect 22308 10310 22354 10362
rect 22058 10308 22114 10310
rect 22138 10308 22194 10310
rect 22218 10308 22274 10310
rect 22298 10308 22354 10310
rect 26278 9818 26334 9820
rect 26358 9818 26414 9820
rect 26438 9818 26494 9820
rect 26518 9818 26574 9820
rect 26278 9766 26324 9818
rect 26324 9766 26334 9818
rect 26358 9766 26388 9818
rect 26388 9766 26400 9818
rect 26400 9766 26414 9818
rect 26438 9766 26452 9818
rect 26452 9766 26464 9818
rect 26464 9766 26494 9818
rect 26518 9766 26528 9818
rect 26528 9766 26574 9818
rect 26278 9764 26334 9766
rect 26358 9764 26414 9766
rect 26438 9764 26494 9766
rect 26518 9764 26574 9766
rect 22058 9274 22114 9276
rect 22138 9274 22194 9276
rect 22218 9274 22274 9276
rect 22298 9274 22354 9276
rect 22058 9222 22104 9274
rect 22104 9222 22114 9274
rect 22138 9222 22168 9274
rect 22168 9222 22180 9274
rect 22180 9222 22194 9274
rect 22218 9222 22232 9274
rect 22232 9222 22244 9274
rect 22244 9222 22274 9274
rect 22298 9222 22308 9274
rect 22308 9222 22354 9274
rect 22058 9220 22114 9222
rect 22138 9220 22194 9222
rect 22218 9220 22274 9222
rect 22298 9220 22354 9222
rect 26278 8730 26334 8732
rect 26358 8730 26414 8732
rect 26438 8730 26494 8732
rect 26518 8730 26574 8732
rect 26278 8678 26324 8730
rect 26324 8678 26334 8730
rect 26358 8678 26388 8730
rect 26388 8678 26400 8730
rect 26400 8678 26414 8730
rect 26438 8678 26452 8730
rect 26452 8678 26464 8730
rect 26464 8678 26494 8730
rect 26518 8678 26528 8730
rect 26528 8678 26574 8730
rect 26278 8676 26334 8678
rect 26358 8676 26414 8678
rect 26438 8676 26494 8678
rect 26518 8676 26574 8678
rect 22058 8186 22114 8188
rect 22138 8186 22194 8188
rect 22218 8186 22274 8188
rect 22298 8186 22354 8188
rect 22058 8134 22104 8186
rect 22104 8134 22114 8186
rect 22138 8134 22168 8186
rect 22168 8134 22180 8186
rect 22180 8134 22194 8186
rect 22218 8134 22232 8186
rect 22232 8134 22244 8186
rect 22244 8134 22274 8186
rect 22298 8134 22308 8186
rect 22308 8134 22354 8186
rect 22058 8132 22114 8134
rect 22138 8132 22194 8134
rect 22218 8132 22274 8134
rect 22298 8132 22354 8134
rect 26278 7642 26334 7644
rect 26358 7642 26414 7644
rect 26438 7642 26494 7644
rect 26518 7642 26574 7644
rect 26278 7590 26324 7642
rect 26324 7590 26334 7642
rect 26358 7590 26388 7642
rect 26388 7590 26400 7642
rect 26400 7590 26414 7642
rect 26438 7590 26452 7642
rect 26452 7590 26464 7642
rect 26464 7590 26494 7642
rect 26518 7590 26528 7642
rect 26528 7590 26574 7642
rect 26278 7588 26334 7590
rect 26358 7588 26414 7590
rect 26438 7588 26494 7590
rect 26518 7588 26574 7590
rect 22058 7098 22114 7100
rect 22138 7098 22194 7100
rect 22218 7098 22274 7100
rect 22298 7098 22354 7100
rect 22058 7046 22104 7098
rect 22104 7046 22114 7098
rect 22138 7046 22168 7098
rect 22168 7046 22180 7098
rect 22180 7046 22194 7098
rect 22218 7046 22232 7098
rect 22232 7046 22244 7098
rect 22244 7046 22274 7098
rect 22298 7046 22308 7098
rect 22308 7046 22354 7098
rect 22058 7044 22114 7046
rect 22138 7044 22194 7046
rect 22218 7044 22274 7046
rect 22298 7044 22354 7046
rect 26278 6554 26334 6556
rect 26358 6554 26414 6556
rect 26438 6554 26494 6556
rect 26518 6554 26574 6556
rect 26278 6502 26324 6554
rect 26324 6502 26334 6554
rect 26358 6502 26388 6554
rect 26388 6502 26400 6554
rect 26400 6502 26414 6554
rect 26438 6502 26452 6554
rect 26452 6502 26464 6554
rect 26464 6502 26494 6554
rect 26518 6502 26528 6554
rect 26528 6502 26574 6554
rect 26278 6500 26334 6502
rect 26358 6500 26414 6502
rect 26438 6500 26494 6502
rect 26518 6500 26574 6502
rect 22058 6010 22114 6012
rect 22138 6010 22194 6012
rect 22218 6010 22274 6012
rect 22298 6010 22354 6012
rect 22058 5958 22104 6010
rect 22104 5958 22114 6010
rect 22138 5958 22168 6010
rect 22168 5958 22180 6010
rect 22180 5958 22194 6010
rect 22218 5958 22232 6010
rect 22232 5958 22244 6010
rect 22244 5958 22274 6010
rect 22298 5958 22308 6010
rect 22308 5958 22354 6010
rect 22058 5956 22114 5958
rect 22138 5956 22194 5958
rect 22218 5956 22274 5958
rect 22298 5956 22354 5958
rect 26278 5466 26334 5468
rect 26358 5466 26414 5468
rect 26438 5466 26494 5468
rect 26518 5466 26574 5468
rect 26278 5414 26324 5466
rect 26324 5414 26334 5466
rect 26358 5414 26388 5466
rect 26388 5414 26400 5466
rect 26400 5414 26414 5466
rect 26438 5414 26452 5466
rect 26452 5414 26464 5466
rect 26464 5414 26494 5466
rect 26518 5414 26528 5466
rect 26528 5414 26574 5466
rect 26278 5412 26334 5414
rect 26358 5412 26414 5414
rect 26438 5412 26494 5414
rect 26518 5412 26574 5414
rect 22058 4922 22114 4924
rect 22138 4922 22194 4924
rect 22218 4922 22274 4924
rect 22298 4922 22354 4924
rect 22058 4870 22104 4922
rect 22104 4870 22114 4922
rect 22138 4870 22168 4922
rect 22168 4870 22180 4922
rect 22180 4870 22194 4922
rect 22218 4870 22232 4922
rect 22232 4870 22244 4922
rect 22244 4870 22274 4922
rect 22298 4870 22308 4922
rect 22308 4870 22354 4922
rect 22058 4868 22114 4870
rect 22138 4868 22194 4870
rect 22218 4868 22274 4870
rect 22298 4868 22354 4870
rect 26278 4378 26334 4380
rect 26358 4378 26414 4380
rect 26438 4378 26494 4380
rect 26518 4378 26574 4380
rect 26278 4326 26324 4378
rect 26324 4326 26334 4378
rect 26358 4326 26388 4378
rect 26388 4326 26400 4378
rect 26400 4326 26414 4378
rect 26438 4326 26452 4378
rect 26452 4326 26464 4378
rect 26464 4326 26494 4378
rect 26518 4326 26528 4378
rect 26528 4326 26574 4378
rect 26278 4324 26334 4326
rect 26358 4324 26414 4326
rect 26438 4324 26494 4326
rect 26518 4324 26574 4326
rect 22058 3834 22114 3836
rect 22138 3834 22194 3836
rect 22218 3834 22274 3836
rect 22298 3834 22354 3836
rect 22058 3782 22104 3834
rect 22104 3782 22114 3834
rect 22138 3782 22168 3834
rect 22168 3782 22180 3834
rect 22180 3782 22194 3834
rect 22218 3782 22232 3834
rect 22232 3782 22244 3834
rect 22244 3782 22274 3834
rect 22298 3782 22308 3834
rect 22308 3782 22354 3834
rect 22058 3780 22114 3782
rect 22138 3780 22194 3782
rect 22218 3780 22274 3782
rect 22298 3780 22354 3782
rect 26278 3290 26334 3292
rect 26358 3290 26414 3292
rect 26438 3290 26494 3292
rect 26518 3290 26574 3292
rect 26278 3238 26324 3290
rect 26324 3238 26334 3290
rect 26358 3238 26388 3290
rect 26388 3238 26400 3290
rect 26400 3238 26414 3290
rect 26438 3238 26452 3290
rect 26452 3238 26464 3290
rect 26464 3238 26494 3290
rect 26518 3238 26528 3290
rect 26528 3238 26574 3290
rect 26278 3236 26334 3238
rect 26358 3236 26414 3238
rect 26438 3236 26494 3238
rect 26518 3236 26574 3238
rect 22058 2746 22114 2748
rect 22138 2746 22194 2748
rect 22218 2746 22274 2748
rect 22298 2746 22354 2748
rect 22058 2694 22104 2746
rect 22104 2694 22114 2746
rect 22138 2694 22168 2746
rect 22168 2694 22180 2746
rect 22180 2694 22194 2746
rect 22218 2694 22232 2746
rect 22232 2694 22244 2746
rect 22244 2694 22274 2746
rect 22298 2694 22308 2746
rect 22308 2694 22354 2746
rect 22058 2692 22114 2694
rect 22138 2692 22194 2694
rect 22218 2692 22274 2694
rect 22298 2692 22354 2694
rect 30499 14714 30555 14716
rect 30579 14714 30635 14716
rect 30659 14714 30715 14716
rect 30739 14714 30795 14716
rect 30499 14662 30545 14714
rect 30545 14662 30555 14714
rect 30579 14662 30609 14714
rect 30609 14662 30621 14714
rect 30621 14662 30635 14714
rect 30659 14662 30673 14714
rect 30673 14662 30685 14714
rect 30685 14662 30715 14714
rect 30739 14662 30749 14714
rect 30749 14662 30795 14714
rect 30499 14660 30555 14662
rect 30579 14660 30635 14662
rect 30659 14660 30715 14662
rect 30739 14660 30795 14662
rect 31298 18420 31354 18456
rect 31298 18400 31300 18420
rect 31300 18400 31352 18420
rect 31352 18400 31354 18420
rect 31206 16532 31208 16552
rect 31208 16532 31260 16552
rect 31260 16532 31262 16552
rect 31206 16496 31262 16532
rect 30499 13626 30555 13628
rect 30579 13626 30635 13628
rect 30659 13626 30715 13628
rect 30739 13626 30795 13628
rect 30499 13574 30545 13626
rect 30545 13574 30555 13626
rect 30579 13574 30609 13626
rect 30609 13574 30621 13626
rect 30621 13574 30635 13626
rect 30659 13574 30673 13626
rect 30673 13574 30685 13626
rect 30685 13574 30715 13626
rect 30739 13574 30749 13626
rect 30749 13574 30795 13626
rect 30499 13572 30555 13574
rect 30579 13572 30635 13574
rect 30659 13572 30715 13574
rect 30739 13572 30795 13574
rect 32034 27512 32090 27568
rect 32494 28328 32550 28384
rect 32034 25472 32090 25528
rect 32034 25064 32090 25120
rect 31758 24656 31814 24712
rect 31574 21004 31630 21040
rect 31574 20984 31576 21004
rect 31576 20984 31628 21004
rect 31628 20984 31630 21004
rect 33230 33768 33286 33824
rect 34334 34620 34336 34640
rect 34336 34620 34388 34640
rect 34388 34620 34390 34640
rect 34334 34584 34390 34620
rect 34426 34040 34482 34096
rect 34334 33360 34390 33416
rect 34719 34842 34775 34844
rect 34799 34842 34855 34844
rect 34879 34842 34935 34844
rect 34959 34842 35015 34844
rect 34719 34790 34765 34842
rect 34765 34790 34775 34842
rect 34799 34790 34829 34842
rect 34829 34790 34841 34842
rect 34841 34790 34855 34842
rect 34879 34790 34893 34842
rect 34893 34790 34905 34842
rect 34905 34790 34935 34842
rect 34959 34790 34969 34842
rect 34969 34790 35015 34842
rect 34719 34788 34775 34790
rect 34799 34788 34855 34790
rect 34879 34788 34935 34790
rect 34959 34788 35015 34790
rect 34719 33754 34775 33756
rect 34799 33754 34855 33756
rect 34879 33754 34935 33756
rect 34959 33754 35015 33756
rect 34719 33702 34765 33754
rect 34765 33702 34775 33754
rect 34799 33702 34829 33754
rect 34829 33702 34841 33754
rect 34841 33702 34855 33754
rect 34879 33702 34893 33754
rect 34893 33702 34905 33754
rect 34905 33702 34935 33754
rect 34959 33702 34969 33754
rect 34969 33702 35015 33754
rect 34719 33700 34775 33702
rect 34799 33700 34855 33702
rect 34879 33700 34935 33702
rect 34959 33700 35015 33702
rect 34610 32816 34666 32872
rect 33230 29824 33286 29880
rect 33322 29588 33324 29608
rect 33324 29588 33376 29608
rect 33376 29588 33378 29608
rect 33322 29552 33378 29588
rect 32770 28600 32826 28656
rect 32678 28464 32734 28520
rect 33874 29688 33930 29744
rect 33414 29008 33470 29064
rect 34719 32666 34775 32668
rect 34799 32666 34855 32668
rect 34879 32666 34935 32668
rect 34959 32666 35015 32668
rect 34719 32614 34765 32666
rect 34765 32614 34775 32666
rect 34799 32614 34829 32666
rect 34829 32614 34841 32666
rect 34841 32614 34855 32666
rect 34879 32614 34893 32666
rect 34893 32614 34905 32666
rect 34905 32614 34935 32666
rect 34959 32614 34969 32666
rect 34969 32614 35015 32666
rect 34719 32612 34775 32614
rect 34799 32612 34855 32614
rect 34879 32612 34935 32614
rect 34959 32612 35015 32614
rect 34334 32000 34390 32056
rect 34719 31578 34775 31580
rect 34799 31578 34855 31580
rect 34879 31578 34935 31580
rect 34959 31578 35015 31580
rect 34719 31526 34765 31578
rect 34765 31526 34775 31578
rect 34799 31526 34829 31578
rect 34829 31526 34841 31578
rect 34841 31526 34855 31578
rect 34879 31526 34893 31578
rect 34893 31526 34905 31578
rect 34905 31526 34935 31578
rect 34959 31526 34969 31578
rect 34969 31526 35015 31578
rect 34719 31524 34775 31526
rect 34799 31524 34855 31526
rect 34879 31524 34935 31526
rect 34959 31524 35015 31526
rect 34334 31340 34390 31376
rect 34334 31320 34336 31340
rect 34336 31320 34388 31340
rect 34388 31320 34390 31340
rect 34719 30490 34775 30492
rect 34799 30490 34855 30492
rect 34879 30490 34935 30492
rect 34959 30490 35015 30492
rect 34719 30438 34765 30490
rect 34765 30438 34775 30490
rect 34799 30438 34829 30490
rect 34829 30438 34841 30490
rect 34841 30438 34855 30490
rect 34879 30438 34893 30490
rect 34893 30438 34905 30490
rect 34905 30438 34935 30490
rect 34959 30438 34969 30490
rect 34969 30438 35015 30490
rect 34719 30436 34775 30438
rect 34799 30436 34855 30438
rect 34879 30436 34935 30438
rect 34959 30436 35015 30438
rect 34719 29402 34775 29404
rect 34799 29402 34855 29404
rect 34879 29402 34935 29404
rect 34959 29402 35015 29404
rect 34719 29350 34765 29402
rect 34765 29350 34775 29402
rect 34799 29350 34829 29402
rect 34829 29350 34841 29402
rect 34841 29350 34855 29402
rect 34879 29350 34893 29402
rect 34893 29350 34905 29402
rect 34905 29350 34935 29402
rect 34959 29350 34969 29402
rect 34969 29350 35015 29402
rect 34719 29348 34775 29350
rect 34799 29348 34855 29350
rect 34879 29348 34935 29350
rect 34959 29348 35015 29350
rect 34719 28314 34775 28316
rect 34799 28314 34855 28316
rect 34879 28314 34935 28316
rect 34959 28314 35015 28316
rect 34719 28262 34765 28314
rect 34765 28262 34775 28314
rect 34799 28262 34829 28314
rect 34829 28262 34841 28314
rect 34841 28262 34855 28314
rect 34879 28262 34893 28314
rect 34893 28262 34905 28314
rect 34905 28262 34935 28314
rect 34959 28262 34969 28314
rect 34969 28262 35015 28314
rect 34719 28260 34775 28262
rect 34799 28260 34855 28262
rect 34879 28260 34935 28262
rect 34959 28260 35015 28262
rect 34334 27956 34336 27976
rect 34336 27956 34388 27976
rect 34388 27956 34390 27976
rect 34334 27920 34390 27956
rect 34719 27226 34775 27228
rect 34799 27226 34855 27228
rect 34879 27226 34935 27228
rect 34959 27226 35015 27228
rect 34719 27174 34765 27226
rect 34765 27174 34775 27226
rect 34799 27174 34829 27226
rect 34829 27174 34841 27226
rect 34841 27174 34855 27226
rect 34879 27174 34893 27226
rect 34893 27174 34905 27226
rect 34905 27174 34935 27226
rect 34959 27174 34969 27226
rect 34969 27174 35015 27226
rect 34719 27172 34775 27174
rect 34799 27172 34855 27174
rect 34879 27172 34935 27174
rect 34959 27172 35015 27174
rect 32494 23840 32550 23896
rect 32494 23432 32550 23488
rect 32494 22616 32550 22672
rect 32678 24656 32734 24712
rect 32678 23704 32734 23760
rect 32678 23604 32680 23624
rect 32680 23604 32732 23624
rect 32732 23604 32734 23624
rect 32678 23568 32734 23604
rect 33322 25336 33378 25392
rect 31850 20848 31906 20904
rect 31482 16768 31538 16824
rect 31758 18808 31814 18864
rect 31666 18400 31722 18456
rect 31758 17040 31814 17096
rect 31574 13932 31630 13968
rect 31574 13912 31576 13932
rect 31576 13912 31628 13932
rect 31628 13912 31630 13932
rect 30499 12538 30555 12540
rect 30579 12538 30635 12540
rect 30659 12538 30715 12540
rect 30739 12538 30795 12540
rect 30499 12486 30545 12538
rect 30545 12486 30555 12538
rect 30579 12486 30609 12538
rect 30609 12486 30621 12538
rect 30621 12486 30635 12538
rect 30659 12486 30673 12538
rect 30673 12486 30685 12538
rect 30685 12486 30715 12538
rect 30739 12486 30749 12538
rect 30749 12486 30795 12538
rect 30499 12484 30555 12486
rect 30579 12484 30635 12486
rect 30659 12484 30715 12486
rect 30739 12484 30795 12486
rect 30499 11450 30555 11452
rect 30579 11450 30635 11452
rect 30659 11450 30715 11452
rect 30739 11450 30795 11452
rect 30499 11398 30545 11450
rect 30545 11398 30555 11450
rect 30579 11398 30609 11450
rect 30609 11398 30621 11450
rect 30621 11398 30635 11450
rect 30659 11398 30673 11450
rect 30673 11398 30685 11450
rect 30685 11398 30715 11450
rect 30739 11398 30749 11450
rect 30749 11398 30795 11450
rect 30499 11396 30555 11398
rect 30579 11396 30635 11398
rect 30659 11396 30715 11398
rect 30739 11396 30795 11398
rect 30499 10362 30555 10364
rect 30579 10362 30635 10364
rect 30659 10362 30715 10364
rect 30739 10362 30795 10364
rect 30499 10310 30545 10362
rect 30545 10310 30555 10362
rect 30579 10310 30609 10362
rect 30609 10310 30621 10362
rect 30621 10310 30635 10362
rect 30659 10310 30673 10362
rect 30673 10310 30685 10362
rect 30685 10310 30715 10362
rect 30739 10310 30749 10362
rect 30749 10310 30795 10362
rect 30499 10308 30555 10310
rect 30579 10308 30635 10310
rect 30659 10308 30715 10310
rect 30739 10308 30795 10310
rect 30499 9274 30555 9276
rect 30579 9274 30635 9276
rect 30659 9274 30715 9276
rect 30739 9274 30795 9276
rect 30499 9222 30545 9274
rect 30545 9222 30555 9274
rect 30579 9222 30609 9274
rect 30609 9222 30621 9274
rect 30621 9222 30635 9274
rect 30659 9222 30673 9274
rect 30673 9222 30685 9274
rect 30685 9222 30715 9274
rect 30739 9222 30749 9274
rect 30749 9222 30795 9274
rect 30499 9220 30555 9222
rect 30579 9220 30635 9222
rect 30659 9220 30715 9222
rect 30739 9220 30795 9222
rect 30499 8186 30555 8188
rect 30579 8186 30635 8188
rect 30659 8186 30715 8188
rect 30739 8186 30795 8188
rect 30499 8134 30545 8186
rect 30545 8134 30555 8186
rect 30579 8134 30609 8186
rect 30609 8134 30621 8186
rect 30621 8134 30635 8186
rect 30659 8134 30673 8186
rect 30673 8134 30685 8186
rect 30685 8134 30715 8186
rect 30739 8134 30749 8186
rect 30749 8134 30795 8186
rect 30499 8132 30555 8134
rect 30579 8132 30635 8134
rect 30659 8132 30715 8134
rect 30739 8132 30795 8134
rect 30499 7098 30555 7100
rect 30579 7098 30635 7100
rect 30659 7098 30715 7100
rect 30739 7098 30795 7100
rect 30499 7046 30545 7098
rect 30545 7046 30555 7098
rect 30579 7046 30609 7098
rect 30609 7046 30621 7098
rect 30621 7046 30635 7098
rect 30659 7046 30673 7098
rect 30673 7046 30685 7098
rect 30685 7046 30715 7098
rect 30739 7046 30749 7098
rect 30749 7046 30795 7098
rect 30499 7044 30555 7046
rect 30579 7044 30635 7046
rect 30659 7044 30715 7046
rect 30739 7044 30795 7046
rect 32402 18944 32458 19000
rect 32402 16244 32458 16280
rect 32402 16224 32404 16244
rect 32404 16224 32456 16244
rect 32456 16224 32458 16244
rect 31850 13524 31906 13560
rect 31850 13504 31852 13524
rect 31852 13504 31904 13524
rect 31904 13504 31906 13524
rect 30499 6010 30555 6012
rect 30579 6010 30635 6012
rect 30659 6010 30715 6012
rect 30739 6010 30795 6012
rect 30499 5958 30545 6010
rect 30545 5958 30555 6010
rect 30579 5958 30609 6010
rect 30609 5958 30621 6010
rect 30621 5958 30635 6010
rect 30659 5958 30673 6010
rect 30673 5958 30685 6010
rect 30685 5958 30715 6010
rect 30739 5958 30749 6010
rect 30749 5958 30795 6010
rect 30499 5956 30555 5958
rect 30579 5956 30635 5958
rect 30659 5956 30715 5958
rect 30739 5956 30795 5958
rect 30499 4922 30555 4924
rect 30579 4922 30635 4924
rect 30659 4922 30715 4924
rect 30739 4922 30795 4924
rect 30499 4870 30545 4922
rect 30545 4870 30555 4922
rect 30579 4870 30609 4922
rect 30609 4870 30621 4922
rect 30621 4870 30635 4922
rect 30659 4870 30673 4922
rect 30673 4870 30685 4922
rect 30685 4870 30715 4922
rect 30739 4870 30749 4922
rect 30749 4870 30795 4922
rect 30499 4868 30555 4870
rect 30579 4868 30635 4870
rect 30659 4868 30715 4870
rect 30739 4868 30795 4870
rect 30499 3834 30555 3836
rect 30579 3834 30635 3836
rect 30659 3834 30715 3836
rect 30739 3834 30795 3836
rect 30499 3782 30545 3834
rect 30545 3782 30555 3834
rect 30579 3782 30609 3834
rect 30609 3782 30621 3834
rect 30621 3782 30635 3834
rect 30659 3782 30673 3834
rect 30673 3782 30685 3834
rect 30685 3782 30715 3834
rect 30739 3782 30749 3834
rect 30749 3782 30795 3834
rect 30499 3780 30555 3782
rect 30579 3780 30635 3782
rect 30659 3780 30715 3782
rect 30739 3780 30795 3782
rect 26278 2202 26334 2204
rect 26358 2202 26414 2204
rect 26438 2202 26494 2204
rect 26518 2202 26574 2204
rect 26278 2150 26324 2202
rect 26324 2150 26334 2202
rect 26358 2150 26388 2202
rect 26388 2150 26400 2202
rect 26400 2150 26414 2202
rect 26438 2150 26452 2202
rect 26452 2150 26464 2202
rect 26464 2150 26494 2202
rect 26518 2150 26528 2202
rect 26528 2150 26574 2202
rect 26278 2148 26334 2150
rect 26358 2148 26414 2150
rect 26438 2148 26494 2150
rect 26518 2148 26574 2150
rect 30499 2746 30555 2748
rect 30579 2746 30635 2748
rect 30659 2746 30715 2748
rect 30739 2746 30795 2748
rect 30499 2694 30545 2746
rect 30545 2694 30555 2746
rect 30579 2694 30609 2746
rect 30609 2694 30621 2746
rect 30621 2694 30635 2746
rect 30659 2694 30673 2746
rect 30673 2694 30685 2746
rect 30685 2694 30715 2746
rect 30739 2694 30749 2746
rect 30749 2694 30795 2746
rect 30499 2692 30555 2694
rect 30579 2692 30635 2694
rect 30659 2692 30715 2694
rect 30739 2692 30795 2694
rect 32678 20712 32734 20768
rect 33046 21120 33102 21176
rect 33046 17992 33102 18048
rect 33598 25200 33654 25256
rect 33690 15544 33746 15600
rect 34719 26138 34775 26140
rect 34799 26138 34855 26140
rect 34879 26138 34935 26140
rect 34959 26138 35015 26140
rect 34719 26086 34765 26138
rect 34765 26086 34775 26138
rect 34799 26086 34829 26138
rect 34829 26086 34841 26138
rect 34841 26086 34855 26138
rect 34879 26086 34893 26138
rect 34893 26086 34905 26138
rect 34905 26086 34935 26138
rect 34959 26086 34969 26138
rect 34969 26086 35015 26138
rect 34719 26084 34775 26086
rect 34799 26084 34855 26086
rect 34879 26084 34935 26086
rect 34959 26084 35015 26086
rect 34334 25900 34390 25936
rect 34334 25880 34336 25900
rect 34336 25880 34388 25900
rect 34388 25880 34390 25900
rect 34334 25220 34390 25256
rect 34334 25200 34336 25220
rect 34336 25200 34388 25220
rect 34388 25200 34390 25220
rect 34719 25050 34775 25052
rect 34799 25050 34855 25052
rect 34879 25050 34935 25052
rect 34959 25050 35015 25052
rect 34719 24998 34765 25050
rect 34765 24998 34775 25050
rect 34799 24998 34829 25050
rect 34829 24998 34841 25050
rect 34841 24998 34855 25050
rect 34879 24998 34893 25050
rect 34893 24998 34905 25050
rect 34905 24998 34935 25050
rect 34959 24998 34969 25050
rect 34969 24998 35015 25050
rect 34719 24996 34775 24998
rect 34799 24996 34855 24998
rect 34879 24996 34935 24998
rect 34959 24996 35015 24998
rect 34426 24520 34482 24576
rect 34719 23962 34775 23964
rect 34799 23962 34855 23964
rect 34879 23962 34935 23964
rect 34959 23962 35015 23964
rect 34719 23910 34765 23962
rect 34765 23910 34775 23962
rect 34799 23910 34829 23962
rect 34829 23910 34841 23962
rect 34841 23910 34855 23962
rect 34879 23910 34893 23962
rect 34893 23910 34905 23962
rect 34905 23910 34935 23962
rect 34959 23910 34969 23962
rect 34969 23910 35015 23962
rect 34719 23908 34775 23910
rect 34799 23908 34855 23910
rect 34879 23908 34935 23910
rect 34959 23908 35015 23910
rect 34334 23704 34390 23760
rect 34334 23180 34390 23216
rect 34334 23160 34336 23180
rect 34336 23160 34388 23180
rect 34388 23160 34390 23180
rect 34334 22752 34390 22808
rect 34242 20596 34298 20632
rect 34242 20576 34244 20596
rect 34244 20576 34296 20596
rect 34296 20576 34298 20596
rect 34334 20440 34390 20496
rect 34334 19796 34336 19816
rect 34336 19796 34388 19816
rect 34388 19796 34390 19816
rect 34334 19760 34390 19796
rect 34334 19080 34390 19136
rect 34334 17740 34390 17776
rect 34334 17720 34336 17740
rect 34336 17720 34388 17740
rect 34388 17720 34390 17740
rect 34334 17076 34336 17096
rect 34336 17076 34388 17096
rect 34388 17076 34390 17096
rect 34334 17040 34390 17076
rect 34719 22874 34775 22876
rect 34799 22874 34855 22876
rect 34879 22874 34935 22876
rect 34959 22874 35015 22876
rect 34719 22822 34765 22874
rect 34765 22822 34775 22874
rect 34799 22822 34829 22874
rect 34829 22822 34841 22874
rect 34841 22822 34855 22874
rect 34879 22822 34893 22874
rect 34893 22822 34905 22874
rect 34905 22822 34935 22874
rect 34959 22822 34969 22874
rect 34969 22822 35015 22874
rect 34719 22820 34775 22822
rect 34799 22820 34855 22822
rect 34879 22820 34935 22822
rect 34959 22820 35015 22822
rect 34719 21786 34775 21788
rect 34799 21786 34855 21788
rect 34879 21786 34935 21788
rect 34959 21786 35015 21788
rect 34719 21734 34765 21786
rect 34765 21734 34775 21786
rect 34799 21734 34829 21786
rect 34829 21734 34841 21786
rect 34841 21734 34855 21786
rect 34879 21734 34893 21786
rect 34893 21734 34905 21786
rect 34905 21734 34935 21786
rect 34959 21734 34969 21786
rect 34969 21734 35015 21786
rect 34719 21732 34775 21734
rect 34799 21732 34855 21734
rect 34879 21732 34935 21734
rect 34959 21732 35015 21734
rect 34719 20698 34775 20700
rect 34799 20698 34855 20700
rect 34879 20698 34935 20700
rect 34959 20698 35015 20700
rect 34719 20646 34765 20698
rect 34765 20646 34775 20698
rect 34799 20646 34829 20698
rect 34829 20646 34841 20698
rect 34841 20646 34855 20698
rect 34879 20646 34893 20698
rect 34893 20646 34905 20698
rect 34905 20646 34935 20698
rect 34959 20646 34969 20698
rect 34969 20646 35015 20698
rect 34719 20644 34775 20646
rect 34799 20644 34855 20646
rect 34879 20644 34935 20646
rect 34959 20644 35015 20646
rect 34719 19610 34775 19612
rect 34799 19610 34855 19612
rect 34879 19610 34935 19612
rect 34959 19610 35015 19612
rect 34719 19558 34765 19610
rect 34765 19558 34775 19610
rect 34799 19558 34829 19610
rect 34829 19558 34841 19610
rect 34841 19558 34855 19610
rect 34879 19558 34893 19610
rect 34893 19558 34905 19610
rect 34905 19558 34935 19610
rect 34959 19558 34969 19610
rect 34969 19558 35015 19610
rect 34719 19556 34775 19558
rect 34799 19556 34855 19558
rect 34879 19556 34935 19558
rect 34959 19556 35015 19558
rect 34719 18522 34775 18524
rect 34799 18522 34855 18524
rect 34879 18522 34935 18524
rect 34959 18522 35015 18524
rect 34719 18470 34765 18522
rect 34765 18470 34775 18522
rect 34799 18470 34829 18522
rect 34829 18470 34841 18522
rect 34841 18470 34855 18522
rect 34879 18470 34893 18522
rect 34893 18470 34905 18522
rect 34905 18470 34935 18522
rect 34959 18470 34969 18522
rect 34969 18470 35015 18522
rect 34719 18468 34775 18470
rect 34799 18468 34855 18470
rect 34879 18468 34935 18470
rect 34959 18468 35015 18470
rect 34719 17434 34775 17436
rect 34799 17434 34855 17436
rect 34879 17434 34935 17436
rect 34959 17434 35015 17436
rect 34719 17382 34765 17434
rect 34765 17382 34775 17434
rect 34799 17382 34829 17434
rect 34829 17382 34841 17434
rect 34841 17382 34855 17434
rect 34879 17382 34893 17434
rect 34893 17382 34905 17434
rect 34905 17382 34935 17434
rect 34959 17382 34969 17434
rect 34969 17382 35015 17434
rect 34719 17380 34775 17382
rect 34799 17380 34855 17382
rect 34879 17380 34935 17382
rect 34959 17380 35015 17382
rect 35162 16360 35218 16416
rect 34719 16346 34775 16348
rect 34799 16346 34855 16348
rect 34879 16346 34935 16348
rect 34959 16346 35015 16348
rect 34719 16294 34765 16346
rect 34765 16294 34775 16346
rect 34799 16294 34829 16346
rect 34829 16294 34841 16346
rect 34841 16294 34855 16346
rect 34879 16294 34893 16346
rect 34893 16294 34905 16346
rect 34905 16294 34935 16346
rect 34959 16294 34969 16346
rect 34969 16294 35015 16346
rect 34719 16292 34775 16294
rect 34799 16292 34855 16294
rect 34879 16292 34935 16294
rect 34959 16292 35015 16294
rect 33782 15020 33838 15056
rect 33782 15000 33784 15020
rect 33784 15000 33836 15020
rect 33836 15000 33838 15020
rect 33598 13524 33654 13560
rect 33598 13504 33600 13524
rect 33600 13504 33652 13524
rect 33652 13504 33654 13524
rect 33782 13368 33838 13424
rect 33966 11756 34022 11792
rect 33966 11736 33968 11756
rect 33968 11736 34020 11756
rect 34020 11736 34022 11756
rect 33046 4120 33102 4176
rect 34719 15258 34775 15260
rect 34799 15258 34855 15260
rect 34879 15258 34935 15260
rect 34959 15258 35015 15260
rect 34719 15206 34765 15258
rect 34765 15206 34775 15258
rect 34799 15206 34829 15258
rect 34829 15206 34841 15258
rect 34841 15206 34855 15258
rect 34879 15206 34893 15258
rect 34893 15206 34905 15258
rect 34905 15206 34935 15258
rect 34959 15206 34969 15258
rect 34969 15206 35015 15258
rect 34719 15204 34775 15206
rect 34799 15204 34855 15206
rect 34879 15204 34935 15206
rect 34959 15204 35015 15206
rect 34334 14356 34336 14376
rect 34336 14356 34388 14376
rect 34388 14356 34390 14376
rect 34334 14320 34390 14356
rect 34719 14170 34775 14172
rect 34799 14170 34855 14172
rect 34879 14170 34935 14172
rect 34959 14170 35015 14172
rect 34719 14118 34765 14170
rect 34765 14118 34775 14170
rect 34799 14118 34829 14170
rect 34829 14118 34841 14170
rect 34841 14118 34855 14170
rect 34879 14118 34893 14170
rect 34893 14118 34905 14170
rect 34905 14118 34935 14170
rect 34959 14118 34969 14170
rect 34969 14118 35015 14170
rect 34719 14116 34775 14118
rect 34799 14116 34855 14118
rect 34879 14116 34935 14118
rect 34959 14116 35015 14118
rect 34334 13640 34390 13696
rect 34719 13082 34775 13084
rect 34799 13082 34855 13084
rect 34879 13082 34935 13084
rect 34959 13082 35015 13084
rect 34719 13030 34765 13082
rect 34765 13030 34775 13082
rect 34799 13030 34829 13082
rect 34829 13030 34841 13082
rect 34841 13030 34855 13082
rect 34879 13030 34893 13082
rect 34893 13030 34905 13082
rect 34905 13030 34935 13082
rect 34959 13030 34969 13082
rect 34969 13030 35015 13082
rect 34719 13028 34775 13030
rect 34799 13028 34855 13030
rect 34879 13028 34935 13030
rect 34959 13028 35015 13030
rect 34334 12860 34336 12880
rect 34336 12860 34388 12880
rect 34388 12860 34390 12880
rect 34334 12824 34390 12860
rect 34334 12300 34390 12336
rect 34334 12280 34336 12300
rect 34336 12280 34388 12300
rect 34388 12280 34390 12300
rect 34719 11994 34775 11996
rect 34799 11994 34855 11996
rect 34879 11994 34935 11996
rect 34959 11994 35015 11996
rect 34719 11942 34765 11994
rect 34765 11942 34775 11994
rect 34799 11942 34829 11994
rect 34829 11942 34841 11994
rect 34841 11942 34855 11994
rect 34879 11942 34893 11994
rect 34893 11942 34905 11994
rect 34905 11942 34935 11994
rect 34959 11942 34969 11994
rect 34969 11942 35015 11994
rect 34719 11940 34775 11942
rect 34799 11940 34855 11942
rect 34879 11940 34935 11942
rect 34959 11940 35015 11942
rect 34719 10906 34775 10908
rect 34799 10906 34855 10908
rect 34879 10906 34935 10908
rect 34959 10906 35015 10908
rect 34719 10854 34765 10906
rect 34765 10854 34775 10906
rect 34799 10854 34829 10906
rect 34829 10854 34841 10906
rect 34841 10854 34855 10906
rect 34879 10854 34893 10906
rect 34893 10854 34905 10906
rect 34905 10854 34935 10906
rect 34959 10854 34969 10906
rect 34969 10854 35015 10906
rect 34719 10852 34775 10854
rect 34799 10852 34855 10854
rect 34879 10852 34935 10854
rect 34959 10852 35015 10854
rect 34719 9818 34775 9820
rect 34799 9818 34855 9820
rect 34879 9818 34935 9820
rect 34959 9818 35015 9820
rect 34719 9766 34765 9818
rect 34765 9766 34775 9818
rect 34799 9766 34829 9818
rect 34829 9766 34841 9818
rect 34841 9766 34855 9818
rect 34879 9766 34893 9818
rect 34893 9766 34905 9818
rect 34905 9766 34935 9818
rect 34959 9766 34969 9818
rect 34969 9766 35015 9818
rect 34719 9764 34775 9766
rect 34799 9764 34855 9766
rect 34879 9764 34935 9766
rect 34959 9764 35015 9766
rect 34058 9560 34114 9616
rect 34334 8880 34390 8936
rect 34719 8730 34775 8732
rect 34799 8730 34855 8732
rect 34879 8730 34935 8732
rect 34959 8730 35015 8732
rect 34719 8678 34765 8730
rect 34765 8678 34775 8730
rect 34799 8678 34829 8730
rect 34829 8678 34841 8730
rect 34841 8678 34855 8730
rect 34879 8678 34893 8730
rect 34893 8678 34905 8730
rect 34905 8678 34935 8730
rect 34959 8678 34969 8730
rect 34969 8678 35015 8730
rect 34719 8676 34775 8678
rect 34799 8676 34855 8678
rect 34879 8676 34935 8678
rect 34959 8676 35015 8678
rect 34719 7642 34775 7644
rect 34799 7642 34855 7644
rect 34879 7642 34935 7644
rect 34959 7642 35015 7644
rect 34719 7590 34765 7642
rect 34765 7590 34775 7642
rect 34799 7590 34829 7642
rect 34829 7590 34841 7642
rect 34841 7590 34855 7642
rect 34879 7590 34893 7642
rect 34893 7590 34905 7642
rect 34905 7590 34935 7642
rect 34959 7590 34969 7642
rect 34969 7590 35015 7642
rect 34719 7588 34775 7590
rect 34799 7588 34855 7590
rect 34879 7588 34935 7590
rect 34959 7588 35015 7590
rect 34334 6860 34390 6896
rect 34334 6840 34336 6860
rect 34336 6840 34388 6860
rect 34388 6840 34390 6860
rect 34719 6554 34775 6556
rect 34799 6554 34855 6556
rect 34879 6554 34935 6556
rect 34959 6554 35015 6556
rect 34719 6502 34765 6554
rect 34765 6502 34775 6554
rect 34799 6502 34829 6554
rect 34829 6502 34841 6554
rect 34841 6502 34855 6554
rect 34879 6502 34893 6554
rect 34893 6502 34905 6554
rect 34905 6502 34935 6554
rect 34959 6502 34969 6554
rect 34969 6502 35015 6554
rect 34719 6500 34775 6502
rect 34799 6500 34855 6502
rect 34879 6500 34935 6502
rect 34959 6500 35015 6502
rect 34334 4800 34390 4856
rect 34334 3440 34390 3496
rect 34719 5466 34775 5468
rect 34799 5466 34855 5468
rect 34879 5466 34935 5468
rect 34959 5466 35015 5468
rect 34719 5414 34765 5466
rect 34765 5414 34775 5466
rect 34799 5414 34829 5466
rect 34829 5414 34841 5466
rect 34841 5414 34855 5466
rect 34879 5414 34893 5466
rect 34893 5414 34905 5466
rect 34905 5414 34935 5466
rect 34959 5414 34969 5466
rect 34969 5414 35015 5466
rect 34719 5412 34775 5414
rect 34799 5412 34855 5414
rect 34879 5412 34935 5414
rect 34959 5412 35015 5414
rect 34719 4378 34775 4380
rect 34799 4378 34855 4380
rect 34879 4378 34935 4380
rect 34959 4378 35015 4380
rect 34719 4326 34765 4378
rect 34765 4326 34775 4378
rect 34799 4326 34829 4378
rect 34829 4326 34841 4378
rect 34841 4326 34855 4378
rect 34879 4326 34893 4378
rect 34893 4326 34905 4378
rect 34905 4326 34935 4378
rect 34959 4326 34969 4378
rect 34969 4326 35015 4378
rect 34719 4324 34775 4326
rect 34799 4324 34855 4326
rect 34879 4324 34935 4326
rect 34959 4324 35015 4326
rect 34719 3290 34775 3292
rect 34799 3290 34855 3292
rect 34879 3290 34935 3292
rect 34959 3290 35015 3292
rect 34719 3238 34765 3290
rect 34765 3238 34775 3290
rect 34799 3238 34829 3290
rect 34829 3238 34841 3290
rect 34841 3238 34855 3290
rect 34879 3238 34893 3290
rect 34893 3238 34905 3290
rect 34905 3238 34935 3290
rect 34959 3238 34969 3290
rect 34969 3238 35015 3290
rect 34719 3236 34775 3238
rect 34799 3236 34855 3238
rect 34879 3236 34935 3238
rect 34959 3236 35015 3238
rect 34719 2202 34775 2204
rect 34799 2202 34855 2204
rect 34879 2202 34935 2204
rect 34959 2202 35015 2204
rect 34719 2150 34765 2202
rect 34765 2150 34775 2202
rect 34799 2150 34829 2202
rect 34829 2150 34841 2202
rect 34841 2150 34855 2202
rect 34879 2150 34893 2202
rect 34893 2150 34905 2202
rect 34905 2150 34935 2202
rect 34959 2150 34969 2202
rect 34969 2150 35015 2202
rect 34719 2148 34775 2150
rect 34799 2148 34855 2150
rect 34879 2148 34935 2150
rect 34959 2148 35015 2150
rect 34610 856 34666 912
rect 35898 2080 35954 2136
rect 31850 40 31906 96
<< metal3 >>
rect 200 41578 800 41668
rect 2773 41578 2839 41581
rect 200 41576 2839 41578
rect 200 41520 2778 41576
rect 2834 41520 2839 41576
rect 200 41518 2839 41520
rect 200 41428 800 41518
rect 2773 41515 2839 41518
rect 200 40898 800 40988
rect 3417 40898 3483 40901
rect 200 40896 3483 40898
rect 200 40840 3422 40896
rect 3478 40840 3483 40896
rect 200 40838 3483 40840
rect 200 40748 800 40838
rect 3417 40835 3483 40838
rect 33041 40898 33107 40901
rect 35200 40898 35800 40988
rect 33041 40896 35800 40898
rect 33041 40840 33046 40896
rect 33102 40840 35800 40896
rect 33041 40838 35800 40840
rect 33041 40835 33107 40838
rect 35200 40748 35800 40838
rect 35200 40068 35800 40308
rect 5166 39744 5482 39745
rect 5166 39680 5172 39744
rect 5236 39680 5252 39744
rect 5316 39680 5332 39744
rect 5396 39680 5412 39744
rect 5476 39680 5482 39744
rect 5166 39679 5482 39680
rect 13607 39744 13923 39745
rect 13607 39680 13613 39744
rect 13677 39680 13693 39744
rect 13757 39680 13773 39744
rect 13837 39680 13853 39744
rect 13917 39680 13923 39744
rect 13607 39679 13923 39680
rect 22048 39744 22364 39745
rect 22048 39680 22054 39744
rect 22118 39680 22134 39744
rect 22198 39680 22214 39744
rect 22278 39680 22294 39744
rect 22358 39680 22364 39744
rect 22048 39679 22364 39680
rect 30489 39744 30805 39745
rect 30489 39680 30495 39744
rect 30559 39680 30575 39744
rect 30639 39680 30655 39744
rect 30719 39680 30735 39744
rect 30799 39680 30805 39744
rect 30489 39679 30805 39680
rect 200 39388 800 39628
rect 32213 39538 32279 39541
rect 35200 39538 35800 39628
rect 32213 39536 35800 39538
rect 32213 39480 32218 39536
rect 32274 39480 35800 39536
rect 32213 39478 35800 39480
rect 32213 39475 32279 39478
rect 13721 39402 13787 39405
rect 30966 39402 30972 39404
rect 13721 39400 30972 39402
rect 13721 39344 13726 39400
rect 13782 39344 30972 39400
rect 13721 39342 30972 39344
rect 13721 39339 13787 39342
rect 30966 39340 30972 39342
rect 31036 39340 31042 39404
rect 35200 39388 35800 39478
rect 9386 39200 9702 39201
rect 9386 39136 9392 39200
rect 9456 39136 9472 39200
rect 9536 39136 9552 39200
rect 9616 39136 9632 39200
rect 9696 39136 9702 39200
rect 9386 39135 9702 39136
rect 17827 39200 18143 39201
rect 17827 39136 17833 39200
rect 17897 39136 17913 39200
rect 17977 39136 17993 39200
rect 18057 39136 18073 39200
rect 18137 39136 18143 39200
rect 17827 39135 18143 39136
rect 26268 39200 26584 39201
rect 26268 39136 26274 39200
rect 26338 39136 26354 39200
rect 26418 39136 26434 39200
rect 26498 39136 26514 39200
rect 26578 39136 26584 39200
rect 26268 39135 26584 39136
rect 34709 39200 35025 39201
rect 34709 39136 34715 39200
rect 34779 39136 34795 39200
rect 34859 39136 34875 39200
rect 34939 39136 34955 39200
rect 35019 39136 35025 39200
rect 34709 39135 35025 39136
rect 21449 38994 21515 38997
rect 27613 38994 27679 38997
rect 21449 38992 27679 38994
rect 200 38858 800 38948
rect 21449 38936 21454 38992
rect 21510 38936 27618 38992
rect 27674 38936 27679 38992
rect 21449 38934 27679 38936
rect 21449 38931 21515 38934
rect 27613 38931 27679 38934
rect 3509 38858 3575 38861
rect 200 38856 3575 38858
rect 200 38800 3514 38856
rect 3570 38800 3575 38856
rect 200 38798 3575 38800
rect 200 38708 800 38798
rect 3509 38795 3575 38798
rect 34329 38858 34395 38861
rect 35200 38858 35800 38948
rect 34329 38856 35800 38858
rect 34329 38800 34334 38856
rect 34390 38800 35800 38856
rect 34329 38798 35800 38800
rect 34329 38795 34395 38798
rect 35200 38708 35800 38798
rect 5166 38656 5482 38657
rect 5166 38592 5172 38656
rect 5236 38592 5252 38656
rect 5316 38592 5332 38656
rect 5396 38592 5412 38656
rect 5476 38592 5482 38656
rect 5166 38591 5482 38592
rect 13607 38656 13923 38657
rect 13607 38592 13613 38656
rect 13677 38592 13693 38656
rect 13757 38592 13773 38656
rect 13837 38592 13853 38656
rect 13917 38592 13923 38656
rect 13607 38591 13923 38592
rect 22048 38656 22364 38657
rect 22048 38592 22054 38656
rect 22118 38592 22134 38656
rect 22198 38592 22214 38656
rect 22278 38592 22294 38656
rect 22358 38592 22364 38656
rect 22048 38591 22364 38592
rect 30489 38656 30805 38657
rect 30489 38592 30495 38656
rect 30559 38592 30575 38656
rect 30639 38592 30655 38656
rect 30719 38592 30735 38656
rect 30799 38592 30805 38656
rect 30489 38591 30805 38592
rect 21357 38314 21423 38317
rect 26417 38314 26483 38317
rect 21357 38312 26483 38314
rect 200 38028 800 38268
rect 21357 38256 21362 38312
rect 21418 38256 26422 38312
rect 26478 38256 26483 38312
rect 21357 38254 26483 38256
rect 21357 38251 21423 38254
rect 26417 38251 26483 38254
rect 35200 38178 35800 38268
rect 9386 38112 9702 38113
rect 9386 38048 9392 38112
rect 9456 38048 9472 38112
rect 9536 38048 9552 38112
rect 9616 38048 9632 38112
rect 9696 38048 9702 38112
rect 9386 38047 9702 38048
rect 17827 38112 18143 38113
rect 17827 38048 17833 38112
rect 17897 38048 17913 38112
rect 17977 38048 17993 38112
rect 18057 38048 18073 38112
rect 18137 38048 18143 38112
rect 17827 38047 18143 38048
rect 26268 38112 26584 38113
rect 26268 38048 26274 38112
rect 26338 38048 26354 38112
rect 26418 38048 26434 38112
rect 26498 38048 26514 38112
rect 26578 38048 26584 38112
rect 26268 38047 26584 38048
rect 34709 38112 35025 38113
rect 34709 38048 34715 38112
rect 34779 38048 34795 38112
rect 34859 38048 34875 38112
rect 34939 38048 34955 38112
rect 35019 38048 35025 38112
rect 34709 38047 35025 38048
rect 35160 38028 35800 38178
rect 35160 37982 35266 38028
rect 23749 37906 23815 37909
rect 25313 37906 25379 37909
rect 23749 37904 25379 37906
rect 23749 37848 23754 37904
rect 23810 37848 25318 37904
rect 25374 37848 25379 37904
rect 23749 37846 25379 37848
rect 23749 37843 23815 37846
rect 25313 37843 25379 37846
rect 30005 37906 30071 37909
rect 32213 37906 32279 37909
rect 30005 37904 32279 37906
rect 30005 37848 30010 37904
rect 30066 37848 32218 37904
rect 32274 37848 32279 37904
rect 30005 37846 32279 37848
rect 30005 37843 30071 37846
rect 32213 37843 32279 37846
rect 34329 37906 34395 37909
rect 35206 37906 35266 37982
rect 34329 37904 35266 37906
rect 34329 37848 34334 37904
rect 34390 37848 35266 37904
rect 34329 37846 35266 37848
rect 34329 37843 34395 37846
rect 25037 37770 25103 37773
rect 27153 37770 27219 37773
rect 25037 37768 27219 37770
rect 25037 37712 25042 37768
rect 25098 37712 27158 37768
rect 27214 37712 27219 37768
rect 25037 37710 27219 37712
rect 25037 37707 25103 37710
rect 27153 37707 27219 37710
rect 29913 37770 29979 37773
rect 32121 37770 32187 37773
rect 29913 37768 32187 37770
rect 29913 37712 29918 37768
rect 29974 37712 32126 37768
rect 32182 37712 32187 37768
rect 29913 37710 32187 37712
rect 29913 37707 29979 37710
rect 32121 37707 32187 37710
rect 28073 37634 28139 37637
rect 28758 37634 28764 37636
rect 28073 37632 28764 37634
rect 200 37498 800 37588
rect 28073 37576 28078 37632
rect 28134 37576 28764 37632
rect 28073 37574 28764 37576
rect 28073 37571 28139 37574
rect 28758 37572 28764 37574
rect 28828 37572 28834 37636
rect 5166 37568 5482 37569
rect 5166 37504 5172 37568
rect 5236 37504 5252 37568
rect 5316 37504 5332 37568
rect 5396 37504 5412 37568
rect 5476 37504 5482 37568
rect 5166 37503 5482 37504
rect 13607 37568 13923 37569
rect 13607 37504 13613 37568
rect 13677 37504 13693 37568
rect 13757 37504 13773 37568
rect 13837 37504 13853 37568
rect 13917 37504 13923 37568
rect 13607 37503 13923 37504
rect 22048 37568 22364 37569
rect 22048 37504 22054 37568
rect 22118 37504 22134 37568
rect 22198 37504 22214 37568
rect 22278 37504 22294 37568
rect 22358 37504 22364 37568
rect 22048 37503 22364 37504
rect 30489 37568 30805 37569
rect 30489 37504 30495 37568
rect 30559 37504 30575 37568
rect 30639 37504 30655 37568
rect 30719 37504 30735 37568
rect 30799 37504 30805 37568
rect 30489 37503 30805 37504
rect 2037 37498 2103 37501
rect 200 37496 2103 37498
rect 200 37440 2042 37496
rect 2098 37440 2103 37496
rect 200 37438 2103 37440
rect 200 37348 800 37438
rect 2037 37435 2103 37438
rect 24025 37498 24091 37501
rect 28942 37498 28948 37500
rect 24025 37496 28948 37498
rect 24025 37440 24030 37496
rect 24086 37440 28948 37496
rect 24025 37438 28948 37440
rect 24025 37435 24091 37438
rect 28942 37436 28948 37438
rect 29012 37436 29018 37500
rect 29085 37498 29151 37501
rect 29310 37498 29316 37500
rect 29085 37496 29316 37498
rect 29085 37440 29090 37496
rect 29146 37440 29316 37496
rect 29085 37438 29316 37440
rect 29085 37435 29151 37438
rect 29310 37436 29316 37438
rect 29380 37436 29386 37500
rect 31937 37498 32003 37501
rect 30928 37496 32003 37498
rect 30928 37440 31942 37496
rect 31998 37440 32003 37496
rect 30928 37438 32003 37440
rect 25681 37362 25747 37365
rect 29729 37362 29795 37365
rect 25681 37360 29795 37362
rect 25681 37304 25686 37360
rect 25742 37304 29734 37360
rect 29790 37304 29795 37360
rect 25681 37302 29795 37304
rect 25681 37299 25747 37302
rect 29729 37299 29795 37302
rect 30005 37362 30071 37365
rect 30928 37362 30988 37438
rect 31937 37435 32003 37438
rect 30005 37360 30988 37362
rect 30005 37304 30010 37360
rect 30066 37304 30988 37360
rect 35200 37348 35800 37588
rect 30005 37302 30988 37304
rect 30005 37299 30071 37302
rect 18873 37226 18939 37229
rect 31017 37226 31083 37229
rect 18873 37224 31083 37226
rect 18873 37168 18878 37224
rect 18934 37168 31022 37224
rect 31078 37168 31083 37224
rect 18873 37166 31083 37168
rect 18873 37163 18939 37166
rect 31017 37163 31083 37166
rect 31293 37226 31359 37229
rect 31518 37226 31524 37228
rect 31293 37224 31524 37226
rect 31293 37168 31298 37224
rect 31354 37168 31524 37224
rect 31293 37166 31524 37168
rect 31293 37163 31359 37166
rect 31518 37164 31524 37166
rect 31588 37164 31594 37228
rect 23473 37090 23539 37093
rect 24669 37092 24735 37093
rect 30925 37092 30991 37093
rect 24669 37090 24716 37092
rect 23473 37088 24716 37090
rect 23473 37032 23478 37088
rect 23534 37032 24674 37088
rect 23473 37030 24716 37032
rect 23473 37027 23539 37030
rect 24669 37028 24716 37030
rect 24780 37028 24786 37092
rect 30925 37090 30972 37092
rect 30880 37088 30972 37090
rect 30880 37032 30930 37088
rect 30880 37030 30972 37032
rect 30925 37028 30972 37030
rect 31036 37028 31042 37092
rect 24669 37027 24735 37028
rect 30925 37027 30991 37028
rect 9386 37024 9702 37025
rect 9386 36960 9392 37024
rect 9456 36960 9472 37024
rect 9536 36960 9552 37024
rect 9616 36960 9632 37024
rect 9696 36960 9702 37024
rect 9386 36959 9702 36960
rect 17827 37024 18143 37025
rect 17827 36960 17833 37024
rect 17897 36960 17913 37024
rect 17977 36960 17993 37024
rect 18057 36960 18073 37024
rect 18137 36960 18143 37024
rect 17827 36959 18143 36960
rect 26268 37024 26584 37025
rect 26268 36960 26274 37024
rect 26338 36960 26354 37024
rect 26418 36960 26434 37024
rect 26498 36960 26514 37024
rect 26578 36960 26584 37024
rect 26268 36959 26584 36960
rect 34709 37024 35025 37025
rect 34709 36960 34715 37024
rect 34779 36960 34795 37024
rect 34859 36960 34875 37024
rect 34939 36960 34955 37024
rect 35019 36960 35025 37024
rect 34709 36959 35025 36960
rect 27153 36954 27219 36957
rect 32305 36954 32371 36957
rect 27153 36952 32371 36954
rect 200 36818 800 36908
rect 27153 36896 27158 36952
rect 27214 36896 32310 36952
rect 32366 36896 32371 36952
rect 27153 36894 32371 36896
rect 27153 36891 27219 36894
rect 32305 36891 32371 36894
rect 2773 36818 2839 36821
rect 200 36816 2839 36818
rect 200 36760 2778 36816
rect 2834 36760 2839 36816
rect 200 36758 2839 36760
rect 200 36668 800 36758
rect 2773 36755 2839 36758
rect 17585 36818 17651 36821
rect 32029 36818 32095 36821
rect 17585 36816 32095 36818
rect 17585 36760 17590 36816
rect 17646 36760 32034 36816
rect 32090 36760 32095 36816
rect 17585 36758 32095 36760
rect 17585 36755 17651 36758
rect 32029 36755 32095 36758
rect 34329 36818 34395 36821
rect 35200 36818 35800 36908
rect 34329 36816 35800 36818
rect 34329 36760 34334 36816
rect 34390 36760 35800 36816
rect 34329 36758 35800 36760
rect 34329 36755 34395 36758
rect 20621 36682 20687 36685
rect 32489 36682 32555 36685
rect 20621 36680 32555 36682
rect 20621 36624 20626 36680
rect 20682 36624 32494 36680
rect 32550 36624 32555 36680
rect 35200 36668 35800 36758
rect 20621 36622 32555 36624
rect 20621 36619 20687 36622
rect 32489 36619 32555 36622
rect 29177 36548 29243 36549
rect 29126 36546 29132 36548
rect 29086 36486 29132 36546
rect 29196 36544 29243 36548
rect 29238 36488 29243 36544
rect 29126 36484 29132 36486
rect 29196 36484 29243 36488
rect 29177 36483 29243 36484
rect 29453 36548 29519 36549
rect 29453 36544 29500 36548
rect 29564 36546 29570 36548
rect 29453 36488 29458 36544
rect 29453 36484 29500 36488
rect 29564 36486 29610 36546
rect 29564 36484 29570 36486
rect 29453 36483 29519 36484
rect 5166 36480 5482 36481
rect 5166 36416 5172 36480
rect 5236 36416 5252 36480
rect 5316 36416 5332 36480
rect 5396 36416 5412 36480
rect 5476 36416 5482 36480
rect 5166 36415 5482 36416
rect 13607 36480 13923 36481
rect 13607 36416 13613 36480
rect 13677 36416 13693 36480
rect 13757 36416 13773 36480
rect 13837 36416 13853 36480
rect 13917 36416 13923 36480
rect 13607 36415 13923 36416
rect 22048 36480 22364 36481
rect 22048 36416 22054 36480
rect 22118 36416 22134 36480
rect 22198 36416 22214 36480
rect 22278 36416 22294 36480
rect 22358 36416 22364 36480
rect 22048 36415 22364 36416
rect 30489 36480 30805 36481
rect 30489 36416 30495 36480
rect 30559 36416 30575 36480
rect 30639 36416 30655 36480
rect 30719 36416 30735 36480
rect 30799 36416 30805 36480
rect 30489 36415 30805 36416
rect 22461 36410 22527 36413
rect 29085 36410 29151 36413
rect 22461 36408 29151 36410
rect 22461 36352 22466 36408
rect 22522 36352 29090 36408
rect 29146 36352 29151 36408
rect 22461 36350 29151 36352
rect 22461 36347 22527 36350
rect 29085 36347 29151 36350
rect 29913 36410 29979 36413
rect 31109 36412 31175 36413
rect 30230 36410 30236 36412
rect 29913 36408 30236 36410
rect 29913 36352 29918 36408
rect 29974 36352 30236 36408
rect 29913 36350 30236 36352
rect 29913 36347 29979 36350
rect 30230 36348 30236 36350
rect 30300 36348 30306 36412
rect 31109 36408 31156 36412
rect 31220 36410 31226 36412
rect 31109 36352 31114 36408
rect 31109 36348 31156 36352
rect 31220 36350 31266 36410
rect 31220 36348 31226 36350
rect 31109 36347 31175 36348
rect 23289 36274 23355 36277
rect 24945 36274 25011 36277
rect 29177 36274 29243 36277
rect 23289 36272 29243 36274
rect 200 36138 800 36228
rect 23289 36216 23294 36272
rect 23350 36216 24950 36272
rect 25006 36216 29182 36272
rect 29238 36216 29243 36272
rect 23289 36214 29243 36216
rect 23289 36211 23355 36214
rect 24945 36211 25011 36214
rect 29177 36211 29243 36214
rect 2865 36138 2931 36141
rect 200 36136 2931 36138
rect 200 36080 2870 36136
rect 2926 36080 2931 36136
rect 200 36078 2931 36080
rect 200 35988 800 36078
rect 2865 36075 2931 36078
rect 25313 36138 25379 36141
rect 27153 36138 27219 36141
rect 25313 36136 27219 36138
rect 25313 36080 25318 36136
rect 25374 36080 27158 36136
rect 27214 36080 27219 36136
rect 25313 36078 27219 36080
rect 25313 36075 25379 36078
rect 27153 36075 27219 36078
rect 30925 36138 30991 36141
rect 32213 36138 32279 36141
rect 35200 36138 35800 36228
rect 30925 36136 32279 36138
rect 30925 36080 30930 36136
rect 30986 36080 32218 36136
rect 32274 36080 32279 36136
rect 30925 36078 32279 36080
rect 30925 36075 30991 36078
rect 32213 36075 32279 36078
rect 32400 36078 35800 36138
rect 27654 35940 27660 36004
rect 27724 36002 27730 36004
rect 28257 36002 28323 36005
rect 27724 36000 28323 36002
rect 27724 35944 28262 36000
rect 28318 35944 28323 36000
rect 27724 35942 28323 35944
rect 27724 35940 27730 35942
rect 28257 35939 28323 35942
rect 28809 36002 28875 36005
rect 32400 36002 32460 36078
rect 28809 36000 32460 36002
rect 28809 35944 28814 36000
rect 28870 35944 32460 36000
rect 35200 35988 35800 36078
rect 28809 35942 32460 35944
rect 28809 35939 28875 35942
rect 9386 35936 9702 35937
rect 9386 35872 9392 35936
rect 9456 35872 9472 35936
rect 9536 35872 9552 35936
rect 9616 35872 9632 35936
rect 9696 35872 9702 35936
rect 9386 35871 9702 35872
rect 17827 35936 18143 35937
rect 17827 35872 17833 35936
rect 17897 35872 17913 35936
rect 17977 35872 17993 35936
rect 18057 35872 18073 35936
rect 18137 35872 18143 35936
rect 17827 35871 18143 35872
rect 26268 35936 26584 35937
rect 26268 35872 26274 35936
rect 26338 35872 26354 35936
rect 26418 35872 26434 35936
rect 26498 35872 26514 35936
rect 26578 35872 26584 35936
rect 26268 35871 26584 35872
rect 34709 35936 35025 35937
rect 34709 35872 34715 35936
rect 34779 35872 34795 35936
rect 34859 35872 34875 35936
rect 34939 35872 34955 35936
rect 35019 35872 35025 35936
rect 34709 35871 35025 35872
rect 22277 35866 22343 35869
rect 24485 35866 24551 35869
rect 29177 35868 29243 35869
rect 22277 35864 24551 35866
rect 22277 35808 22282 35864
rect 22338 35808 24490 35864
rect 24546 35808 24551 35864
rect 22277 35806 24551 35808
rect 22277 35803 22343 35806
rect 24485 35803 24551 35806
rect 29126 35804 29132 35868
rect 29196 35866 29243 35868
rect 29913 35866 29979 35869
rect 31293 35866 31359 35869
rect 29196 35864 29288 35866
rect 29238 35808 29288 35864
rect 29196 35806 29288 35808
rect 29913 35864 31359 35866
rect 29913 35808 29918 35864
rect 29974 35808 31298 35864
rect 31354 35808 31359 35864
rect 29913 35806 31359 35808
rect 29196 35804 29243 35806
rect 29177 35803 29243 35804
rect 29913 35803 29979 35806
rect 31293 35803 31359 35806
rect 20621 35730 20687 35733
rect 27153 35730 27219 35733
rect 20621 35728 27219 35730
rect 20621 35672 20626 35728
rect 20682 35672 27158 35728
rect 27214 35672 27219 35728
rect 20621 35670 27219 35672
rect 20621 35667 20687 35670
rect 27153 35667 27219 35670
rect 28165 35730 28231 35733
rect 28625 35730 28691 35733
rect 31753 35730 31819 35733
rect 28165 35728 31819 35730
rect 28165 35672 28170 35728
rect 28226 35672 28630 35728
rect 28686 35672 31758 35728
rect 31814 35672 31819 35728
rect 28165 35670 31819 35672
rect 28165 35667 28231 35670
rect 28625 35667 28691 35670
rect 31753 35667 31819 35670
rect 19793 35594 19859 35597
rect 19793 35592 32322 35594
rect 200 35458 800 35548
rect 19793 35536 19798 35592
rect 19854 35536 32322 35592
rect 19793 35534 32322 35536
rect 19793 35531 19859 35534
rect 2773 35458 2839 35461
rect 200 35456 2839 35458
rect 200 35400 2778 35456
rect 2834 35400 2839 35456
rect 200 35398 2839 35400
rect 200 35308 800 35398
rect 2773 35395 2839 35398
rect 30925 35458 30991 35461
rect 31753 35458 31819 35461
rect 32262 35460 32322 35534
rect 30925 35456 31819 35458
rect 30925 35400 30930 35456
rect 30986 35400 31758 35456
rect 31814 35400 31819 35456
rect 30925 35398 31819 35400
rect 30925 35395 30991 35398
rect 31753 35395 31819 35398
rect 32254 35396 32260 35460
rect 32324 35458 32330 35460
rect 32765 35458 32831 35461
rect 32324 35456 32831 35458
rect 32324 35400 32770 35456
rect 32826 35400 32831 35456
rect 32324 35398 32831 35400
rect 32324 35396 32330 35398
rect 32765 35395 32831 35398
rect 5166 35392 5482 35393
rect 5166 35328 5172 35392
rect 5236 35328 5252 35392
rect 5316 35328 5332 35392
rect 5396 35328 5412 35392
rect 5476 35328 5482 35392
rect 5166 35327 5482 35328
rect 13607 35392 13923 35393
rect 13607 35328 13613 35392
rect 13677 35328 13693 35392
rect 13757 35328 13773 35392
rect 13837 35328 13853 35392
rect 13917 35328 13923 35392
rect 13607 35327 13923 35328
rect 22048 35392 22364 35393
rect 22048 35328 22054 35392
rect 22118 35328 22134 35392
rect 22198 35328 22214 35392
rect 22278 35328 22294 35392
rect 22358 35328 22364 35392
rect 22048 35327 22364 35328
rect 30489 35392 30805 35393
rect 30489 35328 30495 35392
rect 30559 35328 30575 35392
rect 30639 35328 30655 35392
rect 30719 35328 30735 35392
rect 30799 35328 30805 35392
rect 30489 35327 30805 35328
rect 19333 35186 19399 35189
rect 27613 35186 27679 35189
rect 19333 35184 27679 35186
rect 19333 35128 19338 35184
rect 19394 35128 27618 35184
rect 27674 35128 27679 35184
rect 19333 35126 27679 35128
rect 19333 35123 19399 35126
rect 27613 35123 27679 35126
rect 28942 35124 28948 35188
rect 29012 35186 29018 35188
rect 32489 35186 32555 35189
rect 29012 35184 32555 35186
rect 29012 35128 32494 35184
rect 32550 35128 32555 35184
rect 29012 35126 32555 35128
rect 29012 35124 29018 35126
rect 32489 35123 32555 35126
rect 21449 35050 21515 35053
rect 22737 35050 22803 35053
rect 21449 35048 22803 35050
rect 21449 34992 21454 35048
rect 21510 34992 22742 35048
rect 22798 34992 22803 35048
rect 21449 34990 22803 34992
rect 21449 34987 21515 34990
rect 22737 34987 22803 34990
rect 24117 35050 24183 35053
rect 29361 35050 29427 35053
rect 24117 35048 29427 35050
rect 24117 34992 24122 35048
rect 24178 34992 29366 35048
rect 29422 34992 29427 35048
rect 24117 34990 29427 34992
rect 24117 34987 24183 34990
rect 29361 34987 29427 34990
rect 200 34628 800 34868
rect 9386 34848 9702 34849
rect 9386 34784 9392 34848
rect 9456 34784 9472 34848
rect 9536 34784 9552 34848
rect 9616 34784 9632 34848
rect 9696 34784 9702 34848
rect 9386 34783 9702 34784
rect 17827 34848 18143 34849
rect 17827 34784 17833 34848
rect 17897 34784 17913 34848
rect 17977 34784 17993 34848
rect 18057 34784 18073 34848
rect 18137 34784 18143 34848
rect 17827 34783 18143 34784
rect 26268 34848 26584 34849
rect 26268 34784 26274 34848
rect 26338 34784 26354 34848
rect 26418 34784 26434 34848
rect 26498 34784 26514 34848
rect 26578 34784 26584 34848
rect 26268 34783 26584 34784
rect 34709 34848 35025 34849
rect 34709 34784 34715 34848
rect 34779 34784 34795 34848
rect 34859 34784 34875 34848
rect 34939 34784 34955 34848
rect 35019 34784 35025 34848
rect 34709 34783 35025 34784
rect 35200 34778 35800 34868
rect 17585 34642 17651 34645
rect 23422 34642 23428 34644
rect 17585 34640 23428 34642
rect 17585 34584 17590 34640
rect 17646 34584 23428 34640
rect 17585 34582 23428 34584
rect 17585 34579 17651 34582
rect 23422 34580 23428 34582
rect 23492 34580 23498 34644
rect 34329 34642 34395 34645
rect 35160 34642 35800 34778
rect 34329 34640 35800 34642
rect 34329 34584 34334 34640
rect 34390 34628 35800 34640
rect 34390 34584 35220 34628
rect 34329 34582 35220 34584
rect 34329 34579 34395 34582
rect 27613 34506 27679 34509
rect 30189 34506 30255 34509
rect 27613 34504 30255 34506
rect 27613 34448 27618 34504
rect 27674 34448 30194 34504
rect 30250 34448 30255 34504
rect 27613 34446 30255 34448
rect 27613 34443 27679 34446
rect 30189 34443 30255 34446
rect 5166 34304 5482 34305
rect 5166 34240 5172 34304
rect 5236 34240 5252 34304
rect 5316 34240 5332 34304
rect 5396 34240 5412 34304
rect 5476 34240 5482 34304
rect 5166 34239 5482 34240
rect 13607 34304 13923 34305
rect 13607 34240 13613 34304
rect 13677 34240 13693 34304
rect 13757 34240 13773 34304
rect 13837 34240 13853 34304
rect 13917 34240 13923 34304
rect 13607 34239 13923 34240
rect 22048 34304 22364 34305
rect 22048 34240 22054 34304
rect 22118 34240 22134 34304
rect 22198 34240 22214 34304
rect 22278 34240 22294 34304
rect 22358 34240 22364 34304
rect 22048 34239 22364 34240
rect 30489 34304 30805 34305
rect 30489 34240 30495 34304
rect 30559 34240 30575 34304
rect 30639 34240 30655 34304
rect 30719 34240 30735 34304
rect 30799 34240 30805 34304
rect 30489 34239 30805 34240
rect 23473 34234 23539 34237
rect 23473 34232 29010 34234
rect 200 34098 800 34188
rect 23473 34176 23478 34232
rect 23534 34176 29010 34232
rect 23473 34174 29010 34176
rect 23473 34171 23539 34174
rect 2773 34098 2839 34101
rect 200 34096 2839 34098
rect 200 34040 2778 34096
rect 2834 34040 2839 34096
rect 200 34038 2839 34040
rect 200 33948 800 34038
rect 2773 34035 2839 34038
rect 24761 34098 24827 34101
rect 28533 34098 28599 34101
rect 24761 34096 28599 34098
rect 24761 34040 24766 34096
rect 24822 34040 28538 34096
rect 28594 34040 28599 34096
rect 24761 34038 28599 34040
rect 28950 34098 29010 34174
rect 32029 34098 32095 34101
rect 28950 34096 32095 34098
rect 28950 34040 32034 34096
rect 32090 34040 32095 34096
rect 28950 34038 32095 34040
rect 24761 34035 24827 34038
rect 28533 34035 28599 34038
rect 32029 34035 32095 34038
rect 34421 34098 34487 34101
rect 35200 34098 35800 34188
rect 34421 34096 35800 34098
rect 34421 34040 34426 34096
rect 34482 34040 35800 34096
rect 34421 34038 35800 34040
rect 34421 34035 34487 34038
rect 21173 33962 21239 33965
rect 21173 33960 31770 33962
rect 21173 33904 21178 33960
rect 21234 33904 31770 33960
rect 35200 33948 35800 34038
rect 21173 33902 31770 33904
rect 21173 33899 21239 33902
rect 31710 33826 31770 33902
rect 33225 33826 33291 33829
rect 31710 33824 33291 33826
rect 31710 33768 33230 33824
rect 33286 33768 33291 33824
rect 31710 33766 33291 33768
rect 33225 33763 33291 33766
rect 9386 33760 9702 33761
rect 9386 33696 9392 33760
rect 9456 33696 9472 33760
rect 9536 33696 9552 33760
rect 9616 33696 9632 33760
rect 9696 33696 9702 33760
rect 9386 33695 9702 33696
rect 17827 33760 18143 33761
rect 17827 33696 17833 33760
rect 17897 33696 17913 33760
rect 17977 33696 17993 33760
rect 18057 33696 18073 33760
rect 18137 33696 18143 33760
rect 17827 33695 18143 33696
rect 26268 33760 26584 33761
rect 26268 33696 26274 33760
rect 26338 33696 26354 33760
rect 26418 33696 26434 33760
rect 26498 33696 26514 33760
rect 26578 33696 26584 33760
rect 26268 33695 26584 33696
rect 34709 33760 35025 33761
rect 34709 33696 34715 33760
rect 34779 33696 34795 33760
rect 34859 33696 34875 33760
rect 34939 33696 34955 33760
rect 35019 33696 35025 33760
rect 34709 33695 35025 33696
rect 19977 33690 20043 33693
rect 21725 33690 21791 33693
rect 19977 33688 21791 33690
rect 19977 33632 19982 33688
rect 20038 33632 21730 33688
rect 21786 33632 21791 33688
rect 19977 33630 21791 33632
rect 19977 33627 20043 33630
rect 21725 33627 21791 33630
rect 31518 33628 31524 33692
rect 31588 33690 31594 33692
rect 31661 33690 31727 33693
rect 31588 33688 31727 33690
rect 31588 33632 31666 33688
rect 31722 33632 31727 33688
rect 31588 33630 31727 33632
rect 31588 33628 31594 33630
rect 31661 33627 31727 33630
rect 21265 33554 21331 33557
rect 23657 33554 23723 33557
rect 26693 33554 26759 33557
rect 21265 33552 26759 33554
rect 21265 33496 21270 33552
rect 21326 33496 23662 33552
rect 23718 33496 26698 33552
rect 26754 33496 26759 33552
rect 21265 33494 26759 33496
rect 21265 33491 21331 33494
rect 23657 33491 23723 33494
rect 26693 33491 26759 33494
rect 28758 33492 28764 33556
rect 28828 33554 28834 33556
rect 31845 33554 31911 33557
rect 28828 33552 31911 33554
rect 28828 33496 31850 33552
rect 31906 33496 31911 33552
rect 28828 33494 31911 33496
rect 28828 33492 28834 33494
rect 31845 33491 31911 33494
rect 34329 33418 34395 33421
rect 35200 33418 35800 33508
rect 34329 33416 35800 33418
rect 34329 33360 34334 33416
rect 34390 33360 35800 33416
rect 34329 33358 35800 33360
rect 34329 33355 34395 33358
rect 27613 33282 27679 33285
rect 28809 33282 28875 33285
rect 27613 33280 28875 33282
rect 27613 33224 27618 33280
rect 27674 33224 28814 33280
rect 28870 33224 28875 33280
rect 35200 33268 35800 33358
rect 27613 33222 28875 33224
rect 27613 33219 27679 33222
rect 28809 33219 28875 33222
rect 5166 33216 5482 33217
rect 5166 33152 5172 33216
rect 5236 33152 5252 33216
rect 5316 33152 5332 33216
rect 5396 33152 5412 33216
rect 5476 33152 5482 33216
rect 5166 33151 5482 33152
rect 13607 33216 13923 33217
rect 13607 33152 13613 33216
rect 13677 33152 13693 33216
rect 13757 33152 13773 33216
rect 13837 33152 13853 33216
rect 13917 33152 13923 33216
rect 13607 33151 13923 33152
rect 22048 33216 22364 33217
rect 22048 33152 22054 33216
rect 22118 33152 22134 33216
rect 22198 33152 22214 33216
rect 22278 33152 22294 33216
rect 22358 33152 22364 33216
rect 22048 33151 22364 33152
rect 30489 33216 30805 33217
rect 30489 33152 30495 33216
rect 30559 33152 30575 33216
rect 30639 33152 30655 33216
rect 30719 33152 30735 33216
rect 30799 33152 30805 33216
rect 30489 33151 30805 33152
rect 28533 33146 28599 33149
rect 28809 33146 28875 33149
rect 28533 33144 28875 33146
rect 28533 33088 28538 33144
rect 28594 33088 28814 33144
rect 28870 33088 28875 33144
rect 28533 33086 28875 33088
rect 28533 33083 28599 33086
rect 28809 33083 28875 33086
rect 19425 33010 19491 33013
rect 20621 33010 20687 33013
rect 19425 33008 20687 33010
rect 19425 32952 19430 33008
rect 19486 32952 20626 33008
rect 20682 32952 20687 33008
rect 19425 32950 20687 32952
rect 19425 32947 19491 32950
rect 20621 32947 20687 32950
rect 25497 32874 25563 32877
rect 29177 32874 29243 32877
rect 25497 32872 29243 32874
rect 200 32588 800 32828
rect 25497 32816 25502 32872
rect 25558 32816 29182 32872
rect 29238 32816 29243 32872
rect 25497 32814 29243 32816
rect 25497 32811 25563 32814
rect 28398 32741 28458 32814
rect 29177 32811 29243 32814
rect 34605 32874 34671 32877
rect 34605 32872 35220 32874
rect 34605 32816 34610 32872
rect 34666 32828 35220 32872
rect 34666 32816 35800 32828
rect 34605 32814 35800 32816
rect 34605 32811 34671 32814
rect 28398 32736 28507 32741
rect 28398 32680 28446 32736
rect 28502 32680 28507 32736
rect 28398 32678 28507 32680
rect 35160 32678 35800 32814
rect 28441 32675 28507 32678
rect 9386 32672 9702 32673
rect 9386 32608 9392 32672
rect 9456 32608 9472 32672
rect 9536 32608 9552 32672
rect 9616 32608 9632 32672
rect 9696 32608 9702 32672
rect 9386 32607 9702 32608
rect 17827 32672 18143 32673
rect 17827 32608 17833 32672
rect 17897 32608 17913 32672
rect 17977 32608 17993 32672
rect 18057 32608 18073 32672
rect 18137 32608 18143 32672
rect 17827 32607 18143 32608
rect 26268 32672 26584 32673
rect 26268 32608 26274 32672
rect 26338 32608 26354 32672
rect 26418 32608 26434 32672
rect 26498 32608 26514 32672
rect 26578 32608 26584 32672
rect 26268 32607 26584 32608
rect 34709 32672 35025 32673
rect 34709 32608 34715 32672
rect 34779 32608 34795 32672
rect 34859 32608 34875 32672
rect 34939 32608 34955 32672
rect 35019 32608 35025 32672
rect 34709 32607 35025 32608
rect 31150 32540 31156 32604
rect 31220 32602 31226 32604
rect 31293 32602 31359 32605
rect 31220 32600 31359 32602
rect 31220 32544 31298 32600
rect 31354 32544 31359 32600
rect 35200 32588 35800 32678
rect 31220 32542 31359 32544
rect 31220 32540 31226 32542
rect 31293 32539 31359 32542
rect 25129 32466 25195 32469
rect 29453 32466 29519 32469
rect 25129 32464 29519 32466
rect 25129 32408 25134 32464
rect 25190 32408 29458 32464
rect 29514 32408 29519 32464
rect 25129 32406 29519 32408
rect 25129 32403 25195 32406
rect 29453 32403 29519 32406
rect 22645 32330 22711 32333
rect 24577 32330 24643 32333
rect 22645 32328 24643 32330
rect 22645 32272 22650 32328
rect 22706 32272 24582 32328
rect 24638 32272 24643 32328
rect 22645 32270 24643 32272
rect 22645 32267 22711 32270
rect 24577 32267 24643 32270
rect 200 32058 800 32148
rect 5166 32128 5482 32129
rect 5166 32064 5172 32128
rect 5236 32064 5252 32128
rect 5316 32064 5332 32128
rect 5396 32064 5412 32128
rect 5476 32064 5482 32128
rect 5166 32063 5482 32064
rect 13607 32128 13923 32129
rect 13607 32064 13613 32128
rect 13677 32064 13693 32128
rect 13757 32064 13773 32128
rect 13837 32064 13853 32128
rect 13917 32064 13923 32128
rect 13607 32063 13923 32064
rect 22048 32128 22364 32129
rect 22048 32064 22054 32128
rect 22118 32064 22134 32128
rect 22198 32064 22214 32128
rect 22278 32064 22294 32128
rect 22358 32064 22364 32128
rect 22048 32063 22364 32064
rect 30489 32128 30805 32129
rect 30489 32064 30495 32128
rect 30559 32064 30575 32128
rect 30639 32064 30655 32128
rect 30719 32064 30735 32128
rect 30799 32064 30805 32128
rect 30489 32063 30805 32064
rect 3509 32058 3575 32061
rect 200 32056 3575 32058
rect 200 32000 3514 32056
rect 3570 32000 3575 32056
rect 200 31998 3575 32000
rect 200 31908 800 31998
rect 3509 31995 3575 31998
rect 34329 32058 34395 32061
rect 35200 32058 35800 32148
rect 34329 32056 35800 32058
rect 34329 32000 34334 32056
rect 34390 32000 35800 32056
rect 34329 31998 35800 32000
rect 34329 31995 34395 31998
rect 22737 31922 22803 31925
rect 22921 31922 22987 31925
rect 22737 31920 22987 31922
rect 22737 31864 22742 31920
rect 22798 31864 22926 31920
rect 22982 31864 22987 31920
rect 22737 31862 22987 31864
rect 22737 31859 22803 31862
rect 22921 31859 22987 31862
rect 25129 31922 25195 31925
rect 25773 31922 25839 31925
rect 25129 31920 25839 31922
rect 25129 31864 25134 31920
rect 25190 31864 25778 31920
rect 25834 31864 25839 31920
rect 25129 31862 25839 31864
rect 25129 31859 25195 31862
rect 25773 31859 25839 31862
rect 28901 31922 28967 31925
rect 32581 31922 32647 31925
rect 28901 31920 32647 31922
rect 28901 31864 28906 31920
rect 28962 31864 32586 31920
rect 32642 31864 32647 31920
rect 35200 31908 35800 31998
rect 28901 31862 32647 31864
rect 28901 31859 28967 31862
rect 32581 31859 32647 31862
rect 24117 31786 24183 31789
rect 30925 31786 30991 31789
rect 24117 31784 30991 31786
rect 24117 31728 24122 31784
rect 24178 31728 30930 31784
rect 30986 31728 30991 31784
rect 24117 31726 30991 31728
rect 24117 31723 24183 31726
rect 30925 31723 30991 31726
rect 27889 31650 27955 31653
rect 28809 31650 28875 31653
rect 27889 31648 28875 31650
rect 27889 31592 27894 31648
rect 27950 31592 28814 31648
rect 28870 31592 28875 31648
rect 27889 31590 28875 31592
rect 27889 31587 27955 31590
rect 28809 31587 28875 31590
rect 9386 31584 9702 31585
rect 9386 31520 9392 31584
rect 9456 31520 9472 31584
rect 9536 31520 9552 31584
rect 9616 31520 9632 31584
rect 9696 31520 9702 31584
rect 9386 31519 9702 31520
rect 17827 31584 18143 31585
rect 17827 31520 17833 31584
rect 17897 31520 17913 31584
rect 17977 31520 17993 31584
rect 18057 31520 18073 31584
rect 18137 31520 18143 31584
rect 17827 31519 18143 31520
rect 26268 31584 26584 31585
rect 26268 31520 26274 31584
rect 26338 31520 26354 31584
rect 26418 31520 26434 31584
rect 26498 31520 26514 31584
rect 26578 31520 26584 31584
rect 26268 31519 26584 31520
rect 34709 31584 35025 31585
rect 34709 31520 34715 31584
rect 34779 31520 34795 31584
rect 34859 31520 34875 31584
rect 34939 31520 34955 31584
rect 35019 31520 35025 31584
rect 34709 31519 35025 31520
rect 29729 31514 29795 31517
rect 32213 31514 32279 31517
rect 29729 31512 32279 31514
rect 200 31378 800 31468
rect 29729 31456 29734 31512
rect 29790 31456 32218 31512
rect 32274 31456 32279 31512
rect 29729 31454 32279 31456
rect 29729 31451 29795 31454
rect 32213 31451 32279 31454
rect 2773 31378 2839 31381
rect 200 31376 2839 31378
rect 200 31320 2778 31376
rect 2834 31320 2839 31376
rect 200 31318 2839 31320
rect 200 31228 800 31318
rect 2773 31315 2839 31318
rect 20621 31378 20687 31381
rect 27613 31378 27679 31381
rect 20621 31376 27679 31378
rect 20621 31320 20626 31376
rect 20682 31320 27618 31376
rect 27674 31320 27679 31376
rect 20621 31318 27679 31320
rect 20621 31315 20687 31318
rect 27613 31315 27679 31318
rect 34329 31378 34395 31381
rect 35200 31378 35800 31468
rect 34329 31376 35800 31378
rect 34329 31320 34334 31376
rect 34390 31320 35800 31376
rect 34329 31318 35800 31320
rect 34329 31315 34395 31318
rect 35200 31228 35800 31318
rect 29453 31108 29519 31109
rect 29453 31106 29500 31108
rect 29408 31104 29500 31106
rect 29408 31048 29458 31104
rect 29408 31046 29500 31048
rect 29453 31044 29500 31046
rect 29564 31044 29570 31108
rect 29453 31043 29519 31044
rect 5166 31040 5482 31041
rect 5166 30976 5172 31040
rect 5236 30976 5252 31040
rect 5316 30976 5332 31040
rect 5396 30976 5412 31040
rect 5476 30976 5482 31040
rect 5166 30975 5482 30976
rect 13607 31040 13923 31041
rect 13607 30976 13613 31040
rect 13677 30976 13693 31040
rect 13757 30976 13773 31040
rect 13837 30976 13853 31040
rect 13917 30976 13923 31040
rect 13607 30975 13923 30976
rect 22048 31040 22364 31041
rect 22048 30976 22054 31040
rect 22118 30976 22134 31040
rect 22198 30976 22214 31040
rect 22278 30976 22294 31040
rect 22358 30976 22364 31040
rect 22048 30975 22364 30976
rect 30489 31040 30805 31041
rect 30489 30976 30495 31040
rect 30559 30976 30575 31040
rect 30639 30976 30655 31040
rect 30719 30976 30735 31040
rect 30799 30976 30805 31040
rect 30489 30975 30805 30976
rect 200 30548 800 30788
rect 29085 30698 29151 30701
rect 31017 30698 31083 30701
rect 29085 30696 31083 30698
rect 29085 30640 29090 30696
rect 29146 30640 31022 30696
rect 31078 30640 31083 30696
rect 29085 30638 31083 30640
rect 29085 30635 29151 30638
rect 31017 30635 31083 30638
rect 35200 30548 35800 30788
rect 9386 30496 9702 30497
rect 9386 30432 9392 30496
rect 9456 30432 9472 30496
rect 9536 30432 9552 30496
rect 9616 30432 9632 30496
rect 9696 30432 9702 30496
rect 9386 30431 9702 30432
rect 17827 30496 18143 30497
rect 17827 30432 17833 30496
rect 17897 30432 17913 30496
rect 17977 30432 17993 30496
rect 18057 30432 18073 30496
rect 18137 30432 18143 30496
rect 17827 30431 18143 30432
rect 26268 30496 26584 30497
rect 26268 30432 26274 30496
rect 26338 30432 26354 30496
rect 26418 30432 26434 30496
rect 26498 30432 26514 30496
rect 26578 30432 26584 30496
rect 26268 30431 26584 30432
rect 34709 30496 35025 30497
rect 34709 30432 34715 30496
rect 34779 30432 34795 30496
rect 34859 30432 34875 30496
rect 34939 30432 34955 30496
rect 35019 30432 35025 30496
rect 34709 30431 35025 30432
rect 19609 30290 19675 30293
rect 21909 30290 21975 30293
rect 19609 30288 21975 30290
rect 19609 30232 19614 30288
rect 19670 30232 21914 30288
rect 21970 30232 21975 30288
rect 19609 30230 21975 30232
rect 19609 30227 19675 30230
rect 21909 30227 21975 30230
rect 19609 30154 19675 30157
rect 28993 30154 29059 30157
rect 19609 30152 29059 30154
rect 200 29868 800 30108
rect 19609 30096 19614 30152
rect 19670 30096 28998 30152
rect 29054 30096 29059 30152
rect 19609 30094 29059 30096
rect 19609 30091 19675 30094
rect 28993 30091 29059 30094
rect 5166 29952 5482 29953
rect 5166 29888 5172 29952
rect 5236 29888 5252 29952
rect 5316 29888 5332 29952
rect 5396 29888 5412 29952
rect 5476 29888 5482 29952
rect 5166 29887 5482 29888
rect 13607 29952 13923 29953
rect 13607 29888 13613 29952
rect 13677 29888 13693 29952
rect 13757 29888 13773 29952
rect 13837 29888 13853 29952
rect 13917 29888 13923 29952
rect 13607 29887 13923 29888
rect 22048 29952 22364 29953
rect 22048 29888 22054 29952
rect 22118 29888 22134 29952
rect 22198 29888 22214 29952
rect 22278 29888 22294 29952
rect 22358 29888 22364 29952
rect 22048 29887 22364 29888
rect 30489 29952 30805 29953
rect 30489 29888 30495 29952
rect 30559 29888 30575 29952
rect 30639 29888 30655 29952
rect 30719 29888 30735 29952
rect 30799 29888 30805 29952
rect 30489 29887 30805 29888
rect 27337 29882 27403 29885
rect 27654 29882 27660 29884
rect 27337 29880 27660 29882
rect 27337 29824 27342 29880
rect 27398 29824 27660 29880
rect 27337 29822 27660 29824
rect 27337 29819 27403 29822
rect 27654 29820 27660 29822
rect 27724 29820 27730 29884
rect 31937 29882 32003 29885
rect 33225 29882 33291 29885
rect 31937 29880 33291 29882
rect 31937 29824 31942 29880
rect 31998 29824 33230 29880
rect 33286 29824 33291 29880
rect 35200 29868 35800 30108
rect 31937 29822 33291 29824
rect 31937 29819 32003 29822
rect 33225 29819 33291 29822
rect 17861 29746 17927 29749
rect 33869 29746 33935 29749
rect 17861 29744 33935 29746
rect 17861 29688 17866 29744
rect 17922 29688 33874 29744
rect 33930 29688 33935 29744
rect 17861 29686 33935 29688
rect 17861 29683 17927 29686
rect 33869 29683 33935 29686
rect 18689 29610 18755 29613
rect 19241 29610 19307 29613
rect 18689 29608 19307 29610
rect 18689 29552 18694 29608
rect 18750 29552 19246 29608
rect 19302 29552 19307 29608
rect 18689 29550 19307 29552
rect 18689 29547 18755 29550
rect 19241 29547 19307 29550
rect 22921 29610 22987 29613
rect 27797 29610 27863 29613
rect 29637 29610 29703 29613
rect 22921 29608 27722 29610
rect 22921 29552 22926 29608
rect 22982 29552 27722 29608
rect 22921 29550 27722 29552
rect 22921 29547 22987 29550
rect 18597 29474 18663 29477
rect 25037 29474 25103 29477
rect 18597 29472 25103 29474
rect 200 29188 800 29428
rect 18597 29416 18602 29472
rect 18658 29416 25042 29472
rect 25098 29416 25103 29472
rect 18597 29414 25103 29416
rect 18597 29411 18663 29414
rect 25037 29411 25103 29414
rect 9386 29408 9702 29409
rect 9386 29344 9392 29408
rect 9456 29344 9472 29408
rect 9536 29344 9552 29408
rect 9616 29344 9632 29408
rect 9696 29344 9702 29408
rect 9386 29343 9702 29344
rect 17827 29408 18143 29409
rect 17827 29344 17833 29408
rect 17897 29344 17913 29408
rect 17977 29344 17993 29408
rect 18057 29344 18073 29408
rect 18137 29344 18143 29408
rect 17827 29343 18143 29344
rect 26268 29408 26584 29409
rect 26268 29344 26274 29408
rect 26338 29344 26354 29408
rect 26418 29344 26434 29408
rect 26498 29344 26514 29408
rect 26578 29344 26584 29408
rect 26268 29343 26584 29344
rect 27662 29338 27722 29550
rect 27797 29608 29703 29610
rect 27797 29552 27802 29608
rect 27858 29552 29642 29608
rect 29698 29552 29703 29608
rect 27797 29550 29703 29552
rect 27797 29547 27863 29550
rect 29637 29547 29703 29550
rect 30230 29548 30236 29612
rect 30300 29610 30306 29612
rect 30833 29610 30899 29613
rect 30300 29608 30899 29610
rect 30300 29552 30838 29608
rect 30894 29552 30899 29608
rect 30300 29550 30899 29552
rect 30300 29548 30306 29550
rect 30833 29547 30899 29550
rect 31753 29610 31819 29613
rect 33317 29610 33383 29613
rect 31753 29608 33383 29610
rect 31753 29552 31758 29608
rect 31814 29552 33322 29608
rect 33378 29552 33383 29608
rect 31753 29550 33383 29552
rect 31753 29547 31819 29550
rect 33317 29547 33383 29550
rect 29269 29474 29335 29477
rect 31569 29474 31635 29477
rect 29269 29472 31635 29474
rect 29269 29416 29274 29472
rect 29330 29416 31574 29472
rect 31630 29416 31635 29472
rect 29269 29414 31635 29416
rect 29269 29411 29335 29414
rect 31569 29411 31635 29414
rect 34709 29408 35025 29409
rect 34709 29344 34715 29408
rect 34779 29344 34795 29408
rect 34859 29344 34875 29408
rect 34939 29344 34955 29408
rect 35019 29344 35025 29408
rect 34709 29343 35025 29344
rect 35200 29338 35800 29428
rect 27662 29278 32644 29338
rect 16849 29202 16915 29205
rect 18321 29202 18387 29205
rect 16849 29200 18387 29202
rect 16849 29144 16854 29200
rect 16910 29144 18326 29200
rect 18382 29144 18387 29200
rect 16849 29142 18387 29144
rect 16849 29139 16915 29142
rect 18321 29139 18387 29142
rect 22001 29202 22067 29205
rect 22461 29202 22527 29205
rect 22001 29200 22527 29202
rect 22001 29144 22006 29200
rect 22062 29144 22466 29200
rect 22522 29144 22527 29200
rect 22001 29142 22527 29144
rect 22001 29139 22067 29142
rect 22461 29139 22527 29142
rect 23473 29202 23539 29205
rect 27705 29202 27771 29205
rect 23473 29200 27771 29202
rect 23473 29144 23478 29200
rect 23534 29144 27710 29200
rect 27766 29144 27771 29200
rect 23473 29142 27771 29144
rect 23473 29139 23539 29142
rect 27705 29139 27771 29142
rect 30925 29202 30991 29205
rect 31845 29202 31911 29205
rect 30925 29200 31911 29202
rect 30925 29144 30930 29200
rect 30986 29144 31850 29200
rect 31906 29144 31911 29200
rect 30925 29142 31911 29144
rect 30925 29139 30991 29142
rect 31845 29139 31911 29142
rect 32254 29140 32260 29204
rect 32324 29202 32330 29204
rect 32397 29202 32463 29205
rect 32324 29200 32463 29202
rect 32324 29144 32402 29200
rect 32458 29144 32463 29200
rect 32324 29142 32463 29144
rect 32584 29202 32644 29278
rect 35160 29202 35800 29338
rect 32584 29188 35800 29202
rect 32584 29142 35220 29188
rect 32324 29140 32330 29142
rect 32397 29139 32463 29142
rect 22277 29066 22343 29069
rect 26877 29066 26943 29069
rect 33409 29066 33475 29069
rect 22277 29064 26943 29066
rect 22277 29008 22282 29064
rect 22338 29008 26882 29064
rect 26938 29008 26943 29064
rect 22277 29006 26943 29008
rect 22277 29003 22343 29006
rect 26877 29003 26943 29006
rect 28950 29064 33475 29066
rect 28950 29008 33414 29064
rect 33470 29008 33475 29064
rect 28950 29006 33475 29008
rect 17585 28930 17651 28933
rect 18965 28930 19031 28933
rect 17585 28928 19031 28930
rect 17585 28872 17590 28928
rect 17646 28872 18970 28928
rect 19026 28872 19031 28928
rect 17585 28870 19031 28872
rect 17585 28867 17651 28870
rect 18965 28867 19031 28870
rect 27797 28930 27863 28933
rect 28950 28930 29010 29006
rect 33409 29003 33475 29006
rect 27797 28928 29010 28930
rect 27797 28872 27802 28928
rect 27858 28872 29010 28928
rect 27797 28870 29010 28872
rect 27797 28867 27863 28870
rect 5166 28864 5482 28865
rect 5166 28800 5172 28864
rect 5236 28800 5252 28864
rect 5316 28800 5332 28864
rect 5396 28800 5412 28864
rect 5476 28800 5482 28864
rect 5166 28799 5482 28800
rect 13607 28864 13923 28865
rect 13607 28800 13613 28864
rect 13677 28800 13693 28864
rect 13757 28800 13773 28864
rect 13837 28800 13853 28864
rect 13917 28800 13923 28864
rect 13607 28799 13923 28800
rect 22048 28864 22364 28865
rect 22048 28800 22054 28864
rect 22118 28800 22134 28864
rect 22198 28800 22214 28864
rect 22278 28800 22294 28864
rect 22358 28800 22364 28864
rect 22048 28799 22364 28800
rect 30489 28864 30805 28865
rect 30489 28800 30495 28864
rect 30559 28800 30575 28864
rect 30639 28800 30655 28864
rect 30719 28800 30735 28864
rect 30799 28800 30805 28864
rect 30489 28799 30805 28800
rect 200 28508 800 28748
rect 18321 28658 18387 28661
rect 18965 28658 19031 28661
rect 18321 28656 19031 28658
rect 18321 28600 18326 28656
rect 18382 28600 18970 28656
rect 19026 28600 19031 28656
rect 18321 28598 19031 28600
rect 18321 28595 18387 28598
rect 18965 28595 19031 28598
rect 23422 28596 23428 28660
rect 23492 28658 23498 28660
rect 32765 28658 32831 28661
rect 23492 28656 32831 28658
rect 23492 28600 32770 28656
rect 32826 28600 32831 28656
rect 23492 28598 32831 28600
rect 23492 28596 23498 28598
rect 32765 28595 32831 28598
rect 16113 28522 16179 28525
rect 23473 28522 23539 28525
rect 16113 28520 23539 28522
rect 16113 28464 16118 28520
rect 16174 28464 23478 28520
rect 23534 28464 23539 28520
rect 16113 28462 23539 28464
rect 16113 28459 16179 28462
rect 23473 28459 23539 28462
rect 27613 28522 27679 28525
rect 32673 28522 32739 28525
rect 27613 28520 32739 28522
rect 27613 28464 27618 28520
rect 27674 28464 32678 28520
rect 32734 28464 32739 28520
rect 27613 28462 32739 28464
rect 27613 28459 27679 28462
rect 32673 28459 32739 28462
rect 28901 28386 28967 28389
rect 32489 28386 32555 28389
rect 28901 28384 32555 28386
rect 28901 28328 28906 28384
rect 28962 28328 32494 28384
rect 32550 28328 32555 28384
rect 28901 28326 32555 28328
rect 28901 28323 28967 28326
rect 32489 28323 32555 28326
rect 9386 28320 9702 28321
rect 9386 28256 9392 28320
rect 9456 28256 9472 28320
rect 9536 28256 9552 28320
rect 9616 28256 9632 28320
rect 9696 28256 9702 28320
rect 9386 28255 9702 28256
rect 17827 28320 18143 28321
rect 17827 28256 17833 28320
rect 17897 28256 17913 28320
rect 17977 28256 17993 28320
rect 18057 28256 18073 28320
rect 18137 28256 18143 28320
rect 17827 28255 18143 28256
rect 26268 28320 26584 28321
rect 26268 28256 26274 28320
rect 26338 28256 26354 28320
rect 26418 28256 26434 28320
rect 26498 28256 26514 28320
rect 26578 28256 26584 28320
rect 26268 28255 26584 28256
rect 34709 28320 35025 28321
rect 34709 28256 34715 28320
rect 34779 28256 34795 28320
rect 34859 28256 34875 28320
rect 34939 28256 34955 28320
rect 35019 28256 35025 28320
rect 34709 28255 35025 28256
rect 29637 28250 29703 28253
rect 31017 28250 31083 28253
rect 29637 28248 31083 28250
rect 29637 28192 29642 28248
rect 29698 28192 31022 28248
rect 31078 28192 31083 28248
rect 29637 28190 31083 28192
rect 29637 28187 29703 28190
rect 31017 28187 31083 28190
rect 20437 28114 20503 28117
rect 24209 28114 24275 28117
rect 29085 28116 29151 28117
rect 29085 28114 29132 28116
rect 20437 28112 24275 28114
rect 200 27828 800 28068
rect 20437 28056 20442 28112
rect 20498 28056 24214 28112
rect 24270 28056 24275 28112
rect 20437 28054 24275 28056
rect 29040 28112 29132 28114
rect 29040 28056 29090 28112
rect 29040 28054 29132 28056
rect 20437 28051 20503 28054
rect 24209 28051 24275 28054
rect 29085 28052 29132 28054
rect 29196 28052 29202 28116
rect 29085 28051 29151 28052
rect 28073 27978 28139 27981
rect 28993 27978 29059 27981
rect 31753 27978 31819 27981
rect 28073 27976 31819 27978
rect 28073 27920 28078 27976
rect 28134 27920 28998 27976
rect 29054 27920 31758 27976
rect 31814 27920 31819 27976
rect 28073 27918 31819 27920
rect 28073 27915 28139 27918
rect 28993 27915 29059 27918
rect 31753 27915 31819 27918
rect 34329 27978 34395 27981
rect 35200 27978 35800 28068
rect 34329 27976 35800 27978
rect 34329 27920 34334 27976
rect 34390 27920 35800 27976
rect 34329 27918 35800 27920
rect 34329 27915 34395 27918
rect 35200 27828 35800 27918
rect 5166 27776 5482 27777
rect 5166 27712 5172 27776
rect 5236 27712 5252 27776
rect 5316 27712 5332 27776
rect 5396 27712 5412 27776
rect 5476 27712 5482 27776
rect 5166 27711 5482 27712
rect 13607 27776 13923 27777
rect 13607 27712 13613 27776
rect 13677 27712 13693 27776
rect 13757 27712 13773 27776
rect 13837 27712 13853 27776
rect 13917 27712 13923 27776
rect 13607 27711 13923 27712
rect 22048 27776 22364 27777
rect 22048 27712 22054 27776
rect 22118 27712 22134 27776
rect 22198 27712 22214 27776
rect 22278 27712 22294 27776
rect 22358 27712 22364 27776
rect 22048 27711 22364 27712
rect 30489 27776 30805 27777
rect 30489 27712 30495 27776
rect 30559 27712 30575 27776
rect 30639 27712 30655 27776
rect 30719 27712 30735 27776
rect 30799 27712 30805 27776
rect 30489 27711 30805 27712
rect 28809 27706 28875 27709
rect 29637 27706 29703 27709
rect 28809 27704 29703 27706
rect 28809 27648 28814 27704
rect 28870 27648 29642 27704
rect 29698 27648 29703 27704
rect 28809 27646 29703 27648
rect 28809 27643 28875 27646
rect 29637 27643 29703 27646
rect 18689 27570 18755 27573
rect 30925 27570 30991 27573
rect 32029 27572 32095 27573
rect 32029 27570 32076 27572
rect 18689 27568 32076 27570
rect 18689 27512 18694 27568
rect 18750 27512 30930 27568
rect 30986 27512 32034 27568
rect 18689 27510 32076 27512
rect 18689 27507 18755 27510
rect 30925 27507 30991 27510
rect 32029 27508 32076 27510
rect 32140 27508 32146 27572
rect 32029 27507 32095 27508
rect 200 27148 800 27388
rect 9386 27232 9702 27233
rect 9386 27168 9392 27232
rect 9456 27168 9472 27232
rect 9536 27168 9552 27232
rect 9616 27168 9632 27232
rect 9696 27168 9702 27232
rect 9386 27167 9702 27168
rect 17827 27232 18143 27233
rect 17827 27168 17833 27232
rect 17897 27168 17913 27232
rect 17977 27168 17993 27232
rect 18057 27168 18073 27232
rect 18137 27168 18143 27232
rect 17827 27167 18143 27168
rect 26268 27232 26584 27233
rect 26268 27168 26274 27232
rect 26338 27168 26354 27232
rect 26418 27168 26434 27232
rect 26498 27168 26514 27232
rect 26578 27168 26584 27232
rect 26268 27167 26584 27168
rect 34709 27232 35025 27233
rect 34709 27168 34715 27232
rect 34779 27168 34795 27232
rect 34859 27168 34875 27232
rect 34939 27168 34955 27232
rect 35019 27168 35025 27232
rect 34709 27167 35025 27168
rect 35200 27148 35800 27388
rect 19057 26890 19123 26893
rect 26325 26890 26391 26893
rect 19057 26888 26391 26890
rect 19057 26832 19062 26888
rect 19118 26832 26330 26888
rect 26386 26832 26391 26888
rect 19057 26830 26391 26832
rect 19057 26827 19123 26830
rect 26325 26827 26391 26830
rect 5166 26688 5482 26689
rect 5166 26624 5172 26688
rect 5236 26624 5252 26688
rect 5316 26624 5332 26688
rect 5396 26624 5412 26688
rect 5476 26624 5482 26688
rect 5166 26623 5482 26624
rect 13607 26688 13923 26689
rect 13607 26624 13613 26688
rect 13677 26624 13693 26688
rect 13757 26624 13773 26688
rect 13837 26624 13853 26688
rect 13917 26624 13923 26688
rect 13607 26623 13923 26624
rect 22048 26688 22364 26689
rect 22048 26624 22054 26688
rect 22118 26624 22134 26688
rect 22198 26624 22214 26688
rect 22278 26624 22294 26688
rect 22358 26624 22364 26688
rect 22048 26623 22364 26624
rect 30489 26688 30805 26689
rect 30489 26624 30495 26688
rect 30559 26624 30575 26688
rect 30639 26624 30655 26688
rect 30719 26624 30735 26688
rect 30799 26624 30805 26688
rect 30489 26623 30805 26624
rect 18965 26482 19031 26485
rect 18965 26480 27630 26482
rect 18965 26424 18970 26480
rect 19026 26424 27630 26480
rect 35200 26468 35800 26708
rect 18965 26422 27630 26424
rect 18965 26419 19031 26422
rect 19241 26346 19307 26349
rect 23381 26346 23447 26349
rect 19241 26344 23447 26346
rect 19241 26288 19246 26344
rect 19302 26288 23386 26344
rect 23442 26288 23447 26344
rect 19241 26286 23447 26288
rect 27570 26346 27630 26422
rect 31293 26346 31359 26349
rect 27570 26344 31359 26346
rect 27570 26288 31298 26344
rect 31354 26288 31359 26344
rect 27570 26286 31359 26288
rect 19241 26283 19307 26286
rect 23381 26283 23447 26286
rect 31293 26283 31359 26286
rect 9386 26144 9702 26145
rect 9386 26080 9392 26144
rect 9456 26080 9472 26144
rect 9536 26080 9552 26144
rect 9616 26080 9632 26144
rect 9696 26080 9702 26144
rect 9386 26079 9702 26080
rect 17827 26144 18143 26145
rect 17827 26080 17833 26144
rect 17897 26080 17913 26144
rect 17977 26080 17993 26144
rect 18057 26080 18073 26144
rect 18137 26080 18143 26144
rect 17827 26079 18143 26080
rect 26268 26144 26584 26145
rect 26268 26080 26274 26144
rect 26338 26080 26354 26144
rect 26418 26080 26434 26144
rect 26498 26080 26514 26144
rect 26578 26080 26584 26144
rect 26268 26079 26584 26080
rect 34709 26144 35025 26145
rect 34709 26080 34715 26144
rect 34779 26080 34795 26144
rect 34859 26080 34875 26144
rect 34939 26080 34955 26144
rect 35019 26080 35025 26144
rect 34709 26079 35025 26080
rect 200 25788 800 26028
rect 20069 25938 20135 25941
rect 24945 25938 25011 25941
rect 25957 25938 26023 25941
rect 28165 25938 28231 25941
rect 20069 25936 28231 25938
rect 20069 25880 20074 25936
rect 20130 25880 24950 25936
rect 25006 25880 25962 25936
rect 26018 25880 28170 25936
rect 28226 25880 28231 25936
rect 20069 25878 28231 25880
rect 20069 25875 20135 25878
rect 24945 25875 25011 25878
rect 25957 25875 26023 25878
rect 28165 25875 28231 25878
rect 34329 25938 34395 25941
rect 35200 25938 35800 26028
rect 34329 25936 35800 25938
rect 34329 25880 34334 25936
rect 34390 25880 35800 25936
rect 34329 25878 35800 25880
rect 34329 25875 34395 25878
rect 25773 25802 25839 25805
rect 27429 25802 27495 25805
rect 25773 25800 27495 25802
rect 25773 25744 25778 25800
rect 25834 25744 27434 25800
rect 27490 25744 27495 25800
rect 35200 25788 35800 25878
rect 25773 25742 27495 25744
rect 25773 25739 25839 25742
rect 27429 25739 27495 25742
rect 25681 25666 25747 25669
rect 27429 25666 27495 25669
rect 25681 25664 27495 25666
rect 25681 25608 25686 25664
rect 25742 25608 27434 25664
rect 27490 25608 27495 25664
rect 25681 25606 27495 25608
rect 25681 25603 25747 25606
rect 27429 25603 27495 25606
rect 5166 25600 5482 25601
rect 5166 25536 5172 25600
rect 5236 25536 5252 25600
rect 5316 25536 5332 25600
rect 5396 25536 5412 25600
rect 5476 25536 5482 25600
rect 5166 25535 5482 25536
rect 13607 25600 13923 25601
rect 13607 25536 13613 25600
rect 13677 25536 13693 25600
rect 13757 25536 13773 25600
rect 13837 25536 13853 25600
rect 13917 25536 13923 25600
rect 13607 25535 13923 25536
rect 22048 25600 22364 25601
rect 22048 25536 22054 25600
rect 22118 25536 22134 25600
rect 22198 25536 22214 25600
rect 22278 25536 22294 25600
rect 22358 25536 22364 25600
rect 22048 25535 22364 25536
rect 30489 25600 30805 25601
rect 30489 25536 30495 25600
rect 30559 25536 30575 25600
rect 30639 25536 30655 25600
rect 30719 25536 30735 25600
rect 30799 25536 30805 25600
rect 30489 25535 30805 25536
rect 27337 25530 27403 25533
rect 32029 25530 32095 25533
rect 22510 25528 27403 25530
rect 22510 25472 27342 25528
rect 27398 25472 27403 25528
rect 22510 25470 27403 25472
rect 20621 25394 20687 25397
rect 22510 25394 22570 25470
rect 27337 25467 27403 25470
rect 30928 25528 32095 25530
rect 30928 25472 32034 25528
rect 32090 25472 32095 25528
rect 30928 25470 32095 25472
rect 20621 25392 22570 25394
rect 200 25258 800 25348
rect 20621 25336 20626 25392
rect 20682 25336 22570 25392
rect 20621 25334 22570 25336
rect 26509 25394 26575 25397
rect 26877 25394 26943 25397
rect 26509 25392 26943 25394
rect 26509 25336 26514 25392
rect 26570 25336 26882 25392
rect 26938 25336 26943 25392
rect 26509 25334 26943 25336
rect 20621 25331 20687 25334
rect 26509 25331 26575 25334
rect 26877 25331 26943 25334
rect 28993 25394 29059 25397
rect 30928 25394 30988 25470
rect 32029 25467 32095 25470
rect 28993 25392 30988 25394
rect 28993 25336 28998 25392
rect 29054 25336 30988 25392
rect 28993 25334 30988 25336
rect 31109 25394 31175 25397
rect 33317 25394 33383 25397
rect 31109 25392 33383 25394
rect 31109 25336 31114 25392
rect 31170 25336 33322 25392
rect 33378 25336 33383 25392
rect 31109 25334 33383 25336
rect 28993 25331 29059 25334
rect 31109 25331 31175 25334
rect 33317 25331 33383 25334
rect 2773 25258 2839 25261
rect 200 25256 2839 25258
rect 200 25200 2778 25256
rect 2834 25200 2839 25256
rect 200 25198 2839 25200
rect 200 25108 800 25198
rect 2773 25195 2839 25198
rect 18045 25258 18111 25261
rect 26417 25258 26483 25261
rect 18045 25256 26483 25258
rect 18045 25200 18050 25256
rect 18106 25200 26422 25256
rect 26478 25200 26483 25256
rect 18045 25198 26483 25200
rect 18045 25195 18111 25198
rect 26417 25195 26483 25198
rect 31569 25258 31635 25261
rect 33593 25258 33659 25261
rect 31569 25256 33659 25258
rect 31569 25200 31574 25256
rect 31630 25200 33598 25256
rect 33654 25200 33659 25256
rect 31569 25198 33659 25200
rect 31569 25195 31635 25198
rect 33593 25195 33659 25198
rect 34329 25258 34395 25261
rect 35200 25258 35800 25348
rect 34329 25256 35800 25258
rect 34329 25200 34334 25256
rect 34390 25200 35800 25256
rect 34329 25198 35800 25200
rect 34329 25195 34395 25198
rect 31569 25122 31635 25125
rect 32029 25122 32095 25125
rect 31569 25120 32095 25122
rect 31569 25064 31574 25120
rect 31630 25064 32034 25120
rect 32090 25064 32095 25120
rect 35200 25108 35800 25198
rect 31569 25062 32095 25064
rect 31569 25059 31635 25062
rect 32029 25059 32095 25062
rect 9386 25056 9702 25057
rect 9386 24992 9392 25056
rect 9456 24992 9472 25056
rect 9536 24992 9552 25056
rect 9616 24992 9632 25056
rect 9696 24992 9702 25056
rect 9386 24991 9702 24992
rect 17827 25056 18143 25057
rect 17827 24992 17833 25056
rect 17897 24992 17913 25056
rect 17977 24992 17993 25056
rect 18057 24992 18073 25056
rect 18137 24992 18143 25056
rect 17827 24991 18143 24992
rect 26268 25056 26584 25057
rect 26268 24992 26274 25056
rect 26338 24992 26354 25056
rect 26418 24992 26434 25056
rect 26498 24992 26514 25056
rect 26578 24992 26584 25056
rect 26268 24991 26584 24992
rect 34709 25056 35025 25057
rect 34709 24992 34715 25056
rect 34779 24992 34795 25056
rect 34859 24992 34875 25056
rect 34939 24992 34955 25056
rect 35019 24992 35025 25056
rect 34709 24991 35025 24992
rect 21173 24986 21239 24989
rect 24393 24986 24459 24989
rect 21173 24984 24459 24986
rect 21173 24928 21178 24984
rect 21234 24928 24398 24984
rect 24454 24928 24459 24984
rect 21173 24926 24459 24928
rect 21173 24923 21239 24926
rect 24393 24923 24459 24926
rect 31477 24988 31543 24989
rect 31477 24984 31524 24988
rect 31588 24986 31594 24988
rect 31477 24928 31482 24984
rect 31477 24924 31524 24928
rect 31588 24926 31634 24986
rect 31588 24924 31594 24926
rect 31477 24923 31543 24924
rect 19333 24850 19399 24853
rect 27521 24850 27587 24853
rect 19333 24848 27587 24850
rect 19333 24792 19338 24848
rect 19394 24792 27526 24848
rect 27582 24792 27587 24848
rect 19333 24790 27587 24792
rect 19333 24787 19399 24790
rect 27521 24787 27587 24790
rect 200 24428 800 24668
rect 31334 24652 31340 24716
rect 31404 24714 31410 24716
rect 31753 24714 31819 24717
rect 31404 24712 31819 24714
rect 31404 24656 31758 24712
rect 31814 24656 31819 24712
rect 31404 24654 31819 24656
rect 31404 24652 31410 24654
rect 31753 24651 31819 24654
rect 32673 24714 32739 24717
rect 32806 24714 32812 24716
rect 32673 24712 32812 24714
rect 32673 24656 32678 24712
rect 32734 24656 32812 24712
rect 32673 24654 32812 24656
rect 32673 24651 32739 24654
rect 32806 24652 32812 24654
rect 32876 24652 32882 24716
rect 34421 24578 34487 24581
rect 35200 24578 35800 24668
rect 34421 24576 35800 24578
rect 34421 24520 34426 24576
rect 34482 24520 35800 24576
rect 34421 24518 35800 24520
rect 34421 24515 34487 24518
rect 5166 24512 5482 24513
rect 5166 24448 5172 24512
rect 5236 24448 5252 24512
rect 5316 24448 5332 24512
rect 5396 24448 5412 24512
rect 5476 24448 5482 24512
rect 5166 24447 5482 24448
rect 13607 24512 13923 24513
rect 13607 24448 13613 24512
rect 13677 24448 13693 24512
rect 13757 24448 13773 24512
rect 13837 24448 13853 24512
rect 13917 24448 13923 24512
rect 13607 24447 13923 24448
rect 22048 24512 22364 24513
rect 22048 24448 22054 24512
rect 22118 24448 22134 24512
rect 22198 24448 22214 24512
rect 22278 24448 22294 24512
rect 22358 24448 22364 24512
rect 22048 24447 22364 24448
rect 30489 24512 30805 24513
rect 30489 24448 30495 24512
rect 30559 24448 30575 24512
rect 30639 24448 30655 24512
rect 30719 24448 30735 24512
rect 30799 24448 30805 24512
rect 30489 24447 30805 24448
rect 35200 24428 35800 24518
rect 22277 24306 22343 24309
rect 24577 24306 24643 24309
rect 22277 24304 24643 24306
rect 22277 24248 22282 24304
rect 22338 24248 24582 24304
rect 24638 24248 24643 24304
rect 22277 24246 24643 24248
rect 22277 24243 22343 24246
rect 24577 24243 24643 24246
rect 15745 24170 15811 24173
rect 17125 24170 17191 24173
rect 15745 24168 17191 24170
rect 15745 24112 15750 24168
rect 15806 24112 17130 24168
rect 17186 24112 17191 24168
rect 15745 24110 17191 24112
rect 15745 24107 15811 24110
rect 17125 24107 17191 24110
rect 200 23748 800 23988
rect 9386 23968 9702 23969
rect 9386 23904 9392 23968
rect 9456 23904 9472 23968
rect 9536 23904 9552 23968
rect 9616 23904 9632 23968
rect 9696 23904 9702 23968
rect 9386 23903 9702 23904
rect 17827 23968 18143 23969
rect 17827 23904 17833 23968
rect 17897 23904 17913 23968
rect 17977 23904 17993 23968
rect 18057 23904 18073 23968
rect 18137 23904 18143 23968
rect 17827 23903 18143 23904
rect 26268 23968 26584 23969
rect 26268 23904 26274 23968
rect 26338 23904 26354 23968
rect 26418 23904 26434 23968
rect 26498 23904 26514 23968
rect 26578 23904 26584 23968
rect 26268 23903 26584 23904
rect 34709 23968 35025 23969
rect 34709 23904 34715 23968
rect 34779 23904 34795 23968
rect 34859 23904 34875 23968
rect 34939 23904 34955 23968
rect 35019 23904 35025 23968
rect 34709 23903 35025 23904
rect 32489 23898 32555 23901
rect 33726 23898 33732 23900
rect 32489 23896 33732 23898
rect 32489 23840 32494 23896
rect 32550 23840 33732 23896
rect 32489 23838 33732 23840
rect 32489 23835 32555 23838
rect 33726 23836 33732 23838
rect 33796 23836 33802 23900
rect 35200 23898 35800 23988
rect 17953 23762 18019 23765
rect 19241 23762 19307 23765
rect 17953 23760 19307 23762
rect 17953 23704 17958 23760
rect 18014 23704 19246 23760
rect 19302 23704 19307 23760
rect 17953 23702 19307 23704
rect 17953 23699 18019 23702
rect 19241 23699 19307 23702
rect 31886 23700 31892 23764
rect 31956 23762 31962 23764
rect 32673 23762 32739 23765
rect 31956 23760 32739 23762
rect 31956 23704 32678 23760
rect 32734 23704 32739 23760
rect 31956 23702 32739 23704
rect 31956 23700 31962 23702
rect 32673 23699 32739 23702
rect 34329 23762 34395 23765
rect 35160 23762 35800 23898
rect 34329 23760 35800 23762
rect 34329 23704 34334 23760
rect 34390 23748 35800 23760
rect 34390 23704 35220 23748
rect 34329 23702 35220 23704
rect 34329 23699 34395 23702
rect 29494 23564 29500 23628
rect 29564 23626 29570 23628
rect 32673 23626 32739 23629
rect 29564 23624 32739 23626
rect 29564 23568 32678 23624
rect 32734 23568 32739 23624
rect 29564 23566 32739 23568
rect 29564 23564 29570 23566
rect 32673 23563 32739 23566
rect 22829 23490 22895 23493
rect 26734 23490 26740 23492
rect 22829 23488 26740 23490
rect 22829 23432 22834 23488
rect 22890 23432 26740 23488
rect 22829 23430 26740 23432
rect 22829 23427 22895 23430
rect 26734 23428 26740 23430
rect 26804 23428 26810 23492
rect 32489 23490 32555 23493
rect 33910 23490 33916 23492
rect 32489 23488 33916 23490
rect 32489 23432 32494 23488
rect 32550 23432 33916 23488
rect 32489 23430 33916 23432
rect 32489 23427 32555 23430
rect 33910 23428 33916 23430
rect 33980 23428 33986 23492
rect 5166 23424 5482 23425
rect 5166 23360 5172 23424
rect 5236 23360 5252 23424
rect 5316 23360 5332 23424
rect 5396 23360 5412 23424
rect 5476 23360 5482 23424
rect 5166 23359 5482 23360
rect 13607 23424 13923 23425
rect 13607 23360 13613 23424
rect 13677 23360 13693 23424
rect 13757 23360 13773 23424
rect 13837 23360 13853 23424
rect 13917 23360 13923 23424
rect 13607 23359 13923 23360
rect 22048 23424 22364 23425
rect 22048 23360 22054 23424
rect 22118 23360 22134 23424
rect 22198 23360 22214 23424
rect 22278 23360 22294 23424
rect 22358 23360 22364 23424
rect 22048 23359 22364 23360
rect 30489 23424 30805 23425
rect 30489 23360 30495 23424
rect 30559 23360 30575 23424
rect 30639 23360 30655 23424
rect 30719 23360 30735 23424
rect 30799 23360 30805 23424
rect 30489 23359 30805 23360
rect 200 23068 800 23308
rect 34329 23218 34395 23221
rect 35200 23218 35800 23308
rect 34329 23216 35800 23218
rect 34329 23160 34334 23216
rect 34390 23160 35800 23216
rect 34329 23158 35800 23160
rect 34329 23155 34395 23158
rect 27613 23082 27679 23085
rect 28809 23082 28875 23085
rect 27613 23080 28875 23082
rect 27613 23024 27618 23080
rect 27674 23024 28814 23080
rect 28870 23024 28875 23080
rect 35200 23068 35800 23158
rect 27613 23022 28875 23024
rect 27613 23019 27679 23022
rect 28809 23019 28875 23022
rect 9386 22880 9702 22881
rect 9386 22816 9392 22880
rect 9456 22816 9472 22880
rect 9536 22816 9552 22880
rect 9616 22816 9632 22880
rect 9696 22816 9702 22880
rect 9386 22815 9702 22816
rect 17827 22880 18143 22881
rect 17827 22816 17833 22880
rect 17897 22816 17913 22880
rect 17977 22816 17993 22880
rect 18057 22816 18073 22880
rect 18137 22816 18143 22880
rect 17827 22815 18143 22816
rect 26268 22880 26584 22881
rect 26268 22816 26274 22880
rect 26338 22816 26354 22880
rect 26418 22816 26434 22880
rect 26498 22816 26514 22880
rect 26578 22816 26584 22880
rect 26268 22815 26584 22816
rect 34709 22880 35025 22881
rect 34709 22816 34715 22880
rect 34779 22816 34795 22880
rect 34859 22816 34875 22880
rect 34939 22816 34955 22880
rect 35019 22816 35025 22880
rect 34709 22815 35025 22816
rect 28993 22810 29059 22813
rect 34329 22810 34395 22813
rect 28993 22808 34395 22810
rect 28993 22752 28998 22808
rect 29054 22752 34334 22808
rect 34390 22752 34395 22808
rect 28993 22750 34395 22752
rect 28993 22747 29059 22750
rect 34329 22747 34395 22750
rect 32489 22674 32555 22677
rect 34094 22674 34100 22676
rect 32489 22672 34100 22674
rect 200 22388 800 22628
rect 32489 22616 32494 22672
rect 32550 22616 34100 22672
rect 32489 22614 34100 22616
rect 32489 22611 32555 22614
rect 34094 22612 34100 22614
rect 34164 22612 34170 22676
rect 35200 22388 35800 22628
rect 5166 22336 5482 22337
rect 5166 22272 5172 22336
rect 5236 22272 5252 22336
rect 5316 22272 5332 22336
rect 5396 22272 5412 22336
rect 5476 22272 5482 22336
rect 5166 22271 5482 22272
rect 13607 22336 13923 22337
rect 13607 22272 13613 22336
rect 13677 22272 13693 22336
rect 13757 22272 13773 22336
rect 13837 22272 13853 22336
rect 13917 22272 13923 22336
rect 13607 22271 13923 22272
rect 22048 22336 22364 22337
rect 22048 22272 22054 22336
rect 22118 22272 22134 22336
rect 22198 22272 22214 22336
rect 22278 22272 22294 22336
rect 22358 22272 22364 22336
rect 22048 22271 22364 22272
rect 30489 22336 30805 22337
rect 30489 22272 30495 22336
rect 30559 22272 30575 22336
rect 30639 22272 30655 22336
rect 30719 22272 30735 22336
rect 30799 22272 30805 22336
rect 30489 22271 30805 22272
rect 28717 22266 28783 22269
rect 29678 22266 29684 22268
rect 28717 22264 29684 22266
rect 28717 22208 28722 22264
rect 28778 22208 29684 22264
rect 28717 22206 29684 22208
rect 28717 22203 28783 22206
rect 29678 22204 29684 22206
rect 29748 22204 29754 22268
rect 20529 21994 20595 21997
rect 25129 21994 25195 21997
rect 20529 21992 25195 21994
rect 200 21708 800 21948
rect 20529 21936 20534 21992
rect 20590 21936 25134 21992
rect 25190 21936 25195 21992
rect 20529 21934 25195 21936
rect 20529 21931 20595 21934
rect 25129 21931 25195 21934
rect 28993 21858 29059 21861
rect 29126 21858 29132 21860
rect 28993 21856 29132 21858
rect 28993 21800 28998 21856
rect 29054 21800 29132 21856
rect 28993 21798 29132 21800
rect 28993 21795 29059 21798
rect 29126 21796 29132 21798
rect 29196 21796 29202 21860
rect 9386 21792 9702 21793
rect 9386 21728 9392 21792
rect 9456 21728 9472 21792
rect 9536 21728 9552 21792
rect 9616 21728 9632 21792
rect 9696 21728 9702 21792
rect 9386 21727 9702 21728
rect 17827 21792 18143 21793
rect 17827 21728 17833 21792
rect 17897 21728 17913 21792
rect 17977 21728 17993 21792
rect 18057 21728 18073 21792
rect 18137 21728 18143 21792
rect 17827 21727 18143 21728
rect 26268 21792 26584 21793
rect 26268 21728 26274 21792
rect 26338 21728 26354 21792
rect 26418 21728 26434 21792
rect 26498 21728 26514 21792
rect 26578 21728 26584 21792
rect 26268 21727 26584 21728
rect 34709 21792 35025 21793
rect 34709 21728 34715 21792
rect 34779 21728 34795 21792
rect 34859 21728 34875 21792
rect 34939 21728 34955 21792
rect 35019 21728 35025 21792
rect 34709 21727 35025 21728
rect 20989 21586 21055 21589
rect 23289 21586 23355 21589
rect 20989 21584 23355 21586
rect 20989 21528 20994 21584
rect 21050 21528 23294 21584
rect 23350 21528 23355 21584
rect 20989 21526 23355 21528
rect 20989 21523 21055 21526
rect 23289 21523 23355 21526
rect 21357 21450 21423 21453
rect 22001 21450 22067 21453
rect 21357 21448 22067 21450
rect 21357 21392 21362 21448
rect 21418 21392 22006 21448
rect 22062 21392 22067 21448
rect 21357 21390 22067 21392
rect 21357 21387 21423 21390
rect 22001 21387 22067 21390
rect 200 21028 800 21268
rect 5166 21248 5482 21249
rect 5166 21184 5172 21248
rect 5236 21184 5252 21248
rect 5316 21184 5332 21248
rect 5396 21184 5412 21248
rect 5476 21184 5482 21248
rect 5166 21183 5482 21184
rect 13607 21248 13923 21249
rect 13607 21184 13613 21248
rect 13677 21184 13693 21248
rect 13757 21184 13773 21248
rect 13837 21184 13853 21248
rect 13917 21184 13923 21248
rect 13607 21183 13923 21184
rect 22048 21248 22364 21249
rect 22048 21184 22054 21248
rect 22118 21184 22134 21248
rect 22198 21184 22214 21248
rect 22278 21184 22294 21248
rect 22358 21184 22364 21248
rect 22048 21183 22364 21184
rect 30489 21248 30805 21249
rect 30489 21184 30495 21248
rect 30559 21184 30575 21248
rect 30639 21184 30655 21248
rect 30719 21184 30735 21248
rect 30799 21184 30805 21248
rect 30489 21183 30805 21184
rect 33041 21178 33107 21181
rect 35200 21178 35800 21268
rect 33041 21176 35800 21178
rect 33041 21120 33046 21176
rect 33102 21120 35800 21176
rect 33041 21118 35800 21120
rect 33041 21115 33107 21118
rect 30465 21042 30531 21045
rect 31569 21042 31635 21045
rect 30465 21040 31635 21042
rect 30465 20984 30470 21040
rect 30526 20984 31574 21040
rect 31630 20984 31635 21040
rect 35200 21028 35800 21118
rect 30465 20982 31635 20984
rect 30465 20979 30531 20982
rect 31569 20979 31635 20982
rect 22093 20906 22159 20909
rect 24209 20906 24275 20909
rect 22093 20904 24275 20906
rect 22093 20848 22098 20904
rect 22154 20848 24214 20904
rect 24270 20848 24275 20904
rect 22093 20846 24275 20848
rect 22093 20843 22159 20846
rect 24209 20843 24275 20846
rect 31845 20906 31911 20909
rect 32254 20906 32260 20908
rect 31845 20904 32260 20906
rect 31845 20848 31850 20904
rect 31906 20848 32260 20904
rect 31845 20846 32260 20848
rect 31845 20843 31911 20846
rect 32254 20844 32260 20846
rect 32324 20844 32330 20908
rect 25681 20772 25747 20773
rect 25630 20770 25636 20772
rect 25590 20710 25636 20770
rect 25700 20768 25747 20772
rect 25742 20712 25747 20768
rect 25630 20708 25636 20710
rect 25700 20708 25747 20712
rect 25681 20707 25747 20708
rect 30373 20770 30439 20773
rect 30966 20770 30972 20772
rect 30373 20768 30972 20770
rect 30373 20712 30378 20768
rect 30434 20712 30972 20768
rect 30373 20710 30972 20712
rect 30373 20707 30439 20710
rect 30966 20708 30972 20710
rect 31036 20708 31042 20772
rect 31150 20708 31156 20772
rect 31220 20770 31226 20772
rect 32673 20770 32739 20773
rect 31220 20768 32739 20770
rect 31220 20712 32678 20768
rect 32734 20712 32739 20768
rect 31220 20710 32739 20712
rect 31220 20708 31226 20710
rect 32673 20707 32739 20710
rect 9386 20704 9702 20705
rect 9386 20640 9392 20704
rect 9456 20640 9472 20704
rect 9536 20640 9552 20704
rect 9616 20640 9632 20704
rect 9696 20640 9702 20704
rect 9386 20639 9702 20640
rect 17827 20704 18143 20705
rect 17827 20640 17833 20704
rect 17897 20640 17913 20704
rect 17977 20640 17993 20704
rect 18057 20640 18073 20704
rect 18137 20640 18143 20704
rect 17827 20639 18143 20640
rect 26268 20704 26584 20705
rect 26268 20640 26274 20704
rect 26338 20640 26354 20704
rect 26418 20640 26434 20704
rect 26498 20640 26514 20704
rect 26578 20640 26584 20704
rect 26268 20639 26584 20640
rect 34709 20704 35025 20705
rect 34709 20640 34715 20704
rect 34779 20640 34795 20704
rect 34859 20640 34875 20704
rect 34939 20640 34955 20704
rect 35019 20640 35025 20704
rect 34709 20639 35025 20640
rect 29729 20634 29795 20637
rect 34237 20634 34303 20637
rect 29729 20632 34303 20634
rect 200 20348 800 20588
rect 29729 20576 29734 20632
rect 29790 20576 34242 20632
rect 34298 20576 34303 20632
rect 29729 20574 34303 20576
rect 29729 20571 29795 20574
rect 34237 20571 34303 20574
rect 34329 20498 34395 20501
rect 35200 20498 35800 20588
rect 34329 20496 35800 20498
rect 34329 20440 34334 20496
rect 34390 20440 35800 20496
rect 34329 20438 35800 20440
rect 34329 20435 34395 20438
rect 35200 20348 35800 20438
rect 5166 20160 5482 20161
rect 5166 20096 5172 20160
rect 5236 20096 5252 20160
rect 5316 20096 5332 20160
rect 5396 20096 5412 20160
rect 5476 20096 5482 20160
rect 5166 20095 5482 20096
rect 13607 20160 13923 20161
rect 13607 20096 13613 20160
rect 13677 20096 13693 20160
rect 13757 20096 13773 20160
rect 13837 20096 13853 20160
rect 13917 20096 13923 20160
rect 13607 20095 13923 20096
rect 22048 20160 22364 20161
rect 22048 20096 22054 20160
rect 22118 20096 22134 20160
rect 22198 20096 22214 20160
rect 22278 20096 22294 20160
rect 22358 20096 22364 20160
rect 22048 20095 22364 20096
rect 30489 20160 30805 20161
rect 30489 20096 30495 20160
rect 30559 20096 30575 20160
rect 30639 20096 30655 20160
rect 30719 20096 30735 20160
rect 30799 20096 30805 20160
rect 30489 20095 30805 20096
rect 34329 19818 34395 19821
rect 35200 19818 35800 19908
rect 34329 19816 35800 19818
rect 34329 19760 34334 19816
rect 34390 19760 35800 19816
rect 34329 19758 35800 19760
rect 34329 19755 34395 19758
rect 27705 19682 27771 19685
rect 29361 19682 29427 19685
rect 27705 19680 29427 19682
rect 27705 19624 27710 19680
rect 27766 19624 29366 19680
rect 29422 19624 29427 19680
rect 35200 19668 35800 19758
rect 27705 19622 29427 19624
rect 27705 19619 27771 19622
rect 29361 19619 29427 19622
rect 9386 19616 9702 19617
rect 9386 19552 9392 19616
rect 9456 19552 9472 19616
rect 9536 19552 9552 19616
rect 9616 19552 9632 19616
rect 9696 19552 9702 19616
rect 9386 19551 9702 19552
rect 17827 19616 18143 19617
rect 17827 19552 17833 19616
rect 17897 19552 17913 19616
rect 17977 19552 17993 19616
rect 18057 19552 18073 19616
rect 18137 19552 18143 19616
rect 17827 19551 18143 19552
rect 26268 19616 26584 19617
rect 26268 19552 26274 19616
rect 26338 19552 26354 19616
rect 26418 19552 26434 19616
rect 26498 19552 26514 19616
rect 26578 19552 26584 19616
rect 26268 19551 26584 19552
rect 34709 19616 35025 19617
rect 34709 19552 34715 19616
rect 34779 19552 34795 19616
rect 34859 19552 34875 19616
rect 34939 19552 34955 19616
rect 35019 19552 35025 19616
rect 34709 19551 35025 19552
rect 200 19138 800 19228
rect 2221 19138 2287 19141
rect 200 19136 2287 19138
rect 200 19080 2226 19136
rect 2282 19080 2287 19136
rect 200 19078 2287 19080
rect 200 18988 800 19078
rect 2221 19075 2287 19078
rect 34329 19138 34395 19141
rect 35200 19138 35800 19228
rect 34329 19136 35800 19138
rect 34329 19080 34334 19136
rect 34390 19080 35800 19136
rect 34329 19078 35800 19080
rect 34329 19075 34395 19078
rect 5166 19072 5482 19073
rect 5166 19008 5172 19072
rect 5236 19008 5252 19072
rect 5316 19008 5332 19072
rect 5396 19008 5412 19072
rect 5476 19008 5482 19072
rect 5166 19007 5482 19008
rect 13607 19072 13923 19073
rect 13607 19008 13613 19072
rect 13677 19008 13693 19072
rect 13757 19008 13773 19072
rect 13837 19008 13853 19072
rect 13917 19008 13923 19072
rect 13607 19007 13923 19008
rect 22048 19072 22364 19073
rect 22048 19008 22054 19072
rect 22118 19008 22134 19072
rect 22198 19008 22214 19072
rect 22278 19008 22294 19072
rect 22358 19008 22364 19072
rect 22048 19007 22364 19008
rect 30489 19072 30805 19073
rect 30489 19008 30495 19072
rect 30559 19008 30575 19072
rect 30639 19008 30655 19072
rect 30719 19008 30735 19072
rect 30799 19008 30805 19072
rect 30489 19007 30805 19008
rect 32254 18940 32260 19004
rect 32324 19002 32330 19004
rect 32397 19002 32463 19005
rect 32324 19000 32463 19002
rect 32324 18944 32402 19000
rect 32458 18944 32463 19000
rect 35200 18988 35800 19078
rect 32324 18942 32463 18944
rect 32324 18940 32330 18942
rect 32397 18939 32463 18942
rect 29729 18866 29795 18869
rect 31753 18866 31819 18869
rect 29729 18864 31819 18866
rect 29729 18808 29734 18864
rect 29790 18808 31758 18864
rect 31814 18808 31819 18864
rect 29729 18806 31819 18808
rect 29729 18803 29795 18806
rect 31753 18803 31819 18806
rect 19517 18730 19583 18733
rect 27654 18730 27660 18732
rect 19517 18728 27660 18730
rect 19517 18672 19522 18728
rect 19578 18672 27660 18728
rect 19517 18670 27660 18672
rect 19517 18667 19583 18670
rect 27654 18668 27660 18670
rect 27724 18730 27730 18732
rect 28257 18730 28323 18733
rect 27724 18728 28323 18730
rect 27724 18672 28262 18728
rect 28318 18672 28323 18728
rect 27724 18670 28323 18672
rect 27724 18668 27730 18670
rect 28257 18667 28323 18670
rect 24577 18596 24643 18597
rect 24526 18594 24532 18596
rect 200 18458 800 18548
rect 24486 18534 24532 18594
rect 24596 18592 24643 18596
rect 24638 18536 24643 18592
rect 24526 18532 24532 18534
rect 24596 18532 24643 18536
rect 24577 18531 24643 18532
rect 9386 18528 9702 18529
rect 9386 18464 9392 18528
rect 9456 18464 9472 18528
rect 9536 18464 9552 18528
rect 9616 18464 9632 18528
rect 9696 18464 9702 18528
rect 9386 18463 9702 18464
rect 17827 18528 18143 18529
rect 17827 18464 17833 18528
rect 17897 18464 17913 18528
rect 17977 18464 17993 18528
rect 18057 18464 18073 18528
rect 18137 18464 18143 18528
rect 17827 18463 18143 18464
rect 26268 18528 26584 18529
rect 26268 18464 26274 18528
rect 26338 18464 26354 18528
rect 26418 18464 26434 18528
rect 26498 18464 26514 18528
rect 26578 18464 26584 18528
rect 26268 18463 26584 18464
rect 34709 18528 35025 18529
rect 34709 18464 34715 18528
rect 34779 18464 34795 18528
rect 34859 18464 34875 18528
rect 34939 18464 34955 18528
rect 35019 18464 35025 18528
rect 34709 18463 35025 18464
rect 2773 18458 2839 18461
rect 200 18456 2839 18458
rect 200 18400 2778 18456
rect 2834 18400 2839 18456
rect 200 18398 2839 18400
rect 200 18308 800 18398
rect 2773 18395 2839 18398
rect 31293 18458 31359 18461
rect 31661 18458 31727 18461
rect 31293 18456 31727 18458
rect 31293 18400 31298 18456
rect 31354 18400 31666 18456
rect 31722 18400 31727 18456
rect 31293 18398 31727 18400
rect 31293 18395 31359 18398
rect 31661 18395 31727 18398
rect 35200 18308 35800 18548
rect 32806 17988 32812 18052
rect 32876 18050 32882 18052
rect 33041 18050 33107 18053
rect 32876 18048 33107 18050
rect 32876 17992 33046 18048
rect 33102 17992 33107 18048
rect 32876 17990 33107 17992
rect 32876 17988 32882 17990
rect 33041 17987 33107 17990
rect 5166 17984 5482 17985
rect 5166 17920 5172 17984
rect 5236 17920 5252 17984
rect 5316 17920 5332 17984
rect 5396 17920 5412 17984
rect 5476 17920 5482 17984
rect 5166 17919 5482 17920
rect 13607 17984 13923 17985
rect 13607 17920 13613 17984
rect 13677 17920 13693 17984
rect 13757 17920 13773 17984
rect 13837 17920 13853 17984
rect 13917 17920 13923 17984
rect 13607 17919 13923 17920
rect 22048 17984 22364 17985
rect 22048 17920 22054 17984
rect 22118 17920 22134 17984
rect 22198 17920 22214 17984
rect 22278 17920 22294 17984
rect 22358 17920 22364 17984
rect 22048 17919 22364 17920
rect 30489 17984 30805 17985
rect 30489 17920 30495 17984
rect 30559 17920 30575 17984
rect 30639 17920 30655 17984
rect 30719 17920 30735 17984
rect 30799 17920 30805 17984
rect 30489 17919 30805 17920
rect 200 17628 800 17868
rect 34329 17778 34395 17781
rect 35200 17778 35800 17868
rect 34329 17776 35800 17778
rect 34329 17720 34334 17776
rect 34390 17720 35800 17776
rect 34329 17718 35800 17720
rect 34329 17715 34395 17718
rect 35200 17628 35800 17718
rect 9386 17440 9702 17441
rect 9386 17376 9392 17440
rect 9456 17376 9472 17440
rect 9536 17376 9552 17440
rect 9616 17376 9632 17440
rect 9696 17376 9702 17440
rect 9386 17375 9702 17376
rect 17827 17440 18143 17441
rect 17827 17376 17833 17440
rect 17897 17376 17913 17440
rect 17977 17376 17993 17440
rect 18057 17376 18073 17440
rect 18137 17376 18143 17440
rect 17827 17375 18143 17376
rect 26268 17440 26584 17441
rect 26268 17376 26274 17440
rect 26338 17376 26354 17440
rect 26418 17376 26434 17440
rect 26498 17376 26514 17440
rect 26578 17376 26584 17440
rect 26268 17375 26584 17376
rect 34709 17440 35025 17441
rect 34709 17376 34715 17440
rect 34779 17376 34795 17440
rect 34859 17376 34875 17440
rect 34939 17376 34955 17440
rect 35019 17376 35025 17440
rect 34709 17375 35025 17376
rect 200 17098 800 17188
rect 2773 17098 2839 17101
rect 200 17096 2839 17098
rect 200 17040 2778 17096
rect 2834 17040 2839 17096
rect 200 17038 2839 17040
rect 200 16948 800 17038
rect 2773 17035 2839 17038
rect 30465 17098 30531 17101
rect 31753 17098 31819 17101
rect 30465 17096 31819 17098
rect 30465 17040 30470 17096
rect 30526 17040 31758 17096
rect 31814 17040 31819 17096
rect 30465 17038 31819 17040
rect 30465 17035 30531 17038
rect 31753 17035 31819 17038
rect 34329 17098 34395 17101
rect 35200 17098 35800 17188
rect 34329 17096 35800 17098
rect 34329 17040 34334 17096
rect 34390 17040 35800 17096
rect 34329 17038 35800 17040
rect 34329 17035 34395 17038
rect 35200 16948 35800 17038
rect 5166 16896 5482 16897
rect 5166 16832 5172 16896
rect 5236 16832 5252 16896
rect 5316 16832 5332 16896
rect 5396 16832 5412 16896
rect 5476 16832 5482 16896
rect 5166 16831 5482 16832
rect 13607 16896 13923 16897
rect 13607 16832 13613 16896
rect 13677 16832 13693 16896
rect 13757 16832 13773 16896
rect 13837 16832 13853 16896
rect 13917 16832 13923 16896
rect 13607 16831 13923 16832
rect 22048 16896 22364 16897
rect 22048 16832 22054 16896
rect 22118 16832 22134 16896
rect 22198 16832 22214 16896
rect 22278 16832 22294 16896
rect 22358 16832 22364 16896
rect 22048 16831 22364 16832
rect 30489 16896 30805 16897
rect 30489 16832 30495 16896
rect 30559 16832 30575 16896
rect 30639 16832 30655 16896
rect 30719 16832 30735 16896
rect 30799 16832 30805 16896
rect 30489 16831 30805 16832
rect 30925 16826 30991 16829
rect 31150 16826 31156 16828
rect 30925 16824 31156 16826
rect 30925 16768 30930 16824
rect 30986 16768 31156 16824
rect 30925 16766 31156 16768
rect 30925 16763 30991 16766
rect 31150 16764 31156 16766
rect 31220 16764 31226 16828
rect 31334 16764 31340 16828
rect 31404 16826 31410 16828
rect 31477 16826 31543 16829
rect 31404 16824 31543 16826
rect 31404 16768 31482 16824
rect 31538 16768 31543 16824
rect 31404 16766 31543 16768
rect 31404 16764 31410 16766
rect 31477 16763 31543 16766
rect 29545 16690 29611 16693
rect 30465 16690 30531 16693
rect 29545 16688 30531 16690
rect 29545 16632 29550 16688
rect 29606 16632 30470 16688
rect 30526 16632 30531 16688
rect 29545 16630 30531 16632
rect 29545 16627 29611 16630
rect 30465 16627 30531 16630
rect 30649 16690 30715 16693
rect 32070 16690 32076 16692
rect 30649 16688 32076 16690
rect 30649 16632 30654 16688
rect 30710 16632 32076 16688
rect 30649 16630 32076 16632
rect 30649 16627 30715 16630
rect 32070 16628 32076 16630
rect 32140 16628 32146 16692
rect 200 16268 800 16508
rect 24526 16492 24532 16556
rect 24596 16554 24602 16556
rect 25865 16554 25931 16557
rect 24596 16552 25931 16554
rect 24596 16496 25870 16552
rect 25926 16496 25931 16552
rect 24596 16494 25931 16496
rect 24596 16492 24602 16494
rect 25865 16491 25931 16494
rect 29678 16492 29684 16556
rect 29748 16554 29754 16556
rect 31201 16554 31267 16557
rect 29748 16552 31267 16554
rect 29748 16496 31206 16552
rect 31262 16496 31267 16552
rect 29748 16494 31267 16496
rect 29748 16492 29754 16494
rect 31201 16491 31267 16494
rect 35200 16421 35800 16508
rect 35157 16416 35800 16421
rect 35157 16360 35162 16416
rect 35218 16360 35800 16416
rect 35157 16355 35800 16360
rect 9386 16352 9702 16353
rect 9386 16288 9392 16352
rect 9456 16288 9472 16352
rect 9536 16288 9552 16352
rect 9616 16288 9632 16352
rect 9696 16288 9702 16352
rect 9386 16287 9702 16288
rect 17827 16352 18143 16353
rect 17827 16288 17833 16352
rect 17897 16288 17913 16352
rect 17977 16288 17993 16352
rect 18057 16288 18073 16352
rect 18137 16288 18143 16352
rect 17827 16287 18143 16288
rect 26268 16352 26584 16353
rect 26268 16288 26274 16352
rect 26338 16288 26354 16352
rect 26418 16288 26434 16352
rect 26498 16288 26514 16352
rect 26578 16288 26584 16352
rect 26268 16287 26584 16288
rect 34709 16352 35025 16353
rect 34709 16288 34715 16352
rect 34779 16288 34795 16352
rect 34859 16288 34875 16352
rect 34939 16288 34955 16352
rect 35019 16288 35025 16352
rect 34709 16287 35025 16288
rect 30741 16282 30807 16285
rect 30966 16282 30972 16284
rect 30741 16280 30972 16282
rect 30741 16224 30746 16280
rect 30802 16224 30972 16280
rect 30741 16222 30972 16224
rect 30741 16219 30807 16222
rect 30966 16220 30972 16222
rect 31036 16220 31042 16284
rect 31518 16220 31524 16284
rect 31588 16282 31594 16284
rect 32397 16282 32463 16285
rect 31588 16280 32463 16282
rect 31588 16224 32402 16280
rect 32458 16224 32463 16280
rect 35200 16268 35800 16355
rect 31588 16222 32463 16224
rect 31588 16220 31594 16222
rect 32397 16219 32463 16222
rect 29085 16146 29151 16149
rect 29361 16146 29427 16149
rect 29085 16144 29427 16146
rect 29085 16088 29090 16144
rect 29146 16088 29366 16144
rect 29422 16088 29427 16144
rect 29085 16086 29427 16088
rect 29085 16083 29151 16086
rect 29361 16083 29427 16086
rect 29085 16010 29151 16013
rect 29821 16010 29887 16013
rect 29085 16008 29887 16010
rect 29085 15952 29090 16008
rect 29146 15952 29826 16008
rect 29882 15952 29887 16008
rect 29085 15950 29887 15952
rect 29085 15947 29151 15950
rect 29821 15947 29887 15950
rect 200 15738 800 15828
rect 5166 15808 5482 15809
rect 5166 15744 5172 15808
rect 5236 15744 5252 15808
rect 5316 15744 5332 15808
rect 5396 15744 5412 15808
rect 5476 15744 5482 15808
rect 5166 15743 5482 15744
rect 13607 15808 13923 15809
rect 13607 15744 13613 15808
rect 13677 15744 13693 15808
rect 13757 15744 13773 15808
rect 13837 15744 13853 15808
rect 13917 15744 13923 15808
rect 13607 15743 13923 15744
rect 22048 15808 22364 15809
rect 22048 15744 22054 15808
rect 22118 15744 22134 15808
rect 22198 15744 22214 15808
rect 22278 15744 22294 15808
rect 22358 15744 22364 15808
rect 22048 15743 22364 15744
rect 30489 15808 30805 15809
rect 30489 15744 30495 15808
rect 30559 15744 30575 15808
rect 30639 15744 30655 15808
rect 30719 15744 30735 15808
rect 30799 15744 30805 15808
rect 30489 15743 30805 15744
rect 2773 15738 2839 15741
rect 200 15736 2839 15738
rect 200 15680 2778 15736
rect 2834 15680 2839 15736
rect 200 15678 2839 15680
rect 200 15588 800 15678
rect 2773 15675 2839 15678
rect 28993 15602 29059 15605
rect 30833 15602 30899 15605
rect 33685 15602 33751 15605
rect 28993 15600 33751 15602
rect 28993 15544 28998 15600
rect 29054 15544 30838 15600
rect 30894 15544 33690 15600
rect 33746 15544 33751 15600
rect 35200 15588 35800 15828
rect 28993 15542 33751 15544
rect 28993 15539 29059 15542
rect 30833 15539 30899 15542
rect 33685 15539 33751 15542
rect 23565 15466 23631 15469
rect 26417 15466 26483 15469
rect 23565 15464 26483 15466
rect 23565 15408 23570 15464
rect 23626 15408 26422 15464
rect 26478 15408 26483 15464
rect 23565 15406 26483 15408
rect 23565 15403 23631 15406
rect 26417 15403 26483 15406
rect 25589 15332 25655 15333
rect 25589 15330 25636 15332
rect 25544 15328 25636 15330
rect 25544 15272 25594 15328
rect 25544 15270 25636 15272
rect 25589 15268 25636 15270
rect 25700 15268 25706 15332
rect 25589 15267 25655 15268
rect 9386 15264 9702 15265
rect 9386 15200 9392 15264
rect 9456 15200 9472 15264
rect 9536 15200 9552 15264
rect 9616 15200 9632 15264
rect 9696 15200 9702 15264
rect 9386 15199 9702 15200
rect 17827 15264 18143 15265
rect 17827 15200 17833 15264
rect 17897 15200 17913 15264
rect 17977 15200 17993 15264
rect 18057 15200 18073 15264
rect 18137 15200 18143 15264
rect 17827 15199 18143 15200
rect 26268 15264 26584 15265
rect 26268 15200 26274 15264
rect 26338 15200 26354 15264
rect 26418 15200 26434 15264
rect 26498 15200 26514 15264
rect 26578 15200 26584 15264
rect 26268 15199 26584 15200
rect 34709 15264 35025 15265
rect 34709 15200 34715 15264
rect 34779 15200 34795 15264
rect 34859 15200 34875 15264
rect 34939 15200 34955 15264
rect 35019 15200 35025 15264
rect 34709 15199 35025 15200
rect 29361 15194 29427 15197
rect 29494 15194 29500 15196
rect 29361 15192 29500 15194
rect 200 14908 800 15148
rect 29361 15136 29366 15192
rect 29422 15136 29500 15192
rect 29361 15134 29500 15136
rect 29361 15131 29427 15134
rect 29494 15132 29500 15134
rect 29564 15132 29570 15196
rect 22001 15058 22067 15061
rect 24710 15058 24716 15060
rect 22001 15056 24716 15058
rect 22001 15000 22006 15056
rect 22062 15000 24716 15056
rect 22001 14998 24716 15000
rect 22001 14995 22067 14998
rect 24710 14996 24716 14998
rect 24780 14996 24786 15060
rect 25589 15058 25655 15061
rect 27654 15058 27660 15060
rect 25589 15056 27660 15058
rect 25589 15000 25594 15056
rect 25650 15000 27660 15056
rect 25589 14998 27660 15000
rect 25589 14995 25655 14998
rect 27654 14996 27660 14998
rect 27724 14996 27730 15060
rect 33777 15058 33843 15061
rect 33910 15058 33916 15060
rect 33777 15056 33916 15058
rect 33777 15000 33782 15056
rect 33838 15000 33916 15056
rect 33777 14998 33916 15000
rect 33777 14995 33843 14998
rect 33910 14996 33916 14998
rect 33980 14996 33986 15060
rect 5166 14720 5482 14721
rect 5166 14656 5172 14720
rect 5236 14656 5252 14720
rect 5316 14656 5332 14720
rect 5396 14656 5412 14720
rect 5476 14656 5482 14720
rect 5166 14655 5482 14656
rect 13607 14720 13923 14721
rect 13607 14656 13613 14720
rect 13677 14656 13693 14720
rect 13757 14656 13773 14720
rect 13837 14656 13853 14720
rect 13917 14656 13923 14720
rect 13607 14655 13923 14656
rect 22048 14720 22364 14721
rect 22048 14656 22054 14720
rect 22118 14656 22134 14720
rect 22198 14656 22214 14720
rect 22278 14656 22294 14720
rect 22358 14656 22364 14720
rect 22048 14655 22364 14656
rect 30489 14720 30805 14721
rect 30489 14656 30495 14720
rect 30559 14656 30575 14720
rect 30639 14656 30655 14720
rect 30719 14656 30735 14720
rect 30799 14656 30805 14720
rect 30489 14655 30805 14656
rect 200 14378 800 14468
rect 2773 14378 2839 14381
rect 200 14376 2839 14378
rect 200 14320 2778 14376
rect 2834 14320 2839 14376
rect 200 14318 2839 14320
rect 200 14228 800 14318
rect 2773 14315 2839 14318
rect 34329 14378 34395 14381
rect 35200 14378 35800 14468
rect 34329 14376 35800 14378
rect 34329 14320 34334 14376
rect 34390 14320 35800 14376
rect 34329 14318 35800 14320
rect 34329 14315 34395 14318
rect 35200 14228 35800 14318
rect 9386 14176 9702 14177
rect 9386 14112 9392 14176
rect 9456 14112 9472 14176
rect 9536 14112 9552 14176
rect 9616 14112 9632 14176
rect 9696 14112 9702 14176
rect 9386 14111 9702 14112
rect 17827 14176 18143 14177
rect 17827 14112 17833 14176
rect 17897 14112 17913 14176
rect 17977 14112 17993 14176
rect 18057 14112 18073 14176
rect 18137 14112 18143 14176
rect 17827 14111 18143 14112
rect 26268 14176 26584 14177
rect 26268 14112 26274 14176
rect 26338 14112 26354 14176
rect 26418 14112 26434 14176
rect 26498 14112 26514 14176
rect 26578 14112 26584 14176
rect 26268 14111 26584 14112
rect 34709 14176 35025 14177
rect 34709 14112 34715 14176
rect 34779 14112 34795 14176
rect 34859 14112 34875 14176
rect 34939 14112 34955 14176
rect 35019 14112 35025 14176
rect 34709 14111 35025 14112
rect 26734 13908 26740 13972
rect 26804 13970 26810 13972
rect 31569 13970 31635 13973
rect 26804 13968 31635 13970
rect 26804 13912 31574 13968
rect 31630 13912 31635 13968
rect 26804 13910 31635 13912
rect 26804 13908 26810 13910
rect 31569 13907 31635 13910
rect 200 13698 800 13788
rect 2773 13698 2839 13701
rect 200 13696 2839 13698
rect 200 13640 2778 13696
rect 2834 13640 2839 13696
rect 200 13638 2839 13640
rect 200 13548 800 13638
rect 2773 13635 2839 13638
rect 34329 13698 34395 13701
rect 35200 13698 35800 13788
rect 34329 13696 35800 13698
rect 34329 13640 34334 13696
rect 34390 13640 35800 13696
rect 34329 13638 35800 13640
rect 34329 13635 34395 13638
rect 5166 13632 5482 13633
rect 5166 13568 5172 13632
rect 5236 13568 5252 13632
rect 5316 13568 5332 13632
rect 5396 13568 5412 13632
rect 5476 13568 5482 13632
rect 5166 13567 5482 13568
rect 13607 13632 13923 13633
rect 13607 13568 13613 13632
rect 13677 13568 13693 13632
rect 13757 13568 13773 13632
rect 13837 13568 13853 13632
rect 13917 13568 13923 13632
rect 13607 13567 13923 13568
rect 22048 13632 22364 13633
rect 22048 13568 22054 13632
rect 22118 13568 22134 13632
rect 22198 13568 22214 13632
rect 22278 13568 22294 13632
rect 22358 13568 22364 13632
rect 22048 13567 22364 13568
rect 30489 13632 30805 13633
rect 30489 13568 30495 13632
rect 30559 13568 30575 13632
rect 30639 13568 30655 13632
rect 30719 13568 30735 13632
rect 30799 13568 30805 13632
rect 30489 13567 30805 13568
rect 31845 13564 31911 13565
rect 31845 13562 31892 13564
rect 31800 13560 31892 13562
rect 31800 13504 31850 13560
rect 31800 13502 31892 13504
rect 31845 13500 31892 13502
rect 31956 13500 31962 13564
rect 33593 13562 33659 13565
rect 33726 13562 33732 13564
rect 33593 13560 33732 13562
rect 33593 13504 33598 13560
rect 33654 13504 33732 13560
rect 33593 13502 33732 13504
rect 31845 13499 31911 13500
rect 33593 13499 33659 13502
rect 33726 13500 33732 13502
rect 33796 13500 33802 13564
rect 35200 13548 35800 13638
rect 29126 13364 29132 13428
rect 29196 13426 29202 13428
rect 33777 13426 33843 13429
rect 29196 13424 33843 13426
rect 29196 13368 33782 13424
rect 33838 13368 33843 13424
rect 29196 13366 33843 13368
rect 29196 13364 29202 13366
rect 33777 13363 33843 13366
rect 9386 13088 9702 13089
rect 9386 13024 9392 13088
rect 9456 13024 9472 13088
rect 9536 13024 9552 13088
rect 9616 13024 9632 13088
rect 9696 13024 9702 13088
rect 9386 13023 9702 13024
rect 17827 13088 18143 13089
rect 17827 13024 17833 13088
rect 17897 13024 17913 13088
rect 17977 13024 17993 13088
rect 18057 13024 18073 13088
rect 18137 13024 18143 13088
rect 17827 13023 18143 13024
rect 26268 13088 26584 13089
rect 26268 13024 26274 13088
rect 26338 13024 26354 13088
rect 26418 13024 26434 13088
rect 26498 13024 26514 13088
rect 26578 13024 26584 13088
rect 26268 13023 26584 13024
rect 34709 13088 35025 13089
rect 34709 13024 34715 13088
rect 34779 13024 34795 13088
rect 34859 13024 34875 13088
rect 34939 13024 34955 13088
rect 35019 13024 35025 13088
rect 34709 13023 35025 13024
rect 35200 13018 35800 13108
rect 34329 12882 34395 12885
rect 35160 12882 35800 13018
rect 34329 12880 35800 12882
rect 34329 12824 34334 12880
rect 34390 12868 35800 12880
rect 34390 12824 35220 12868
rect 34329 12822 35220 12824
rect 34329 12819 34395 12822
rect 5166 12544 5482 12545
rect 5166 12480 5172 12544
rect 5236 12480 5252 12544
rect 5316 12480 5332 12544
rect 5396 12480 5412 12544
rect 5476 12480 5482 12544
rect 5166 12479 5482 12480
rect 13607 12544 13923 12545
rect 13607 12480 13613 12544
rect 13677 12480 13693 12544
rect 13757 12480 13773 12544
rect 13837 12480 13853 12544
rect 13917 12480 13923 12544
rect 13607 12479 13923 12480
rect 22048 12544 22364 12545
rect 22048 12480 22054 12544
rect 22118 12480 22134 12544
rect 22198 12480 22214 12544
rect 22278 12480 22294 12544
rect 22358 12480 22364 12544
rect 22048 12479 22364 12480
rect 30489 12544 30805 12545
rect 30489 12480 30495 12544
rect 30559 12480 30575 12544
rect 30639 12480 30655 12544
rect 30719 12480 30735 12544
rect 30799 12480 30805 12544
rect 30489 12479 30805 12480
rect 200 12188 800 12428
rect 34329 12338 34395 12341
rect 35200 12338 35800 12428
rect 34329 12336 35800 12338
rect 34329 12280 34334 12336
rect 34390 12280 35800 12336
rect 34329 12278 35800 12280
rect 34329 12275 34395 12278
rect 35200 12188 35800 12278
rect 9386 12000 9702 12001
rect 9386 11936 9392 12000
rect 9456 11936 9472 12000
rect 9536 11936 9552 12000
rect 9616 11936 9632 12000
rect 9696 11936 9702 12000
rect 9386 11935 9702 11936
rect 17827 12000 18143 12001
rect 17827 11936 17833 12000
rect 17897 11936 17913 12000
rect 17977 11936 17993 12000
rect 18057 11936 18073 12000
rect 18137 11936 18143 12000
rect 17827 11935 18143 11936
rect 26268 12000 26584 12001
rect 26268 11936 26274 12000
rect 26338 11936 26354 12000
rect 26418 11936 26434 12000
rect 26498 11936 26514 12000
rect 26578 11936 26584 12000
rect 26268 11935 26584 11936
rect 34709 12000 35025 12001
rect 34709 11936 34715 12000
rect 34779 11936 34795 12000
rect 34859 11936 34875 12000
rect 34939 11936 34955 12000
rect 35019 11936 35025 12000
rect 34709 11935 35025 11936
rect 33961 11794 34027 11797
rect 34094 11794 34100 11796
rect 33961 11792 34100 11794
rect 200 11658 800 11748
rect 33961 11736 33966 11792
rect 34022 11736 34100 11792
rect 33961 11734 34100 11736
rect 33961 11731 34027 11734
rect 34094 11732 34100 11734
rect 34164 11732 34170 11796
rect 2773 11658 2839 11661
rect 200 11656 2839 11658
rect 200 11600 2778 11656
rect 2834 11600 2839 11656
rect 200 11598 2839 11600
rect 200 11508 800 11598
rect 2773 11595 2839 11598
rect 35200 11508 35800 11748
rect 5166 11456 5482 11457
rect 5166 11392 5172 11456
rect 5236 11392 5252 11456
rect 5316 11392 5332 11456
rect 5396 11392 5412 11456
rect 5476 11392 5482 11456
rect 5166 11391 5482 11392
rect 13607 11456 13923 11457
rect 13607 11392 13613 11456
rect 13677 11392 13693 11456
rect 13757 11392 13773 11456
rect 13837 11392 13853 11456
rect 13917 11392 13923 11456
rect 13607 11391 13923 11392
rect 22048 11456 22364 11457
rect 22048 11392 22054 11456
rect 22118 11392 22134 11456
rect 22198 11392 22214 11456
rect 22278 11392 22294 11456
rect 22358 11392 22364 11456
rect 22048 11391 22364 11392
rect 30489 11456 30805 11457
rect 30489 11392 30495 11456
rect 30559 11392 30575 11456
rect 30639 11392 30655 11456
rect 30719 11392 30735 11456
rect 30799 11392 30805 11456
rect 30489 11391 30805 11392
rect 200 10978 800 11068
rect 2773 10978 2839 10981
rect 200 10976 2839 10978
rect 200 10920 2778 10976
rect 2834 10920 2839 10976
rect 200 10918 2839 10920
rect 200 10828 800 10918
rect 2773 10915 2839 10918
rect 9386 10912 9702 10913
rect 9386 10848 9392 10912
rect 9456 10848 9472 10912
rect 9536 10848 9552 10912
rect 9616 10848 9632 10912
rect 9696 10848 9702 10912
rect 9386 10847 9702 10848
rect 17827 10912 18143 10913
rect 17827 10848 17833 10912
rect 17897 10848 17913 10912
rect 17977 10848 17993 10912
rect 18057 10848 18073 10912
rect 18137 10848 18143 10912
rect 17827 10847 18143 10848
rect 26268 10912 26584 10913
rect 26268 10848 26274 10912
rect 26338 10848 26354 10912
rect 26418 10848 26434 10912
rect 26498 10848 26514 10912
rect 26578 10848 26584 10912
rect 26268 10847 26584 10848
rect 34709 10912 35025 10913
rect 34709 10848 34715 10912
rect 34779 10848 34795 10912
rect 34859 10848 34875 10912
rect 34939 10848 34955 10912
rect 35019 10848 35025 10912
rect 34709 10847 35025 10848
rect 35200 10828 35800 11068
rect 200 10148 800 10388
rect 5166 10368 5482 10369
rect 5166 10304 5172 10368
rect 5236 10304 5252 10368
rect 5316 10304 5332 10368
rect 5396 10304 5412 10368
rect 5476 10304 5482 10368
rect 5166 10303 5482 10304
rect 13607 10368 13923 10369
rect 13607 10304 13613 10368
rect 13677 10304 13693 10368
rect 13757 10304 13773 10368
rect 13837 10304 13853 10368
rect 13917 10304 13923 10368
rect 13607 10303 13923 10304
rect 22048 10368 22364 10369
rect 22048 10304 22054 10368
rect 22118 10304 22134 10368
rect 22198 10304 22214 10368
rect 22278 10304 22294 10368
rect 22358 10304 22364 10368
rect 22048 10303 22364 10304
rect 30489 10368 30805 10369
rect 30489 10304 30495 10368
rect 30559 10304 30575 10368
rect 30639 10304 30655 10368
rect 30719 10304 30735 10368
rect 30799 10304 30805 10368
rect 30489 10303 30805 10304
rect 35200 10148 35800 10388
rect 9386 9824 9702 9825
rect 9386 9760 9392 9824
rect 9456 9760 9472 9824
rect 9536 9760 9552 9824
rect 9616 9760 9632 9824
rect 9696 9760 9702 9824
rect 9386 9759 9702 9760
rect 17827 9824 18143 9825
rect 17827 9760 17833 9824
rect 17897 9760 17913 9824
rect 17977 9760 17993 9824
rect 18057 9760 18073 9824
rect 18137 9760 18143 9824
rect 17827 9759 18143 9760
rect 26268 9824 26584 9825
rect 26268 9760 26274 9824
rect 26338 9760 26354 9824
rect 26418 9760 26434 9824
rect 26498 9760 26514 9824
rect 26578 9760 26584 9824
rect 26268 9759 26584 9760
rect 34709 9824 35025 9825
rect 34709 9760 34715 9824
rect 34779 9760 34795 9824
rect 34859 9760 34875 9824
rect 34939 9760 34955 9824
rect 35019 9760 35025 9824
rect 34709 9759 35025 9760
rect 200 9468 800 9708
rect 34053 9618 34119 9621
rect 35200 9618 35800 9708
rect 34053 9616 35800 9618
rect 34053 9560 34058 9616
rect 34114 9560 35800 9616
rect 34053 9558 35800 9560
rect 34053 9555 34119 9558
rect 35200 9468 35800 9558
rect 5166 9280 5482 9281
rect 5166 9216 5172 9280
rect 5236 9216 5252 9280
rect 5316 9216 5332 9280
rect 5396 9216 5412 9280
rect 5476 9216 5482 9280
rect 5166 9215 5482 9216
rect 13607 9280 13923 9281
rect 13607 9216 13613 9280
rect 13677 9216 13693 9280
rect 13757 9216 13773 9280
rect 13837 9216 13853 9280
rect 13917 9216 13923 9280
rect 13607 9215 13923 9216
rect 22048 9280 22364 9281
rect 22048 9216 22054 9280
rect 22118 9216 22134 9280
rect 22198 9216 22214 9280
rect 22278 9216 22294 9280
rect 22358 9216 22364 9280
rect 22048 9215 22364 9216
rect 30489 9280 30805 9281
rect 30489 9216 30495 9280
rect 30559 9216 30575 9280
rect 30639 9216 30655 9280
rect 30719 9216 30735 9280
rect 30799 9216 30805 9280
rect 30489 9215 30805 9216
rect 200 8938 800 9028
rect 2773 8938 2839 8941
rect 200 8936 2839 8938
rect 200 8880 2778 8936
rect 2834 8880 2839 8936
rect 200 8878 2839 8880
rect 200 8788 800 8878
rect 2773 8875 2839 8878
rect 34329 8938 34395 8941
rect 35200 8938 35800 9028
rect 34329 8936 35800 8938
rect 34329 8880 34334 8936
rect 34390 8880 35800 8936
rect 34329 8878 35800 8880
rect 34329 8875 34395 8878
rect 35200 8788 35800 8878
rect 9386 8736 9702 8737
rect 9386 8672 9392 8736
rect 9456 8672 9472 8736
rect 9536 8672 9552 8736
rect 9616 8672 9632 8736
rect 9696 8672 9702 8736
rect 9386 8671 9702 8672
rect 17827 8736 18143 8737
rect 17827 8672 17833 8736
rect 17897 8672 17913 8736
rect 17977 8672 17993 8736
rect 18057 8672 18073 8736
rect 18137 8672 18143 8736
rect 17827 8671 18143 8672
rect 26268 8736 26584 8737
rect 26268 8672 26274 8736
rect 26338 8672 26354 8736
rect 26418 8672 26434 8736
rect 26498 8672 26514 8736
rect 26578 8672 26584 8736
rect 26268 8671 26584 8672
rect 34709 8736 35025 8737
rect 34709 8672 34715 8736
rect 34779 8672 34795 8736
rect 34859 8672 34875 8736
rect 34939 8672 34955 8736
rect 35019 8672 35025 8736
rect 34709 8671 35025 8672
rect 200 8258 800 8348
rect 2773 8258 2839 8261
rect 200 8256 2839 8258
rect 200 8200 2778 8256
rect 2834 8200 2839 8256
rect 200 8198 2839 8200
rect 200 8108 800 8198
rect 2773 8195 2839 8198
rect 5166 8192 5482 8193
rect 5166 8128 5172 8192
rect 5236 8128 5252 8192
rect 5316 8128 5332 8192
rect 5396 8128 5412 8192
rect 5476 8128 5482 8192
rect 5166 8127 5482 8128
rect 13607 8192 13923 8193
rect 13607 8128 13613 8192
rect 13677 8128 13693 8192
rect 13757 8128 13773 8192
rect 13837 8128 13853 8192
rect 13917 8128 13923 8192
rect 13607 8127 13923 8128
rect 22048 8192 22364 8193
rect 22048 8128 22054 8192
rect 22118 8128 22134 8192
rect 22198 8128 22214 8192
rect 22278 8128 22294 8192
rect 22358 8128 22364 8192
rect 22048 8127 22364 8128
rect 30489 8192 30805 8193
rect 30489 8128 30495 8192
rect 30559 8128 30575 8192
rect 30639 8128 30655 8192
rect 30719 8128 30735 8192
rect 30799 8128 30805 8192
rect 30489 8127 30805 8128
rect 200 7578 800 7668
rect 9386 7648 9702 7649
rect 9386 7584 9392 7648
rect 9456 7584 9472 7648
rect 9536 7584 9552 7648
rect 9616 7584 9632 7648
rect 9696 7584 9702 7648
rect 9386 7583 9702 7584
rect 17827 7648 18143 7649
rect 17827 7584 17833 7648
rect 17897 7584 17913 7648
rect 17977 7584 17993 7648
rect 18057 7584 18073 7648
rect 18137 7584 18143 7648
rect 17827 7583 18143 7584
rect 26268 7648 26584 7649
rect 26268 7584 26274 7648
rect 26338 7584 26354 7648
rect 26418 7584 26434 7648
rect 26498 7584 26514 7648
rect 26578 7584 26584 7648
rect 26268 7583 26584 7584
rect 34709 7648 35025 7649
rect 34709 7584 34715 7648
rect 34779 7584 34795 7648
rect 34859 7584 34875 7648
rect 34939 7584 34955 7648
rect 35019 7584 35025 7648
rect 34709 7583 35025 7584
rect 2773 7578 2839 7581
rect 200 7576 2839 7578
rect 200 7520 2778 7576
rect 2834 7520 2839 7576
rect 200 7518 2839 7520
rect 200 7428 800 7518
rect 2773 7515 2839 7518
rect 35200 7428 35800 7668
rect 5166 7104 5482 7105
rect 5166 7040 5172 7104
rect 5236 7040 5252 7104
rect 5316 7040 5332 7104
rect 5396 7040 5412 7104
rect 5476 7040 5482 7104
rect 5166 7039 5482 7040
rect 13607 7104 13923 7105
rect 13607 7040 13613 7104
rect 13677 7040 13693 7104
rect 13757 7040 13773 7104
rect 13837 7040 13853 7104
rect 13917 7040 13923 7104
rect 13607 7039 13923 7040
rect 22048 7104 22364 7105
rect 22048 7040 22054 7104
rect 22118 7040 22134 7104
rect 22198 7040 22214 7104
rect 22278 7040 22294 7104
rect 22358 7040 22364 7104
rect 22048 7039 22364 7040
rect 30489 7104 30805 7105
rect 30489 7040 30495 7104
rect 30559 7040 30575 7104
rect 30639 7040 30655 7104
rect 30719 7040 30735 7104
rect 30799 7040 30805 7104
rect 30489 7039 30805 7040
rect 200 6748 800 6988
rect 34329 6898 34395 6901
rect 35200 6898 35800 6988
rect 34329 6896 35800 6898
rect 34329 6840 34334 6896
rect 34390 6840 35800 6896
rect 34329 6838 35800 6840
rect 34329 6835 34395 6838
rect 35200 6748 35800 6838
rect 9386 6560 9702 6561
rect 9386 6496 9392 6560
rect 9456 6496 9472 6560
rect 9536 6496 9552 6560
rect 9616 6496 9632 6560
rect 9696 6496 9702 6560
rect 9386 6495 9702 6496
rect 17827 6560 18143 6561
rect 17827 6496 17833 6560
rect 17897 6496 17913 6560
rect 17977 6496 17993 6560
rect 18057 6496 18073 6560
rect 18137 6496 18143 6560
rect 17827 6495 18143 6496
rect 26268 6560 26584 6561
rect 26268 6496 26274 6560
rect 26338 6496 26354 6560
rect 26418 6496 26434 6560
rect 26498 6496 26514 6560
rect 26578 6496 26584 6560
rect 26268 6495 26584 6496
rect 34709 6560 35025 6561
rect 34709 6496 34715 6560
rect 34779 6496 34795 6560
rect 34859 6496 34875 6560
rect 34939 6496 34955 6560
rect 35019 6496 35025 6560
rect 34709 6495 35025 6496
rect 35200 6068 35800 6308
rect 5166 6016 5482 6017
rect 5166 5952 5172 6016
rect 5236 5952 5252 6016
rect 5316 5952 5332 6016
rect 5396 5952 5412 6016
rect 5476 5952 5482 6016
rect 5166 5951 5482 5952
rect 13607 6016 13923 6017
rect 13607 5952 13613 6016
rect 13677 5952 13693 6016
rect 13757 5952 13773 6016
rect 13837 5952 13853 6016
rect 13917 5952 13923 6016
rect 13607 5951 13923 5952
rect 22048 6016 22364 6017
rect 22048 5952 22054 6016
rect 22118 5952 22134 6016
rect 22198 5952 22214 6016
rect 22278 5952 22294 6016
rect 22358 5952 22364 6016
rect 22048 5951 22364 5952
rect 30489 6016 30805 6017
rect 30489 5952 30495 6016
rect 30559 5952 30575 6016
rect 30639 5952 30655 6016
rect 30719 5952 30735 6016
rect 30799 5952 30805 6016
rect 30489 5951 30805 5952
rect 200 5538 800 5628
rect 3417 5538 3483 5541
rect 200 5536 3483 5538
rect 200 5480 3422 5536
rect 3478 5480 3483 5536
rect 200 5478 3483 5480
rect 200 5388 800 5478
rect 3417 5475 3483 5478
rect 9386 5472 9702 5473
rect 9386 5408 9392 5472
rect 9456 5408 9472 5472
rect 9536 5408 9552 5472
rect 9616 5408 9632 5472
rect 9696 5408 9702 5472
rect 9386 5407 9702 5408
rect 17827 5472 18143 5473
rect 17827 5408 17833 5472
rect 17897 5408 17913 5472
rect 17977 5408 17993 5472
rect 18057 5408 18073 5472
rect 18137 5408 18143 5472
rect 17827 5407 18143 5408
rect 26268 5472 26584 5473
rect 26268 5408 26274 5472
rect 26338 5408 26354 5472
rect 26418 5408 26434 5472
rect 26498 5408 26514 5472
rect 26578 5408 26584 5472
rect 26268 5407 26584 5408
rect 34709 5472 35025 5473
rect 34709 5408 34715 5472
rect 34779 5408 34795 5472
rect 34859 5408 34875 5472
rect 34939 5408 34955 5472
rect 35019 5408 35025 5472
rect 34709 5407 35025 5408
rect 35200 5388 35800 5628
rect 200 4858 800 4948
rect 5166 4928 5482 4929
rect 5166 4864 5172 4928
rect 5236 4864 5252 4928
rect 5316 4864 5332 4928
rect 5396 4864 5412 4928
rect 5476 4864 5482 4928
rect 5166 4863 5482 4864
rect 13607 4928 13923 4929
rect 13607 4864 13613 4928
rect 13677 4864 13693 4928
rect 13757 4864 13773 4928
rect 13837 4864 13853 4928
rect 13917 4864 13923 4928
rect 13607 4863 13923 4864
rect 22048 4928 22364 4929
rect 22048 4864 22054 4928
rect 22118 4864 22134 4928
rect 22198 4864 22214 4928
rect 22278 4864 22294 4928
rect 22358 4864 22364 4928
rect 22048 4863 22364 4864
rect 30489 4928 30805 4929
rect 30489 4864 30495 4928
rect 30559 4864 30575 4928
rect 30639 4864 30655 4928
rect 30719 4864 30735 4928
rect 30799 4864 30805 4928
rect 30489 4863 30805 4864
rect 2773 4858 2839 4861
rect 200 4856 2839 4858
rect 200 4800 2778 4856
rect 2834 4800 2839 4856
rect 200 4798 2839 4800
rect 200 4708 800 4798
rect 2773 4795 2839 4798
rect 34329 4858 34395 4861
rect 35200 4858 35800 4948
rect 34329 4856 35800 4858
rect 34329 4800 34334 4856
rect 34390 4800 35800 4856
rect 34329 4798 35800 4800
rect 34329 4795 34395 4798
rect 35200 4708 35800 4798
rect 9386 4384 9702 4385
rect 9386 4320 9392 4384
rect 9456 4320 9472 4384
rect 9536 4320 9552 4384
rect 9616 4320 9632 4384
rect 9696 4320 9702 4384
rect 9386 4319 9702 4320
rect 17827 4384 18143 4385
rect 17827 4320 17833 4384
rect 17897 4320 17913 4384
rect 17977 4320 17993 4384
rect 18057 4320 18073 4384
rect 18137 4320 18143 4384
rect 17827 4319 18143 4320
rect 26268 4384 26584 4385
rect 26268 4320 26274 4384
rect 26338 4320 26354 4384
rect 26418 4320 26434 4384
rect 26498 4320 26514 4384
rect 26578 4320 26584 4384
rect 26268 4319 26584 4320
rect 34709 4384 35025 4385
rect 34709 4320 34715 4384
rect 34779 4320 34795 4384
rect 34859 4320 34875 4384
rect 34939 4320 34955 4384
rect 35019 4320 35025 4384
rect 34709 4319 35025 4320
rect 200 4178 800 4268
rect 2773 4178 2839 4181
rect 200 4176 2839 4178
rect 200 4120 2778 4176
rect 2834 4120 2839 4176
rect 200 4118 2839 4120
rect 200 4028 800 4118
rect 2773 4115 2839 4118
rect 33041 4178 33107 4181
rect 35200 4178 35800 4268
rect 33041 4176 35800 4178
rect 33041 4120 33046 4176
rect 33102 4120 35800 4176
rect 33041 4118 35800 4120
rect 33041 4115 33107 4118
rect 35200 4028 35800 4118
rect 5166 3840 5482 3841
rect 5166 3776 5172 3840
rect 5236 3776 5252 3840
rect 5316 3776 5332 3840
rect 5396 3776 5412 3840
rect 5476 3776 5482 3840
rect 5166 3775 5482 3776
rect 13607 3840 13923 3841
rect 13607 3776 13613 3840
rect 13677 3776 13693 3840
rect 13757 3776 13773 3840
rect 13837 3776 13853 3840
rect 13917 3776 13923 3840
rect 13607 3775 13923 3776
rect 22048 3840 22364 3841
rect 22048 3776 22054 3840
rect 22118 3776 22134 3840
rect 22198 3776 22214 3840
rect 22278 3776 22294 3840
rect 22358 3776 22364 3840
rect 22048 3775 22364 3776
rect 30489 3840 30805 3841
rect 30489 3776 30495 3840
rect 30559 3776 30575 3840
rect 30639 3776 30655 3840
rect 30719 3776 30735 3840
rect 30799 3776 30805 3840
rect 30489 3775 30805 3776
rect 200 3498 800 3588
rect 2865 3498 2931 3501
rect 200 3496 2931 3498
rect 200 3440 2870 3496
rect 2926 3440 2931 3496
rect 200 3438 2931 3440
rect 200 3348 800 3438
rect 2865 3435 2931 3438
rect 34329 3498 34395 3501
rect 35200 3498 35800 3588
rect 34329 3496 35800 3498
rect 34329 3440 34334 3496
rect 34390 3440 35800 3496
rect 34329 3438 35800 3440
rect 34329 3435 34395 3438
rect 35200 3348 35800 3438
rect 9386 3296 9702 3297
rect 9386 3232 9392 3296
rect 9456 3232 9472 3296
rect 9536 3232 9552 3296
rect 9616 3232 9632 3296
rect 9696 3232 9702 3296
rect 9386 3231 9702 3232
rect 17827 3296 18143 3297
rect 17827 3232 17833 3296
rect 17897 3232 17913 3296
rect 17977 3232 17993 3296
rect 18057 3232 18073 3296
rect 18137 3232 18143 3296
rect 17827 3231 18143 3232
rect 26268 3296 26584 3297
rect 26268 3232 26274 3296
rect 26338 3232 26354 3296
rect 26418 3232 26434 3296
rect 26498 3232 26514 3296
rect 26578 3232 26584 3296
rect 26268 3231 26584 3232
rect 34709 3296 35025 3297
rect 34709 3232 34715 3296
rect 34779 3232 34795 3296
rect 34859 3232 34875 3296
rect 34939 3232 34955 3296
rect 35019 3232 35025 3296
rect 34709 3231 35025 3232
rect 200 2818 800 2908
rect 3969 2818 4035 2821
rect 200 2816 4035 2818
rect 200 2760 3974 2816
rect 4030 2760 4035 2816
rect 200 2758 4035 2760
rect 200 2668 800 2758
rect 3969 2755 4035 2758
rect 5166 2752 5482 2753
rect 5166 2688 5172 2752
rect 5236 2688 5252 2752
rect 5316 2688 5332 2752
rect 5396 2688 5412 2752
rect 5476 2688 5482 2752
rect 5166 2687 5482 2688
rect 13607 2752 13923 2753
rect 13607 2688 13613 2752
rect 13677 2688 13693 2752
rect 13757 2688 13773 2752
rect 13837 2688 13853 2752
rect 13917 2688 13923 2752
rect 13607 2687 13923 2688
rect 22048 2752 22364 2753
rect 22048 2688 22054 2752
rect 22118 2688 22134 2752
rect 22198 2688 22214 2752
rect 22278 2688 22294 2752
rect 22358 2688 22364 2752
rect 22048 2687 22364 2688
rect 30489 2752 30805 2753
rect 30489 2688 30495 2752
rect 30559 2688 30575 2752
rect 30639 2688 30655 2752
rect 30719 2688 30735 2752
rect 30799 2688 30805 2752
rect 30489 2687 30805 2688
rect 35200 2668 35800 2908
rect 200 2138 800 2228
rect 9386 2208 9702 2209
rect 9386 2144 9392 2208
rect 9456 2144 9472 2208
rect 9536 2144 9552 2208
rect 9616 2144 9632 2208
rect 9696 2144 9702 2208
rect 9386 2143 9702 2144
rect 17827 2208 18143 2209
rect 17827 2144 17833 2208
rect 17897 2144 17913 2208
rect 17977 2144 17993 2208
rect 18057 2144 18073 2208
rect 18137 2144 18143 2208
rect 17827 2143 18143 2144
rect 26268 2208 26584 2209
rect 26268 2144 26274 2208
rect 26338 2144 26354 2208
rect 26418 2144 26434 2208
rect 26498 2144 26514 2208
rect 26578 2144 26584 2208
rect 26268 2143 26584 2144
rect 34709 2208 35025 2209
rect 34709 2144 34715 2208
rect 34779 2144 34795 2208
rect 34859 2144 34875 2208
rect 34939 2144 34955 2208
rect 35019 2144 35025 2208
rect 34709 2143 35025 2144
rect 2773 2138 2839 2141
rect 200 2136 2839 2138
rect 200 2080 2778 2136
rect 2834 2080 2839 2136
rect 200 2078 2839 2080
rect 200 1988 800 2078
rect 2773 2075 2839 2078
rect 35200 2138 35800 2228
rect 35893 2138 35959 2141
rect 35200 2136 35959 2138
rect 35200 2080 35898 2136
rect 35954 2080 35959 2136
rect 35200 2078 35959 2080
rect 35200 1988 35800 2078
rect 35893 2075 35959 2078
rect 200 1458 800 1548
rect 4061 1458 4127 1461
rect 200 1456 4127 1458
rect 200 1400 4066 1456
rect 4122 1400 4127 1456
rect 200 1398 4127 1400
rect 200 1308 800 1398
rect 4061 1395 4127 1398
rect 34605 914 34671 917
rect 34605 912 34714 914
rect 200 628 800 868
rect 34605 856 34610 912
rect 34666 856 34714 912
rect 34605 851 34714 856
rect 34654 778 34714 851
rect 35200 778 35800 868
rect 34654 718 35800 778
rect 35200 628 35800 718
rect 31845 98 31911 101
rect 35200 98 35800 188
rect 31845 96 35800 98
rect 31845 40 31850 96
rect 31906 40 35800 96
rect 31845 38 35800 40
rect 31845 35 31911 38
rect 35200 -52 35800 38
<< via3 >>
rect 5172 39740 5236 39744
rect 5172 39684 5176 39740
rect 5176 39684 5232 39740
rect 5232 39684 5236 39740
rect 5172 39680 5236 39684
rect 5252 39740 5316 39744
rect 5252 39684 5256 39740
rect 5256 39684 5312 39740
rect 5312 39684 5316 39740
rect 5252 39680 5316 39684
rect 5332 39740 5396 39744
rect 5332 39684 5336 39740
rect 5336 39684 5392 39740
rect 5392 39684 5396 39740
rect 5332 39680 5396 39684
rect 5412 39740 5476 39744
rect 5412 39684 5416 39740
rect 5416 39684 5472 39740
rect 5472 39684 5476 39740
rect 5412 39680 5476 39684
rect 13613 39740 13677 39744
rect 13613 39684 13617 39740
rect 13617 39684 13673 39740
rect 13673 39684 13677 39740
rect 13613 39680 13677 39684
rect 13693 39740 13757 39744
rect 13693 39684 13697 39740
rect 13697 39684 13753 39740
rect 13753 39684 13757 39740
rect 13693 39680 13757 39684
rect 13773 39740 13837 39744
rect 13773 39684 13777 39740
rect 13777 39684 13833 39740
rect 13833 39684 13837 39740
rect 13773 39680 13837 39684
rect 13853 39740 13917 39744
rect 13853 39684 13857 39740
rect 13857 39684 13913 39740
rect 13913 39684 13917 39740
rect 13853 39680 13917 39684
rect 22054 39740 22118 39744
rect 22054 39684 22058 39740
rect 22058 39684 22114 39740
rect 22114 39684 22118 39740
rect 22054 39680 22118 39684
rect 22134 39740 22198 39744
rect 22134 39684 22138 39740
rect 22138 39684 22194 39740
rect 22194 39684 22198 39740
rect 22134 39680 22198 39684
rect 22214 39740 22278 39744
rect 22214 39684 22218 39740
rect 22218 39684 22274 39740
rect 22274 39684 22278 39740
rect 22214 39680 22278 39684
rect 22294 39740 22358 39744
rect 22294 39684 22298 39740
rect 22298 39684 22354 39740
rect 22354 39684 22358 39740
rect 22294 39680 22358 39684
rect 30495 39740 30559 39744
rect 30495 39684 30499 39740
rect 30499 39684 30555 39740
rect 30555 39684 30559 39740
rect 30495 39680 30559 39684
rect 30575 39740 30639 39744
rect 30575 39684 30579 39740
rect 30579 39684 30635 39740
rect 30635 39684 30639 39740
rect 30575 39680 30639 39684
rect 30655 39740 30719 39744
rect 30655 39684 30659 39740
rect 30659 39684 30715 39740
rect 30715 39684 30719 39740
rect 30655 39680 30719 39684
rect 30735 39740 30799 39744
rect 30735 39684 30739 39740
rect 30739 39684 30795 39740
rect 30795 39684 30799 39740
rect 30735 39680 30799 39684
rect 30972 39340 31036 39404
rect 9392 39196 9456 39200
rect 9392 39140 9396 39196
rect 9396 39140 9452 39196
rect 9452 39140 9456 39196
rect 9392 39136 9456 39140
rect 9472 39196 9536 39200
rect 9472 39140 9476 39196
rect 9476 39140 9532 39196
rect 9532 39140 9536 39196
rect 9472 39136 9536 39140
rect 9552 39196 9616 39200
rect 9552 39140 9556 39196
rect 9556 39140 9612 39196
rect 9612 39140 9616 39196
rect 9552 39136 9616 39140
rect 9632 39196 9696 39200
rect 9632 39140 9636 39196
rect 9636 39140 9692 39196
rect 9692 39140 9696 39196
rect 9632 39136 9696 39140
rect 17833 39196 17897 39200
rect 17833 39140 17837 39196
rect 17837 39140 17893 39196
rect 17893 39140 17897 39196
rect 17833 39136 17897 39140
rect 17913 39196 17977 39200
rect 17913 39140 17917 39196
rect 17917 39140 17973 39196
rect 17973 39140 17977 39196
rect 17913 39136 17977 39140
rect 17993 39196 18057 39200
rect 17993 39140 17997 39196
rect 17997 39140 18053 39196
rect 18053 39140 18057 39196
rect 17993 39136 18057 39140
rect 18073 39196 18137 39200
rect 18073 39140 18077 39196
rect 18077 39140 18133 39196
rect 18133 39140 18137 39196
rect 18073 39136 18137 39140
rect 26274 39196 26338 39200
rect 26274 39140 26278 39196
rect 26278 39140 26334 39196
rect 26334 39140 26338 39196
rect 26274 39136 26338 39140
rect 26354 39196 26418 39200
rect 26354 39140 26358 39196
rect 26358 39140 26414 39196
rect 26414 39140 26418 39196
rect 26354 39136 26418 39140
rect 26434 39196 26498 39200
rect 26434 39140 26438 39196
rect 26438 39140 26494 39196
rect 26494 39140 26498 39196
rect 26434 39136 26498 39140
rect 26514 39196 26578 39200
rect 26514 39140 26518 39196
rect 26518 39140 26574 39196
rect 26574 39140 26578 39196
rect 26514 39136 26578 39140
rect 34715 39196 34779 39200
rect 34715 39140 34719 39196
rect 34719 39140 34775 39196
rect 34775 39140 34779 39196
rect 34715 39136 34779 39140
rect 34795 39196 34859 39200
rect 34795 39140 34799 39196
rect 34799 39140 34855 39196
rect 34855 39140 34859 39196
rect 34795 39136 34859 39140
rect 34875 39196 34939 39200
rect 34875 39140 34879 39196
rect 34879 39140 34935 39196
rect 34935 39140 34939 39196
rect 34875 39136 34939 39140
rect 34955 39196 35019 39200
rect 34955 39140 34959 39196
rect 34959 39140 35015 39196
rect 35015 39140 35019 39196
rect 34955 39136 35019 39140
rect 5172 38652 5236 38656
rect 5172 38596 5176 38652
rect 5176 38596 5232 38652
rect 5232 38596 5236 38652
rect 5172 38592 5236 38596
rect 5252 38652 5316 38656
rect 5252 38596 5256 38652
rect 5256 38596 5312 38652
rect 5312 38596 5316 38652
rect 5252 38592 5316 38596
rect 5332 38652 5396 38656
rect 5332 38596 5336 38652
rect 5336 38596 5392 38652
rect 5392 38596 5396 38652
rect 5332 38592 5396 38596
rect 5412 38652 5476 38656
rect 5412 38596 5416 38652
rect 5416 38596 5472 38652
rect 5472 38596 5476 38652
rect 5412 38592 5476 38596
rect 13613 38652 13677 38656
rect 13613 38596 13617 38652
rect 13617 38596 13673 38652
rect 13673 38596 13677 38652
rect 13613 38592 13677 38596
rect 13693 38652 13757 38656
rect 13693 38596 13697 38652
rect 13697 38596 13753 38652
rect 13753 38596 13757 38652
rect 13693 38592 13757 38596
rect 13773 38652 13837 38656
rect 13773 38596 13777 38652
rect 13777 38596 13833 38652
rect 13833 38596 13837 38652
rect 13773 38592 13837 38596
rect 13853 38652 13917 38656
rect 13853 38596 13857 38652
rect 13857 38596 13913 38652
rect 13913 38596 13917 38652
rect 13853 38592 13917 38596
rect 22054 38652 22118 38656
rect 22054 38596 22058 38652
rect 22058 38596 22114 38652
rect 22114 38596 22118 38652
rect 22054 38592 22118 38596
rect 22134 38652 22198 38656
rect 22134 38596 22138 38652
rect 22138 38596 22194 38652
rect 22194 38596 22198 38652
rect 22134 38592 22198 38596
rect 22214 38652 22278 38656
rect 22214 38596 22218 38652
rect 22218 38596 22274 38652
rect 22274 38596 22278 38652
rect 22214 38592 22278 38596
rect 22294 38652 22358 38656
rect 22294 38596 22298 38652
rect 22298 38596 22354 38652
rect 22354 38596 22358 38652
rect 22294 38592 22358 38596
rect 30495 38652 30559 38656
rect 30495 38596 30499 38652
rect 30499 38596 30555 38652
rect 30555 38596 30559 38652
rect 30495 38592 30559 38596
rect 30575 38652 30639 38656
rect 30575 38596 30579 38652
rect 30579 38596 30635 38652
rect 30635 38596 30639 38652
rect 30575 38592 30639 38596
rect 30655 38652 30719 38656
rect 30655 38596 30659 38652
rect 30659 38596 30715 38652
rect 30715 38596 30719 38652
rect 30655 38592 30719 38596
rect 30735 38652 30799 38656
rect 30735 38596 30739 38652
rect 30739 38596 30795 38652
rect 30795 38596 30799 38652
rect 30735 38592 30799 38596
rect 9392 38108 9456 38112
rect 9392 38052 9396 38108
rect 9396 38052 9452 38108
rect 9452 38052 9456 38108
rect 9392 38048 9456 38052
rect 9472 38108 9536 38112
rect 9472 38052 9476 38108
rect 9476 38052 9532 38108
rect 9532 38052 9536 38108
rect 9472 38048 9536 38052
rect 9552 38108 9616 38112
rect 9552 38052 9556 38108
rect 9556 38052 9612 38108
rect 9612 38052 9616 38108
rect 9552 38048 9616 38052
rect 9632 38108 9696 38112
rect 9632 38052 9636 38108
rect 9636 38052 9692 38108
rect 9692 38052 9696 38108
rect 9632 38048 9696 38052
rect 17833 38108 17897 38112
rect 17833 38052 17837 38108
rect 17837 38052 17893 38108
rect 17893 38052 17897 38108
rect 17833 38048 17897 38052
rect 17913 38108 17977 38112
rect 17913 38052 17917 38108
rect 17917 38052 17973 38108
rect 17973 38052 17977 38108
rect 17913 38048 17977 38052
rect 17993 38108 18057 38112
rect 17993 38052 17997 38108
rect 17997 38052 18053 38108
rect 18053 38052 18057 38108
rect 17993 38048 18057 38052
rect 18073 38108 18137 38112
rect 18073 38052 18077 38108
rect 18077 38052 18133 38108
rect 18133 38052 18137 38108
rect 18073 38048 18137 38052
rect 26274 38108 26338 38112
rect 26274 38052 26278 38108
rect 26278 38052 26334 38108
rect 26334 38052 26338 38108
rect 26274 38048 26338 38052
rect 26354 38108 26418 38112
rect 26354 38052 26358 38108
rect 26358 38052 26414 38108
rect 26414 38052 26418 38108
rect 26354 38048 26418 38052
rect 26434 38108 26498 38112
rect 26434 38052 26438 38108
rect 26438 38052 26494 38108
rect 26494 38052 26498 38108
rect 26434 38048 26498 38052
rect 26514 38108 26578 38112
rect 26514 38052 26518 38108
rect 26518 38052 26574 38108
rect 26574 38052 26578 38108
rect 26514 38048 26578 38052
rect 34715 38108 34779 38112
rect 34715 38052 34719 38108
rect 34719 38052 34775 38108
rect 34775 38052 34779 38108
rect 34715 38048 34779 38052
rect 34795 38108 34859 38112
rect 34795 38052 34799 38108
rect 34799 38052 34855 38108
rect 34855 38052 34859 38108
rect 34795 38048 34859 38052
rect 34875 38108 34939 38112
rect 34875 38052 34879 38108
rect 34879 38052 34935 38108
rect 34935 38052 34939 38108
rect 34875 38048 34939 38052
rect 34955 38108 35019 38112
rect 34955 38052 34959 38108
rect 34959 38052 35015 38108
rect 35015 38052 35019 38108
rect 34955 38048 35019 38052
rect 28764 37572 28828 37636
rect 5172 37564 5236 37568
rect 5172 37508 5176 37564
rect 5176 37508 5232 37564
rect 5232 37508 5236 37564
rect 5172 37504 5236 37508
rect 5252 37564 5316 37568
rect 5252 37508 5256 37564
rect 5256 37508 5312 37564
rect 5312 37508 5316 37564
rect 5252 37504 5316 37508
rect 5332 37564 5396 37568
rect 5332 37508 5336 37564
rect 5336 37508 5392 37564
rect 5392 37508 5396 37564
rect 5332 37504 5396 37508
rect 5412 37564 5476 37568
rect 5412 37508 5416 37564
rect 5416 37508 5472 37564
rect 5472 37508 5476 37564
rect 5412 37504 5476 37508
rect 13613 37564 13677 37568
rect 13613 37508 13617 37564
rect 13617 37508 13673 37564
rect 13673 37508 13677 37564
rect 13613 37504 13677 37508
rect 13693 37564 13757 37568
rect 13693 37508 13697 37564
rect 13697 37508 13753 37564
rect 13753 37508 13757 37564
rect 13693 37504 13757 37508
rect 13773 37564 13837 37568
rect 13773 37508 13777 37564
rect 13777 37508 13833 37564
rect 13833 37508 13837 37564
rect 13773 37504 13837 37508
rect 13853 37564 13917 37568
rect 13853 37508 13857 37564
rect 13857 37508 13913 37564
rect 13913 37508 13917 37564
rect 13853 37504 13917 37508
rect 22054 37564 22118 37568
rect 22054 37508 22058 37564
rect 22058 37508 22114 37564
rect 22114 37508 22118 37564
rect 22054 37504 22118 37508
rect 22134 37564 22198 37568
rect 22134 37508 22138 37564
rect 22138 37508 22194 37564
rect 22194 37508 22198 37564
rect 22134 37504 22198 37508
rect 22214 37564 22278 37568
rect 22214 37508 22218 37564
rect 22218 37508 22274 37564
rect 22274 37508 22278 37564
rect 22214 37504 22278 37508
rect 22294 37564 22358 37568
rect 22294 37508 22298 37564
rect 22298 37508 22354 37564
rect 22354 37508 22358 37564
rect 22294 37504 22358 37508
rect 30495 37564 30559 37568
rect 30495 37508 30499 37564
rect 30499 37508 30555 37564
rect 30555 37508 30559 37564
rect 30495 37504 30559 37508
rect 30575 37564 30639 37568
rect 30575 37508 30579 37564
rect 30579 37508 30635 37564
rect 30635 37508 30639 37564
rect 30575 37504 30639 37508
rect 30655 37564 30719 37568
rect 30655 37508 30659 37564
rect 30659 37508 30715 37564
rect 30715 37508 30719 37564
rect 30655 37504 30719 37508
rect 30735 37564 30799 37568
rect 30735 37508 30739 37564
rect 30739 37508 30795 37564
rect 30795 37508 30799 37564
rect 30735 37504 30799 37508
rect 28948 37436 29012 37500
rect 29316 37436 29380 37500
rect 31524 37164 31588 37228
rect 24716 37088 24780 37092
rect 24716 37032 24730 37088
rect 24730 37032 24780 37088
rect 24716 37028 24780 37032
rect 30972 37088 31036 37092
rect 30972 37032 30986 37088
rect 30986 37032 31036 37088
rect 30972 37028 31036 37032
rect 9392 37020 9456 37024
rect 9392 36964 9396 37020
rect 9396 36964 9452 37020
rect 9452 36964 9456 37020
rect 9392 36960 9456 36964
rect 9472 37020 9536 37024
rect 9472 36964 9476 37020
rect 9476 36964 9532 37020
rect 9532 36964 9536 37020
rect 9472 36960 9536 36964
rect 9552 37020 9616 37024
rect 9552 36964 9556 37020
rect 9556 36964 9612 37020
rect 9612 36964 9616 37020
rect 9552 36960 9616 36964
rect 9632 37020 9696 37024
rect 9632 36964 9636 37020
rect 9636 36964 9692 37020
rect 9692 36964 9696 37020
rect 9632 36960 9696 36964
rect 17833 37020 17897 37024
rect 17833 36964 17837 37020
rect 17837 36964 17893 37020
rect 17893 36964 17897 37020
rect 17833 36960 17897 36964
rect 17913 37020 17977 37024
rect 17913 36964 17917 37020
rect 17917 36964 17973 37020
rect 17973 36964 17977 37020
rect 17913 36960 17977 36964
rect 17993 37020 18057 37024
rect 17993 36964 17997 37020
rect 17997 36964 18053 37020
rect 18053 36964 18057 37020
rect 17993 36960 18057 36964
rect 18073 37020 18137 37024
rect 18073 36964 18077 37020
rect 18077 36964 18133 37020
rect 18133 36964 18137 37020
rect 18073 36960 18137 36964
rect 26274 37020 26338 37024
rect 26274 36964 26278 37020
rect 26278 36964 26334 37020
rect 26334 36964 26338 37020
rect 26274 36960 26338 36964
rect 26354 37020 26418 37024
rect 26354 36964 26358 37020
rect 26358 36964 26414 37020
rect 26414 36964 26418 37020
rect 26354 36960 26418 36964
rect 26434 37020 26498 37024
rect 26434 36964 26438 37020
rect 26438 36964 26494 37020
rect 26494 36964 26498 37020
rect 26434 36960 26498 36964
rect 26514 37020 26578 37024
rect 26514 36964 26518 37020
rect 26518 36964 26574 37020
rect 26574 36964 26578 37020
rect 26514 36960 26578 36964
rect 34715 37020 34779 37024
rect 34715 36964 34719 37020
rect 34719 36964 34775 37020
rect 34775 36964 34779 37020
rect 34715 36960 34779 36964
rect 34795 37020 34859 37024
rect 34795 36964 34799 37020
rect 34799 36964 34855 37020
rect 34855 36964 34859 37020
rect 34795 36960 34859 36964
rect 34875 37020 34939 37024
rect 34875 36964 34879 37020
rect 34879 36964 34935 37020
rect 34935 36964 34939 37020
rect 34875 36960 34939 36964
rect 34955 37020 35019 37024
rect 34955 36964 34959 37020
rect 34959 36964 35015 37020
rect 35015 36964 35019 37020
rect 34955 36960 35019 36964
rect 29132 36544 29196 36548
rect 29132 36488 29182 36544
rect 29182 36488 29196 36544
rect 29132 36484 29196 36488
rect 29500 36544 29564 36548
rect 29500 36488 29514 36544
rect 29514 36488 29564 36544
rect 29500 36484 29564 36488
rect 5172 36476 5236 36480
rect 5172 36420 5176 36476
rect 5176 36420 5232 36476
rect 5232 36420 5236 36476
rect 5172 36416 5236 36420
rect 5252 36476 5316 36480
rect 5252 36420 5256 36476
rect 5256 36420 5312 36476
rect 5312 36420 5316 36476
rect 5252 36416 5316 36420
rect 5332 36476 5396 36480
rect 5332 36420 5336 36476
rect 5336 36420 5392 36476
rect 5392 36420 5396 36476
rect 5332 36416 5396 36420
rect 5412 36476 5476 36480
rect 5412 36420 5416 36476
rect 5416 36420 5472 36476
rect 5472 36420 5476 36476
rect 5412 36416 5476 36420
rect 13613 36476 13677 36480
rect 13613 36420 13617 36476
rect 13617 36420 13673 36476
rect 13673 36420 13677 36476
rect 13613 36416 13677 36420
rect 13693 36476 13757 36480
rect 13693 36420 13697 36476
rect 13697 36420 13753 36476
rect 13753 36420 13757 36476
rect 13693 36416 13757 36420
rect 13773 36476 13837 36480
rect 13773 36420 13777 36476
rect 13777 36420 13833 36476
rect 13833 36420 13837 36476
rect 13773 36416 13837 36420
rect 13853 36476 13917 36480
rect 13853 36420 13857 36476
rect 13857 36420 13913 36476
rect 13913 36420 13917 36476
rect 13853 36416 13917 36420
rect 22054 36476 22118 36480
rect 22054 36420 22058 36476
rect 22058 36420 22114 36476
rect 22114 36420 22118 36476
rect 22054 36416 22118 36420
rect 22134 36476 22198 36480
rect 22134 36420 22138 36476
rect 22138 36420 22194 36476
rect 22194 36420 22198 36476
rect 22134 36416 22198 36420
rect 22214 36476 22278 36480
rect 22214 36420 22218 36476
rect 22218 36420 22274 36476
rect 22274 36420 22278 36476
rect 22214 36416 22278 36420
rect 22294 36476 22358 36480
rect 22294 36420 22298 36476
rect 22298 36420 22354 36476
rect 22354 36420 22358 36476
rect 22294 36416 22358 36420
rect 30495 36476 30559 36480
rect 30495 36420 30499 36476
rect 30499 36420 30555 36476
rect 30555 36420 30559 36476
rect 30495 36416 30559 36420
rect 30575 36476 30639 36480
rect 30575 36420 30579 36476
rect 30579 36420 30635 36476
rect 30635 36420 30639 36476
rect 30575 36416 30639 36420
rect 30655 36476 30719 36480
rect 30655 36420 30659 36476
rect 30659 36420 30715 36476
rect 30715 36420 30719 36476
rect 30655 36416 30719 36420
rect 30735 36476 30799 36480
rect 30735 36420 30739 36476
rect 30739 36420 30795 36476
rect 30795 36420 30799 36476
rect 30735 36416 30799 36420
rect 30236 36348 30300 36412
rect 31156 36408 31220 36412
rect 31156 36352 31170 36408
rect 31170 36352 31220 36408
rect 31156 36348 31220 36352
rect 27660 35940 27724 36004
rect 9392 35932 9456 35936
rect 9392 35876 9396 35932
rect 9396 35876 9452 35932
rect 9452 35876 9456 35932
rect 9392 35872 9456 35876
rect 9472 35932 9536 35936
rect 9472 35876 9476 35932
rect 9476 35876 9532 35932
rect 9532 35876 9536 35932
rect 9472 35872 9536 35876
rect 9552 35932 9616 35936
rect 9552 35876 9556 35932
rect 9556 35876 9612 35932
rect 9612 35876 9616 35932
rect 9552 35872 9616 35876
rect 9632 35932 9696 35936
rect 9632 35876 9636 35932
rect 9636 35876 9692 35932
rect 9692 35876 9696 35932
rect 9632 35872 9696 35876
rect 17833 35932 17897 35936
rect 17833 35876 17837 35932
rect 17837 35876 17893 35932
rect 17893 35876 17897 35932
rect 17833 35872 17897 35876
rect 17913 35932 17977 35936
rect 17913 35876 17917 35932
rect 17917 35876 17973 35932
rect 17973 35876 17977 35932
rect 17913 35872 17977 35876
rect 17993 35932 18057 35936
rect 17993 35876 17997 35932
rect 17997 35876 18053 35932
rect 18053 35876 18057 35932
rect 17993 35872 18057 35876
rect 18073 35932 18137 35936
rect 18073 35876 18077 35932
rect 18077 35876 18133 35932
rect 18133 35876 18137 35932
rect 18073 35872 18137 35876
rect 26274 35932 26338 35936
rect 26274 35876 26278 35932
rect 26278 35876 26334 35932
rect 26334 35876 26338 35932
rect 26274 35872 26338 35876
rect 26354 35932 26418 35936
rect 26354 35876 26358 35932
rect 26358 35876 26414 35932
rect 26414 35876 26418 35932
rect 26354 35872 26418 35876
rect 26434 35932 26498 35936
rect 26434 35876 26438 35932
rect 26438 35876 26494 35932
rect 26494 35876 26498 35932
rect 26434 35872 26498 35876
rect 26514 35932 26578 35936
rect 26514 35876 26518 35932
rect 26518 35876 26574 35932
rect 26574 35876 26578 35932
rect 26514 35872 26578 35876
rect 34715 35932 34779 35936
rect 34715 35876 34719 35932
rect 34719 35876 34775 35932
rect 34775 35876 34779 35932
rect 34715 35872 34779 35876
rect 34795 35932 34859 35936
rect 34795 35876 34799 35932
rect 34799 35876 34855 35932
rect 34855 35876 34859 35932
rect 34795 35872 34859 35876
rect 34875 35932 34939 35936
rect 34875 35876 34879 35932
rect 34879 35876 34935 35932
rect 34935 35876 34939 35932
rect 34875 35872 34939 35876
rect 34955 35932 35019 35936
rect 34955 35876 34959 35932
rect 34959 35876 35015 35932
rect 35015 35876 35019 35932
rect 34955 35872 35019 35876
rect 29132 35864 29196 35868
rect 29132 35808 29182 35864
rect 29182 35808 29196 35864
rect 29132 35804 29196 35808
rect 32260 35396 32324 35460
rect 5172 35388 5236 35392
rect 5172 35332 5176 35388
rect 5176 35332 5232 35388
rect 5232 35332 5236 35388
rect 5172 35328 5236 35332
rect 5252 35388 5316 35392
rect 5252 35332 5256 35388
rect 5256 35332 5312 35388
rect 5312 35332 5316 35388
rect 5252 35328 5316 35332
rect 5332 35388 5396 35392
rect 5332 35332 5336 35388
rect 5336 35332 5392 35388
rect 5392 35332 5396 35388
rect 5332 35328 5396 35332
rect 5412 35388 5476 35392
rect 5412 35332 5416 35388
rect 5416 35332 5472 35388
rect 5472 35332 5476 35388
rect 5412 35328 5476 35332
rect 13613 35388 13677 35392
rect 13613 35332 13617 35388
rect 13617 35332 13673 35388
rect 13673 35332 13677 35388
rect 13613 35328 13677 35332
rect 13693 35388 13757 35392
rect 13693 35332 13697 35388
rect 13697 35332 13753 35388
rect 13753 35332 13757 35388
rect 13693 35328 13757 35332
rect 13773 35388 13837 35392
rect 13773 35332 13777 35388
rect 13777 35332 13833 35388
rect 13833 35332 13837 35388
rect 13773 35328 13837 35332
rect 13853 35388 13917 35392
rect 13853 35332 13857 35388
rect 13857 35332 13913 35388
rect 13913 35332 13917 35388
rect 13853 35328 13917 35332
rect 22054 35388 22118 35392
rect 22054 35332 22058 35388
rect 22058 35332 22114 35388
rect 22114 35332 22118 35388
rect 22054 35328 22118 35332
rect 22134 35388 22198 35392
rect 22134 35332 22138 35388
rect 22138 35332 22194 35388
rect 22194 35332 22198 35388
rect 22134 35328 22198 35332
rect 22214 35388 22278 35392
rect 22214 35332 22218 35388
rect 22218 35332 22274 35388
rect 22274 35332 22278 35388
rect 22214 35328 22278 35332
rect 22294 35388 22358 35392
rect 22294 35332 22298 35388
rect 22298 35332 22354 35388
rect 22354 35332 22358 35388
rect 22294 35328 22358 35332
rect 30495 35388 30559 35392
rect 30495 35332 30499 35388
rect 30499 35332 30555 35388
rect 30555 35332 30559 35388
rect 30495 35328 30559 35332
rect 30575 35388 30639 35392
rect 30575 35332 30579 35388
rect 30579 35332 30635 35388
rect 30635 35332 30639 35388
rect 30575 35328 30639 35332
rect 30655 35388 30719 35392
rect 30655 35332 30659 35388
rect 30659 35332 30715 35388
rect 30715 35332 30719 35388
rect 30655 35328 30719 35332
rect 30735 35388 30799 35392
rect 30735 35332 30739 35388
rect 30739 35332 30795 35388
rect 30795 35332 30799 35388
rect 30735 35328 30799 35332
rect 28948 35124 29012 35188
rect 9392 34844 9456 34848
rect 9392 34788 9396 34844
rect 9396 34788 9452 34844
rect 9452 34788 9456 34844
rect 9392 34784 9456 34788
rect 9472 34844 9536 34848
rect 9472 34788 9476 34844
rect 9476 34788 9532 34844
rect 9532 34788 9536 34844
rect 9472 34784 9536 34788
rect 9552 34844 9616 34848
rect 9552 34788 9556 34844
rect 9556 34788 9612 34844
rect 9612 34788 9616 34844
rect 9552 34784 9616 34788
rect 9632 34844 9696 34848
rect 9632 34788 9636 34844
rect 9636 34788 9692 34844
rect 9692 34788 9696 34844
rect 9632 34784 9696 34788
rect 17833 34844 17897 34848
rect 17833 34788 17837 34844
rect 17837 34788 17893 34844
rect 17893 34788 17897 34844
rect 17833 34784 17897 34788
rect 17913 34844 17977 34848
rect 17913 34788 17917 34844
rect 17917 34788 17973 34844
rect 17973 34788 17977 34844
rect 17913 34784 17977 34788
rect 17993 34844 18057 34848
rect 17993 34788 17997 34844
rect 17997 34788 18053 34844
rect 18053 34788 18057 34844
rect 17993 34784 18057 34788
rect 18073 34844 18137 34848
rect 18073 34788 18077 34844
rect 18077 34788 18133 34844
rect 18133 34788 18137 34844
rect 18073 34784 18137 34788
rect 26274 34844 26338 34848
rect 26274 34788 26278 34844
rect 26278 34788 26334 34844
rect 26334 34788 26338 34844
rect 26274 34784 26338 34788
rect 26354 34844 26418 34848
rect 26354 34788 26358 34844
rect 26358 34788 26414 34844
rect 26414 34788 26418 34844
rect 26354 34784 26418 34788
rect 26434 34844 26498 34848
rect 26434 34788 26438 34844
rect 26438 34788 26494 34844
rect 26494 34788 26498 34844
rect 26434 34784 26498 34788
rect 26514 34844 26578 34848
rect 26514 34788 26518 34844
rect 26518 34788 26574 34844
rect 26574 34788 26578 34844
rect 26514 34784 26578 34788
rect 34715 34844 34779 34848
rect 34715 34788 34719 34844
rect 34719 34788 34775 34844
rect 34775 34788 34779 34844
rect 34715 34784 34779 34788
rect 34795 34844 34859 34848
rect 34795 34788 34799 34844
rect 34799 34788 34855 34844
rect 34855 34788 34859 34844
rect 34795 34784 34859 34788
rect 34875 34844 34939 34848
rect 34875 34788 34879 34844
rect 34879 34788 34935 34844
rect 34935 34788 34939 34844
rect 34875 34784 34939 34788
rect 34955 34844 35019 34848
rect 34955 34788 34959 34844
rect 34959 34788 35015 34844
rect 35015 34788 35019 34844
rect 34955 34784 35019 34788
rect 23428 34580 23492 34644
rect 5172 34300 5236 34304
rect 5172 34244 5176 34300
rect 5176 34244 5232 34300
rect 5232 34244 5236 34300
rect 5172 34240 5236 34244
rect 5252 34300 5316 34304
rect 5252 34244 5256 34300
rect 5256 34244 5312 34300
rect 5312 34244 5316 34300
rect 5252 34240 5316 34244
rect 5332 34300 5396 34304
rect 5332 34244 5336 34300
rect 5336 34244 5392 34300
rect 5392 34244 5396 34300
rect 5332 34240 5396 34244
rect 5412 34300 5476 34304
rect 5412 34244 5416 34300
rect 5416 34244 5472 34300
rect 5472 34244 5476 34300
rect 5412 34240 5476 34244
rect 13613 34300 13677 34304
rect 13613 34244 13617 34300
rect 13617 34244 13673 34300
rect 13673 34244 13677 34300
rect 13613 34240 13677 34244
rect 13693 34300 13757 34304
rect 13693 34244 13697 34300
rect 13697 34244 13753 34300
rect 13753 34244 13757 34300
rect 13693 34240 13757 34244
rect 13773 34300 13837 34304
rect 13773 34244 13777 34300
rect 13777 34244 13833 34300
rect 13833 34244 13837 34300
rect 13773 34240 13837 34244
rect 13853 34300 13917 34304
rect 13853 34244 13857 34300
rect 13857 34244 13913 34300
rect 13913 34244 13917 34300
rect 13853 34240 13917 34244
rect 22054 34300 22118 34304
rect 22054 34244 22058 34300
rect 22058 34244 22114 34300
rect 22114 34244 22118 34300
rect 22054 34240 22118 34244
rect 22134 34300 22198 34304
rect 22134 34244 22138 34300
rect 22138 34244 22194 34300
rect 22194 34244 22198 34300
rect 22134 34240 22198 34244
rect 22214 34300 22278 34304
rect 22214 34244 22218 34300
rect 22218 34244 22274 34300
rect 22274 34244 22278 34300
rect 22214 34240 22278 34244
rect 22294 34300 22358 34304
rect 22294 34244 22298 34300
rect 22298 34244 22354 34300
rect 22354 34244 22358 34300
rect 22294 34240 22358 34244
rect 30495 34300 30559 34304
rect 30495 34244 30499 34300
rect 30499 34244 30555 34300
rect 30555 34244 30559 34300
rect 30495 34240 30559 34244
rect 30575 34300 30639 34304
rect 30575 34244 30579 34300
rect 30579 34244 30635 34300
rect 30635 34244 30639 34300
rect 30575 34240 30639 34244
rect 30655 34300 30719 34304
rect 30655 34244 30659 34300
rect 30659 34244 30715 34300
rect 30715 34244 30719 34300
rect 30655 34240 30719 34244
rect 30735 34300 30799 34304
rect 30735 34244 30739 34300
rect 30739 34244 30795 34300
rect 30795 34244 30799 34300
rect 30735 34240 30799 34244
rect 9392 33756 9456 33760
rect 9392 33700 9396 33756
rect 9396 33700 9452 33756
rect 9452 33700 9456 33756
rect 9392 33696 9456 33700
rect 9472 33756 9536 33760
rect 9472 33700 9476 33756
rect 9476 33700 9532 33756
rect 9532 33700 9536 33756
rect 9472 33696 9536 33700
rect 9552 33756 9616 33760
rect 9552 33700 9556 33756
rect 9556 33700 9612 33756
rect 9612 33700 9616 33756
rect 9552 33696 9616 33700
rect 9632 33756 9696 33760
rect 9632 33700 9636 33756
rect 9636 33700 9692 33756
rect 9692 33700 9696 33756
rect 9632 33696 9696 33700
rect 17833 33756 17897 33760
rect 17833 33700 17837 33756
rect 17837 33700 17893 33756
rect 17893 33700 17897 33756
rect 17833 33696 17897 33700
rect 17913 33756 17977 33760
rect 17913 33700 17917 33756
rect 17917 33700 17973 33756
rect 17973 33700 17977 33756
rect 17913 33696 17977 33700
rect 17993 33756 18057 33760
rect 17993 33700 17997 33756
rect 17997 33700 18053 33756
rect 18053 33700 18057 33756
rect 17993 33696 18057 33700
rect 18073 33756 18137 33760
rect 18073 33700 18077 33756
rect 18077 33700 18133 33756
rect 18133 33700 18137 33756
rect 18073 33696 18137 33700
rect 26274 33756 26338 33760
rect 26274 33700 26278 33756
rect 26278 33700 26334 33756
rect 26334 33700 26338 33756
rect 26274 33696 26338 33700
rect 26354 33756 26418 33760
rect 26354 33700 26358 33756
rect 26358 33700 26414 33756
rect 26414 33700 26418 33756
rect 26354 33696 26418 33700
rect 26434 33756 26498 33760
rect 26434 33700 26438 33756
rect 26438 33700 26494 33756
rect 26494 33700 26498 33756
rect 26434 33696 26498 33700
rect 26514 33756 26578 33760
rect 26514 33700 26518 33756
rect 26518 33700 26574 33756
rect 26574 33700 26578 33756
rect 26514 33696 26578 33700
rect 34715 33756 34779 33760
rect 34715 33700 34719 33756
rect 34719 33700 34775 33756
rect 34775 33700 34779 33756
rect 34715 33696 34779 33700
rect 34795 33756 34859 33760
rect 34795 33700 34799 33756
rect 34799 33700 34855 33756
rect 34855 33700 34859 33756
rect 34795 33696 34859 33700
rect 34875 33756 34939 33760
rect 34875 33700 34879 33756
rect 34879 33700 34935 33756
rect 34935 33700 34939 33756
rect 34875 33696 34939 33700
rect 34955 33756 35019 33760
rect 34955 33700 34959 33756
rect 34959 33700 35015 33756
rect 35015 33700 35019 33756
rect 34955 33696 35019 33700
rect 31524 33628 31588 33692
rect 28764 33492 28828 33556
rect 5172 33212 5236 33216
rect 5172 33156 5176 33212
rect 5176 33156 5232 33212
rect 5232 33156 5236 33212
rect 5172 33152 5236 33156
rect 5252 33212 5316 33216
rect 5252 33156 5256 33212
rect 5256 33156 5312 33212
rect 5312 33156 5316 33212
rect 5252 33152 5316 33156
rect 5332 33212 5396 33216
rect 5332 33156 5336 33212
rect 5336 33156 5392 33212
rect 5392 33156 5396 33212
rect 5332 33152 5396 33156
rect 5412 33212 5476 33216
rect 5412 33156 5416 33212
rect 5416 33156 5472 33212
rect 5472 33156 5476 33212
rect 5412 33152 5476 33156
rect 13613 33212 13677 33216
rect 13613 33156 13617 33212
rect 13617 33156 13673 33212
rect 13673 33156 13677 33212
rect 13613 33152 13677 33156
rect 13693 33212 13757 33216
rect 13693 33156 13697 33212
rect 13697 33156 13753 33212
rect 13753 33156 13757 33212
rect 13693 33152 13757 33156
rect 13773 33212 13837 33216
rect 13773 33156 13777 33212
rect 13777 33156 13833 33212
rect 13833 33156 13837 33212
rect 13773 33152 13837 33156
rect 13853 33212 13917 33216
rect 13853 33156 13857 33212
rect 13857 33156 13913 33212
rect 13913 33156 13917 33212
rect 13853 33152 13917 33156
rect 22054 33212 22118 33216
rect 22054 33156 22058 33212
rect 22058 33156 22114 33212
rect 22114 33156 22118 33212
rect 22054 33152 22118 33156
rect 22134 33212 22198 33216
rect 22134 33156 22138 33212
rect 22138 33156 22194 33212
rect 22194 33156 22198 33212
rect 22134 33152 22198 33156
rect 22214 33212 22278 33216
rect 22214 33156 22218 33212
rect 22218 33156 22274 33212
rect 22274 33156 22278 33212
rect 22214 33152 22278 33156
rect 22294 33212 22358 33216
rect 22294 33156 22298 33212
rect 22298 33156 22354 33212
rect 22354 33156 22358 33212
rect 22294 33152 22358 33156
rect 30495 33212 30559 33216
rect 30495 33156 30499 33212
rect 30499 33156 30555 33212
rect 30555 33156 30559 33212
rect 30495 33152 30559 33156
rect 30575 33212 30639 33216
rect 30575 33156 30579 33212
rect 30579 33156 30635 33212
rect 30635 33156 30639 33212
rect 30575 33152 30639 33156
rect 30655 33212 30719 33216
rect 30655 33156 30659 33212
rect 30659 33156 30715 33212
rect 30715 33156 30719 33212
rect 30655 33152 30719 33156
rect 30735 33212 30799 33216
rect 30735 33156 30739 33212
rect 30739 33156 30795 33212
rect 30795 33156 30799 33212
rect 30735 33152 30799 33156
rect 9392 32668 9456 32672
rect 9392 32612 9396 32668
rect 9396 32612 9452 32668
rect 9452 32612 9456 32668
rect 9392 32608 9456 32612
rect 9472 32668 9536 32672
rect 9472 32612 9476 32668
rect 9476 32612 9532 32668
rect 9532 32612 9536 32668
rect 9472 32608 9536 32612
rect 9552 32668 9616 32672
rect 9552 32612 9556 32668
rect 9556 32612 9612 32668
rect 9612 32612 9616 32668
rect 9552 32608 9616 32612
rect 9632 32668 9696 32672
rect 9632 32612 9636 32668
rect 9636 32612 9692 32668
rect 9692 32612 9696 32668
rect 9632 32608 9696 32612
rect 17833 32668 17897 32672
rect 17833 32612 17837 32668
rect 17837 32612 17893 32668
rect 17893 32612 17897 32668
rect 17833 32608 17897 32612
rect 17913 32668 17977 32672
rect 17913 32612 17917 32668
rect 17917 32612 17973 32668
rect 17973 32612 17977 32668
rect 17913 32608 17977 32612
rect 17993 32668 18057 32672
rect 17993 32612 17997 32668
rect 17997 32612 18053 32668
rect 18053 32612 18057 32668
rect 17993 32608 18057 32612
rect 18073 32668 18137 32672
rect 18073 32612 18077 32668
rect 18077 32612 18133 32668
rect 18133 32612 18137 32668
rect 18073 32608 18137 32612
rect 26274 32668 26338 32672
rect 26274 32612 26278 32668
rect 26278 32612 26334 32668
rect 26334 32612 26338 32668
rect 26274 32608 26338 32612
rect 26354 32668 26418 32672
rect 26354 32612 26358 32668
rect 26358 32612 26414 32668
rect 26414 32612 26418 32668
rect 26354 32608 26418 32612
rect 26434 32668 26498 32672
rect 26434 32612 26438 32668
rect 26438 32612 26494 32668
rect 26494 32612 26498 32668
rect 26434 32608 26498 32612
rect 26514 32668 26578 32672
rect 26514 32612 26518 32668
rect 26518 32612 26574 32668
rect 26574 32612 26578 32668
rect 26514 32608 26578 32612
rect 34715 32668 34779 32672
rect 34715 32612 34719 32668
rect 34719 32612 34775 32668
rect 34775 32612 34779 32668
rect 34715 32608 34779 32612
rect 34795 32668 34859 32672
rect 34795 32612 34799 32668
rect 34799 32612 34855 32668
rect 34855 32612 34859 32668
rect 34795 32608 34859 32612
rect 34875 32668 34939 32672
rect 34875 32612 34879 32668
rect 34879 32612 34935 32668
rect 34935 32612 34939 32668
rect 34875 32608 34939 32612
rect 34955 32668 35019 32672
rect 34955 32612 34959 32668
rect 34959 32612 35015 32668
rect 35015 32612 35019 32668
rect 34955 32608 35019 32612
rect 31156 32540 31220 32604
rect 5172 32124 5236 32128
rect 5172 32068 5176 32124
rect 5176 32068 5232 32124
rect 5232 32068 5236 32124
rect 5172 32064 5236 32068
rect 5252 32124 5316 32128
rect 5252 32068 5256 32124
rect 5256 32068 5312 32124
rect 5312 32068 5316 32124
rect 5252 32064 5316 32068
rect 5332 32124 5396 32128
rect 5332 32068 5336 32124
rect 5336 32068 5392 32124
rect 5392 32068 5396 32124
rect 5332 32064 5396 32068
rect 5412 32124 5476 32128
rect 5412 32068 5416 32124
rect 5416 32068 5472 32124
rect 5472 32068 5476 32124
rect 5412 32064 5476 32068
rect 13613 32124 13677 32128
rect 13613 32068 13617 32124
rect 13617 32068 13673 32124
rect 13673 32068 13677 32124
rect 13613 32064 13677 32068
rect 13693 32124 13757 32128
rect 13693 32068 13697 32124
rect 13697 32068 13753 32124
rect 13753 32068 13757 32124
rect 13693 32064 13757 32068
rect 13773 32124 13837 32128
rect 13773 32068 13777 32124
rect 13777 32068 13833 32124
rect 13833 32068 13837 32124
rect 13773 32064 13837 32068
rect 13853 32124 13917 32128
rect 13853 32068 13857 32124
rect 13857 32068 13913 32124
rect 13913 32068 13917 32124
rect 13853 32064 13917 32068
rect 22054 32124 22118 32128
rect 22054 32068 22058 32124
rect 22058 32068 22114 32124
rect 22114 32068 22118 32124
rect 22054 32064 22118 32068
rect 22134 32124 22198 32128
rect 22134 32068 22138 32124
rect 22138 32068 22194 32124
rect 22194 32068 22198 32124
rect 22134 32064 22198 32068
rect 22214 32124 22278 32128
rect 22214 32068 22218 32124
rect 22218 32068 22274 32124
rect 22274 32068 22278 32124
rect 22214 32064 22278 32068
rect 22294 32124 22358 32128
rect 22294 32068 22298 32124
rect 22298 32068 22354 32124
rect 22354 32068 22358 32124
rect 22294 32064 22358 32068
rect 30495 32124 30559 32128
rect 30495 32068 30499 32124
rect 30499 32068 30555 32124
rect 30555 32068 30559 32124
rect 30495 32064 30559 32068
rect 30575 32124 30639 32128
rect 30575 32068 30579 32124
rect 30579 32068 30635 32124
rect 30635 32068 30639 32124
rect 30575 32064 30639 32068
rect 30655 32124 30719 32128
rect 30655 32068 30659 32124
rect 30659 32068 30715 32124
rect 30715 32068 30719 32124
rect 30655 32064 30719 32068
rect 30735 32124 30799 32128
rect 30735 32068 30739 32124
rect 30739 32068 30795 32124
rect 30795 32068 30799 32124
rect 30735 32064 30799 32068
rect 9392 31580 9456 31584
rect 9392 31524 9396 31580
rect 9396 31524 9452 31580
rect 9452 31524 9456 31580
rect 9392 31520 9456 31524
rect 9472 31580 9536 31584
rect 9472 31524 9476 31580
rect 9476 31524 9532 31580
rect 9532 31524 9536 31580
rect 9472 31520 9536 31524
rect 9552 31580 9616 31584
rect 9552 31524 9556 31580
rect 9556 31524 9612 31580
rect 9612 31524 9616 31580
rect 9552 31520 9616 31524
rect 9632 31580 9696 31584
rect 9632 31524 9636 31580
rect 9636 31524 9692 31580
rect 9692 31524 9696 31580
rect 9632 31520 9696 31524
rect 17833 31580 17897 31584
rect 17833 31524 17837 31580
rect 17837 31524 17893 31580
rect 17893 31524 17897 31580
rect 17833 31520 17897 31524
rect 17913 31580 17977 31584
rect 17913 31524 17917 31580
rect 17917 31524 17973 31580
rect 17973 31524 17977 31580
rect 17913 31520 17977 31524
rect 17993 31580 18057 31584
rect 17993 31524 17997 31580
rect 17997 31524 18053 31580
rect 18053 31524 18057 31580
rect 17993 31520 18057 31524
rect 18073 31580 18137 31584
rect 18073 31524 18077 31580
rect 18077 31524 18133 31580
rect 18133 31524 18137 31580
rect 18073 31520 18137 31524
rect 26274 31580 26338 31584
rect 26274 31524 26278 31580
rect 26278 31524 26334 31580
rect 26334 31524 26338 31580
rect 26274 31520 26338 31524
rect 26354 31580 26418 31584
rect 26354 31524 26358 31580
rect 26358 31524 26414 31580
rect 26414 31524 26418 31580
rect 26354 31520 26418 31524
rect 26434 31580 26498 31584
rect 26434 31524 26438 31580
rect 26438 31524 26494 31580
rect 26494 31524 26498 31580
rect 26434 31520 26498 31524
rect 26514 31580 26578 31584
rect 26514 31524 26518 31580
rect 26518 31524 26574 31580
rect 26574 31524 26578 31580
rect 26514 31520 26578 31524
rect 34715 31580 34779 31584
rect 34715 31524 34719 31580
rect 34719 31524 34775 31580
rect 34775 31524 34779 31580
rect 34715 31520 34779 31524
rect 34795 31580 34859 31584
rect 34795 31524 34799 31580
rect 34799 31524 34855 31580
rect 34855 31524 34859 31580
rect 34795 31520 34859 31524
rect 34875 31580 34939 31584
rect 34875 31524 34879 31580
rect 34879 31524 34935 31580
rect 34935 31524 34939 31580
rect 34875 31520 34939 31524
rect 34955 31580 35019 31584
rect 34955 31524 34959 31580
rect 34959 31524 35015 31580
rect 35015 31524 35019 31580
rect 34955 31520 35019 31524
rect 29500 31104 29564 31108
rect 29500 31048 29514 31104
rect 29514 31048 29564 31104
rect 29500 31044 29564 31048
rect 5172 31036 5236 31040
rect 5172 30980 5176 31036
rect 5176 30980 5232 31036
rect 5232 30980 5236 31036
rect 5172 30976 5236 30980
rect 5252 31036 5316 31040
rect 5252 30980 5256 31036
rect 5256 30980 5312 31036
rect 5312 30980 5316 31036
rect 5252 30976 5316 30980
rect 5332 31036 5396 31040
rect 5332 30980 5336 31036
rect 5336 30980 5392 31036
rect 5392 30980 5396 31036
rect 5332 30976 5396 30980
rect 5412 31036 5476 31040
rect 5412 30980 5416 31036
rect 5416 30980 5472 31036
rect 5472 30980 5476 31036
rect 5412 30976 5476 30980
rect 13613 31036 13677 31040
rect 13613 30980 13617 31036
rect 13617 30980 13673 31036
rect 13673 30980 13677 31036
rect 13613 30976 13677 30980
rect 13693 31036 13757 31040
rect 13693 30980 13697 31036
rect 13697 30980 13753 31036
rect 13753 30980 13757 31036
rect 13693 30976 13757 30980
rect 13773 31036 13837 31040
rect 13773 30980 13777 31036
rect 13777 30980 13833 31036
rect 13833 30980 13837 31036
rect 13773 30976 13837 30980
rect 13853 31036 13917 31040
rect 13853 30980 13857 31036
rect 13857 30980 13913 31036
rect 13913 30980 13917 31036
rect 13853 30976 13917 30980
rect 22054 31036 22118 31040
rect 22054 30980 22058 31036
rect 22058 30980 22114 31036
rect 22114 30980 22118 31036
rect 22054 30976 22118 30980
rect 22134 31036 22198 31040
rect 22134 30980 22138 31036
rect 22138 30980 22194 31036
rect 22194 30980 22198 31036
rect 22134 30976 22198 30980
rect 22214 31036 22278 31040
rect 22214 30980 22218 31036
rect 22218 30980 22274 31036
rect 22274 30980 22278 31036
rect 22214 30976 22278 30980
rect 22294 31036 22358 31040
rect 22294 30980 22298 31036
rect 22298 30980 22354 31036
rect 22354 30980 22358 31036
rect 22294 30976 22358 30980
rect 30495 31036 30559 31040
rect 30495 30980 30499 31036
rect 30499 30980 30555 31036
rect 30555 30980 30559 31036
rect 30495 30976 30559 30980
rect 30575 31036 30639 31040
rect 30575 30980 30579 31036
rect 30579 30980 30635 31036
rect 30635 30980 30639 31036
rect 30575 30976 30639 30980
rect 30655 31036 30719 31040
rect 30655 30980 30659 31036
rect 30659 30980 30715 31036
rect 30715 30980 30719 31036
rect 30655 30976 30719 30980
rect 30735 31036 30799 31040
rect 30735 30980 30739 31036
rect 30739 30980 30795 31036
rect 30795 30980 30799 31036
rect 30735 30976 30799 30980
rect 9392 30492 9456 30496
rect 9392 30436 9396 30492
rect 9396 30436 9452 30492
rect 9452 30436 9456 30492
rect 9392 30432 9456 30436
rect 9472 30492 9536 30496
rect 9472 30436 9476 30492
rect 9476 30436 9532 30492
rect 9532 30436 9536 30492
rect 9472 30432 9536 30436
rect 9552 30492 9616 30496
rect 9552 30436 9556 30492
rect 9556 30436 9612 30492
rect 9612 30436 9616 30492
rect 9552 30432 9616 30436
rect 9632 30492 9696 30496
rect 9632 30436 9636 30492
rect 9636 30436 9692 30492
rect 9692 30436 9696 30492
rect 9632 30432 9696 30436
rect 17833 30492 17897 30496
rect 17833 30436 17837 30492
rect 17837 30436 17893 30492
rect 17893 30436 17897 30492
rect 17833 30432 17897 30436
rect 17913 30492 17977 30496
rect 17913 30436 17917 30492
rect 17917 30436 17973 30492
rect 17973 30436 17977 30492
rect 17913 30432 17977 30436
rect 17993 30492 18057 30496
rect 17993 30436 17997 30492
rect 17997 30436 18053 30492
rect 18053 30436 18057 30492
rect 17993 30432 18057 30436
rect 18073 30492 18137 30496
rect 18073 30436 18077 30492
rect 18077 30436 18133 30492
rect 18133 30436 18137 30492
rect 18073 30432 18137 30436
rect 26274 30492 26338 30496
rect 26274 30436 26278 30492
rect 26278 30436 26334 30492
rect 26334 30436 26338 30492
rect 26274 30432 26338 30436
rect 26354 30492 26418 30496
rect 26354 30436 26358 30492
rect 26358 30436 26414 30492
rect 26414 30436 26418 30492
rect 26354 30432 26418 30436
rect 26434 30492 26498 30496
rect 26434 30436 26438 30492
rect 26438 30436 26494 30492
rect 26494 30436 26498 30492
rect 26434 30432 26498 30436
rect 26514 30492 26578 30496
rect 26514 30436 26518 30492
rect 26518 30436 26574 30492
rect 26574 30436 26578 30492
rect 26514 30432 26578 30436
rect 34715 30492 34779 30496
rect 34715 30436 34719 30492
rect 34719 30436 34775 30492
rect 34775 30436 34779 30492
rect 34715 30432 34779 30436
rect 34795 30492 34859 30496
rect 34795 30436 34799 30492
rect 34799 30436 34855 30492
rect 34855 30436 34859 30492
rect 34795 30432 34859 30436
rect 34875 30492 34939 30496
rect 34875 30436 34879 30492
rect 34879 30436 34935 30492
rect 34935 30436 34939 30492
rect 34875 30432 34939 30436
rect 34955 30492 35019 30496
rect 34955 30436 34959 30492
rect 34959 30436 35015 30492
rect 35015 30436 35019 30492
rect 34955 30432 35019 30436
rect 5172 29948 5236 29952
rect 5172 29892 5176 29948
rect 5176 29892 5232 29948
rect 5232 29892 5236 29948
rect 5172 29888 5236 29892
rect 5252 29948 5316 29952
rect 5252 29892 5256 29948
rect 5256 29892 5312 29948
rect 5312 29892 5316 29948
rect 5252 29888 5316 29892
rect 5332 29948 5396 29952
rect 5332 29892 5336 29948
rect 5336 29892 5392 29948
rect 5392 29892 5396 29948
rect 5332 29888 5396 29892
rect 5412 29948 5476 29952
rect 5412 29892 5416 29948
rect 5416 29892 5472 29948
rect 5472 29892 5476 29948
rect 5412 29888 5476 29892
rect 13613 29948 13677 29952
rect 13613 29892 13617 29948
rect 13617 29892 13673 29948
rect 13673 29892 13677 29948
rect 13613 29888 13677 29892
rect 13693 29948 13757 29952
rect 13693 29892 13697 29948
rect 13697 29892 13753 29948
rect 13753 29892 13757 29948
rect 13693 29888 13757 29892
rect 13773 29948 13837 29952
rect 13773 29892 13777 29948
rect 13777 29892 13833 29948
rect 13833 29892 13837 29948
rect 13773 29888 13837 29892
rect 13853 29948 13917 29952
rect 13853 29892 13857 29948
rect 13857 29892 13913 29948
rect 13913 29892 13917 29948
rect 13853 29888 13917 29892
rect 22054 29948 22118 29952
rect 22054 29892 22058 29948
rect 22058 29892 22114 29948
rect 22114 29892 22118 29948
rect 22054 29888 22118 29892
rect 22134 29948 22198 29952
rect 22134 29892 22138 29948
rect 22138 29892 22194 29948
rect 22194 29892 22198 29948
rect 22134 29888 22198 29892
rect 22214 29948 22278 29952
rect 22214 29892 22218 29948
rect 22218 29892 22274 29948
rect 22274 29892 22278 29948
rect 22214 29888 22278 29892
rect 22294 29948 22358 29952
rect 22294 29892 22298 29948
rect 22298 29892 22354 29948
rect 22354 29892 22358 29948
rect 22294 29888 22358 29892
rect 30495 29948 30559 29952
rect 30495 29892 30499 29948
rect 30499 29892 30555 29948
rect 30555 29892 30559 29948
rect 30495 29888 30559 29892
rect 30575 29948 30639 29952
rect 30575 29892 30579 29948
rect 30579 29892 30635 29948
rect 30635 29892 30639 29948
rect 30575 29888 30639 29892
rect 30655 29948 30719 29952
rect 30655 29892 30659 29948
rect 30659 29892 30715 29948
rect 30715 29892 30719 29948
rect 30655 29888 30719 29892
rect 30735 29948 30799 29952
rect 30735 29892 30739 29948
rect 30739 29892 30795 29948
rect 30795 29892 30799 29948
rect 30735 29888 30799 29892
rect 27660 29820 27724 29884
rect 9392 29404 9456 29408
rect 9392 29348 9396 29404
rect 9396 29348 9452 29404
rect 9452 29348 9456 29404
rect 9392 29344 9456 29348
rect 9472 29404 9536 29408
rect 9472 29348 9476 29404
rect 9476 29348 9532 29404
rect 9532 29348 9536 29404
rect 9472 29344 9536 29348
rect 9552 29404 9616 29408
rect 9552 29348 9556 29404
rect 9556 29348 9612 29404
rect 9612 29348 9616 29404
rect 9552 29344 9616 29348
rect 9632 29404 9696 29408
rect 9632 29348 9636 29404
rect 9636 29348 9692 29404
rect 9692 29348 9696 29404
rect 9632 29344 9696 29348
rect 17833 29404 17897 29408
rect 17833 29348 17837 29404
rect 17837 29348 17893 29404
rect 17893 29348 17897 29404
rect 17833 29344 17897 29348
rect 17913 29404 17977 29408
rect 17913 29348 17917 29404
rect 17917 29348 17973 29404
rect 17973 29348 17977 29404
rect 17913 29344 17977 29348
rect 17993 29404 18057 29408
rect 17993 29348 17997 29404
rect 17997 29348 18053 29404
rect 18053 29348 18057 29404
rect 17993 29344 18057 29348
rect 18073 29404 18137 29408
rect 18073 29348 18077 29404
rect 18077 29348 18133 29404
rect 18133 29348 18137 29404
rect 18073 29344 18137 29348
rect 26274 29404 26338 29408
rect 26274 29348 26278 29404
rect 26278 29348 26334 29404
rect 26334 29348 26338 29404
rect 26274 29344 26338 29348
rect 26354 29404 26418 29408
rect 26354 29348 26358 29404
rect 26358 29348 26414 29404
rect 26414 29348 26418 29404
rect 26354 29344 26418 29348
rect 26434 29404 26498 29408
rect 26434 29348 26438 29404
rect 26438 29348 26494 29404
rect 26494 29348 26498 29404
rect 26434 29344 26498 29348
rect 26514 29404 26578 29408
rect 26514 29348 26518 29404
rect 26518 29348 26574 29404
rect 26574 29348 26578 29404
rect 26514 29344 26578 29348
rect 30236 29548 30300 29612
rect 34715 29404 34779 29408
rect 34715 29348 34719 29404
rect 34719 29348 34775 29404
rect 34775 29348 34779 29404
rect 34715 29344 34779 29348
rect 34795 29404 34859 29408
rect 34795 29348 34799 29404
rect 34799 29348 34855 29404
rect 34855 29348 34859 29404
rect 34795 29344 34859 29348
rect 34875 29404 34939 29408
rect 34875 29348 34879 29404
rect 34879 29348 34935 29404
rect 34935 29348 34939 29404
rect 34875 29344 34939 29348
rect 34955 29404 35019 29408
rect 34955 29348 34959 29404
rect 34959 29348 35015 29404
rect 35015 29348 35019 29404
rect 34955 29344 35019 29348
rect 32260 29140 32324 29204
rect 5172 28860 5236 28864
rect 5172 28804 5176 28860
rect 5176 28804 5232 28860
rect 5232 28804 5236 28860
rect 5172 28800 5236 28804
rect 5252 28860 5316 28864
rect 5252 28804 5256 28860
rect 5256 28804 5312 28860
rect 5312 28804 5316 28860
rect 5252 28800 5316 28804
rect 5332 28860 5396 28864
rect 5332 28804 5336 28860
rect 5336 28804 5392 28860
rect 5392 28804 5396 28860
rect 5332 28800 5396 28804
rect 5412 28860 5476 28864
rect 5412 28804 5416 28860
rect 5416 28804 5472 28860
rect 5472 28804 5476 28860
rect 5412 28800 5476 28804
rect 13613 28860 13677 28864
rect 13613 28804 13617 28860
rect 13617 28804 13673 28860
rect 13673 28804 13677 28860
rect 13613 28800 13677 28804
rect 13693 28860 13757 28864
rect 13693 28804 13697 28860
rect 13697 28804 13753 28860
rect 13753 28804 13757 28860
rect 13693 28800 13757 28804
rect 13773 28860 13837 28864
rect 13773 28804 13777 28860
rect 13777 28804 13833 28860
rect 13833 28804 13837 28860
rect 13773 28800 13837 28804
rect 13853 28860 13917 28864
rect 13853 28804 13857 28860
rect 13857 28804 13913 28860
rect 13913 28804 13917 28860
rect 13853 28800 13917 28804
rect 22054 28860 22118 28864
rect 22054 28804 22058 28860
rect 22058 28804 22114 28860
rect 22114 28804 22118 28860
rect 22054 28800 22118 28804
rect 22134 28860 22198 28864
rect 22134 28804 22138 28860
rect 22138 28804 22194 28860
rect 22194 28804 22198 28860
rect 22134 28800 22198 28804
rect 22214 28860 22278 28864
rect 22214 28804 22218 28860
rect 22218 28804 22274 28860
rect 22274 28804 22278 28860
rect 22214 28800 22278 28804
rect 22294 28860 22358 28864
rect 22294 28804 22298 28860
rect 22298 28804 22354 28860
rect 22354 28804 22358 28860
rect 22294 28800 22358 28804
rect 30495 28860 30559 28864
rect 30495 28804 30499 28860
rect 30499 28804 30555 28860
rect 30555 28804 30559 28860
rect 30495 28800 30559 28804
rect 30575 28860 30639 28864
rect 30575 28804 30579 28860
rect 30579 28804 30635 28860
rect 30635 28804 30639 28860
rect 30575 28800 30639 28804
rect 30655 28860 30719 28864
rect 30655 28804 30659 28860
rect 30659 28804 30715 28860
rect 30715 28804 30719 28860
rect 30655 28800 30719 28804
rect 30735 28860 30799 28864
rect 30735 28804 30739 28860
rect 30739 28804 30795 28860
rect 30795 28804 30799 28860
rect 30735 28800 30799 28804
rect 23428 28596 23492 28660
rect 9392 28316 9456 28320
rect 9392 28260 9396 28316
rect 9396 28260 9452 28316
rect 9452 28260 9456 28316
rect 9392 28256 9456 28260
rect 9472 28316 9536 28320
rect 9472 28260 9476 28316
rect 9476 28260 9532 28316
rect 9532 28260 9536 28316
rect 9472 28256 9536 28260
rect 9552 28316 9616 28320
rect 9552 28260 9556 28316
rect 9556 28260 9612 28316
rect 9612 28260 9616 28316
rect 9552 28256 9616 28260
rect 9632 28316 9696 28320
rect 9632 28260 9636 28316
rect 9636 28260 9692 28316
rect 9692 28260 9696 28316
rect 9632 28256 9696 28260
rect 17833 28316 17897 28320
rect 17833 28260 17837 28316
rect 17837 28260 17893 28316
rect 17893 28260 17897 28316
rect 17833 28256 17897 28260
rect 17913 28316 17977 28320
rect 17913 28260 17917 28316
rect 17917 28260 17973 28316
rect 17973 28260 17977 28316
rect 17913 28256 17977 28260
rect 17993 28316 18057 28320
rect 17993 28260 17997 28316
rect 17997 28260 18053 28316
rect 18053 28260 18057 28316
rect 17993 28256 18057 28260
rect 18073 28316 18137 28320
rect 18073 28260 18077 28316
rect 18077 28260 18133 28316
rect 18133 28260 18137 28316
rect 18073 28256 18137 28260
rect 26274 28316 26338 28320
rect 26274 28260 26278 28316
rect 26278 28260 26334 28316
rect 26334 28260 26338 28316
rect 26274 28256 26338 28260
rect 26354 28316 26418 28320
rect 26354 28260 26358 28316
rect 26358 28260 26414 28316
rect 26414 28260 26418 28316
rect 26354 28256 26418 28260
rect 26434 28316 26498 28320
rect 26434 28260 26438 28316
rect 26438 28260 26494 28316
rect 26494 28260 26498 28316
rect 26434 28256 26498 28260
rect 26514 28316 26578 28320
rect 26514 28260 26518 28316
rect 26518 28260 26574 28316
rect 26574 28260 26578 28316
rect 26514 28256 26578 28260
rect 34715 28316 34779 28320
rect 34715 28260 34719 28316
rect 34719 28260 34775 28316
rect 34775 28260 34779 28316
rect 34715 28256 34779 28260
rect 34795 28316 34859 28320
rect 34795 28260 34799 28316
rect 34799 28260 34855 28316
rect 34855 28260 34859 28316
rect 34795 28256 34859 28260
rect 34875 28316 34939 28320
rect 34875 28260 34879 28316
rect 34879 28260 34935 28316
rect 34935 28260 34939 28316
rect 34875 28256 34939 28260
rect 34955 28316 35019 28320
rect 34955 28260 34959 28316
rect 34959 28260 35015 28316
rect 35015 28260 35019 28316
rect 34955 28256 35019 28260
rect 29132 28112 29196 28116
rect 29132 28056 29146 28112
rect 29146 28056 29196 28112
rect 29132 28052 29196 28056
rect 5172 27772 5236 27776
rect 5172 27716 5176 27772
rect 5176 27716 5232 27772
rect 5232 27716 5236 27772
rect 5172 27712 5236 27716
rect 5252 27772 5316 27776
rect 5252 27716 5256 27772
rect 5256 27716 5312 27772
rect 5312 27716 5316 27772
rect 5252 27712 5316 27716
rect 5332 27772 5396 27776
rect 5332 27716 5336 27772
rect 5336 27716 5392 27772
rect 5392 27716 5396 27772
rect 5332 27712 5396 27716
rect 5412 27772 5476 27776
rect 5412 27716 5416 27772
rect 5416 27716 5472 27772
rect 5472 27716 5476 27772
rect 5412 27712 5476 27716
rect 13613 27772 13677 27776
rect 13613 27716 13617 27772
rect 13617 27716 13673 27772
rect 13673 27716 13677 27772
rect 13613 27712 13677 27716
rect 13693 27772 13757 27776
rect 13693 27716 13697 27772
rect 13697 27716 13753 27772
rect 13753 27716 13757 27772
rect 13693 27712 13757 27716
rect 13773 27772 13837 27776
rect 13773 27716 13777 27772
rect 13777 27716 13833 27772
rect 13833 27716 13837 27772
rect 13773 27712 13837 27716
rect 13853 27772 13917 27776
rect 13853 27716 13857 27772
rect 13857 27716 13913 27772
rect 13913 27716 13917 27772
rect 13853 27712 13917 27716
rect 22054 27772 22118 27776
rect 22054 27716 22058 27772
rect 22058 27716 22114 27772
rect 22114 27716 22118 27772
rect 22054 27712 22118 27716
rect 22134 27772 22198 27776
rect 22134 27716 22138 27772
rect 22138 27716 22194 27772
rect 22194 27716 22198 27772
rect 22134 27712 22198 27716
rect 22214 27772 22278 27776
rect 22214 27716 22218 27772
rect 22218 27716 22274 27772
rect 22274 27716 22278 27772
rect 22214 27712 22278 27716
rect 22294 27772 22358 27776
rect 22294 27716 22298 27772
rect 22298 27716 22354 27772
rect 22354 27716 22358 27772
rect 22294 27712 22358 27716
rect 30495 27772 30559 27776
rect 30495 27716 30499 27772
rect 30499 27716 30555 27772
rect 30555 27716 30559 27772
rect 30495 27712 30559 27716
rect 30575 27772 30639 27776
rect 30575 27716 30579 27772
rect 30579 27716 30635 27772
rect 30635 27716 30639 27772
rect 30575 27712 30639 27716
rect 30655 27772 30719 27776
rect 30655 27716 30659 27772
rect 30659 27716 30715 27772
rect 30715 27716 30719 27772
rect 30655 27712 30719 27716
rect 30735 27772 30799 27776
rect 30735 27716 30739 27772
rect 30739 27716 30795 27772
rect 30795 27716 30799 27772
rect 30735 27712 30799 27716
rect 32076 27568 32140 27572
rect 32076 27512 32090 27568
rect 32090 27512 32140 27568
rect 32076 27508 32140 27512
rect 9392 27228 9456 27232
rect 9392 27172 9396 27228
rect 9396 27172 9452 27228
rect 9452 27172 9456 27228
rect 9392 27168 9456 27172
rect 9472 27228 9536 27232
rect 9472 27172 9476 27228
rect 9476 27172 9532 27228
rect 9532 27172 9536 27228
rect 9472 27168 9536 27172
rect 9552 27228 9616 27232
rect 9552 27172 9556 27228
rect 9556 27172 9612 27228
rect 9612 27172 9616 27228
rect 9552 27168 9616 27172
rect 9632 27228 9696 27232
rect 9632 27172 9636 27228
rect 9636 27172 9692 27228
rect 9692 27172 9696 27228
rect 9632 27168 9696 27172
rect 17833 27228 17897 27232
rect 17833 27172 17837 27228
rect 17837 27172 17893 27228
rect 17893 27172 17897 27228
rect 17833 27168 17897 27172
rect 17913 27228 17977 27232
rect 17913 27172 17917 27228
rect 17917 27172 17973 27228
rect 17973 27172 17977 27228
rect 17913 27168 17977 27172
rect 17993 27228 18057 27232
rect 17993 27172 17997 27228
rect 17997 27172 18053 27228
rect 18053 27172 18057 27228
rect 17993 27168 18057 27172
rect 18073 27228 18137 27232
rect 18073 27172 18077 27228
rect 18077 27172 18133 27228
rect 18133 27172 18137 27228
rect 18073 27168 18137 27172
rect 26274 27228 26338 27232
rect 26274 27172 26278 27228
rect 26278 27172 26334 27228
rect 26334 27172 26338 27228
rect 26274 27168 26338 27172
rect 26354 27228 26418 27232
rect 26354 27172 26358 27228
rect 26358 27172 26414 27228
rect 26414 27172 26418 27228
rect 26354 27168 26418 27172
rect 26434 27228 26498 27232
rect 26434 27172 26438 27228
rect 26438 27172 26494 27228
rect 26494 27172 26498 27228
rect 26434 27168 26498 27172
rect 26514 27228 26578 27232
rect 26514 27172 26518 27228
rect 26518 27172 26574 27228
rect 26574 27172 26578 27228
rect 26514 27168 26578 27172
rect 34715 27228 34779 27232
rect 34715 27172 34719 27228
rect 34719 27172 34775 27228
rect 34775 27172 34779 27228
rect 34715 27168 34779 27172
rect 34795 27228 34859 27232
rect 34795 27172 34799 27228
rect 34799 27172 34855 27228
rect 34855 27172 34859 27228
rect 34795 27168 34859 27172
rect 34875 27228 34939 27232
rect 34875 27172 34879 27228
rect 34879 27172 34935 27228
rect 34935 27172 34939 27228
rect 34875 27168 34939 27172
rect 34955 27228 35019 27232
rect 34955 27172 34959 27228
rect 34959 27172 35015 27228
rect 35015 27172 35019 27228
rect 34955 27168 35019 27172
rect 5172 26684 5236 26688
rect 5172 26628 5176 26684
rect 5176 26628 5232 26684
rect 5232 26628 5236 26684
rect 5172 26624 5236 26628
rect 5252 26684 5316 26688
rect 5252 26628 5256 26684
rect 5256 26628 5312 26684
rect 5312 26628 5316 26684
rect 5252 26624 5316 26628
rect 5332 26684 5396 26688
rect 5332 26628 5336 26684
rect 5336 26628 5392 26684
rect 5392 26628 5396 26684
rect 5332 26624 5396 26628
rect 5412 26684 5476 26688
rect 5412 26628 5416 26684
rect 5416 26628 5472 26684
rect 5472 26628 5476 26684
rect 5412 26624 5476 26628
rect 13613 26684 13677 26688
rect 13613 26628 13617 26684
rect 13617 26628 13673 26684
rect 13673 26628 13677 26684
rect 13613 26624 13677 26628
rect 13693 26684 13757 26688
rect 13693 26628 13697 26684
rect 13697 26628 13753 26684
rect 13753 26628 13757 26684
rect 13693 26624 13757 26628
rect 13773 26684 13837 26688
rect 13773 26628 13777 26684
rect 13777 26628 13833 26684
rect 13833 26628 13837 26684
rect 13773 26624 13837 26628
rect 13853 26684 13917 26688
rect 13853 26628 13857 26684
rect 13857 26628 13913 26684
rect 13913 26628 13917 26684
rect 13853 26624 13917 26628
rect 22054 26684 22118 26688
rect 22054 26628 22058 26684
rect 22058 26628 22114 26684
rect 22114 26628 22118 26684
rect 22054 26624 22118 26628
rect 22134 26684 22198 26688
rect 22134 26628 22138 26684
rect 22138 26628 22194 26684
rect 22194 26628 22198 26684
rect 22134 26624 22198 26628
rect 22214 26684 22278 26688
rect 22214 26628 22218 26684
rect 22218 26628 22274 26684
rect 22274 26628 22278 26684
rect 22214 26624 22278 26628
rect 22294 26684 22358 26688
rect 22294 26628 22298 26684
rect 22298 26628 22354 26684
rect 22354 26628 22358 26684
rect 22294 26624 22358 26628
rect 30495 26684 30559 26688
rect 30495 26628 30499 26684
rect 30499 26628 30555 26684
rect 30555 26628 30559 26684
rect 30495 26624 30559 26628
rect 30575 26684 30639 26688
rect 30575 26628 30579 26684
rect 30579 26628 30635 26684
rect 30635 26628 30639 26684
rect 30575 26624 30639 26628
rect 30655 26684 30719 26688
rect 30655 26628 30659 26684
rect 30659 26628 30715 26684
rect 30715 26628 30719 26684
rect 30655 26624 30719 26628
rect 30735 26684 30799 26688
rect 30735 26628 30739 26684
rect 30739 26628 30795 26684
rect 30795 26628 30799 26684
rect 30735 26624 30799 26628
rect 9392 26140 9456 26144
rect 9392 26084 9396 26140
rect 9396 26084 9452 26140
rect 9452 26084 9456 26140
rect 9392 26080 9456 26084
rect 9472 26140 9536 26144
rect 9472 26084 9476 26140
rect 9476 26084 9532 26140
rect 9532 26084 9536 26140
rect 9472 26080 9536 26084
rect 9552 26140 9616 26144
rect 9552 26084 9556 26140
rect 9556 26084 9612 26140
rect 9612 26084 9616 26140
rect 9552 26080 9616 26084
rect 9632 26140 9696 26144
rect 9632 26084 9636 26140
rect 9636 26084 9692 26140
rect 9692 26084 9696 26140
rect 9632 26080 9696 26084
rect 17833 26140 17897 26144
rect 17833 26084 17837 26140
rect 17837 26084 17893 26140
rect 17893 26084 17897 26140
rect 17833 26080 17897 26084
rect 17913 26140 17977 26144
rect 17913 26084 17917 26140
rect 17917 26084 17973 26140
rect 17973 26084 17977 26140
rect 17913 26080 17977 26084
rect 17993 26140 18057 26144
rect 17993 26084 17997 26140
rect 17997 26084 18053 26140
rect 18053 26084 18057 26140
rect 17993 26080 18057 26084
rect 18073 26140 18137 26144
rect 18073 26084 18077 26140
rect 18077 26084 18133 26140
rect 18133 26084 18137 26140
rect 18073 26080 18137 26084
rect 26274 26140 26338 26144
rect 26274 26084 26278 26140
rect 26278 26084 26334 26140
rect 26334 26084 26338 26140
rect 26274 26080 26338 26084
rect 26354 26140 26418 26144
rect 26354 26084 26358 26140
rect 26358 26084 26414 26140
rect 26414 26084 26418 26140
rect 26354 26080 26418 26084
rect 26434 26140 26498 26144
rect 26434 26084 26438 26140
rect 26438 26084 26494 26140
rect 26494 26084 26498 26140
rect 26434 26080 26498 26084
rect 26514 26140 26578 26144
rect 26514 26084 26518 26140
rect 26518 26084 26574 26140
rect 26574 26084 26578 26140
rect 26514 26080 26578 26084
rect 34715 26140 34779 26144
rect 34715 26084 34719 26140
rect 34719 26084 34775 26140
rect 34775 26084 34779 26140
rect 34715 26080 34779 26084
rect 34795 26140 34859 26144
rect 34795 26084 34799 26140
rect 34799 26084 34855 26140
rect 34855 26084 34859 26140
rect 34795 26080 34859 26084
rect 34875 26140 34939 26144
rect 34875 26084 34879 26140
rect 34879 26084 34935 26140
rect 34935 26084 34939 26140
rect 34875 26080 34939 26084
rect 34955 26140 35019 26144
rect 34955 26084 34959 26140
rect 34959 26084 35015 26140
rect 35015 26084 35019 26140
rect 34955 26080 35019 26084
rect 5172 25596 5236 25600
rect 5172 25540 5176 25596
rect 5176 25540 5232 25596
rect 5232 25540 5236 25596
rect 5172 25536 5236 25540
rect 5252 25596 5316 25600
rect 5252 25540 5256 25596
rect 5256 25540 5312 25596
rect 5312 25540 5316 25596
rect 5252 25536 5316 25540
rect 5332 25596 5396 25600
rect 5332 25540 5336 25596
rect 5336 25540 5392 25596
rect 5392 25540 5396 25596
rect 5332 25536 5396 25540
rect 5412 25596 5476 25600
rect 5412 25540 5416 25596
rect 5416 25540 5472 25596
rect 5472 25540 5476 25596
rect 5412 25536 5476 25540
rect 13613 25596 13677 25600
rect 13613 25540 13617 25596
rect 13617 25540 13673 25596
rect 13673 25540 13677 25596
rect 13613 25536 13677 25540
rect 13693 25596 13757 25600
rect 13693 25540 13697 25596
rect 13697 25540 13753 25596
rect 13753 25540 13757 25596
rect 13693 25536 13757 25540
rect 13773 25596 13837 25600
rect 13773 25540 13777 25596
rect 13777 25540 13833 25596
rect 13833 25540 13837 25596
rect 13773 25536 13837 25540
rect 13853 25596 13917 25600
rect 13853 25540 13857 25596
rect 13857 25540 13913 25596
rect 13913 25540 13917 25596
rect 13853 25536 13917 25540
rect 22054 25596 22118 25600
rect 22054 25540 22058 25596
rect 22058 25540 22114 25596
rect 22114 25540 22118 25596
rect 22054 25536 22118 25540
rect 22134 25596 22198 25600
rect 22134 25540 22138 25596
rect 22138 25540 22194 25596
rect 22194 25540 22198 25596
rect 22134 25536 22198 25540
rect 22214 25596 22278 25600
rect 22214 25540 22218 25596
rect 22218 25540 22274 25596
rect 22274 25540 22278 25596
rect 22214 25536 22278 25540
rect 22294 25596 22358 25600
rect 22294 25540 22298 25596
rect 22298 25540 22354 25596
rect 22354 25540 22358 25596
rect 22294 25536 22358 25540
rect 30495 25596 30559 25600
rect 30495 25540 30499 25596
rect 30499 25540 30555 25596
rect 30555 25540 30559 25596
rect 30495 25536 30559 25540
rect 30575 25596 30639 25600
rect 30575 25540 30579 25596
rect 30579 25540 30635 25596
rect 30635 25540 30639 25596
rect 30575 25536 30639 25540
rect 30655 25596 30719 25600
rect 30655 25540 30659 25596
rect 30659 25540 30715 25596
rect 30715 25540 30719 25596
rect 30655 25536 30719 25540
rect 30735 25596 30799 25600
rect 30735 25540 30739 25596
rect 30739 25540 30795 25596
rect 30795 25540 30799 25596
rect 30735 25536 30799 25540
rect 9392 25052 9456 25056
rect 9392 24996 9396 25052
rect 9396 24996 9452 25052
rect 9452 24996 9456 25052
rect 9392 24992 9456 24996
rect 9472 25052 9536 25056
rect 9472 24996 9476 25052
rect 9476 24996 9532 25052
rect 9532 24996 9536 25052
rect 9472 24992 9536 24996
rect 9552 25052 9616 25056
rect 9552 24996 9556 25052
rect 9556 24996 9612 25052
rect 9612 24996 9616 25052
rect 9552 24992 9616 24996
rect 9632 25052 9696 25056
rect 9632 24996 9636 25052
rect 9636 24996 9692 25052
rect 9692 24996 9696 25052
rect 9632 24992 9696 24996
rect 17833 25052 17897 25056
rect 17833 24996 17837 25052
rect 17837 24996 17893 25052
rect 17893 24996 17897 25052
rect 17833 24992 17897 24996
rect 17913 25052 17977 25056
rect 17913 24996 17917 25052
rect 17917 24996 17973 25052
rect 17973 24996 17977 25052
rect 17913 24992 17977 24996
rect 17993 25052 18057 25056
rect 17993 24996 17997 25052
rect 17997 24996 18053 25052
rect 18053 24996 18057 25052
rect 17993 24992 18057 24996
rect 18073 25052 18137 25056
rect 18073 24996 18077 25052
rect 18077 24996 18133 25052
rect 18133 24996 18137 25052
rect 18073 24992 18137 24996
rect 26274 25052 26338 25056
rect 26274 24996 26278 25052
rect 26278 24996 26334 25052
rect 26334 24996 26338 25052
rect 26274 24992 26338 24996
rect 26354 25052 26418 25056
rect 26354 24996 26358 25052
rect 26358 24996 26414 25052
rect 26414 24996 26418 25052
rect 26354 24992 26418 24996
rect 26434 25052 26498 25056
rect 26434 24996 26438 25052
rect 26438 24996 26494 25052
rect 26494 24996 26498 25052
rect 26434 24992 26498 24996
rect 26514 25052 26578 25056
rect 26514 24996 26518 25052
rect 26518 24996 26574 25052
rect 26574 24996 26578 25052
rect 26514 24992 26578 24996
rect 34715 25052 34779 25056
rect 34715 24996 34719 25052
rect 34719 24996 34775 25052
rect 34775 24996 34779 25052
rect 34715 24992 34779 24996
rect 34795 25052 34859 25056
rect 34795 24996 34799 25052
rect 34799 24996 34855 25052
rect 34855 24996 34859 25052
rect 34795 24992 34859 24996
rect 34875 25052 34939 25056
rect 34875 24996 34879 25052
rect 34879 24996 34935 25052
rect 34935 24996 34939 25052
rect 34875 24992 34939 24996
rect 34955 25052 35019 25056
rect 34955 24996 34959 25052
rect 34959 24996 35015 25052
rect 35015 24996 35019 25052
rect 34955 24992 35019 24996
rect 31524 24984 31588 24988
rect 31524 24928 31538 24984
rect 31538 24928 31588 24984
rect 31524 24924 31588 24928
rect 31340 24652 31404 24716
rect 32812 24652 32876 24716
rect 5172 24508 5236 24512
rect 5172 24452 5176 24508
rect 5176 24452 5232 24508
rect 5232 24452 5236 24508
rect 5172 24448 5236 24452
rect 5252 24508 5316 24512
rect 5252 24452 5256 24508
rect 5256 24452 5312 24508
rect 5312 24452 5316 24508
rect 5252 24448 5316 24452
rect 5332 24508 5396 24512
rect 5332 24452 5336 24508
rect 5336 24452 5392 24508
rect 5392 24452 5396 24508
rect 5332 24448 5396 24452
rect 5412 24508 5476 24512
rect 5412 24452 5416 24508
rect 5416 24452 5472 24508
rect 5472 24452 5476 24508
rect 5412 24448 5476 24452
rect 13613 24508 13677 24512
rect 13613 24452 13617 24508
rect 13617 24452 13673 24508
rect 13673 24452 13677 24508
rect 13613 24448 13677 24452
rect 13693 24508 13757 24512
rect 13693 24452 13697 24508
rect 13697 24452 13753 24508
rect 13753 24452 13757 24508
rect 13693 24448 13757 24452
rect 13773 24508 13837 24512
rect 13773 24452 13777 24508
rect 13777 24452 13833 24508
rect 13833 24452 13837 24508
rect 13773 24448 13837 24452
rect 13853 24508 13917 24512
rect 13853 24452 13857 24508
rect 13857 24452 13913 24508
rect 13913 24452 13917 24508
rect 13853 24448 13917 24452
rect 22054 24508 22118 24512
rect 22054 24452 22058 24508
rect 22058 24452 22114 24508
rect 22114 24452 22118 24508
rect 22054 24448 22118 24452
rect 22134 24508 22198 24512
rect 22134 24452 22138 24508
rect 22138 24452 22194 24508
rect 22194 24452 22198 24508
rect 22134 24448 22198 24452
rect 22214 24508 22278 24512
rect 22214 24452 22218 24508
rect 22218 24452 22274 24508
rect 22274 24452 22278 24508
rect 22214 24448 22278 24452
rect 22294 24508 22358 24512
rect 22294 24452 22298 24508
rect 22298 24452 22354 24508
rect 22354 24452 22358 24508
rect 22294 24448 22358 24452
rect 30495 24508 30559 24512
rect 30495 24452 30499 24508
rect 30499 24452 30555 24508
rect 30555 24452 30559 24508
rect 30495 24448 30559 24452
rect 30575 24508 30639 24512
rect 30575 24452 30579 24508
rect 30579 24452 30635 24508
rect 30635 24452 30639 24508
rect 30575 24448 30639 24452
rect 30655 24508 30719 24512
rect 30655 24452 30659 24508
rect 30659 24452 30715 24508
rect 30715 24452 30719 24508
rect 30655 24448 30719 24452
rect 30735 24508 30799 24512
rect 30735 24452 30739 24508
rect 30739 24452 30795 24508
rect 30795 24452 30799 24508
rect 30735 24448 30799 24452
rect 9392 23964 9456 23968
rect 9392 23908 9396 23964
rect 9396 23908 9452 23964
rect 9452 23908 9456 23964
rect 9392 23904 9456 23908
rect 9472 23964 9536 23968
rect 9472 23908 9476 23964
rect 9476 23908 9532 23964
rect 9532 23908 9536 23964
rect 9472 23904 9536 23908
rect 9552 23964 9616 23968
rect 9552 23908 9556 23964
rect 9556 23908 9612 23964
rect 9612 23908 9616 23964
rect 9552 23904 9616 23908
rect 9632 23964 9696 23968
rect 9632 23908 9636 23964
rect 9636 23908 9692 23964
rect 9692 23908 9696 23964
rect 9632 23904 9696 23908
rect 17833 23964 17897 23968
rect 17833 23908 17837 23964
rect 17837 23908 17893 23964
rect 17893 23908 17897 23964
rect 17833 23904 17897 23908
rect 17913 23964 17977 23968
rect 17913 23908 17917 23964
rect 17917 23908 17973 23964
rect 17973 23908 17977 23964
rect 17913 23904 17977 23908
rect 17993 23964 18057 23968
rect 17993 23908 17997 23964
rect 17997 23908 18053 23964
rect 18053 23908 18057 23964
rect 17993 23904 18057 23908
rect 18073 23964 18137 23968
rect 18073 23908 18077 23964
rect 18077 23908 18133 23964
rect 18133 23908 18137 23964
rect 18073 23904 18137 23908
rect 26274 23964 26338 23968
rect 26274 23908 26278 23964
rect 26278 23908 26334 23964
rect 26334 23908 26338 23964
rect 26274 23904 26338 23908
rect 26354 23964 26418 23968
rect 26354 23908 26358 23964
rect 26358 23908 26414 23964
rect 26414 23908 26418 23964
rect 26354 23904 26418 23908
rect 26434 23964 26498 23968
rect 26434 23908 26438 23964
rect 26438 23908 26494 23964
rect 26494 23908 26498 23964
rect 26434 23904 26498 23908
rect 26514 23964 26578 23968
rect 26514 23908 26518 23964
rect 26518 23908 26574 23964
rect 26574 23908 26578 23964
rect 26514 23904 26578 23908
rect 34715 23964 34779 23968
rect 34715 23908 34719 23964
rect 34719 23908 34775 23964
rect 34775 23908 34779 23964
rect 34715 23904 34779 23908
rect 34795 23964 34859 23968
rect 34795 23908 34799 23964
rect 34799 23908 34855 23964
rect 34855 23908 34859 23964
rect 34795 23904 34859 23908
rect 34875 23964 34939 23968
rect 34875 23908 34879 23964
rect 34879 23908 34935 23964
rect 34935 23908 34939 23964
rect 34875 23904 34939 23908
rect 34955 23964 35019 23968
rect 34955 23908 34959 23964
rect 34959 23908 35015 23964
rect 35015 23908 35019 23964
rect 34955 23904 35019 23908
rect 33732 23836 33796 23900
rect 31892 23700 31956 23764
rect 29500 23564 29564 23628
rect 26740 23428 26804 23492
rect 33916 23428 33980 23492
rect 5172 23420 5236 23424
rect 5172 23364 5176 23420
rect 5176 23364 5232 23420
rect 5232 23364 5236 23420
rect 5172 23360 5236 23364
rect 5252 23420 5316 23424
rect 5252 23364 5256 23420
rect 5256 23364 5312 23420
rect 5312 23364 5316 23420
rect 5252 23360 5316 23364
rect 5332 23420 5396 23424
rect 5332 23364 5336 23420
rect 5336 23364 5392 23420
rect 5392 23364 5396 23420
rect 5332 23360 5396 23364
rect 5412 23420 5476 23424
rect 5412 23364 5416 23420
rect 5416 23364 5472 23420
rect 5472 23364 5476 23420
rect 5412 23360 5476 23364
rect 13613 23420 13677 23424
rect 13613 23364 13617 23420
rect 13617 23364 13673 23420
rect 13673 23364 13677 23420
rect 13613 23360 13677 23364
rect 13693 23420 13757 23424
rect 13693 23364 13697 23420
rect 13697 23364 13753 23420
rect 13753 23364 13757 23420
rect 13693 23360 13757 23364
rect 13773 23420 13837 23424
rect 13773 23364 13777 23420
rect 13777 23364 13833 23420
rect 13833 23364 13837 23420
rect 13773 23360 13837 23364
rect 13853 23420 13917 23424
rect 13853 23364 13857 23420
rect 13857 23364 13913 23420
rect 13913 23364 13917 23420
rect 13853 23360 13917 23364
rect 22054 23420 22118 23424
rect 22054 23364 22058 23420
rect 22058 23364 22114 23420
rect 22114 23364 22118 23420
rect 22054 23360 22118 23364
rect 22134 23420 22198 23424
rect 22134 23364 22138 23420
rect 22138 23364 22194 23420
rect 22194 23364 22198 23420
rect 22134 23360 22198 23364
rect 22214 23420 22278 23424
rect 22214 23364 22218 23420
rect 22218 23364 22274 23420
rect 22274 23364 22278 23420
rect 22214 23360 22278 23364
rect 22294 23420 22358 23424
rect 22294 23364 22298 23420
rect 22298 23364 22354 23420
rect 22354 23364 22358 23420
rect 22294 23360 22358 23364
rect 30495 23420 30559 23424
rect 30495 23364 30499 23420
rect 30499 23364 30555 23420
rect 30555 23364 30559 23420
rect 30495 23360 30559 23364
rect 30575 23420 30639 23424
rect 30575 23364 30579 23420
rect 30579 23364 30635 23420
rect 30635 23364 30639 23420
rect 30575 23360 30639 23364
rect 30655 23420 30719 23424
rect 30655 23364 30659 23420
rect 30659 23364 30715 23420
rect 30715 23364 30719 23420
rect 30655 23360 30719 23364
rect 30735 23420 30799 23424
rect 30735 23364 30739 23420
rect 30739 23364 30795 23420
rect 30795 23364 30799 23420
rect 30735 23360 30799 23364
rect 9392 22876 9456 22880
rect 9392 22820 9396 22876
rect 9396 22820 9452 22876
rect 9452 22820 9456 22876
rect 9392 22816 9456 22820
rect 9472 22876 9536 22880
rect 9472 22820 9476 22876
rect 9476 22820 9532 22876
rect 9532 22820 9536 22876
rect 9472 22816 9536 22820
rect 9552 22876 9616 22880
rect 9552 22820 9556 22876
rect 9556 22820 9612 22876
rect 9612 22820 9616 22876
rect 9552 22816 9616 22820
rect 9632 22876 9696 22880
rect 9632 22820 9636 22876
rect 9636 22820 9692 22876
rect 9692 22820 9696 22876
rect 9632 22816 9696 22820
rect 17833 22876 17897 22880
rect 17833 22820 17837 22876
rect 17837 22820 17893 22876
rect 17893 22820 17897 22876
rect 17833 22816 17897 22820
rect 17913 22876 17977 22880
rect 17913 22820 17917 22876
rect 17917 22820 17973 22876
rect 17973 22820 17977 22876
rect 17913 22816 17977 22820
rect 17993 22876 18057 22880
rect 17993 22820 17997 22876
rect 17997 22820 18053 22876
rect 18053 22820 18057 22876
rect 17993 22816 18057 22820
rect 18073 22876 18137 22880
rect 18073 22820 18077 22876
rect 18077 22820 18133 22876
rect 18133 22820 18137 22876
rect 18073 22816 18137 22820
rect 26274 22876 26338 22880
rect 26274 22820 26278 22876
rect 26278 22820 26334 22876
rect 26334 22820 26338 22876
rect 26274 22816 26338 22820
rect 26354 22876 26418 22880
rect 26354 22820 26358 22876
rect 26358 22820 26414 22876
rect 26414 22820 26418 22876
rect 26354 22816 26418 22820
rect 26434 22876 26498 22880
rect 26434 22820 26438 22876
rect 26438 22820 26494 22876
rect 26494 22820 26498 22876
rect 26434 22816 26498 22820
rect 26514 22876 26578 22880
rect 26514 22820 26518 22876
rect 26518 22820 26574 22876
rect 26574 22820 26578 22876
rect 26514 22816 26578 22820
rect 34715 22876 34779 22880
rect 34715 22820 34719 22876
rect 34719 22820 34775 22876
rect 34775 22820 34779 22876
rect 34715 22816 34779 22820
rect 34795 22876 34859 22880
rect 34795 22820 34799 22876
rect 34799 22820 34855 22876
rect 34855 22820 34859 22876
rect 34795 22816 34859 22820
rect 34875 22876 34939 22880
rect 34875 22820 34879 22876
rect 34879 22820 34935 22876
rect 34935 22820 34939 22876
rect 34875 22816 34939 22820
rect 34955 22876 35019 22880
rect 34955 22820 34959 22876
rect 34959 22820 35015 22876
rect 35015 22820 35019 22876
rect 34955 22816 35019 22820
rect 34100 22612 34164 22676
rect 5172 22332 5236 22336
rect 5172 22276 5176 22332
rect 5176 22276 5232 22332
rect 5232 22276 5236 22332
rect 5172 22272 5236 22276
rect 5252 22332 5316 22336
rect 5252 22276 5256 22332
rect 5256 22276 5312 22332
rect 5312 22276 5316 22332
rect 5252 22272 5316 22276
rect 5332 22332 5396 22336
rect 5332 22276 5336 22332
rect 5336 22276 5392 22332
rect 5392 22276 5396 22332
rect 5332 22272 5396 22276
rect 5412 22332 5476 22336
rect 5412 22276 5416 22332
rect 5416 22276 5472 22332
rect 5472 22276 5476 22332
rect 5412 22272 5476 22276
rect 13613 22332 13677 22336
rect 13613 22276 13617 22332
rect 13617 22276 13673 22332
rect 13673 22276 13677 22332
rect 13613 22272 13677 22276
rect 13693 22332 13757 22336
rect 13693 22276 13697 22332
rect 13697 22276 13753 22332
rect 13753 22276 13757 22332
rect 13693 22272 13757 22276
rect 13773 22332 13837 22336
rect 13773 22276 13777 22332
rect 13777 22276 13833 22332
rect 13833 22276 13837 22332
rect 13773 22272 13837 22276
rect 13853 22332 13917 22336
rect 13853 22276 13857 22332
rect 13857 22276 13913 22332
rect 13913 22276 13917 22332
rect 13853 22272 13917 22276
rect 22054 22332 22118 22336
rect 22054 22276 22058 22332
rect 22058 22276 22114 22332
rect 22114 22276 22118 22332
rect 22054 22272 22118 22276
rect 22134 22332 22198 22336
rect 22134 22276 22138 22332
rect 22138 22276 22194 22332
rect 22194 22276 22198 22332
rect 22134 22272 22198 22276
rect 22214 22332 22278 22336
rect 22214 22276 22218 22332
rect 22218 22276 22274 22332
rect 22274 22276 22278 22332
rect 22214 22272 22278 22276
rect 22294 22332 22358 22336
rect 22294 22276 22298 22332
rect 22298 22276 22354 22332
rect 22354 22276 22358 22332
rect 22294 22272 22358 22276
rect 30495 22332 30559 22336
rect 30495 22276 30499 22332
rect 30499 22276 30555 22332
rect 30555 22276 30559 22332
rect 30495 22272 30559 22276
rect 30575 22332 30639 22336
rect 30575 22276 30579 22332
rect 30579 22276 30635 22332
rect 30635 22276 30639 22332
rect 30575 22272 30639 22276
rect 30655 22332 30719 22336
rect 30655 22276 30659 22332
rect 30659 22276 30715 22332
rect 30715 22276 30719 22332
rect 30655 22272 30719 22276
rect 30735 22332 30799 22336
rect 30735 22276 30739 22332
rect 30739 22276 30795 22332
rect 30795 22276 30799 22332
rect 30735 22272 30799 22276
rect 29684 22204 29748 22268
rect 29132 21796 29196 21860
rect 9392 21788 9456 21792
rect 9392 21732 9396 21788
rect 9396 21732 9452 21788
rect 9452 21732 9456 21788
rect 9392 21728 9456 21732
rect 9472 21788 9536 21792
rect 9472 21732 9476 21788
rect 9476 21732 9532 21788
rect 9532 21732 9536 21788
rect 9472 21728 9536 21732
rect 9552 21788 9616 21792
rect 9552 21732 9556 21788
rect 9556 21732 9612 21788
rect 9612 21732 9616 21788
rect 9552 21728 9616 21732
rect 9632 21788 9696 21792
rect 9632 21732 9636 21788
rect 9636 21732 9692 21788
rect 9692 21732 9696 21788
rect 9632 21728 9696 21732
rect 17833 21788 17897 21792
rect 17833 21732 17837 21788
rect 17837 21732 17893 21788
rect 17893 21732 17897 21788
rect 17833 21728 17897 21732
rect 17913 21788 17977 21792
rect 17913 21732 17917 21788
rect 17917 21732 17973 21788
rect 17973 21732 17977 21788
rect 17913 21728 17977 21732
rect 17993 21788 18057 21792
rect 17993 21732 17997 21788
rect 17997 21732 18053 21788
rect 18053 21732 18057 21788
rect 17993 21728 18057 21732
rect 18073 21788 18137 21792
rect 18073 21732 18077 21788
rect 18077 21732 18133 21788
rect 18133 21732 18137 21788
rect 18073 21728 18137 21732
rect 26274 21788 26338 21792
rect 26274 21732 26278 21788
rect 26278 21732 26334 21788
rect 26334 21732 26338 21788
rect 26274 21728 26338 21732
rect 26354 21788 26418 21792
rect 26354 21732 26358 21788
rect 26358 21732 26414 21788
rect 26414 21732 26418 21788
rect 26354 21728 26418 21732
rect 26434 21788 26498 21792
rect 26434 21732 26438 21788
rect 26438 21732 26494 21788
rect 26494 21732 26498 21788
rect 26434 21728 26498 21732
rect 26514 21788 26578 21792
rect 26514 21732 26518 21788
rect 26518 21732 26574 21788
rect 26574 21732 26578 21788
rect 26514 21728 26578 21732
rect 34715 21788 34779 21792
rect 34715 21732 34719 21788
rect 34719 21732 34775 21788
rect 34775 21732 34779 21788
rect 34715 21728 34779 21732
rect 34795 21788 34859 21792
rect 34795 21732 34799 21788
rect 34799 21732 34855 21788
rect 34855 21732 34859 21788
rect 34795 21728 34859 21732
rect 34875 21788 34939 21792
rect 34875 21732 34879 21788
rect 34879 21732 34935 21788
rect 34935 21732 34939 21788
rect 34875 21728 34939 21732
rect 34955 21788 35019 21792
rect 34955 21732 34959 21788
rect 34959 21732 35015 21788
rect 35015 21732 35019 21788
rect 34955 21728 35019 21732
rect 5172 21244 5236 21248
rect 5172 21188 5176 21244
rect 5176 21188 5232 21244
rect 5232 21188 5236 21244
rect 5172 21184 5236 21188
rect 5252 21244 5316 21248
rect 5252 21188 5256 21244
rect 5256 21188 5312 21244
rect 5312 21188 5316 21244
rect 5252 21184 5316 21188
rect 5332 21244 5396 21248
rect 5332 21188 5336 21244
rect 5336 21188 5392 21244
rect 5392 21188 5396 21244
rect 5332 21184 5396 21188
rect 5412 21244 5476 21248
rect 5412 21188 5416 21244
rect 5416 21188 5472 21244
rect 5472 21188 5476 21244
rect 5412 21184 5476 21188
rect 13613 21244 13677 21248
rect 13613 21188 13617 21244
rect 13617 21188 13673 21244
rect 13673 21188 13677 21244
rect 13613 21184 13677 21188
rect 13693 21244 13757 21248
rect 13693 21188 13697 21244
rect 13697 21188 13753 21244
rect 13753 21188 13757 21244
rect 13693 21184 13757 21188
rect 13773 21244 13837 21248
rect 13773 21188 13777 21244
rect 13777 21188 13833 21244
rect 13833 21188 13837 21244
rect 13773 21184 13837 21188
rect 13853 21244 13917 21248
rect 13853 21188 13857 21244
rect 13857 21188 13913 21244
rect 13913 21188 13917 21244
rect 13853 21184 13917 21188
rect 22054 21244 22118 21248
rect 22054 21188 22058 21244
rect 22058 21188 22114 21244
rect 22114 21188 22118 21244
rect 22054 21184 22118 21188
rect 22134 21244 22198 21248
rect 22134 21188 22138 21244
rect 22138 21188 22194 21244
rect 22194 21188 22198 21244
rect 22134 21184 22198 21188
rect 22214 21244 22278 21248
rect 22214 21188 22218 21244
rect 22218 21188 22274 21244
rect 22274 21188 22278 21244
rect 22214 21184 22278 21188
rect 22294 21244 22358 21248
rect 22294 21188 22298 21244
rect 22298 21188 22354 21244
rect 22354 21188 22358 21244
rect 22294 21184 22358 21188
rect 30495 21244 30559 21248
rect 30495 21188 30499 21244
rect 30499 21188 30555 21244
rect 30555 21188 30559 21244
rect 30495 21184 30559 21188
rect 30575 21244 30639 21248
rect 30575 21188 30579 21244
rect 30579 21188 30635 21244
rect 30635 21188 30639 21244
rect 30575 21184 30639 21188
rect 30655 21244 30719 21248
rect 30655 21188 30659 21244
rect 30659 21188 30715 21244
rect 30715 21188 30719 21244
rect 30655 21184 30719 21188
rect 30735 21244 30799 21248
rect 30735 21188 30739 21244
rect 30739 21188 30795 21244
rect 30795 21188 30799 21244
rect 30735 21184 30799 21188
rect 32260 20844 32324 20908
rect 25636 20768 25700 20772
rect 25636 20712 25686 20768
rect 25686 20712 25700 20768
rect 25636 20708 25700 20712
rect 30972 20708 31036 20772
rect 31156 20708 31220 20772
rect 9392 20700 9456 20704
rect 9392 20644 9396 20700
rect 9396 20644 9452 20700
rect 9452 20644 9456 20700
rect 9392 20640 9456 20644
rect 9472 20700 9536 20704
rect 9472 20644 9476 20700
rect 9476 20644 9532 20700
rect 9532 20644 9536 20700
rect 9472 20640 9536 20644
rect 9552 20700 9616 20704
rect 9552 20644 9556 20700
rect 9556 20644 9612 20700
rect 9612 20644 9616 20700
rect 9552 20640 9616 20644
rect 9632 20700 9696 20704
rect 9632 20644 9636 20700
rect 9636 20644 9692 20700
rect 9692 20644 9696 20700
rect 9632 20640 9696 20644
rect 17833 20700 17897 20704
rect 17833 20644 17837 20700
rect 17837 20644 17893 20700
rect 17893 20644 17897 20700
rect 17833 20640 17897 20644
rect 17913 20700 17977 20704
rect 17913 20644 17917 20700
rect 17917 20644 17973 20700
rect 17973 20644 17977 20700
rect 17913 20640 17977 20644
rect 17993 20700 18057 20704
rect 17993 20644 17997 20700
rect 17997 20644 18053 20700
rect 18053 20644 18057 20700
rect 17993 20640 18057 20644
rect 18073 20700 18137 20704
rect 18073 20644 18077 20700
rect 18077 20644 18133 20700
rect 18133 20644 18137 20700
rect 18073 20640 18137 20644
rect 26274 20700 26338 20704
rect 26274 20644 26278 20700
rect 26278 20644 26334 20700
rect 26334 20644 26338 20700
rect 26274 20640 26338 20644
rect 26354 20700 26418 20704
rect 26354 20644 26358 20700
rect 26358 20644 26414 20700
rect 26414 20644 26418 20700
rect 26354 20640 26418 20644
rect 26434 20700 26498 20704
rect 26434 20644 26438 20700
rect 26438 20644 26494 20700
rect 26494 20644 26498 20700
rect 26434 20640 26498 20644
rect 26514 20700 26578 20704
rect 26514 20644 26518 20700
rect 26518 20644 26574 20700
rect 26574 20644 26578 20700
rect 26514 20640 26578 20644
rect 34715 20700 34779 20704
rect 34715 20644 34719 20700
rect 34719 20644 34775 20700
rect 34775 20644 34779 20700
rect 34715 20640 34779 20644
rect 34795 20700 34859 20704
rect 34795 20644 34799 20700
rect 34799 20644 34855 20700
rect 34855 20644 34859 20700
rect 34795 20640 34859 20644
rect 34875 20700 34939 20704
rect 34875 20644 34879 20700
rect 34879 20644 34935 20700
rect 34935 20644 34939 20700
rect 34875 20640 34939 20644
rect 34955 20700 35019 20704
rect 34955 20644 34959 20700
rect 34959 20644 35015 20700
rect 35015 20644 35019 20700
rect 34955 20640 35019 20644
rect 5172 20156 5236 20160
rect 5172 20100 5176 20156
rect 5176 20100 5232 20156
rect 5232 20100 5236 20156
rect 5172 20096 5236 20100
rect 5252 20156 5316 20160
rect 5252 20100 5256 20156
rect 5256 20100 5312 20156
rect 5312 20100 5316 20156
rect 5252 20096 5316 20100
rect 5332 20156 5396 20160
rect 5332 20100 5336 20156
rect 5336 20100 5392 20156
rect 5392 20100 5396 20156
rect 5332 20096 5396 20100
rect 5412 20156 5476 20160
rect 5412 20100 5416 20156
rect 5416 20100 5472 20156
rect 5472 20100 5476 20156
rect 5412 20096 5476 20100
rect 13613 20156 13677 20160
rect 13613 20100 13617 20156
rect 13617 20100 13673 20156
rect 13673 20100 13677 20156
rect 13613 20096 13677 20100
rect 13693 20156 13757 20160
rect 13693 20100 13697 20156
rect 13697 20100 13753 20156
rect 13753 20100 13757 20156
rect 13693 20096 13757 20100
rect 13773 20156 13837 20160
rect 13773 20100 13777 20156
rect 13777 20100 13833 20156
rect 13833 20100 13837 20156
rect 13773 20096 13837 20100
rect 13853 20156 13917 20160
rect 13853 20100 13857 20156
rect 13857 20100 13913 20156
rect 13913 20100 13917 20156
rect 13853 20096 13917 20100
rect 22054 20156 22118 20160
rect 22054 20100 22058 20156
rect 22058 20100 22114 20156
rect 22114 20100 22118 20156
rect 22054 20096 22118 20100
rect 22134 20156 22198 20160
rect 22134 20100 22138 20156
rect 22138 20100 22194 20156
rect 22194 20100 22198 20156
rect 22134 20096 22198 20100
rect 22214 20156 22278 20160
rect 22214 20100 22218 20156
rect 22218 20100 22274 20156
rect 22274 20100 22278 20156
rect 22214 20096 22278 20100
rect 22294 20156 22358 20160
rect 22294 20100 22298 20156
rect 22298 20100 22354 20156
rect 22354 20100 22358 20156
rect 22294 20096 22358 20100
rect 30495 20156 30559 20160
rect 30495 20100 30499 20156
rect 30499 20100 30555 20156
rect 30555 20100 30559 20156
rect 30495 20096 30559 20100
rect 30575 20156 30639 20160
rect 30575 20100 30579 20156
rect 30579 20100 30635 20156
rect 30635 20100 30639 20156
rect 30575 20096 30639 20100
rect 30655 20156 30719 20160
rect 30655 20100 30659 20156
rect 30659 20100 30715 20156
rect 30715 20100 30719 20156
rect 30655 20096 30719 20100
rect 30735 20156 30799 20160
rect 30735 20100 30739 20156
rect 30739 20100 30795 20156
rect 30795 20100 30799 20156
rect 30735 20096 30799 20100
rect 9392 19612 9456 19616
rect 9392 19556 9396 19612
rect 9396 19556 9452 19612
rect 9452 19556 9456 19612
rect 9392 19552 9456 19556
rect 9472 19612 9536 19616
rect 9472 19556 9476 19612
rect 9476 19556 9532 19612
rect 9532 19556 9536 19612
rect 9472 19552 9536 19556
rect 9552 19612 9616 19616
rect 9552 19556 9556 19612
rect 9556 19556 9612 19612
rect 9612 19556 9616 19612
rect 9552 19552 9616 19556
rect 9632 19612 9696 19616
rect 9632 19556 9636 19612
rect 9636 19556 9692 19612
rect 9692 19556 9696 19612
rect 9632 19552 9696 19556
rect 17833 19612 17897 19616
rect 17833 19556 17837 19612
rect 17837 19556 17893 19612
rect 17893 19556 17897 19612
rect 17833 19552 17897 19556
rect 17913 19612 17977 19616
rect 17913 19556 17917 19612
rect 17917 19556 17973 19612
rect 17973 19556 17977 19612
rect 17913 19552 17977 19556
rect 17993 19612 18057 19616
rect 17993 19556 17997 19612
rect 17997 19556 18053 19612
rect 18053 19556 18057 19612
rect 17993 19552 18057 19556
rect 18073 19612 18137 19616
rect 18073 19556 18077 19612
rect 18077 19556 18133 19612
rect 18133 19556 18137 19612
rect 18073 19552 18137 19556
rect 26274 19612 26338 19616
rect 26274 19556 26278 19612
rect 26278 19556 26334 19612
rect 26334 19556 26338 19612
rect 26274 19552 26338 19556
rect 26354 19612 26418 19616
rect 26354 19556 26358 19612
rect 26358 19556 26414 19612
rect 26414 19556 26418 19612
rect 26354 19552 26418 19556
rect 26434 19612 26498 19616
rect 26434 19556 26438 19612
rect 26438 19556 26494 19612
rect 26494 19556 26498 19612
rect 26434 19552 26498 19556
rect 26514 19612 26578 19616
rect 26514 19556 26518 19612
rect 26518 19556 26574 19612
rect 26574 19556 26578 19612
rect 26514 19552 26578 19556
rect 34715 19612 34779 19616
rect 34715 19556 34719 19612
rect 34719 19556 34775 19612
rect 34775 19556 34779 19612
rect 34715 19552 34779 19556
rect 34795 19612 34859 19616
rect 34795 19556 34799 19612
rect 34799 19556 34855 19612
rect 34855 19556 34859 19612
rect 34795 19552 34859 19556
rect 34875 19612 34939 19616
rect 34875 19556 34879 19612
rect 34879 19556 34935 19612
rect 34935 19556 34939 19612
rect 34875 19552 34939 19556
rect 34955 19612 35019 19616
rect 34955 19556 34959 19612
rect 34959 19556 35015 19612
rect 35015 19556 35019 19612
rect 34955 19552 35019 19556
rect 5172 19068 5236 19072
rect 5172 19012 5176 19068
rect 5176 19012 5232 19068
rect 5232 19012 5236 19068
rect 5172 19008 5236 19012
rect 5252 19068 5316 19072
rect 5252 19012 5256 19068
rect 5256 19012 5312 19068
rect 5312 19012 5316 19068
rect 5252 19008 5316 19012
rect 5332 19068 5396 19072
rect 5332 19012 5336 19068
rect 5336 19012 5392 19068
rect 5392 19012 5396 19068
rect 5332 19008 5396 19012
rect 5412 19068 5476 19072
rect 5412 19012 5416 19068
rect 5416 19012 5472 19068
rect 5472 19012 5476 19068
rect 5412 19008 5476 19012
rect 13613 19068 13677 19072
rect 13613 19012 13617 19068
rect 13617 19012 13673 19068
rect 13673 19012 13677 19068
rect 13613 19008 13677 19012
rect 13693 19068 13757 19072
rect 13693 19012 13697 19068
rect 13697 19012 13753 19068
rect 13753 19012 13757 19068
rect 13693 19008 13757 19012
rect 13773 19068 13837 19072
rect 13773 19012 13777 19068
rect 13777 19012 13833 19068
rect 13833 19012 13837 19068
rect 13773 19008 13837 19012
rect 13853 19068 13917 19072
rect 13853 19012 13857 19068
rect 13857 19012 13913 19068
rect 13913 19012 13917 19068
rect 13853 19008 13917 19012
rect 22054 19068 22118 19072
rect 22054 19012 22058 19068
rect 22058 19012 22114 19068
rect 22114 19012 22118 19068
rect 22054 19008 22118 19012
rect 22134 19068 22198 19072
rect 22134 19012 22138 19068
rect 22138 19012 22194 19068
rect 22194 19012 22198 19068
rect 22134 19008 22198 19012
rect 22214 19068 22278 19072
rect 22214 19012 22218 19068
rect 22218 19012 22274 19068
rect 22274 19012 22278 19068
rect 22214 19008 22278 19012
rect 22294 19068 22358 19072
rect 22294 19012 22298 19068
rect 22298 19012 22354 19068
rect 22354 19012 22358 19068
rect 22294 19008 22358 19012
rect 30495 19068 30559 19072
rect 30495 19012 30499 19068
rect 30499 19012 30555 19068
rect 30555 19012 30559 19068
rect 30495 19008 30559 19012
rect 30575 19068 30639 19072
rect 30575 19012 30579 19068
rect 30579 19012 30635 19068
rect 30635 19012 30639 19068
rect 30575 19008 30639 19012
rect 30655 19068 30719 19072
rect 30655 19012 30659 19068
rect 30659 19012 30715 19068
rect 30715 19012 30719 19068
rect 30655 19008 30719 19012
rect 30735 19068 30799 19072
rect 30735 19012 30739 19068
rect 30739 19012 30795 19068
rect 30795 19012 30799 19068
rect 30735 19008 30799 19012
rect 32260 18940 32324 19004
rect 27660 18668 27724 18732
rect 24532 18592 24596 18596
rect 24532 18536 24582 18592
rect 24582 18536 24596 18592
rect 24532 18532 24596 18536
rect 9392 18524 9456 18528
rect 9392 18468 9396 18524
rect 9396 18468 9452 18524
rect 9452 18468 9456 18524
rect 9392 18464 9456 18468
rect 9472 18524 9536 18528
rect 9472 18468 9476 18524
rect 9476 18468 9532 18524
rect 9532 18468 9536 18524
rect 9472 18464 9536 18468
rect 9552 18524 9616 18528
rect 9552 18468 9556 18524
rect 9556 18468 9612 18524
rect 9612 18468 9616 18524
rect 9552 18464 9616 18468
rect 9632 18524 9696 18528
rect 9632 18468 9636 18524
rect 9636 18468 9692 18524
rect 9692 18468 9696 18524
rect 9632 18464 9696 18468
rect 17833 18524 17897 18528
rect 17833 18468 17837 18524
rect 17837 18468 17893 18524
rect 17893 18468 17897 18524
rect 17833 18464 17897 18468
rect 17913 18524 17977 18528
rect 17913 18468 17917 18524
rect 17917 18468 17973 18524
rect 17973 18468 17977 18524
rect 17913 18464 17977 18468
rect 17993 18524 18057 18528
rect 17993 18468 17997 18524
rect 17997 18468 18053 18524
rect 18053 18468 18057 18524
rect 17993 18464 18057 18468
rect 18073 18524 18137 18528
rect 18073 18468 18077 18524
rect 18077 18468 18133 18524
rect 18133 18468 18137 18524
rect 18073 18464 18137 18468
rect 26274 18524 26338 18528
rect 26274 18468 26278 18524
rect 26278 18468 26334 18524
rect 26334 18468 26338 18524
rect 26274 18464 26338 18468
rect 26354 18524 26418 18528
rect 26354 18468 26358 18524
rect 26358 18468 26414 18524
rect 26414 18468 26418 18524
rect 26354 18464 26418 18468
rect 26434 18524 26498 18528
rect 26434 18468 26438 18524
rect 26438 18468 26494 18524
rect 26494 18468 26498 18524
rect 26434 18464 26498 18468
rect 26514 18524 26578 18528
rect 26514 18468 26518 18524
rect 26518 18468 26574 18524
rect 26574 18468 26578 18524
rect 26514 18464 26578 18468
rect 34715 18524 34779 18528
rect 34715 18468 34719 18524
rect 34719 18468 34775 18524
rect 34775 18468 34779 18524
rect 34715 18464 34779 18468
rect 34795 18524 34859 18528
rect 34795 18468 34799 18524
rect 34799 18468 34855 18524
rect 34855 18468 34859 18524
rect 34795 18464 34859 18468
rect 34875 18524 34939 18528
rect 34875 18468 34879 18524
rect 34879 18468 34935 18524
rect 34935 18468 34939 18524
rect 34875 18464 34939 18468
rect 34955 18524 35019 18528
rect 34955 18468 34959 18524
rect 34959 18468 35015 18524
rect 35015 18468 35019 18524
rect 34955 18464 35019 18468
rect 32812 17988 32876 18052
rect 5172 17980 5236 17984
rect 5172 17924 5176 17980
rect 5176 17924 5232 17980
rect 5232 17924 5236 17980
rect 5172 17920 5236 17924
rect 5252 17980 5316 17984
rect 5252 17924 5256 17980
rect 5256 17924 5312 17980
rect 5312 17924 5316 17980
rect 5252 17920 5316 17924
rect 5332 17980 5396 17984
rect 5332 17924 5336 17980
rect 5336 17924 5392 17980
rect 5392 17924 5396 17980
rect 5332 17920 5396 17924
rect 5412 17980 5476 17984
rect 5412 17924 5416 17980
rect 5416 17924 5472 17980
rect 5472 17924 5476 17980
rect 5412 17920 5476 17924
rect 13613 17980 13677 17984
rect 13613 17924 13617 17980
rect 13617 17924 13673 17980
rect 13673 17924 13677 17980
rect 13613 17920 13677 17924
rect 13693 17980 13757 17984
rect 13693 17924 13697 17980
rect 13697 17924 13753 17980
rect 13753 17924 13757 17980
rect 13693 17920 13757 17924
rect 13773 17980 13837 17984
rect 13773 17924 13777 17980
rect 13777 17924 13833 17980
rect 13833 17924 13837 17980
rect 13773 17920 13837 17924
rect 13853 17980 13917 17984
rect 13853 17924 13857 17980
rect 13857 17924 13913 17980
rect 13913 17924 13917 17980
rect 13853 17920 13917 17924
rect 22054 17980 22118 17984
rect 22054 17924 22058 17980
rect 22058 17924 22114 17980
rect 22114 17924 22118 17980
rect 22054 17920 22118 17924
rect 22134 17980 22198 17984
rect 22134 17924 22138 17980
rect 22138 17924 22194 17980
rect 22194 17924 22198 17980
rect 22134 17920 22198 17924
rect 22214 17980 22278 17984
rect 22214 17924 22218 17980
rect 22218 17924 22274 17980
rect 22274 17924 22278 17980
rect 22214 17920 22278 17924
rect 22294 17980 22358 17984
rect 22294 17924 22298 17980
rect 22298 17924 22354 17980
rect 22354 17924 22358 17980
rect 22294 17920 22358 17924
rect 30495 17980 30559 17984
rect 30495 17924 30499 17980
rect 30499 17924 30555 17980
rect 30555 17924 30559 17980
rect 30495 17920 30559 17924
rect 30575 17980 30639 17984
rect 30575 17924 30579 17980
rect 30579 17924 30635 17980
rect 30635 17924 30639 17980
rect 30575 17920 30639 17924
rect 30655 17980 30719 17984
rect 30655 17924 30659 17980
rect 30659 17924 30715 17980
rect 30715 17924 30719 17980
rect 30655 17920 30719 17924
rect 30735 17980 30799 17984
rect 30735 17924 30739 17980
rect 30739 17924 30795 17980
rect 30795 17924 30799 17980
rect 30735 17920 30799 17924
rect 9392 17436 9456 17440
rect 9392 17380 9396 17436
rect 9396 17380 9452 17436
rect 9452 17380 9456 17436
rect 9392 17376 9456 17380
rect 9472 17436 9536 17440
rect 9472 17380 9476 17436
rect 9476 17380 9532 17436
rect 9532 17380 9536 17436
rect 9472 17376 9536 17380
rect 9552 17436 9616 17440
rect 9552 17380 9556 17436
rect 9556 17380 9612 17436
rect 9612 17380 9616 17436
rect 9552 17376 9616 17380
rect 9632 17436 9696 17440
rect 9632 17380 9636 17436
rect 9636 17380 9692 17436
rect 9692 17380 9696 17436
rect 9632 17376 9696 17380
rect 17833 17436 17897 17440
rect 17833 17380 17837 17436
rect 17837 17380 17893 17436
rect 17893 17380 17897 17436
rect 17833 17376 17897 17380
rect 17913 17436 17977 17440
rect 17913 17380 17917 17436
rect 17917 17380 17973 17436
rect 17973 17380 17977 17436
rect 17913 17376 17977 17380
rect 17993 17436 18057 17440
rect 17993 17380 17997 17436
rect 17997 17380 18053 17436
rect 18053 17380 18057 17436
rect 17993 17376 18057 17380
rect 18073 17436 18137 17440
rect 18073 17380 18077 17436
rect 18077 17380 18133 17436
rect 18133 17380 18137 17436
rect 18073 17376 18137 17380
rect 26274 17436 26338 17440
rect 26274 17380 26278 17436
rect 26278 17380 26334 17436
rect 26334 17380 26338 17436
rect 26274 17376 26338 17380
rect 26354 17436 26418 17440
rect 26354 17380 26358 17436
rect 26358 17380 26414 17436
rect 26414 17380 26418 17436
rect 26354 17376 26418 17380
rect 26434 17436 26498 17440
rect 26434 17380 26438 17436
rect 26438 17380 26494 17436
rect 26494 17380 26498 17436
rect 26434 17376 26498 17380
rect 26514 17436 26578 17440
rect 26514 17380 26518 17436
rect 26518 17380 26574 17436
rect 26574 17380 26578 17436
rect 26514 17376 26578 17380
rect 34715 17436 34779 17440
rect 34715 17380 34719 17436
rect 34719 17380 34775 17436
rect 34775 17380 34779 17436
rect 34715 17376 34779 17380
rect 34795 17436 34859 17440
rect 34795 17380 34799 17436
rect 34799 17380 34855 17436
rect 34855 17380 34859 17436
rect 34795 17376 34859 17380
rect 34875 17436 34939 17440
rect 34875 17380 34879 17436
rect 34879 17380 34935 17436
rect 34935 17380 34939 17436
rect 34875 17376 34939 17380
rect 34955 17436 35019 17440
rect 34955 17380 34959 17436
rect 34959 17380 35015 17436
rect 35015 17380 35019 17436
rect 34955 17376 35019 17380
rect 5172 16892 5236 16896
rect 5172 16836 5176 16892
rect 5176 16836 5232 16892
rect 5232 16836 5236 16892
rect 5172 16832 5236 16836
rect 5252 16892 5316 16896
rect 5252 16836 5256 16892
rect 5256 16836 5312 16892
rect 5312 16836 5316 16892
rect 5252 16832 5316 16836
rect 5332 16892 5396 16896
rect 5332 16836 5336 16892
rect 5336 16836 5392 16892
rect 5392 16836 5396 16892
rect 5332 16832 5396 16836
rect 5412 16892 5476 16896
rect 5412 16836 5416 16892
rect 5416 16836 5472 16892
rect 5472 16836 5476 16892
rect 5412 16832 5476 16836
rect 13613 16892 13677 16896
rect 13613 16836 13617 16892
rect 13617 16836 13673 16892
rect 13673 16836 13677 16892
rect 13613 16832 13677 16836
rect 13693 16892 13757 16896
rect 13693 16836 13697 16892
rect 13697 16836 13753 16892
rect 13753 16836 13757 16892
rect 13693 16832 13757 16836
rect 13773 16892 13837 16896
rect 13773 16836 13777 16892
rect 13777 16836 13833 16892
rect 13833 16836 13837 16892
rect 13773 16832 13837 16836
rect 13853 16892 13917 16896
rect 13853 16836 13857 16892
rect 13857 16836 13913 16892
rect 13913 16836 13917 16892
rect 13853 16832 13917 16836
rect 22054 16892 22118 16896
rect 22054 16836 22058 16892
rect 22058 16836 22114 16892
rect 22114 16836 22118 16892
rect 22054 16832 22118 16836
rect 22134 16892 22198 16896
rect 22134 16836 22138 16892
rect 22138 16836 22194 16892
rect 22194 16836 22198 16892
rect 22134 16832 22198 16836
rect 22214 16892 22278 16896
rect 22214 16836 22218 16892
rect 22218 16836 22274 16892
rect 22274 16836 22278 16892
rect 22214 16832 22278 16836
rect 22294 16892 22358 16896
rect 22294 16836 22298 16892
rect 22298 16836 22354 16892
rect 22354 16836 22358 16892
rect 22294 16832 22358 16836
rect 30495 16892 30559 16896
rect 30495 16836 30499 16892
rect 30499 16836 30555 16892
rect 30555 16836 30559 16892
rect 30495 16832 30559 16836
rect 30575 16892 30639 16896
rect 30575 16836 30579 16892
rect 30579 16836 30635 16892
rect 30635 16836 30639 16892
rect 30575 16832 30639 16836
rect 30655 16892 30719 16896
rect 30655 16836 30659 16892
rect 30659 16836 30715 16892
rect 30715 16836 30719 16892
rect 30655 16832 30719 16836
rect 30735 16892 30799 16896
rect 30735 16836 30739 16892
rect 30739 16836 30795 16892
rect 30795 16836 30799 16892
rect 30735 16832 30799 16836
rect 31156 16764 31220 16828
rect 31340 16764 31404 16828
rect 32076 16628 32140 16692
rect 24532 16492 24596 16556
rect 29684 16492 29748 16556
rect 9392 16348 9456 16352
rect 9392 16292 9396 16348
rect 9396 16292 9452 16348
rect 9452 16292 9456 16348
rect 9392 16288 9456 16292
rect 9472 16348 9536 16352
rect 9472 16292 9476 16348
rect 9476 16292 9532 16348
rect 9532 16292 9536 16348
rect 9472 16288 9536 16292
rect 9552 16348 9616 16352
rect 9552 16292 9556 16348
rect 9556 16292 9612 16348
rect 9612 16292 9616 16348
rect 9552 16288 9616 16292
rect 9632 16348 9696 16352
rect 9632 16292 9636 16348
rect 9636 16292 9692 16348
rect 9692 16292 9696 16348
rect 9632 16288 9696 16292
rect 17833 16348 17897 16352
rect 17833 16292 17837 16348
rect 17837 16292 17893 16348
rect 17893 16292 17897 16348
rect 17833 16288 17897 16292
rect 17913 16348 17977 16352
rect 17913 16292 17917 16348
rect 17917 16292 17973 16348
rect 17973 16292 17977 16348
rect 17913 16288 17977 16292
rect 17993 16348 18057 16352
rect 17993 16292 17997 16348
rect 17997 16292 18053 16348
rect 18053 16292 18057 16348
rect 17993 16288 18057 16292
rect 18073 16348 18137 16352
rect 18073 16292 18077 16348
rect 18077 16292 18133 16348
rect 18133 16292 18137 16348
rect 18073 16288 18137 16292
rect 26274 16348 26338 16352
rect 26274 16292 26278 16348
rect 26278 16292 26334 16348
rect 26334 16292 26338 16348
rect 26274 16288 26338 16292
rect 26354 16348 26418 16352
rect 26354 16292 26358 16348
rect 26358 16292 26414 16348
rect 26414 16292 26418 16348
rect 26354 16288 26418 16292
rect 26434 16348 26498 16352
rect 26434 16292 26438 16348
rect 26438 16292 26494 16348
rect 26494 16292 26498 16348
rect 26434 16288 26498 16292
rect 26514 16348 26578 16352
rect 26514 16292 26518 16348
rect 26518 16292 26574 16348
rect 26574 16292 26578 16348
rect 26514 16288 26578 16292
rect 34715 16348 34779 16352
rect 34715 16292 34719 16348
rect 34719 16292 34775 16348
rect 34775 16292 34779 16348
rect 34715 16288 34779 16292
rect 34795 16348 34859 16352
rect 34795 16292 34799 16348
rect 34799 16292 34855 16348
rect 34855 16292 34859 16348
rect 34795 16288 34859 16292
rect 34875 16348 34939 16352
rect 34875 16292 34879 16348
rect 34879 16292 34935 16348
rect 34935 16292 34939 16348
rect 34875 16288 34939 16292
rect 34955 16348 35019 16352
rect 34955 16292 34959 16348
rect 34959 16292 35015 16348
rect 35015 16292 35019 16348
rect 34955 16288 35019 16292
rect 30972 16220 31036 16284
rect 31524 16220 31588 16284
rect 5172 15804 5236 15808
rect 5172 15748 5176 15804
rect 5176 15748 5232 15804
rect 5232 15748 5236 15804
rect 5172 15744 5236 15748
rect 5252 15804 5316 15808
rect 5252 15748 5256 15804
rect 5256 15748 5312 15804
rect 5312 15748 5316 15804
rect 5252 15744 5316 15748
rect 5332 15804 5396 15808
rect 5332 15748 5336 15804
rect 5336 15748 5392 15804
rect 5392 15748 5396 15804
rect 5332 15744 5396 15748
rect 5412 15804 5476 15808
rect 5412 15748 5416 15804
rect 5416 15748 5472 15804
rect 5472 15748 5476 15804
rect 5412 15744 5476 15748
rect 13613 15804 13677 15808
rect 13613 15748 13617 15804
rect 13617 15748 13673 15804
rect 13673 15748 13677 15804
rect 13613 15744 13677 15748
rect 13693 15804 13757 15808
rect 13693 15748 13697 15804
rect 13697 15748 13753 15804
rect 13753 15748 13757 15804
rect 13693 15744 13757 15748
rect 13773 15804 13837 15808
rect 13773 15748 13777 15804
rect 13777 15748 13833 15804
rect 13833 15748 13837 15804
rect 13773 15744 13837 15748
rect 13853 15804 13917 15808
rect 13853 15748 13857 15804
rect 13857 15748 13913 15804
rect 13913 15748 13917 15804
rect 13853 15744 13917 15748
rect 22054 15804 22118 15808
rect 22054 15748 22058 15804
rect 22058 15748 22114 15804
rect 22114 15748 22118 15804
rect 22054 15744 22118 15748
rect 22134 15804 22198 15808
rect 22134 15748 22138 15804
rect 22138 15748 22194 15804
rect 22194 15748 22198 15804
rect 22134 15744 22198 15748
rect 22214 15804 22278 15808
rect 22214 15748 22218 15804
rect 22218 15748 22274 15804
rect 22274 15748 22278 15804
rect 22214 15744 22278 15748
rect 22294 15804 22358 15808
rect 22294 15748 22298 15804
rect 22298 15748 22354 15804
rect 22354 15748 22358 15804
rect 22294 15744 22358 15748
rect 30495 15804 30559 15808
rect 30495 15748 30499 15804
rect 30499 15748 30555 15804
rect 30555 15748 30559 15804
rect 30495 15744 30559 15748
rect 30575 15804 30639 15808
rect 30575 15748 30579 15804
rect 30579 15748 30635 15804
rect 30635 15748 30639 15804
rect 30575 15744 30639 15748
rect 30655 15804 30719 15808
rect 30655 15748 30659 15804
rect 30659 15748 30715 15804
rect 30715 15748 30719 15804
rect 30655 15744 30719 15748
rect 30735 15804 30799 15808
rect 30735 15748 30739 15804
rect 30739 15748 30795 15804
rect 30795 15748 30799 15804
rect 30735 15744 30799 15748
rect 25636 15328 25700 15332
rect 25636 15272 25650 15328
rect 25650 15272 25700 15328
rect 25636 15268 25700 15272
rect 9392 15260 9456 15264
rect 9392 15204 9396 15260
rect 9396 15204 9452 15260
rect 9452 15204 9456 15260
rect 9392 15200 9456 15204
rect 9472 15260 9536 15264
rect 9472 15204 9476 15260
rect 9476 15204 9532 15260
rect 9532 15204 9536 15260
rect 9472 15200 9536 15204
rect 9552 15260 9616 15264
rect 9552 15204 9556 15260
rect 9556 15204 9612 15260
rect 9612 15204 9616 15260
rect 9552 15200 9616 15204
rect 9632 15260 9696 15264
rect 9632 15204 9636 15260
rect 9636 15204 9692 15260
rect 9692 15204 9696 15260
rect 9632 15200 9696 15204
rect 17833 15260 17897 15264
rect 17833 15204 17837 15260
rect 17837 15204 17893 15260
rect 17893 15204 17897 15260
rect 17833 15200 17897 15204
rect 17913 15260 17977 15264
rect 17913 15204 17917 15260
rect 17917 15204 17973 15260
rect 17973 15204 17977 15260
rect 17913 15200 17977 15204
rect 17993 15260 18057 15264
rect 17993 15204 17997 15260
rect 17997 15204 18053 15260
rect 18053 15204 18057 15260
rect 17993 15200 18057 15204
rect 18073 15260 18137 15264
rect 18073 15204 18077 15260
rect 18077 15204 18133 15260
rect 18133 15204 18137 15260
rect 18073 15200 18137 15204
rect 26274 15260 26338 15264
rect 26274 15204 26278 15260
rect 26278 15204 26334 15260
rect 26334 15204 26338 15260
rect 26274 15200 26338 15204
rect 26354 15260 26418 15264
rect 26354 15204 26358 15260
rect 26358 15204 26414 15260
rect 26414 15204 26418 15260
rect 26354 15200 26418 15204
rect 26434 15260 26498 15264
rect 26434 15204 26438 15260
rect 26438 15204 26494 15260
rect 26494 15204 26498 15260
rect 26434 15200 26498 15204
rect 26514 15260 26578 15264
rect 26514 15204 26518 15260
rect 26518 15204 26574 15260
rect 26574 15204 26578 15260
rect 26514 15200 26578 15204
rect 34715 15260 34779 15264
rect 34715 15204 34719 15260
rect 34719 15204 34775 15260
rect 34775 15204 34779 15260
rect 34715 15200 34779 15204
rect 34795 15260 34859 15264
rect 34795 15204 34799 15260
rect 34799 15204 34855 15260
rect 34855 15204 34859 15260
rect 34795 15200 34859 15204
rect 34875 15260 34939 15264
rect 34875 15204 34879 15260
rect 34879 15204 34935 15260
rect 34935 15204 34939 15260
rect 34875 15200 34939 15204
rect 34955 15260 35019 15264
rect 34955 15204 34959 15260
rect 34959 15204 35015 15260
rect 35015 15204 35019 15260
rect 34955 15200 35019 15204
rect 29500 15132 29564 15196
rect 24716 14996 24780 15060
rect 27660 14996 27724 15060
rect 33916 14996 33980 15060
rect 5172 14716 5236 14720
rect 5172 14660 5176 14716
rect 5176 14660 5232 14716
rect 5232 14660 5236 14716
rect 5172 14656 5236 14660
rect 5252 14716 5316 14720
rect 5252 14660 5256 14716
rect 5256 14660 5312 14716
rect 5312 14660 5316 14716
rect 5252 14656 5316 14660
rect 5332 14716 5396 14720
rect 5332 14660 5336 14716
rect 5336 14660 5392 14716
rect 5392 14660 5396 14716
rect 5332 14656 5396 14660
rect 5412 14716 5476 14720
rect 5412 14660 5416 14716
rect 5416 14660 5472 14716
rect 5472 14660 5476 14716
rect 5412 14656 5476 14660
rect 13613 14716 13677 14720
rect 13613 14660 13617 14716
rect 13617 14660 13673 14716
rect 13673 14660 13677 14716
rect 13613 14656 13677 14660
rect 13693 14716 13757 14720
rect 13693 14660 13697 14716
rect 13697 14660 13753 14716
rect 13753 14660 13757 14716
rect 13693 14656 13757 14660
rect 13773 14716 13837 14720
rect 13773 14660 13777 14716
rect 13777 14660 13833 14716
rect 13833 14660 13837 14716
rect 13773 14656 13837 14660
rect 13853 14716 13917 14720
rect 13853 14660 13857 14716
rect 13857 14660 13913 14716
rect 13913 14660 13917 14716
rect 13853 14656 13917 14660
rect 22054 14716 22118 14720
rect 22054 14660 22058 14716
rect 22058 14660 22114 14716
rect 22114 14660 22118 14716
rect 22054 14656 22118 14660
rect 22134 14716 22198 14720
rect 22134 14660 22138 14716
rect 22138 14660 22194 14716
rect 22194 14660 22198 14716
rect 22134 14656 22198 14660
rect 22214 14716 22278 14720
rect 22214 14660 22218 14716
rect 22218 14660 22274 14716
rect 22274 14660 22278 14716
rect 22214 14656 22278 14660
rect 22294 14716 22358 14720
rect 22294 14660 22298 14716
rect 22298 14660 22354 14716
rect 22354 14660 22358 14716
rect 22294 14656 22358 14660
rect 30495 14716 30559 14720
rect 30495 14660 30499 14716
rect 30499 14660 30555 14716
rect 30555 14660 30559 14716
rect 30495 14656 30559 14660
rect 30575 14716 30639 14720
rect 30575 14660 30579 14716
rect 30579 14660 30635 14716
rect 30635 14660 30639 14716
rect 30575 14656 30639 14660
rect 30655 14716 30719 14720
rect 30655 14660 30659 14716
rect 30659 14660 30715 14716
rect 30715 14660 30719 14716
rect 30655 14656 30719 14660
rect 30735 14716 30799 14720
rect 30735 14660 30739 14716
rect 30739 14660 30795 14716
rect 30795 14660 30799 14716
rect 30735 14656 30799 14660
rect 9392 14172 9456 14176
rect 9392 14116 9396 14172
rect 9396 14116 9452 14172
rect 9452 14116 9456 14172
rect 9392 14112 9456 14116
rect 9472 14172 9536 14176
rect 9472 14116 9476 14172
rect 9476 14116 9532 14172
rect 9532 14116 9536 14172
rect 9472 14112 9536 14116
rect 9552 14172 9616 14176
rect 9552 14116 9556 14172
rect 9556 14116 9612 14172
rect 9612 14116 9616 14172
rect 9552 14112 9616 14116
rect 9632 14172 9696 14176
rect 9632 14116 9636 14172
rect 9636 14116 9692 14172
rect 9692 14116 9696 14172
rect 9632 14112 9696 14116
rect 17833 14172 17897 14176
rect 17833 14116 17837 14172
rect 17837 14116 17893 14172
rect 17893 14116 17897 14172
rect 17833 14112 17897 14116
rect 17913 14172 17977 14176
rect 17913 14116 17917 14172
rect 17917 14116 17973 14172
rect 17973 14116 17977 14172
rect 17913 14112 17977 14116
rect 17993 14172 18057 14176
rect 17993 14116 17997 14172
rect 17997 14116 18053 14172
rect 18053 14116 18057 14172
rect 17993 14112 18057 14116
rect 18073 14172 18137 14176
rect 18073 14116 18077 14172
rect 18077 14116 18133 14172
rect 18133 14116 18137 14172
rect 18073 14112 18137 14116
rect 26274 14172 26338 14176
rect 26274 14116 26278 14172
rect 26278 14116 26334 14172
rect 26334 14116 26338 14172
rect 26274 14112 26338 14116
rect 26354 14172 26418 14176
rect 26354 14116 26358 14172
rect 26358 14116 26414 14172
rect 26414 14116 26418 14172
rect 26354 14112 26418 14116
rect 26434 14172 26498 14176
rect 26434 14116 26438 14172
rect 26438 14116 26494 14172
rect 26494 14116 26498 14172
rect 26434 14112 26498 14116
rect 26514 14172 26578 14176
rect 26514 14116 26518 14172
rect 26518 14116 26574 14172
rect 26574 14116 26578 14172
rect 26514 14112 26578 14116
rect 34715 14172 34779 14176
rect 34715 14116 34719 14172
rect 34719 14116 34775 14172
rect 34775 14116 34779 14172
rect 34715 14112 34779 14116
rect 34795 14172 34859 14176
rect 34795 14116 34799 14172
rect 34799 14116 34855 14172
rect 34855 14116 34859 14172
rect 34795 14112 34859 14116
rect 34875 14172 34939 14176
rect 34875 14116 34879 14172
rect 34879 14116 34935 14172
rect 34935 14116 34939 14172
rect 34875 14112 34939 14116
rect 34955 14172 35019 14176
rect 34955 14116 34959 14172
rect 34959 14116 35015 14172
rect 35015 14116 35019 14172
rect 34955 14112 35019 14116
rect 26740 13908 26804 13972
rect 5172 13628 5236 13632
rect 5172 13572 5176 13628
rect 5176 13572 5232 13628
rect 5232 13572 5236 13628
rect 5172 13568 5236 13572
rect 5252 13628 5316 13632
rect 5252 13572 5256 13628
rect 5256 13572 5312 13628
rect 5312 13572 5316 13628
rect 5252 13568 5316 13572
rect 5332 13628 5396 13632
rect 5332 13572 5336 13628
rect 5336 13572 5392 13628
rect 5392 13572 5396 13628
rect 5332 13568 5396 13572
rect 5412 13628 5476 13632
rect 5412 13572 5416 13628
rect 5416 13572 5472 13628
rect 5472 13572 5476 13628
rect 5412 13568 5476 13572
rect 13613 13628 13677 13632
rect 13613 13572 13617 13628
rect 13617 13572 13673 13628
rect 13673 13572 13677 13628
rect 13613 13568 13677 13572
rect 13693 13628 13757 13632
rect 13693 13572 13697 13628
rect 13697 13572 13753 13628
rect 13753 13572 13757 13628
rect 13693 13568 13757 13572
rect 13773 13628 13837 13632
rect 13773 13572 13777 13628
rect 13777 13572 13833 13628
rect 13833 13572 13837 13628
rect 13773 13568 13837 13572
rect 13853 13628 13917 13632
rect 13853 13572 13857 13628
rect 13857 13572 13913 13628
rect 13913 13572 13917 13628
rect 13853 13568 13917 13572
rect 22054 13628 22118 13632
rect 22054 13572 22058 13628
rect 22058 13572 22114 13628
rect 22114 13572 22118 13628
rect 22054 13568 22118 13572
rect 22134 13628 22198 13632
rect 22134 13572 22138 13628
rect 22138 13572 22194 13628
rect 22194 13572 22198 13628
rect 22134 13568 22198 13572
rect 22214 13628 22278 13632
rect 22214 13572 22218 13628
rect 22218 13572 22274 13628
rect 22274 13572 22278 13628
rect 22214 13568 22278 13572
rect 22294 13628 22358 13632
rect 22294 13572 22298 13628
rect 22298 13572 22354 13628
rect 22354 13572 22358 13628
rect 22294 13568 22358 13572
rect 30495 13628 30559 13632
rect 30495 13572 30499 13628
rect 30499 13572 30555 13628
rect 30555 13572 30559 13628
rect 30495 13568 30559 13572
rect 30575 13628 30639 13632
rect 30575 13572 30579 13628
rect 30579 13572 30635 13628
rect 30635 13572 30639 13628
rect 30575 13568 30639 13572
rect 30655 13628 30719 13632
rect 30655 13572 30659 13628
rect 30659 13572 30715 13628
rect 30715 13572 30719 13628
rect 30655 13568 30719 13572
rect 30735 13628 30799 13632
rect 30735 13572 30739 13628
rect 30739 13572 30795 13628
rect 30795 13572 30799 13628
rect 30735 13568 30799 13572
rect 31892 13560 31956 13564
rect 31892 13504 31906 13560
rect 31906 13504 31956 13560
rect 31892 13500 31956 13504
rect 33732 13500 33796 13564
rect 29132 13364 29196 13428
rect 9392 13084 9456 13088
rect 9392 13028 9396 13084
rect 9396 13028 9452 13084
rect 9452 13028 9456 13084
rect 9392 13024 9456 13028
rect 9472 13084 9536 13088
rect 9472 13028 9476 13084
rect 9476 13028 9532 13084
rect 9532 13028 9536 13084
rect 9472 13024 9536 13028
rect 9552 13084 9616 13088
rect 9552 13028 9556 13084
rect 9556 13028 9612 13084
rect 9612 13028 9616 13084
rect 9552 13024 9616 13028
rect 9632 13084 9696 13088
rect 9632 13028 9636 13084
rect 9636 13028 9692 13084
rect 9692 13028 9696 13084
rect 9632 13024 9696 13028
rect 17833 13084 17897 13088
rect 17833 13028 17837 13084
rect 17837 13028 17893 13084
rect 17893 13028 17897 13084
rect 17833 13024 17897 13028
rect 17913 13084 17977 13088
rect 17913 13028 17917 13084
rect 17917 13028 17973 13084
rect 17973 13028 17977 13084
rect 17913 13024 17977 13028
rect 17993 13084 18057 13088
rect 17993 13028 17997 13084
rect 17997 13028 18053 13084
rect 18053 13028 18057 13084
rect 17993 13024 18057 13028
rect 18073 13084 18137 13088
rect 18073 13028 18077 13084
rect 18077 13028 18133 13084
rect 18133 13028 18137 13084
rect 18073 13024 18137 13028
rect 26274 13084 26338 13088
rect 26274 13028 26278 13084
rect 26278 13028 26334 13084
rect 26334 13028 26338 13084
rect 26274 13024 26338 13028
rect 26354 13084 26418 13088
rect 26354 13028 26358 13084
rect 26358 13028 26414 13084
rect 26414 13028 26418 13084
rect 26354 13024 26418 13028
rect 26434 13084 26498 13088
rect 26434 13028 26438 13084
rect 26438 13028 26494 13084
rect 26494 13028 26498 13084
rect 26434 13024 26498 13028
rect 26514 13084 26578 13088
rect 26514 13028 26518 13084
rect 26518 13028 26574 13084
rect 26574 13028 26578 13084
rect 26514 13024 26578 13028
rect 34715 13084 34779 13088
rect 34715 13028 34719 13084
rect 34719 13028 34775 13084
rect 34775 13028 34779 13084
rect 34715 13024 34779 13028
rect 34795 13084 34859 13088
rect 34795 13028 34799 13084
rect 34799 13028 34855 13084
rect 34855 13028 34859 13084
rect 34795 13024 34859 13028
rect 34875 13084 34939 13088
rect 34875 13028 34879 13084
rect 34879 13028 34935 13084
rect 34935 13028 34939 13084
rect 34875 13024 34939 13028
rect 34955 13084 35019 13088
rect 34955 13028 34959 13084
rect 34959 13028 35015 13084
rect 35015 13028 35019 13084
rect 34955 13024 35019 13028
rect 5172 12540 5236 12544
rect 5172 12484 5176 12540
rect 5176 12484 5232 12540
rect 5232 12484 5236 12540
rect 5172 12480 5236 12484
rect 5252 12540 5316 12544
rect 5252 12484 5256 12540
rect 5256 12484 5312 12540
rect 5312 12484 5316 12540
rect 5252 12480 5316 12484
rect 5332 12540 5396 12544
rect 5332 12484 5336 12540
rect 5336 12484 5392 12540
rect 5392 12484 5396 12540
rect 5332 12480 5396 12484
rect 5412 12540 5476 12544
rect 5412 12484 5416 12540
rect 5416 12484 5472 12540
rect 5472 12484 5476 12540
rect 5412 12480 5476 12484
rect 13613 12540 13677 12544
rect 13613 12484 13617 12540
rect 13617 12484 13673 12540
rect 13673 12484 13677 12540
rect 13613 12480 13677 12484
rect 13693 12540 13757 12544
rect 13693 12484 13697 12540
rect 13697 12484 13753 12540
rect 13753 12484 13757 12540
rect 13693 12480 13757 12484
rect 13773 12540 13837 12544
rect 13773 12484 13777 12540
rect 13777 12484 13833 12540
rect 13833 12484 13837 12540
rect 13773 12480 13837 12484
rect 13853 12540 13917 12544
rect 13853 12484 13857 12540
rect 13857 12484 13913 12540
rect 13913 12484 13917 12540
rect 13853 12480 13917 12484
rect 22054 12540 22118 12544
rect 22054 12484 22058 12540
rect 22058 12484 22114 12540
rect 22114 12484 22118 12540
rect 22054 12480 22118 12484
rect 22134 12540 22198 12544
rect 22134 12484 22138 12540
rect 22138 12484 22194 12540
rect 22194 12484 22198 12540
rect 22134 12480 22198 12484
rect 22214 12540 22278 12544
rect 22214 12484 22218 12540
rect 22218 12484 22274 12540
rect 22274 12484 22278 12540
rect 22214 12480 22278 12484
rect 22294 12540 22358 12544
rect 22294 12484 22298 12540
rect 22298 12484 22354 12540
rect 22354 12484 22358 12540
rect 22294 12480 22358 12484
rect 30495 12540 30559 12544
rect 30495 12484 30499 12540
rect 30499 12484 30555 12540
rect 30555 12484 30559 12540
rect 30495 12480 30559 12484
rect 30575 12540 30639 12544
rect 30575 12484 30579 12540
rect 30579 12484 30635 12540
rect 30635 12484 30639 12540
rect 30575 12480 30639 12484
rect 30655 12540 30719 12544
rect 30655 12484 30659 12540
rect 30659 12484 30715 12540
rect 30715 12484 30719 12540
rect 30655 12480 30719 12484
rect 30735 12540 30799 12544
rect 30735 12484 30739 12540
rect 30739 12484 30795 12540
rect 30795 12484 30799 12540
rect 30735 12480 30799 12484
rect 9392 11996 9456 12000
rect 9392 11940 9396 11996
rect 9396 11940 9452 11996
rect 9452 11940 9456 11996
rect 9392 11936 9456 11940
rect 9472 11996 9536 12000
rect 9472 11940 9476 11996
rect 9476 11940 9532 11996
rect 9532 11940 9536 11996
rect 9472 11936 9536 11940
rect 9552 11996 9616 12000
rect 9552 11940 9556 11996
rect 9556 11940 9612 11996
rect 9612 11940 9616 11996
rect 9552 11936 9616 11940
rect 9632 11996 9696 12000
rect 9632 11940 9636 11996
rect 9636 11940 9692 11996
rect 9692 11940 9696 11996
rect 9632 11936 9696 11940
rect 17833 11996 17897 12000
rect 17833 11940 17837 11996
rect 17837 11940 17893 11996
rect 17893 11940 17897 11996
rect 17833 11936 17897 11940
rect 17913 11996 17977 12000
rect 17913 11940 17917 11996
rect 17917 11940 17973 11996
rect 17973 11940 17977 11996
rect 17913 11936 17977 11940
rect 17993 11996 18057 12000
rect 17993 11940 17997 11996
rect 17997 11940 18053 11996
rect 18053 11940 18057 11996
rect 17993 11936 18057 11940
rect 18073 11996 18137 12000
rect 18073 11940 18077 11996
rect 18077 11940 18133 11996
rect 18133 11940 18137 11996
rect 18073 11936 18137 11940
rect 26274 11996 26338 12000
rect 26274 11940 26278 11996
rect 26278 11940 26334 11996
rect 26334 11940 26338 11996
rect 26274 11936 26338 11940
rect 26354 11996 26418 12000
rect 26354 11940 26358 11996
rect 26358 11940 26414 11996
rect 26414 11940 26418 11996
rect 26354 11936 26418 11940
rect 26434 11996 26498 12000
rect 26434 11940 26438 11996
rect 26438 11940 26494 11996
rect 26494 11940 26498 11996
rect 26434 11936 26498 11940
rect 26514 11996 26578 12000
rect 26514 11940 26518 11996
rect 26518 11940 26574 11996
rect 26574 11940 26578 11996
rect 26514 11936 26578 11940
rect 34715 11996 34779 12000
rect 34715 11940 34719 11996
rect 34719 11940 34775 11996
rect 34775 11940 34779 11996
rect 34715 11936 34779 11940
rect 34795 11996 34859 12000
rect 34795 11940 34799 11996
rect 34799 11940 34855 11996
rect 34855 11940 34859 11996
rect 34795 11936 34859 11940
rect 34875 11996 34939 12000
rect 34875 11940 34879 11996
rect 34879 11940 34935 11996
rect 34935 11940 34939 11996
rect 34875 11936 34939 11940
rect 34955 11996 35019 12000
rect 34955 11940 34959 11996
rect 34959 11940 35015 11996
rect 35015 11940 35019 11996
rect 34955 11936 35019 11940
rect 34100 11732 34164 11796
rect 5172 11452 5236 11456
rect 5172 11396 5176 11452
rect 5176 11396 5232 11452
rect 5232 11396 5236 11452
rect 5172 11392 5236 11396
rect 5252 11452 5316 11456
rect 5252 11396 5256 11452
rect 5256 11396 5312 11452
rect 5312 11396 5316 11452
rect 5252 11392 5316 11396
rect 5332 11452 5396 11456
rect 5332 11396 5336 11452
rect 5336 11396 5392 11452
rect 5392 11396 5396 11452
rect 5332 11392 5396 11396
rect 5412 11452 5476 11456
rect 5412 11396 5416 11452
rect 5416 11396 5472 11452
rect 5472 11396 5476 11452
rect 5412 11392 5476 11396
rect 13613 11452 13677 11456
rect 13613 11396 13617 11452
rect 13617 11396 13673 11452
rect 13673 11396 13677 11452
rect 13613 11392 13677 11396
rect 13693 11452 13757 11456
rect 13693 11396 13697 11452
rect 13697 11396 13753 11452
rect 13753 11396 13757 11452
rect 13693 11392 13757 11396
rect 13773 11452 13837 11456
rect 13773 11396 13777 11452
rect 13777 11396 13833 11452
rect 13833 11396 13837 11452
rect 13773 11392 13837 11396
rect 13853 11452 13917 11456
rect 13853 11396 13857 11452
rect 13857 11396 13913 11452
rect 13913 11396 13917 11452
rect 13853 11392 13917 11396
rect 22054 11452 22118 11456
rect 22054 11396 22058 11452
rect 22058 11396 22114 11452
rect 22114 11396 22118 11452
rect 22054 11392 22118 11396
rect 22134 11452 22198 11456
rect 22134 11396 22138 11452
rect 22138 11396 22194 11452
rect 22194 11396 22198 11452
rect 22134 11392 22198 11396
rect 22214 11452 22278 11456
rect 22214 11396 22218 11452
rect 22218 11396 22274 11452
rect 22274 11396 22278 11452
rect 22214 11392 22278 11396
rect 22294 11452 22358 11456
rect 22294 11396 22298 11452
rect 22298 11396 22354 11452
rect 22354 11396 22358 11452
rect 22294 11392 22358 11396
rect 30495 11452 30559 11456
rect 30495 11396 30499 11452
rect 30499 11396 30555 11452
rect 30555 11396 30559 11452
rect 30495 11392 30559 11396
rect 30575 11452 30639 11456
rect 30575 11396 30579 11452
rect 30579 11396 30635 11452
rect 30635 11396 30639 11452
rect 30575 11392 30639 11396
rect 30655 11452 30719 11456
rect 30655 11396 30659 11452
rect 30659 11396 30715 11452
rect 30715 11396 30719 11452
rect 30655 11392 30719 11396
rect 30735 11452 30799 11456
rect 30735 11396 30739 11452
rect 30739 11396 30795 11452
rect 30795 11396 30799 11452
rect 30735 11392 30799 11396
rect 9392 10908 9456 10912
rect 9392 10852 9396 10908
rect 9396 10852 9452 10908
rect 9452 10852 9456 10908
rect 9392 10848 9456 10852
rect 9472 10908 9536 10912
rect 9472 10852 9476 10908
rect 9476 10852 9532 10908
rect 9532 10852 9536 10908
rect 9472 10848 9536 10852
rect 9552 10908 9616 10912
rect 9552 10852 9556 10908
rect 9556 10852 9612 10908
rect 9612 10852 9616 10908
rect 9552 10848 9616 10852
rect 9632 10908 9696 10912
rect 9632 10852 9636 10908
rect 9636 10852 9692 10908
rect 9692 10852 9696 10908
rect 9632 10848 9696 10852
rect 17833 10908 17897 10912
rect 17833 10852 17837 10908
rect 17837 10852 17893 10908
rect 17893 10852 17897 10908
rect 17833 10848 17897 10852
rect 17913 10908 17977 10912
rect 17913 10852 17917 10908
rect 17917 10852 17973 10908
rect 17973 10852 17977 10908
rect 17913 10848 17977 10852
rect 17993 10908 18057 10912
rect 17993 10852 17997 10908
rect 17997 10852 18053 10908
rect 18053 10852 18057 10908
rect 17993 10848 18057 10852
rect 18073 10908 18137 10912
rect 18073 10852 18077 10908
rect 18077 10852 18133 10908
rect 18133 10852 18137 10908
rect 18073 10848 18137 10852
rect 26274 10908 26338 10912
rect 26274 10852 26278 10908
rect 26278 10852 26334 10908
rect 26334 10852 26338 10908
rect 26274 10848 26338 10852
rect 26354 10908 26418 10912
rect 26354 10852 26358 10908
rect 26358 10852 26414 10908
rect 26414 10852 26418 10908
rect 26354 10848 26418 10852
rect 26434 10908 26498 10912
rect 26434 10852 26438 10908
rect 26438 10852 26494 10908
rect 26494 10852 26498 10908
rect 26434 10848 26498 10852
rect 26514 10908 26578 10912
rect 26514 10852 26518 10908
rect 26518 10852 26574 10908
rect 26574 10852 26578 10908
rect 26514 10848 26578 10852
rect 34715 10908 34779 10912
rect 34715 10852 34719 10908
rect 34719 10852 34775 10908
rect 34775 10852 34779 10908
rect 34715 10848 34779 10852
rect 34795 10908 34859 10912
rect 34795 10852 34799 10908
rect 34799 10852 34855 10908
rect 34855 10852 34859 10908
rect 34795 10848 34859 10852
rect 34875 10908 34939 10912
rect 34875 10852 34879 10908
rect 34879 10852 34935 10908
rect 34935 10852 34939 10908
rect 34875 10848 34939 10852
rect 34955 10908 35019 10912
rect 34955 10852 34959 10908
rect 34959 10852 35015 10908
rect 35015 10852 35019 10908
rect 34955 10848 35019 10852
rect 5172 10364 5236 10368
rect 5172 10308 5176 10364
rect 5176 10308 5232 10364
rect 5232 10308 5236 10364
rect 5172 10304 5236 10308
rect 5252 10364 5316 10368
rect 5252 10308 5256 10364
rect 5256 10308 5312 10364
rect 5312 10308 5316 10364
rect 5252 10304 5316 10308
rect 5332 10364 5396 10368
rect 5332 10308 5336 10364
rect 5336 10308 5392 10364
rect 5392 10308 5396 10364
rect 5332 10304 5396 10308
rect 5412 10364 5476 10368
rect 5412 10308 5416 10364
rect 5416 10308 5472 10364
rect 5472 10308 5476 10364
rect 5412 10304 5476 10308
rect 13613 10364 13677 10368
rect 13613 10308 13617 10364
rect 13617 10308 13673 10364
rect 13673 10308 13677 10364
rect 13613 10304 13677 10308
rect 13693 10364 13757 10368
rect 13693 10308 13697 10364
rect 13697 10308 13753 10364
rect 13753 10308 13757 10364
rect 13693 10304 13757 10308
rect 13773 10364 13837 10368
rect 13773 10308 13777 10364
rect 13777 10308 13833 10364
rect 13833 10308 13837 10364
rect 13773 10304 13837 10308
rect 13853 10364 13917 10368
rect 13853 10308 13857 10364
rect 13857 10308 13913 10364
rect 13913 10308 13917 10364
rect 13853 10304 13917 10308
rect 22054 10364 22118 10368
rect 22054 10308 22058 10364
rect 22058 10308 22114 10364
rect 22114 10308 22118 10364
rect 22054 10304 22118 10308
rect 22134 10364 22198 10368
rect 22134 10308 22138 10364
rect 22138 10308 22194 10364
rect 22194 10308 22198 10364
rect 22134 10304 22198 10308
rect 22214 10364 22278 10368
rect 22214 10308 22218 10364
rect 22218 10308 22274 10364
rect 22274 10308 22278 10364
rect 22214 10304 22278 10308
rect 22294 10364 22358 10368
rect 22294 10308 22298 10364
rect 22298 10308 22354 10364
rect 22354 10308 22358 10364
rect 22294 10304 22358 10308
rect 30495 10364 30559 10368
rect 30495 10308 30499 10364
rect 30499 10308 30555 10364
rect 30555 10308 30559 10364
rect 30495 10304 30559 10308
rect 30575 10364 30639 10368
rect 30575 10308 30579 10364
rect 30579 10308 30635 10364
rect 30635 10308 30639 10364
rect 30575 10304 30639 10308
rect 30655 10364 30719 10368
rect 30655 10308 30659 10364
rect 30659 10308 30715 10364
rect 30715 10308 30719 10364
rect 30655 10304 30719 10308
rect 30735 10364 30799 10368
rect 30735 10308 30739 10364
rect 30739 10308 30795 10364
rect 30795 10308 30799 10364
rect 30735 10304 30799 10308
rect 9392 9820 9456 9824
rect 9392 9764 9396 9820
rect 9396 9764 9452 9820
rect 9452 9764 9456 9820
rect 9392 9760 9456 9764
rect 9472 9820 9536 9824
rect 9472 9764 9476 9820
rect 9476 9764 9532 9820
rect 9532 9764 9536 9820
rect 9472 9760 9536 9764
rect 9552 9820 9616 9824
rect 9552 9764 9556 9820
rect 9556 9764 9612 9820
rect 9612 9764 9616 9820
rect 9552 9760 9616 9764
rect 9632 9820 9696 9824
rect 9632 9764 9636 9820
rect 9636 9764 9692 9820
rect 9692 9764 9696 9820
rect 9632 9760 9696 9764
rect 17833 9820 17897 9824
rect 17833 9764 17837 9820
rect 17837 9764 17893 9820
rect 17893 9764 17897 9820
rect 17833 9760 17897 9764
rect 17913 9820 17977 9824
rect 17913 9764 17917 9820
rect 17917 9764 17973 9820
rect 17973 9764 17977 9820
rect 17913 9760 17977 9764
rect 17993 9820 18057 9824
rect 17993 9764 17997 9820
rect 17997 9764 18053 9820
rect 18053 9764 18057 9820
rect 17993 9760 18057 9764
rect 18073 9820 18137 9824
rect 18073 9764 18077 9820
rect 18077 9764 18133 9820
rect 18133 9764 18137 9820
rect 18073 9760 18137 9764
rect 26274 9820 26338 9824
rect 26274 9764 26278 9820
rect 26278 9764 26334 9820
rect 26334 9764 26338 9820
rect 26274 9760 26338 9764
rect 26354 9820 26418 9824
rect 26354 9764 26358 9820
rect 26358 9764 26414 9820
rect 26414 9764 26418 9820
rect 26354 9760 26418 9764
rect 26434 9820 26498 9824
rect 26434 9764 26438 9820
rect 26438 9764 26494 9820
rect 26494 9764 26498 9820
rect 26434 9760 26498 9764
rect 26514 9820 26578 9824
rect 26514 9764 26518 9820
rect 26518 9764 26574 9820
rect 26574 9764 26578 9820
rect 26514 9760 26578 9764
rect 34715 9820 34779 9824
rect 34715 9764 34719 9820
rect 34719 9764 34775 9820
rect 34775 9764 34779 9820
rect 34715 9760 34779 9764
rect 34795 9820 34859 9824
rect 34795 9764 34799 9820
rect 34799 9764 34855 9820
rect 34855 9764 34859 9820
rect 34795 9760 34859 9764
rect 34875 9820 34939 9824
rect 34875 9764 34879 9820
rect 34879 9764 34935 9820
rect 34935 9764 34939 9820
rect 34875 9760 34939 9764
rect 34955 9820 35019 9824
rect 34955 9764 34959 9820
rect 34959 9764 35015 9820
rect 35015 9764 35019 9820
rect 34955 9760 35019 9764
rect 5172 9276 5236 9280
rect 5172 9220 5176 9276
rect 5176 9220 5232 9276
rect 5232 9220 5236 9276
rect 5172 9216 5236 9220
rect 5252 9276 5316 9280
rect 5252 9220 5256 9276
rect 5256 9220 5312 9276
rect 5312 9220 5316 9276
rect 5252 9216 5316 9220
rect 5332 9276 5396 9280
rect 5332 9220 5336 9276
rect 5336 9220 5392 9276
rect 5392 9220 5396 9276
rect 5332 9216 5396 9220
rect 5412 9276 5476 9280
rect 5412 9220 5416 9276
rect 5416 9220 5472 9276
rect 5472 9220 5476 9276
rect 5412 9216 5476 9220
rect 13613 9276 13677 9280
rect 13613 9220 13617 9276
rect 13617 9220 13673 9276
rect 13673 9220 13677 9276
rect 13613 9216 13677 9220
rect 13693 9276 13757 9280
rect 13693 9220 13697 9276
rect 13697 9220 13753 9276
rect 13753 9220 13757 9276
rect 13693 9216 13757 9220
rect 13773 9276 13837 9280
rect 13773 9220 13777 9276
rect 13777 9220 13833 9276
rect 13833 9220 13837 9276
rect 13773 9216 13837 9220
rect 13853 9276 13917 9280
rect 13853 9220 13857 9276
rect 13857 9220 13913 9276
rect 13913 9220 13917 9276
rect 13853 9216 13917 9220
rect 22054 9276 22118 9280
rect 22054 9220 22058 9276
rect 22058 9220 22114 9276
rect 22114 9220 22118 9276
rect 22054 9216 22118 9220
rect 22134 9276 22198 9280
rect 22134 9220 22138 9276
rect 22138 9220 22194 9276
rect 22194 9220 22198 9276
rect 22134 9216 22198 9220
rect 22214 9276 22278 9280
rect 22214 9220 22218 9276
rect 22218 9220 22274 9276
rect 22274 9220 22278 9276
rect 22214 9216 22278 9220
rect 22294 9276 22358 9280
rect 22294 9220 22298 9276
rect 22298 9220 22354 9276
rect 22354 9220 22358 9276
rect 22294 9216 22358 9220
rect 30495 9276 30559 9280
rect 30495 9220 30499 9276
rect 30499 9220 30555 9276
rect 30555 9220 30559 9276
rect 30495 9216 30559 9220
rect 30575 9276 30639 9280
rect 30575 9220 30579 9276
rect 30579 9220 30635 9276
rect 30635 9220 30639 9276
rect 30575 9216 30639 9220
rect 30655 9276 30719 9280
rect 30655 9220 30659 9276
rect 30659 9220 30715 9276
rect 30715 9220 30719 9276
rect 30655 9216 30719 9220
rect 30735 9276 30799 9280
rect 30735 9220 30739 9276
rect 30739 9220 30795 9276
rect 30795 9220 30799 9276
rect 30735 9216 30799 9220
rect 9392 8732 9456 8736
rect 9392 8676 9396 8732
rect 9396 8676 9452 8732
rect 9452 8676 9456 8732
rect 9392 8672 9456 8676
rect 9472 8732 9536 8736
rect 9472 8676 9476 8732
rect 9476 8676 9532 8732
rect 9532 8676 9536 8732
rect 9472 8672 9536 8676
rect 9552 8732 9616 8736
rect 9552 8676 9556 8732
rect 9556 8676 9612 8732
rect 9612 8676 9616 8732
rect 9552 8672 9616 8676
rect 9632 8732 9696 8736
rect 9632 8676 9636 8732
rect 9636 8676 9692 8732
rect 9692 8676 9696 8732
rect 9632 8672 9696 8676
rect 17833 8732 17897 8736
rect 17833 8676 17837 8732
rect 17837 8676 17893 8732
rect 17893 8676 17897 8732
rect 17833 8672 17897 8676
rect 17913 8732 17977 8736
rect 17913 8676 17917 8732
rect 17917 8676 17973 8732
rect 17973 8676 17977 8732
rect 17913 8672 17977 8676
rect 17993 8732 18057 8736
rect 17993 8676 17997 8732
rect 17997 8676 18053 8732
rect 18053 8676 18057 8732
rect 17993 8672 18057 8676
rect 18073 8732 18137 8736
rect 18073 8676 18077 8732
rect 18077 8676 18133 8732
rect 18133 8676 18137 8732
rect 18073 8672 18137 8676
rect 26274 8732 26338 8736
rect 26274 8676 26278 8732
rect 26278 8676 26334 8732
rect 26334 8676 26338 8732
rect 26274 8672 26338 8676
rect 26354 8732 26418 8736
rect 26354 8676 26358 8732
rect 26358 8676 26414 8732
rect 26414 8676 26418 8732
rect 26354 8672 26418 8676
rect 26434 8732 26498 8736
rect 26434 8676 26438 8732
rect 26438 8676 26494 8732
rect 26494 8676 26498 8732
rect 26434 8672 26498 8676
rect 26514 8732 26578 8736
rect 26514 8676 26518 8732
rect 26518 8676 26574 8732
rect 26574 8676 26578 8732
rect 26514 8672 26578 8676
rect 34715 8732 34779 8736
rect 34715 8676 34719 8732
rect 34719 8676 34775 8732
rect 34775 8676 34779 8732
rect 34715 8672 34779 8676
rect 34795 8732 34859 8736
rect 34795 8676 34799 8732
rect 34799 8676 34855 8732
rect 34855 8676 34859 8732
rect 34795 8672 34859 8676
rect 34875 8732 34939 8736
rect 34875 8676 34879 8732
rect 34879 8676 34935 8732
rect 34935 8676 34939 8732
rect 34875 8672 34939 8676
rect 34955 8732 35019 8736
rect 34955 8676 34959 8732
rect 34959 8676 35015 8732
rect 35015 8676 35019 8732
rect 34955 8672 35019 8676
rect 5172 8188 5236 8192
rect 5172 8132 5176 8188
rect 5176 8132 5232 8188
rect 5232 8132 5236 8188
rect 5172 8128 5236 8132
rect 5252 8188 5316 8192
rect 5252 8132 5256 8188
rect 5256 8132 5312 8188
rect 5312 8132 5316 8188
rect 5252 8128 5316 8132
rect 5332 8188 5396 8192
rect 5332 8132 5336 8188
rect 5336 8132 5392 8188
rect 5392 8132 5396 8188
rect 5332 8128 5396 8132
rect 5412 8188 5476 8192
rect 5412 8132 5416 8188
rect 5416 8132 5472 8188
rect 5472 8132 5476 8188
rect 5412 8128 5476 8132
rect 13613 8188 13677 8192
rect 13613 8132 13617 8188
rect 13617 8132 13673 8188
rect 13673 8132 13677 8188
rect 13613 8128 13677 8132
rect 13693 8188 13757 8192
rect 13693 8132 13697 8188
rect 13697 8132 13753 8188
rect 13753 8132 13757 8188
rect 13693 8128 13757 8132
rect 13773 8188 13837 8192
rect 13773 8132 13777 8188
rect 13777 8132 13833 8188
rect 13833 8132 13837 8188
rect 13773 8128 13837 8132
rect 13853 8188 13917 8192
rect 13853 8132 13857 8188
rect 13857 8132 13913 8188
rect 13913 8132 13917 8188
rect 13853 8128 13917 8132
rect 22054 8188 22118 8192
rect 22054 8132 22058 8188
rect 22058 8132 22114 8188
rect 22114 8132 22118 8188
rect 22054 8128 22118 8132
rect 22134 8188 22198 8192
rect 22134 8132 22138 8188
rect 22138 8132 22194 8188
rect 22194 8132 22198 8188
rect 22134 8128 22198 8132
rect 22214 8188 22278 8192
rect 22214 8132 22218 8188
rect 22218 8132 22274 8188
rect 22274 8132 22278 8188
rect 22214 8128 22278 8132
rect 22294 8188 22358 8192
rect 22294 8132 22298 8188
rect 22298 8132 22354 8188
rect 22354 8132 22358 8188
rect 22294 8128 22358 8132
rect 30495 8188 30559 8192
rect 30495 8132 30499 8188
rect 30499 8132 30555 8188
rect 30555 8132 30559 8188
rect 30495 8128 30559 8132
rect 30575 8188 30639 8192
rect 30575 8132 30579 8188
rect 30579 8132 30635 8188
rect 30635 8132 30639 8188
rect 30575 8128 30639 8132
rect 30655 8188 30719 8192
rect 30655 8132 30659 8188
rect 30659 8132 30715 8188
rect 30715 8132 30719 8188
rect 30655 8128 30719 8132
rect 30735 8188 30799 8192
rect 30735 8132 30739 8188
rect 30739 8132 30795 8188
rect 30795 8132 30799 8188
rect 30735 8128 30799 8132
rect 9392 7644 9456 7648
rect 9392 7588 9396 7644
rect 9396 7588 9452 7644
rect 9452 7588 9456 7644
rect 9392 7584 9456 7588
rect 9472 7644 9536 7648
rect 9472 7588 9476 7644
rect 9476 7588 9532 7644
rect 9532 7588 9536 7644
rect 9472 7584 9536 7588
rect 9552 7644 9616 7648
rect 9552 7588 9556 7644
rect 9556 7588 9612 7644
rect 9612 7588 9616 7644
rect 9552 7584 9616 7588
rect 9632 7644 9696 7648
rect 9632 7588 9636 7644
rect 9636 7588 9692 7644
rect 9692 7588 9696 7644
rect 9632 7584 9696 7588
rect 17833 7644 17897 7648
rect 17833 7588 17837 7644
rect 17837 7588 17893 7644
rect 17893 7588 17897 7644
rect 17833 7584 17897 7588
rect 17913 7644 17977 7648
rect 17913 7588 17917 7644
rect 17917 7588 17973 7644
rect 17973 7588 17977 7644
rect 17913 7584 17977 7588
rect 17993 7644 18057 7648
rect 17993 7588 17997 7644
rect 17997 7588 18053 7644
rect 18053 7588 18057 7644
rect 17993 7584 18057 7588
rect 18073 7644 18137 7648
rect 18073 7588 18077 7644
rect 18077 7588 18133 7644
rect 18133 7588 18137 7644
rect 18073 7584 18137 7588
rect 26274 7644 26338 7648
rect 26274 7588 26278 7644
rect 26278 7588 26334 7644
rect 26334 7588 26338 7644
rect 26274 7584 26338 7588
rect 26354 7644 26418 7648
rect 26354 7588 26358 7644
rect 26358 7588 26414 7644
rect 26414 7588 26418 7644
rect 26354 7584 26418 7588
rect 26434 7644 26498 7648
rect 26434 7588 26438 7644
rect 26438 7588 26494 7644
rect 26494 7588 26498 7644
rect 26434 7584 26498 7588
rect 26514 7644 26578 7648
rect 26514 7588 26518 7644
rect 26518 7588 26574 7644
rect 26574 7588 26578 7644
rect 26514 7584 26578 7588
rect 34715 7644 34779 7648
rect 34715 7588 34719 7644
rect 34719 7588 34775 7644
rect 34775 7588 34779 7644
rect 34715 7584 34779 7588
rect 34795 7644 34859 7648
rect 34795 7588 34799 7644
rect 34799 7588 34855 7644
rect 34855 7588 34859 7644
rect 34795 7584 34859 7588
rect 34875 7644 34939 7648
rect 34875 7588 34879 7644
rect 34879 7588 34935 7644
rect 34935 7588 34939 7644
rect 34875 7584 34939 7588
rect 34955 7644 35019 7648
rect 34955 7588 34959 7644
rect 34959 7588 35015 7644
rect 35015 7588 35019 7644
rect 34955 7584 35019 7588
rect 5172 7100 5236 7104
rect 5172 7044 5176 7100
rect 5176 7044 5232 7100
rect 5232 7044 5236 7100
rect 5172 7040 5236 7044
rect 5252 7100 5316 7104
rect 5252 7044 5256 7100
rect 5256 7044 5312 7100
rect 5312 7044 5316 7100
rect 5252 7040 5316 7044
rect 5332 7100 5396 7104
rect 5332 7044 5336 7100
rect 5336 7044 5392 7100
rect 5392 7044 5396 7100
rect 5332 7040 5396 7044
rect 5412 7100 5476 7104
rect 5412 7044 5416 7100
rect 5416 7044 5472 7100
rect 5472 7044 5476 7100
rect 5412 7040 5476 7044
rect 13613 7100 13677 7104
rect 13613 7044 13617 7100
rect 13617 7044 13673 7100
rect 13673 7044 13677 7100
rect 13613 7040 13677 7044
rect 13693 7100 13757 7104
rect 13693 7044 13697 7100
rect 13697 7044 13753 7100
rect 13753 7044 13757 7100
rect 13693 7040 13757 7044
rect 13773 7100 13837 7104
rect 13773 7044 13777 7100
rect 13777 7044 13833 7100
rect 13833 7044 13837 7100
rect 13773 7040 13837 7044
rect 13853 7100 13917 7104
rect 13853 7044 13857 7100
rect 13857 7044 13913 7100
rect 13913 7044 13917 7100
rect 13853 7040 13917 7044
rect 22054 7100 22118 7104
rect 22054 7044 22058 7100
rect 22058 7044 22114 7100
rect 22114 7044 22118 7100
rect 22054 7040 22118 7044
rect 22134 7100 22198 7104
rect 22134 7044 22138 7100
rect 22138 7044 22194 7100
rect 22194 7044 22198 7100
rect 22134 7040 22198 7044
rect 22214 7100 22278 7104
rect 22214 7044 22218 7100
rect 22218 7044 22274 7100
rect 22274 7044 22278 7100
rect 22214 7040 22278 7044
rect 22294 7100 22358 7104
rect 22294 7044 22298 7100
rect 22298 7044 22354 7100
rect 22354 7044 22358 7100
rect 22294 7040 22358 7044
rect 30495 7100 30559 7104
rect 30495 7044 30499 7100
rect 30499 7044 30555 7100
rect 30555 7044 30559 7100
rect 30495 7040 30559 7044
rect 30575 7100 30639 7104
rect 30575 7044 30579 7100
rect 30579 7044 30635 7100
rect 30635 7044 30639 7100
rect 30575 7040 30639 7044
rect 30655 7100 30719 7104
rect 30655 7044 30659 7100
rect 30659 7044 30715 7100
rect 30715 7044 30719 7100
rect 30655 7040 30719 7044
rect 30735 7100 30799 7104
rect 30735 7044 30739 7100
rect 30739 7044 30795 7100
rect 30795 7044 30799 7100
rect 30735 7040 30799 7044
rect 9392 6556 9456 6560
rect 9392 6500 9396 6556
rect 9396 6500 9452 6556
rect 9452 6500 9456 6556
rect 9392 6496 9456 6500
rect 9472 6556 9536 6560
rect 9472 6500 9476 6556
rect 9476 6500 9532 6556
rect 9532 6500 9536 6556
rect 9472 6496 9536 6500
rect 9552 6556 9616 6560
rect 9552 6500 9556 6556
rect 9556 6500 9612 6556
rect 9612 6500 9616 6556
rect 9552 6496 9616 6500
rect 9632 6556 9696 6560
rect 9632 6500 9636 6556
rect 9636 6500 9692 6556
rect 9692 6500 9696 6556
rect 9632 6496 9696 6500
rect 17833 6556 17897 6560
rect 17833 6500 17837 6556
rect 17837 6500 17893 6556
rect 17893 6500 17897 6556
rect 17833 6496 17897 6500
rect 17913 6556 17977 6560
rect 17913 6500 17917 6556
rect 17917 6500 17973 6556
rect 17973 6500 17977 6556
rect 17913 6496 17977 6500
rect 17993 6556 18057 6560
rect 17993 6500 17997 6556
rect 17997 6500 18053 6556
rect 18053 6500 18057 6556
rect 17993 6496 18057 6500
rect 18073 6556 18137 6560
rect 18073 6500 18077 6556
rect 18077 6500 18133 6556
rect 18133 6500 18137 6556
rect 18073 6496 18137 6500
rect 26274 6556 26338 6560
rect 26274 6500 26278 6556
rect 26278 6500 26334 6556
rect 26334 6500 26338 6556
rect 26274 6496 26338 6500
rect 26354 6556 26418 6560
rect 26354 6500 26358 6556
rect 26358 6500 26414 6556
rect 26414 6500 26418 6556
rect 26354 6496 26418 6500
rect 26434 6556 26498 6560
rect 26434 6500 26438 6556
rect 26438 6500 26494 6556
rect 26494 6500 26498 6556
rect 26434 6496 26498 6500
rect 26514 6556 26578 6560
rect 26514 6500 26518 6556
rect 26518 6500 26574 6556
rect 26574 6500 26578 6556
rect 26514 6496 26578 6500
rect 34715 6556 34779 6560
rect 34715 6500 34719 6556
rect 34719 6500 34775 6556
rect 34775 6500 34779 6556
rect 34715 6496 34779 6500
rect 34795 6556 34859 6560
rect 34795 6500 34799 6556
rect 34799 6500 34855 6556
rect 34855 6500 34859 6556
rect 34795 6496 34859 6500
rect 34875 6556 34939 6560
rect 34875 6500 34879 6556
rect 34879 6500 34935 6556
rect 34935 6500 34939 6556
rect 34875 6496 34939 6500
rect 34955 6556 35019 6560
rect 34955 6500 34959 6556
rect 34959 6500 35015 6556
rect 35015 6500 35019 6556
rect 34955 6496 35019 6500
rect 5172 6012 5236 6016
rect 5172 5956 5176 6012
rect 5176 5956 5232 6012
rect 5232 5956 5236 6012
rect 5172 5952 5236 5956
rect 5252 6012 5316 6016
rect 5252 5956 5256 6012
rect 5256 5956 5312 6012
rect 5312 5956 5316 6012
rect 5252 5952 5316 5956
rect 5332 6012 5396 6016
rect 5332 5956 5336 6012
rect 5336 5956 5392 6012
rect 5392 5956 5396 6012
rect 5332 5952 5396 5956
rect 5412 6012 5476 6016
rect 5412 5956 5416 6012
rect 5416 5956 5472 6012
rect 5472 5956 5476 6012
rect 5412 5952 5476 5956
rect 13613 6012 13677 6016
rect 13613 5956 13617 6012
rect 13617 5956 13673 6012
rect 13673 5956 13677 6012
rect 13613 5952 13677 5956
rect 13693 6012 13757 6016
rect 13693 5956 13697 6012
rect 13697 5956 13753 6012
rect 13753 5956 13757 6012
rect 13693 5952 13757 5956
rect 13773 6012 13837 6016
rect 13773 5956 13777 6012
rect 13777 5956 13833 6012
rect 13833 5956 13837 6012
rect 13773 5952 13837 5956
rect 13853 6012 13917 6016
rect 13853 5956 13857 6012
rect 13857 5956 13913 6012
rect 13913 5956 13917 6012
rect 13853 5952 13917 5956
rect 22054 6012 22118 6016
rect 22054 5956 22058 6012
rect 22058 5956 22114 6012
rect 22114 5956 22118 6012
rect 22054 5952 22118 5956
rect 22134 6012 22198 6016
rect 22134 5956 22138 6012
rect 22138 5956 22194 6012
rect 22194 5956 22198 6012
rect 22134 5952 22198 5956
rect 22214 6012 22278 6016
rect 22214 5956 22218 6012
rect 22218 5956 22274 6012
rect 22274 5956 22278 6012
rect 22214 5952 22278 5956
rect 22294 6012 22358 6016
rect 22294 5956 22298 6012
rect 22298 5956 22354 6012
rect 22354 5956 22358 6012
rect 22294 5952 22358 5956
rect 30495 6012 30559 6016
rect 30495 5956 30499 6012
rect 30499 5956 30555 6012
rect 30555 5956 30559 6012
rect 30495 5952 30559 5956
rect 30575 6012 30639 6016
rect 30575 5956 30579 6012
rect 30579 5956 30635 6012
rect 30635 5956 30639 6012
rect 30575 5952 30639 5956
rect 30655 6012 30719 6016
rect 30655 5956 30659 6012
rect 30659 5956 30715 6012
rect 30715 5956 30719 6012
rect 30655 5952 30719 5956
rect 30735 6012 30799 6016
rect 30735 5956 30739 6012
rect 30739 5956 30795 6012
rect 30795 5956 30799 6012
rect 30735 5952 30799 5956
rect 9392 5468 9456 5472
rect 9392 5412 9396 5468
rect 9396 5412 9452 5468
rect 9452 5412 9456 5468
rect 9392 5408 9456 5412
rect 9472 5468 9536 5472
rect 9472 5412 9476 5468
rect 9476 5412 9532 5468
rect 9532 5412 9536 5468
rect 9472 5408 9536 5412
rect 9552 5468 9616 5472
rect 9552 5412 9556 5468
rect 9556 5412 9612 5468
rect 9612 5412 9616 5468
rect 9552 5408 9616 5412
rect 9632 5468 9696 5472
rect 9632 5412 9636 5468
rect 9636 5412 9692 5468
rect 9692 5412 9696 5468
rect 9632 5408 9696 5412
rect 17833 5468 17897 5472
rect 17833 5412 17837 5468
rect 17837 5412 17893 5468
rect 17893 5412 17897 5468
rect 17833 5408 17897 5412
rect 17913 5468 17977 5472
rect 17913 5412 17917 5468
rect 17917 5412 17973 5468
rect 17973 5412 17977 5468
rect 17913 5408 17977 5412
rect 17993 5468 18057 5472
rect 17993 5412 17997 5468
rect 17997 5412 18053 5468
rect 18053 5412 18057 5468
rect 17993 5408 18057 5412
rect 18073 5468 18137 5472
rect 18073 5412 18077 5468
rect 18077 5412 18133 5468
rect 18133 5412 18137 5468
rect 18073 5408 18137 5412
rect 26274 5468 26338 5472
rect 26274 5412 26278 5468
rect 26278 5412 26334 5468
rect 26334 5412 26338 5468
rect 26274 5408 26338 5412
rect 26354 5468 26418 5472
rect 26354 5412 26358 5468
rect 26358 5412 26414 5468
rect 26414 5412 26418 5468
rect 26354 5408 26418 5412
rect 26434 5468 26498 5472
rect 26434 5412 26438 5468
rect 26438 5412 26494 5468
rect 26494 5412 26498 5468
rect 26434 5408 26498 5412
rect 26514 5468 26578 5472
rect 26514 5412 26518 5468
rect 26518 5412 26574 5468
rect 26574 5412 26578 5468
rect 26514 5408 26578 5412
rect 34715 5468 34779 5472
rect 34715 5412 34719 5468
rect 34719 5412 34775 5468
rect 34775 5412 34779 5468
rect 34715 5408 34779 5412
rect 34795 5468 34859 5472
rect 34795 5412 34799 5468
rect 34799 5412 34855 5468
rect 34855 5412 34859 5468
rect 34795 5408 34859 5412
rect 34875 5468 34939 5472
rect 34875 5412 34879 5468
rect 34879 5412 34935 5468
rect 34935 5412 34939 5468
rect 34875 5408 34939 5412
rect 34955 5468 35019 5472
rect 34955 5412 34959 5468
rect 34959 5412 35015 5468
rect 35015 5412 35019 5468
rect 34955 5408 35019 5412
rect 5172 4924 5236 4928
rect 5172 4868 5176 4924
rect 5176 4868 5232 4924
rect 5232 4868 5236 4924
rect 5172 4864 5236 4868
rect 5252 4924 5316 4928
rect 5252 4868 5256 4924
rect 5256 4868 5312 4924
rect 5312 4868 5316 4924
rect 5252 4864 5316 4868
rect 5332 4924 5396 4928
rect 5332 4868 5336 4924
rect 5336 4868 5392 4924
rect 5392 4868 5396 4924
rect 5332 4864 5396 4868
rect 5412 4924 5476 4928
rect 5412 4868 5416 4924
rect 5416 4868 5472 4924
rect 5472 4868 5476 4924
rect 5412 4864 5476 4868
rect 13613 4924 13677 4928
rect 13613 4868 13617 4924
rect 13617 4868 13673 4924
rect 13673 4868 13677 4924
rect 13613 4864 13677 4868
rect 13693 4924 13757 4928
rect 13693 4868 13697 4924
rect 13697 4868 13753 4924
rect 13753 4868 13757 4924
rect 13693 4864 13757 4868
rect 13773 4924 13837 4928
rect 13773 4868 13777 4924
rect 13777 4868 13833 4924
rect 13833 4868 13837 4924
rect 13773 4864 13837 4868
rect 13853 4924 13917 4928
rect 13853 4868 13857 4924
rect 13857 4868 13913 4924
rect 13913 4868 13917 4924
rect 13853 4864 13917 4868
rect 22054 4924 22118 4928
rect 22054 4868 22058 4924
rect 22058 4868 22114 4924
rect 22114 4868 22118 4924
rect 22054 4864 22118 4868
rect 22134 4924 22198 4928
rect 22134 4868 22138 4924
rect 22138 4868 22194 4924
rect 22194 4868 22198 4924
rect 22134 4864 22198 4868
rect 22214 4924 22278 4928
rect 22214 4868 22218 4924
rect 22218 4868 22274 4924
rect 22274 4868 22278 4924
rect 22214 4864 22278 4868
rect 22294 4924 22358 4928
rect 22294 4868 22298 4924
rect 22298 4868 22354 4924
rect 22354 4868 22358 4924
rect 22294 4864 22358 4868
rect 30495 4924 30559 4928
rect 30495 4868 30499 4924
rect 30499 4868 30555 4924
rect 30555 4868 30559 4924
rect 30495 4864 30559 4868
rect 30575 4924 30639 4928
rect 30575 4868 30579 4924
rect 30579 4868 30635 4924
rect 30635 4868 30639 4924
rect 30575 4864 30639 4868
rect 30655 4924 30719 4928
rect 30655 4868 30659 4924
rect 30659 4868 30715 4924
rect 30715 4868 30719 4924
rect 30655 4864 30719 4868
rect 30735 4924 30799 4928
rect 30735 4868 30739 4924
rect 30739 4868 30795 4924
rect 30795 4868 30799 4924
rect 30735 4864 30799 4868
rect 9392 4380 9456 4384
rect 9392 4324 9396 4380
rect 9396 4324 9452 4380
rect 9452 4324 9456 4380
rect 9392 4320 9456 4324
rect 9472 4380 9536 4384
rect 9472 4324 9476 4380
rect 9476 4324 9532 4380
rect 9532 4324 9536 4380
rect 9472 4320 9536 4324
rect 9552 4380 9616 4384
rect 9552 4324 9556 4380
rect 9556 4324 9612 4380
rect 9612 4324 9616 4380
rect 9552 4320 9616 4324
rect 9632 4380 9696 4384
rect 9632 4324 9636 4380
rect 9636 4324 9692 4380
rect 9692 4324 9696 4380
rect 9632 4320 9696 4324
rect 17833 4380 17897 4384
rect 17833 4324 17837 4380
rect 17837 4324 17893 4380
rect 17893 4324 17897 4380
rect 17833 4320 17897 4324
rect 17913 4380 17977 4384
rect 17913 4324 17917 4380
rect 17917 4324 17973 4380
rect 17973 4324 17977 4380
rect 17913 4320 17977 4324
rect 17993 4380 18057 4384
rect 17993 4324 17997 4380
rect 17997 4324 18053 4380
rect 18053 4324 18057 4380
rect 17993 4320 18057 4324
rect 18073 4380 18137 4384
rect 18073 4324 18077 4380
rect 18077 4324 18133 4380
rect 18133 4324 18137 4380
rect 18073 4320 18137 4324
rect 26274 4380 26338 4384
rect 26274 4324 26278 4380
rect 26278 4324 26334 4380
rect 26334 4324 26338 4380
rect 26274 4320 26338 4324
rect 26354 4380 26418 4384
rect 26354 4324 26358 4380
rect 26358 4324 26414 4380
rect 26414 4324 26418 4380
rect 26354 4320 26418 4324
rect 26434 4380 26498 4384
rect 26434 4324 26438 4380
rect 26438 4324 26494 4380
rect 26494 4324 26498 4380
rect 26434 4320 26498 4324
rect 26514 4380 26578 4384
rect 26514 4324 26518 4380
rect 26518 4324 26574 4380
rect 26574 4324 26578 4380
rect 26514 4320 26578 4324
rect 34715 4380 34779 4384
rect 34715 4324 34719 4380
rect 34719 4324 34775 4380
rect 34775 4324 34779 4380
rect 34715 4320 34779 4324
rect 34795 4380 34859 4384
rect 34795 4324 34799 4380
rect 34799 4324 34855 4380
rect 34855 4324 34859 4380
rect 34795 4320 34859 4324
rect 34875 4380 34939 4384
rect 34875 4324 34879 4380
rect 34879 4324 34935 4380
rect 34935 4324 34939 4380
rect 34875 4320 34939 4324
rect 34955 4380 35019 4384
rect 34955 4324 34959 4380
rect 34959 4324 35015 4380
rect 35015 4324 35019 4380
rect 34955 4320 35019 4324
rect 5172 3836 5236 3840
rect 5172 3780 5176 3836
rect 5176 3780 5232 3836
rect 5232 3780 5236 3836
rect 5172 3776 5236 3780
rect 5252 3836 5316 3840
rect 5252 3780 5256 3836
rect 5256 3780 5312 3836
rect 5312 3780 5316 3836
rect 5252 3776 5316 3780
rect 5332 3836 5396 3840
rect 5332 3780 5336 3836
rect 5336 3780 5392 3836
rect 5392 3780 5396 3836
rect 5332 3776 5396 3780
rect 5412 3836 5476 3840
rect 5412 3780 5416 3836
rect 5416 3780 5472 3836
rect 5472 3780 5476 3836
rect 5412 3776 5476 3780
rect 13613 3836 13677 3840
rect 13613 3780 13617 3836
rect 13617 3780 13673 3836
rect 13673 3780 13677 3836
rect 13613 3776 13677 3780
rect 13693 3836 13757 3840
rect 13693 3780 13697 3836
rect 13697 3780 13753 3836
rect 13753 3780 13757 3836
rect 13693 3776 13757 3780
rect 13773 3836 13837 3840
rect 13773 3780 13777 3836
rect 13777 3780 13833 3836
rect 13833 3780 13837 3836
rect 13773 3776 13837 3780
rect 13853 3836 13917 3840
rect 13853 3780 13857 3836
rect 13857 3780 13913 3836
rect 13913 3780 13917 3836
rect 13853 3776 13917 3780
rect 22054 3836 22118 3840
rect 22054 3780 22058 3836
rect 22058 3780 22114 3836
rect 22114 3780 22118 3836
rect 22054 3776 22118 3780
rect 22134 3836 22198 3840
rect 22134 3780 22138 3836
rect 22138 3780 22194 3836
rect 22194 3780 22198 3836
rect 22134 3776 22198 3780
rect 22214 3836 22278 3840
rect 22214 3780 22218 3836
rect 22218 3780 22274 3836
rect 22274 3780 22278 3836
rect 22214 3776 22278 3780
rect 22294 3836 22358 3840
rect 22294 3780 22298 3836
rect 22298 3780 22354 3836
rect 22354 3780 22358 3836
rect 22294 3776 22358 3780
rect 30495 3836 30559 3840
rect 30495 3780 30499 3836
rect 30499 3780 30555 3836
rect 30555 3780 30559 3836
rect 30495 3776 30559 3780
rect 30575 3836 30639 3840
rect 30575 3780 30579 3836
rect 30579 3780 30635 3836
rect 30635 3780 30639 3836
rect 30575 3776 30639 3780
rect 30655 3836 30719 3840
rect 30655 3780 30659 3836
rect 30659 3780 30715 3836
rect 30715 3780 30719 3836
rect 30655 3776 30719 3780
rect 30735 3836 30799 3840
rect 30735 3780 30739 3836
rect 30739 3780 30795 3836
rect 30795 3780 30799 3836
rect 30735 3776 30799 3780
rect 9392 3292 9456 3296
rect 9392 3236 9396 3292
rect 9396 3236 9452 3292
rect 9452 3236 9456 3292
rect 9392 3232 9456 3236
rect 9472 3292 9536 3296
rect 9472 3236 9476 3292
rect 9476 3236 9532 3292
rect 9532 3236 9536 3292
rect 9472 3232 9536 3236
rect 9552 3292 9616 3296
rect 9552 3236 9556 3292
rect 9556 3236 9612 3292
rect 9612 3236 9616 3292
rect 9552 3232 9616 3236
rect 9632 3292 9696 3296
rect 9632 3236 9636 3292
rect 9636 3236 9692 3292
rect 9692 3236 9696 3292
rect 9632 3232 9696 3236
rect 17833 3292 17897 3296
rect 17833 3236 17837 3292
rect 17837 3236 17893 3292
rect 17893 3236 17897 3292
rect 17833 3232 17897 3236
rect 17913 3292 17977 3296
rect 17913 3236 17917 3292
rect 17917 3236 17973 3292
rect 17973 3236 17977 3292
rect 17913 3232 17977 3236
rect 17993 3292 18057 3296
rect 17993 3236 17997 3292
rect 17997 3236 18053 3292
rect 18053 3236 18057 3292
rect 17993 3232 18057 3236
rect 18073 3292 18137 3296
rect 18073 3236 18077 3292
rect 18077 3236 18133 3292
rect 18133 3236 18137 3292
rect 18073 3232 18137 3236
rect 26274 3292 26338 3296
rect 26274 3236 26278 3292
rect 26278 3236 26334 3292
rect 26334 3236 26338 3292
rect 26274 3232 26338 3236
rect 26354 3292 26418 3296
rect 26354 3236 26358 3292
rect 26358 3236 26414 3292
rect 26414 3236 26418 3292
rect 26354 3232 26418 3236
rect 26434 3292 26498 3296
rect 26434 3236 26438 3292
rect 26438 3236 26494 3292
rect 26494 3236 26498 3292
rect 26434 3232 26498 3236
rect 26514 3292 26578 3296
rect 26514 3236 26518 3292
rect 26518 3236 26574 3292
rect 26574 3236 26578 3292
rect 26514 3232 26578 3236
rect 34715 3292 34779 3296
rect 34715 3236 34719 3292
rect 34719 3236 34775 3292
rect 34775 3236 34779 3292
rect 34715 3232 34779 3236
rect 34795 3292 34859 3296
rect 34795 3236 34799 3292
rect 34799 3236 34855 3292
rect 34855 3236 34859 3292
rect 34795 3232 34859 3236
rect 34875 3292 34939 3296
rect 34875 3236 34879 3292
rect 34879 3236 34935 3292
rect 34935 3236 34939 3292
rect 34875 3232 34939 3236
rect 34955 3292 35019 3296
rect 34955 3236 34959 3292
rect 34959 3236 35015 3292
rect 35015 3236 35019 3292
rect 34955 3232 35019 3236
rect 5172 2748 5236 2752
rect 5172 2692 5176 2748
rect 5176 2692 5232 2748
rect 5232 2692 5236 2748
rect 5172 2688 5236 2692
rect 5252 2748 5316 2752
rect 5252 2692 5256 2748
rect 5256 2692 5312 2748
rect 5312 2692 5316 2748
rect 5252 2688 5316 2692
rect 5332 2748 5396 2752
rect 5332 2692 5336 2748
rect 5336 2692 5392 2748
rect 5392 2692 5396 2748
rect 5332 2688 5396 2692
rect 5412 2748 5476 2752
rect 5412 2692 5416 2748
rect 5416 2692 5472 2748
rect 5472 2692 5476 2748
rect 5412 2688 5476 2692
rect 13613 2748 13677 2752
rect 13613 2692 13617 2748
rect 13617 2692 13673 2748
rect 13673 2692 13677 2748
rect 13613 2688 13677 2692
rect 13693 2748 13757 2752
rect 13693 2692 13697 2748
rect 13697 2692 13753 2748
rect 13753 2692 13757 2748
rect 13693 2688 13757 2692
rect 13773 2748 13837 2752
rect 13773 2692 13777 2748
rect 13777 2692 13833 2748
rect 13833 2692 13837 2748
rect 13773 2688 13837 2692
rect 13853 2748 13917 2752
rect 13853 2692 13857 2748
rect 13857 2692 13913 2748
rect 13913 2692 13917 2748
rect 13853 2688 13917 2692
rect 22054 2748 22118 2752
rect 22054 2692 22058 2748
rect 22058 2692 22114 2748
rect 22114 2692 22118 2748
rect 22054 2688 22118 2692
rect 22134 2748 22198 2752
rect 22134 2692 22138 2748
rect 22138 2692 22194 2748
rect 22194 2692 22198 2748
rect 22134 2688 22198 2692
rect 22214 2748 22278 2752
rect 22214 2692 22218 2748
rect 22218 2692 22274 2748
rect 22274 2692 22278 2748
rect 22214 2688 22278 2692
rect 22294 2748 22358 2752
rect 22294 2692 22298 2748
rect 22298 2692 22354 2748
rect 22354 2692 22358 2748
rect 22294 2688 22358 2692
rect 30495 2748 30559 2752
rect 30495 2692 30499 2748
rect 30499 2692 30555 2748
rect 30555 2692 30559 2748
rect 30495 2688 30559 2692
rect 30575 2748 30639 2752
rect 30575 2692 30579 2748
rect 30579 2692 30635 2748
rect 30635 2692 30639 2748
rect 30575 2688 30639 2692
rect 30655 2748 30719 2752
rect 30655 2692 30659 2748
rect 30659 2692 30715 2748
rect 30715 2692 30719 2748
rect 30655 2688 30719 2692
rect 30735 2748 30799 2752
rect 30735 2692 30739 2748
rect 30739 2692 30795 2748
rect 30795 2692 30799 2748
rect 30735 2688 30799 2692
rect 9392 2204 9456 2208
rect 9392 2148 9396 2204
rect 9396 2148 9452 2204
rect 9452 2148 9456 2204
rect 9392 2144 9456 2148
rect 9472 2204 9536 2208
rect 9472 2148 9476 2204
rect 9476 2148 9532 2204
rect 9532 2148 9536 2204
rect 9472 2144 9536 2148
rect 9552 2204 9616 2208
rect 9552 2148 9556 2204
rect 9556 2148 9612 2204
rect 9612 2148 9616 2204
rect 9552 2144 9616 2148
rect 9632 2204 9696 2208
rect 9632 2148 9636 2204
rect 9636 2148 9692 2204
rect 9692 2148 9696 2204
rect 9632 2144 9696 2148
rect 17833 2204 17897 2208
rect 17833 2148 17837 2204
rect 17837 2148 17893 2204
rect 17893 2148 17897 2204
rect 17833 2144 17897 2148
rect 17913 2204 17977 2208
rect 17913 2148 17917 2204
rect 17917 2148 17973 2204
rect 17973 2148 17977 2204
rect 17913 2144 17977 2148
rect 17993 2204 18057 2208
rect 17993 2148 17997 2204
rect 17997 2148 18053 2204
rect 18053 2148 18057 2204
rect 17993 2144 18057 2148
rect 18073 2204 18137 2208
rect 18073 2148 18077 2204
rect 18077 2148 18133 2204
rect 18133 2148 18137 2204
rect 18073 2144 18137 2148
rect 26274 2204 26338 2208
rect 26274 2148 26278 2204
rect 26278 2148 26334 2204
rect 26334 2148 26338 2204
rect 26274 2144 26338 2148
rect 26354 2204 26418 2208
rect 26354 2148 26358 2204
rect 26358 2148 26414 2204
rect 26414 2148 26418 2204
rect 26354 2144 26418 2148
rect 26434 2204 26498 2208
rect 26434 2148 26438 2204
rect 26438 2148 26494 2204
rect 26494 2148 26498 2204
rect 26434 2144 26498 2148
rect 26514 2204 26578 2208
rect 26514 2148 26518 2204
rect 26518 2148 26574 2204
rect 26574 2148 26578 2204
rect 26514 2144 26578 2148
rect 34715 2204 34779 2208
rect 34715 2148 34719 2204
rect 34719 2148 34775 2204
rect 34775 2148 34779 2204
rect 34715 2144 34779 2148
rect 34795 2204 34859 2208
rect 34795 2148 34799 2204
rect 34799 2148 34855 2204
rect 34855 2148 34859 2204
rect 34795 2144 34859 2148
rect 34875 2204 34939 2208
rect 34875 2148 34879 2204
rect 34879 2148 34935 2204
rect 34935 2148 34939 2204
rect 34875 2144 34939 2148
rect 34955 2204 35019 2208
rect 34955 2148 34959 2204
rect 34959 2148 35015 2204
rect 35015 2148 35019 2204
rect 34955 2144 35019 2148
<< metal4 >>
rect 5164 39744 5484 39760
rect 5164 39680 5172 39744
rect 5236 39680 5252 39744
rect 5316 39680 5332 39744
rect 5396 39680 5412 39744
rect 5476 39680 5484 39744
rect 5164 38656 5484 39680
rect 5164 38592 5172 38656
rect 5236 38592 5252 38656
rect 5316 38592 5332 38656
rect 5396 38592 5412 38656
rect 5476 38592 5484 38656
rect 5164 37568 5484 38592
rect 5164 37504 5172 37568
rect 5236 37504 5252 37568
rect 5316 37504 5332 37568
rect 5396 37504 5412 37568
rect 5476 37504 5484 37568
rect 5164 36480 5484 37504
rect 5164 36416 5172 36480
rect 5236 36416 5252 36480
rect 5316 36416 5332 36480
rect 5396 36416 5412 36480
rect 5476 36416 5484 36480
rect 5164 35392 5484 36416
rect 5164 35328 5172 35392
rect 5236 35328 5252 35392
rect 5316 35328 5332 35392
rect 5396 35328 5412 35392
rect 5476 35328 5484 35392
rect 5164 34304 5484 35328
rect 5164 34240 5172 34304
rect 5236 34240 5252 34304
rect 5316 34240 5332 34304
rect 5396 34240 5412 34304
rect 5476 34240 5484 34304
rect 5164 33216 5484 34240
rect 5164 33152 5172 33216
rect 5236 33152 5252 33216
rect 5316 33152 5332 33216
rect 5396 33152 5412 33216
rect 5476 33152 5484 33216
rect 5164 32128 5484 33152
rect 5164 32064 5172 32128
rect 5236 32064 5252 32128
rect 5316 32064 5332 32128
rect 5396 32064 5412 32128
rect 5476 32064 5484 32128
rect 5164 31040 5484 32064
rect 5164 30976 5172 31040
rect 5236 30976 5252 31040
rect 5316 30976 5332 31040
rect 5396 30976 5412 31040
rect 5476 30976 5484 31040
rect 5164 29952 5484 30976
rect 5164 29888 5172 29952
rect 5236 29888 5252 29952
rect 5316 29888 5332 29952
rect 5396 29888 5412 29952
rect 5476 29888 5484 29952
rect 5164 28864 5484 29888
rect 5164 28800 5172 28864
rect 5236 28800 5252 28864
rect 5316 28800 5332 28864
rect 5396 28800 5412 28864
rect 5476 28800 5484 28864
rect 5164 27776 5484 28800
rect 5164 27712 5172 27776
rect 5236 27712 5252 27776
rect 5316 27712 5332 27776
rect 5396 27712 5412 27776
rect 5476 27712 5484 27776
rect 5164 26688 5484 27712
rect 5164 26624 5172 26688
rect 5236 26624 5252 26688
rect 5316 26624 5332 26688
rect 5396 26624 5412 26688
rect 5476 26624 5484 26688
rect 5164 25600 5484 26624
rect 5164 25536 5172 25600
rect 5236 25536 5252 25600
rect 5316 25536 5332 25600
rect 5396 25536 5412 25600
rect 5476 25536 5484 25600
rect 5164 24512 5484 25536
rect 5164 24448 5172 24512
rect 5236 24448 5252 24512
rect 5316 24448 5332 24512
rect 5396 24448 5412 24512
rect 5476 24448 5484 24512
rect 5164 23424 5484 24448
rect 5164 23360 5172 23424
rect 5236 23360 5252 23424
rect 5316 23360 5332 23424
rect 5396 23360 5412 23424
rect 5476 23360 5484 23424
rect 5164 22336 5484 23360
rect 5164 22272 5172 22336
rect 5236 22272 5252 22336
rect 5316 22272 5332 22336
rect 5396 22272 5412 22336
rect 5476 22272 5484 22336
rect 5164 21248 5484 22272
rect 5164 21184 5172 21248
rect 5236 21184 5252 21248
rect 5316 21184 5332 21248
rect 5396 21184 5412 21248
rect 5476 21184 5484 21248
rect 5164 20160 5484 21184
rect 5164 20096 5172 20160
rect 5236 20096 5252 20160
rect 5316 20096 5332 20160
rect 5396 20096 5412 20160
rect 5476 20096 5484 20160
rect 5164 19072 5484 20096
rect 5164 19008 5172 19072
rect 5236 19008 5252 19072
rect 5316 19008 5332 19072
rect 5396 19008 5412 19072
rect 5476 19008 5484 19072
rect 5164 17984 5484 19008
rect 5164 17920 5172 17984
rect 5236 17920 5252 17984
rect 5316 17920 5332 17984
rect 5396 17920 5412 17984
rect 5476 17920 5484 17984
rect 5164 16896 5484 17920
rect 5164 16832 5172 16896
rect 5236 16832 5252 16896
rect 5316 16832 5332 16896
rect 5396 16832 5412 16896
rect 5476 16832 5484 16896
rect 5164 15808 5484 16832
rect 5164 15744 5172 15808
rect 5236 15744 5252 15808
rect 5316 15744 5332 15808
rect 5396 15744 5412 15808
rect 5476 15744 5484 15808
rect 5164 14720 5484 15744
rect 5164 14656 5172 14720
rect 5236 14656 5252 14720
rect 5316 14656 5332 14720
rect 5396 14656 5412 14720
rect 5476 14656 5484 14720
rect 5164 13632 5484 14656
rect 5164 13568 5172 13632
rect 5236 13568 5252 13632
rect 5316 13568 5332 13632
rect 5396 13568 5412 13632
rect 5476 13568 5484 13632
rect 5164 12544 5484 13568
rect 5164 12480 5172 12544
rect 5236 12480 5252 12544
rect 5316 12480 5332 12544
rect 5396 12480 5412 12544
rect 5476 12480 5484 12544
rect 5164 11456 5484 12480
rect 5164 11392 5172 11456
rect 5236 11392 5252 11456
rect 5316 11392 5332 11456
rect 5396 11392 5412 11456
rect 5476 11392 5484 11456
rect 5164 10368 5484 11392
rect 5164 10304 5172 10368
rect 5236 10304 5252 10368
rect 5316 10304 5332 10368
rect 5396 10304 5412 10368
rect 5476 10304 5484 10368
rect 5164 9280 5484 10304
rect 5164 9216 5172 9280
rect 5236 9216 5252 9280
rect 5316 9216 5332 9280
rect 5396 9216 5412 9280
rect 5476 9216 5484 9280
rect 5164 8192 5484 9216
rect 5164 8128 5172 8192
rect 5236 8128 5252 8192
rect 5316 8128 5332 8192
rect 5396 8128 5412 8192
rect 5476 8128 5484 8192
rect 5164 7104 5484 8128
rect 5164 7040 5172 7104
rect 5236 7040 5252 7104
rect 5316 7040 5332 7104
rect 5396 7040 5412 7104
rect 5476 7040 5484 7104
rect 5164 6016 5484 7040
rect 5164 5952 5172 6016
rect 5236 5952 5252 6016
rect 5316 5952 5332 6016
rect 5396 5952 5412 6016
rect 5476 5952 5484 6016
rect 5164 4928 5484 5952
rect 5164 4864 5172 4928
rect 5236 4864 5252 4928
rect 5316 4864 5332 4928
rect 5396 4864 5412 4928
rect 5476 4864 5484 4928
rect 5164 3840 5484 4864
rect 5164 3776 5172 3840
rect 5236 3776 5252 3840
rect 5316 3776 5332 3840
rect 5396 3776 5412 3840
rect 5476 3776 5484 3840
rect 5164 2752 5484 3776
rect 5164 2688 5172 2752
rect 5236 2688 5252 2752
rect 5316 2688 5332 2752
rect 5396 2688 5412 2752
rect 5476 2688 5484 2752
rect 5164 2128 5484 2688
rect 9384 39200 9704 39760
rect 9384 39136 9392 39200
rect 9456 39136 9472 39200
rect 9536 39136 9552 39200
rect 9616 39136 9632 39200
rect 9696 39136 9704 39200
rect 9384 38112 9704 39136
rect 9384 38048 9392 38112
rect 9456 38048 9472 38112
rect 9536 38048 9552 38112
rect 9616 38048 9632 38112
rect 9696 38048 9704 38112
rect 9384 37024 9704 38048
rect 9384 36960 9392 37024
rect 9456 36960 9472 37024
rect 9536 36960 9552 37024
rect 9616 36960 9632 37024
rect 9696 36960 9704 37024
rect 9384 35936 9704 36960
rect 9384 35872 9392 35936
rect 9456 35872 9472 35936
rect 9536 35872 9552 35936
rect 9616 35872 9632 35936
rect 9696 35872 9704 35936
rect 9384 34848 9704 35872
rect 9384 34784 9392 34848
rect 9456 34784 9472 34848
rect 9536 34784 9552 34848
rect 9616 34784 9632 34848
rect 9696 34784 9704 34848
rect 9384 33760 9704 34784
rect 9384 33696 9392 33760
rect 9456 33696 9472 33760
rect 9536 33696 9552 33760
rect 9616 33696 9632 33760
rect 9696 33696 9704 33760
rect 9384 32672 9704 33696
rect 9384 32608 9392 32672
rect 9456 32608 9472 32672
rect 9536 32608 9552 32672
rect 9616 32608 9632 32672
rect 9696 32608 9704 32672
rect 9384 31584 9704 32608
rect 9384 31520 9392 31584
rect 9456 31520 9472 31584
rect 9536 31520 9552 31584
rect 9616 31520 9632 31584
rect 9696 31520 9704 31584
rect 9384 30496 9704 31520
rect 9384 30432 9392 30496
rect 9456 30432 9472 30496
rect 9536 30432 9552 30496
rect 9616 30432 9632 30496
rect 9696 30432 9704 30496
rect 9384 29408 9704 30432
rect 9384 29344 9392 29408
rect 9456 29344 9472 29408
rect 9536 29344 9552 29408
rect 9616 29344 9632 29408
rect 9696 29344 9704 29408
rect 9384 28320 9704 29344
rect 9384 28256 9392 28320
rect 9456 28256 9472 28320
rect 9536 28256 9552 28320
rect 9616 28256 9632 28320
rect 9696 28256 9704 28320
rect 9384 27232 9704 28256
rect 9384 27168 9392 27232
rect 9456 27168 9472 27232
rect 9536 27168 9552 27232
rect 9616 27168 9632 27232
rect 9696 27168 9704 27232
rect 9384 26144 9704 27168
rect 9384 26080 9392 26144
rect 9456 26080 9472 26144
rect 9536 26080 9552 26144
rect 9616 26080 9632 26144
rect 9696 26080 9704 26144
rect 9384 25056 9704 26080
rect 9384 24992 9392 25056
rect 9456 24992 9472 25056
rect 9536 24992 9552 25056
rect 9616 24992 9632 25056
rect 9696 24992 9704 25056
rect 9384 23968 9704 24992
rect 9384 23904 9392 23968
rect 9456 23904 9472 23968
rect 9536 23904 9552 23968
rect 9616 23904 9632 23968
rect 9696 23904 9704 23968
rect 9384 22880 9704 23904
rect 9384 22816 9392 22880
rect 9456 22816 9472 22880
rect 9536 22816 9552 22880
rect 9616 22816 9632 22880
rect 9696 22816 9704 22880
rect 9384 21792 9704 22816
rect 9384 21728 9392 21792
rect 9456 21728 9472 21792
rect 9536 21728 9552 21792
rect 9616 21728 9632 21792
rect 9696 21728 9704 21792
rect 9384 20704 9704 21728
rect 9384 20640 9392 20704
rect 9456 20640 9472 20704
rect 9536 20640 9552 20704
rect 9616 20640 9632 20704
rect 9696 20640 9704 20704
rect 9384 19616 9704 20640
rect 9384 19552 9392 19616
rect 9456 19552 9472 19616
rect 9536 19552 9552 19616
rect 9616 19552 9632 19616
rect 9696 19552 9704 19616
rect 9384 18528 9704 19552
rect 9384 18464 9392 18528
rect 9456 18464 9472 18528
rect 9536 18464 9552 18528
rect 9616 18464 9632 18528
rect 9696 18464 9704 18528
rect 9384 17440 9704 18464
rect 9384 17376 9392 17440
rect 9456 17376 9472 17440
rect 9536 17376 9552 17440
rect 9616 17376 9632 17440
rect 9696 17376 9704 17440
rect 9384 16352 9704 17376
rect 9384 16288 9392 16352
rect 9456 16288 9472 16352
rect 9536 16288 9552 16352
rect 9616 16288 9632 16352
rect 9696 16288 9704 16352
rect 9384 15264 9704 16288
rect 9384 15200 9392 15264
rect 9456 15200 9472 15264
rect 9536 15200 9552 15264
rect 9616 15200 9632 15264
rect 9696 15200 9704 15264
rect 9384 14176 9704 15200
rect 9384 14112 9392 14176
rect 9456 14112 9472 14176
rect 9536 14112 9552 14176
rect 9616 14112 9632 14176
rect 9696 14112 9704 14176
rect 9384 13088 9704 14112
rect 9384 13024 9392 13088
rect 9456 13024 9472 13088
rect 9536 13024 9552 13088
rect 9616 13024 9632 13088
rect 9696 13024 9704 13088
rect 9384 12000 9704 13024
rect 9384 11936 9392 12000
rect 9456 11936 9472 12000
rect 9536 11936 9552 12000
rect 9616 11936 9632 12000
rect 9696 11936 9704 12000
rect 9384 10912 9704 11936
rect 9384 10848 9392 10912
rect 9456 10848 9472 10912
rect 9536 10848 9552 10912
rect 9616 10848 9632 10912
rect 9696 10848 9704 10912
rect 9384 9824 9704 10848
rect 9384 9760 9392 9824
rect 9456 9760 9472 9824
rect 9536 9760 9552 9824
rect 9616 9760 9632 9824
rect 9696 9760 9704 9824
rect 9384 8736 9704 9760
rect 9384 8672 9392 8736
rect 9456 8672 9472 8736
rect 9536 8672 9552 8736
rect 9616 8672 9632 8736
rect 9696 8672 9704 8736
rect 9384 7648 9704 8672
rect 9384 7584 9392 7648
rect 9456 7584 9472 7648
rect 9536 7584 9552 7648
rect 9616 7584 9632 7648
rect 9696 7584 9704 7648
rect 9384 6560 9704 7584
rect 9384 6496 9392 6560
rect 9456 6496 9472 6560
rect 9536 6496 9552 6560
rect 9616 6496 9632 6560
rect 9696 6496 9704 6560
rect 9384 5472 9704 6496
rect 9384 5408 9392 5472
rect 9456 5408 9472 5472
rect 9536 5408 9552 5472
rect 9616 5408 9632 5472
rect 9696 5408 9704 5472
rect 9384 4384 9704 5408
rect 9384 4320 9392 4384
rect 9456 4320 9472 4384
rect 9536 4320 9552 4384
rect 9616 4320 9632 4384
rect 9696 4320 9704 4384
rect 9384 3296 9704 4320
rect 9384 3232 9392 3296
rect 9456 3232 9472 3296
rect 9536 3232 9552 3296
rect 9616 3232 9632 3296
rect 9696 3232 9704 3296
rect 9384 2208 9704 3232
rect 9384 2144 9392 2208
rect 9456 2144 9472 2208
rect 9536 2144 9552 2208
rect 9616 2144 9632 2208
rect 9696 2144 9704 2208
rect 9384 2128 9704 2144
rect 13605 39744 13925 39760
rect 13605 39680 13613 39744
rect 13677 39680 13693 39744
rect 13757 39680 13773 39744
rect 13837 39680 13853 39744
rect 13917 39680 13925 39744
rect 13605 38656 13925 39680
rect 13605 38592 13613 38656
rect 13677 38592 13693 38656
rect 13757 38592 13773 38656
rect 13837 38592 13853 38656
rect 13917 38592 13925 38656
rect 13605 37568 13925 38592
rect 13605 37504 13613 37568
rect 13677 37504 13693 37568
rect 13757 37504 13773 37568
rect 13837 37504 13853 37568
rect 13917 37504 13925 37568
rect 13605 36480 13925 37504
rect 13605 36416 13613 36480
rect 13677 36416 13693 36480
rect 13757 36416 13773 36480
rect 13837 36416 13853 36480
rect 13917 36416 13925 36480
rect 13605 35392 13925 36416
rect 13605 35328 13613 35392
rect 13677 35328 13693 35392
rect 13757 35328 13773 35392
rect 13837 35328 13853 35392
rect 13917 35328 13925 35392
rect 13605 34304 13925 35328
rect 13605 34240 13613 34304
rect 13677 34240 13693 34304
rect 13757 34240 13773 34304
rect 13837 34240 13853 34304
rect 13917 34240 13925 34304
rect 13605 33216 13925 34240
rect 13605 33152 13613 33216
rect 13677 33152 13693 33216
rect 13757 33152 13773 33216
rect 13837 33152 13853 33216
rect 13917 33152 13925 33216
rect 13605 32128 13925 33152
rect 13605 32064 13613 32128
rect 13677 32064 13693 32128
rect 13757 32064 13773 32128
rect 13837 32064 13853 32128
rect 13917 32064 13925 32128
rect 13605 31040 13925 32064
rect 13605 30976 13613 31040
rect 13677 30976 13693 31040
rect 13757 30976 13773 31040
rect 13837 30976 13853 31040
rect 13917 30976 13925 31040
rect 13605 29952 13925 30976
rect 13605 29888 13613 29952
rect 13677 29888 13693 29952
rect 13757 29888 13773 29952
rect 13837 29888 13853 29952
rect 13917 29888 13925 29952
rect 13605 28864 13925 29888
rect 13605 28800 13613 28864
rect 13677 28800 13693 28864
rect 13757 28800 13773 28864
rect 13837 28800 13853 28864
rect 13917 28800 13925 28864
rect 13605 27776 13925 28800
rect 13605 27712 13613 27776
rect 13677 27712 13693 27776
rect 13757 27712 13773 27776
rect 13837 27712 13853 27776
rect 13917 27712 13925 27776
rect 13605 26688 13925 27712
rect 13605 26624 13613 26688
rect 13677 26624 13693 26688
rect 13757 26624 13773 26688
rect 13837 26624 13853 26688
rect 13917 26624 13925 26688
rect 13605 25600 13925 26624
rect 13605 25536 13613 25600
rect 13677 25536 13693 25600
rect 13757 25536 13773 25600
rect 13837 25536 13853 25600
rect 13917 25536 13925 25600
rect 13605 24512 13925 25536
rect 13605 24448 13613 24512
rect 13677 24448 13693 24512
rect 13757 24448 13773 24512
rect 13837 24448 13853 24512
rect 13917 24448 13925 24512
rect 13605 23424 13925 24448
rect 13605 23360 13613 23424
rect 13677 23360 13693 23424
rect 13757 23360 13773 23424
rect 13837 23360 13853 23424
rect 13917 23360 13925 23424
rect 13605 22336 13925 23360
rect 13605 22272 13613 22336
rect 13677 22272 13693 22336
rect 13757 22272 13773 22336
rect 13837 22272 13853 22336
rect 13917 22272 13925 22336
rect 13605 21248 13925 22272
rect 13605 21184 13613 21248
rect 13677 21184 13693 21248
rect 13757 21184 13773 21248
rect 13837 21184 13853 21248
rect 13917 21184 13925 21248
rect 13605 20160 13925 21184
rect 13605 20096 13613 20160
rect 13677 20096 13693 20160
rect 13757 20096 13773 20160
rect 13837 20096 13853 20160
rect 13917 20096 13925 20160
rect 13605 19072 13925 20096
rect 13605 19008 13613 19072
rect 13677 19008 13693 19072
rect 13757 19008 13773 19072
rect 13837 19008 13853 19072
rect 13917 19008 13925 19072
rect 13605 17984 13925 19008
rect 13605 17920 13613 17984
rect 13677 17920 13693 17984
rect 13757 17920 13773 17984
rect 13837 17920 13853 17984
rect 13917 17920 13925 17984
rect 13605 16896 13925 17920
rect 13605 16832 13613 16896
rect 13677 16832 13693 16896
rect 13757 16832 13773 16896
rect 13837 16832 13853 16896
rect 13917 16832 13925 16896
rect 13605 15808 13925 16832
rect 13605 15744 13613 15808
rect 13677 15744 13693 15808
rect 13757 15744 13773 15808
rect 13837 15744 13853 15808
rect 13917 15744 13925 15808
rect 13605 14720 13925 15744
rect 13605 14656 13613 14720
rect 13677 14656 13693 14720
rect 13757 14656 13773 14720
rect 13837 14656 13853 14720
rect 13917 14656 13925 14720
rect 13605 13632 13925 14656
rect 13605 13568 13613 13632
rect 13677 13568 13693 13632
rect 13757 13568 13773 13632
rect 13837 13568 13853 13632
rect 13917 13568 13925 13632
rect 13605 12544 13925 13568
rect 13605 12480 13613 12544
rect 13677 12480 13693 12544
rect 13757 12480 13773 12544
rect 13837 12480 13853 12544
rect 13917 12480 13925 12544
rect 13605 11456 13925 12480
rect 13605 11392 13613 11456
rect 13677 11392 13693 11456
rect 13757 11392 13773 11456
rect 13837 11392 13853 11456
rect 13917 11392 13925 11456
rect 13605 10368 13925 11392
rect 13605 10304 13613 10368
rect 13677 10304 13693 10368
rect 13757 10304 13773 10368
rect 13837 10304 13853 10368
rect 13917 10304 13925 10368
rect 13605 9280 13925 10304
rect 13605 9216 13613 9280
rect 13677 9216 13693 9280
rect 13757 9216 13773 9280
rect 13837 9216 13853 9280
rect 13917 9216 13925 9280
rect 13605 8192 13925 9216
rect 13605 8128 13613 8192
rect 13677 8128 13693 8192
rect 13757 8128 13773 8192
rect 13837 8128 13853 8192
rect 13917 8128 13925 8192
rect 13605 7104 13925 8128
rect 13605 7040 13613 7104
rect 13677 7040 13693 7104
rect 13757 7040 13773 7104
rect 13837 7040 13853 7104
rect 13917 7040 13925 7104
rect 13605 6016 13925 7040
rect 13605 5952 13613 6016
rect 13677 5952 13693 6016
rect 13757 5952 13773 6016
rect 13837 5952 13853 6016
rect 13917 5952 13925 6016
rect 13605 4928 13925 5952
rect 13605 4864 13613 4928
rect 13677 4864 13693 4928
rect 13757 4864 13773 4928
rect 13837 4864 13853 4928
rect 13917 4864 13925 4928
rect 13605 3840 13925 4864
rect 13605 3776 13613 3840
rect 13677 3776 13693 3840
rect 13757 3776 13773 3840
rect 13837 3776 13853 3840
rect 13917 3776 13925 3840
rect 13605 2752 13925 3776
rect 13605 2688 13613 2752
rect 13677 2688 13693 2752
rect 13757 2688 13773 2752
rect 13837 2688 13853 2752
rect 13917 2688 13925 2752
rect 13605 2128 13925 2688
rect 17825 39200 18145 39760
rect 17825 39136 17833 39200
rect 17897 39136 17913 39200
rect 17977 39136 17993 39200
rect 18057 39136 18073 39200
rect 18137 39136 18145 39200
rect 17825 38112 18145 39136
rect 17825 38048 17833 38112
rect 17897 38048 17913 38112
rect 17977 38048 17993 38112
rect 18057 38048 18073 38112
rect 18137 38048 18145 38112
rect 17825 37024 18145 38048
rect 17825 36960 17833 37024
rect 17897 36960 17913 37024
rect 17977 36960 17993 37024
rect 18057 36960 18073 37024
rect 18137 36960 18145 37024
rect 17825 35936 18145 36960
rect 17825 35872 17833 35936
rect 17897 35872 17913 35936
rect 17977 35872 17993 35936
rect 18057 35872 18073 35936
rect 18137 35872 18145 35936
rect 17825 34848 18145 35872
rect 17825 34784 17833 34848
rect 17897 34784 17913 34848
rect 17977 34784 17993 34848
rect 18057 34784 18073 34848
rect 18137 34784 18145 34848
rect 17825 33760 18145 34784
rect 17825 33696 17833 33760
rect 17897 33696 17913 33760
rect 17977 33696 17993 33760
rect 18057 33696 18073 33760
rect 18137 33696 18145 33760
rect 17825 32672 18145 33696
rect 17825 32608 17833 32672
rect 17897 32608 17913 32672
rect 17977 32608 17993 32672
rect 18057 32608 18073 32672
rect 18137 32608 18145 32672
rect 17825 31584 18145 32608
rect 17825 31520 17833 31584
rect 17897 31520 17913 31584
rect 17977 31520 17993 31584
rect 18057 31520 18073 31584
rect 18137 31520 18145 31584
rect 17825 30496 18145 31520
rect 17825 30432 17833 30496
rect 17897 30432 17913 30496
rect 17977 30432 17993 30496
rect 18057 30432 18073 30496
rect 18137 30432 18145 30496
rect 17825 29408 18145 30432
rect 17825 29344 17833 29408
rect 17897 29344 17913 29408
rect 17977 29344 17993 29408
rect 18057 29344 18073 29408
rect 18137 29344 18145 29408
rect 17825 28320 18145 29344
rect 17825 28256 17833 28320
rect 17897 28256 17913 28320
rect 17977 28256 17993 28320
rect 18057 28256 18073 28320
rect 18137 28256 18145 28320
rect 17825 27232 18145 28256
rect 17825 27168 17833 27232
rect 17897 27168 17913 27232
rect 17977 27168 17993 27232
rect 18057 27168 18073 27232
rect 18137 27168 18145 27232
rect 17825 26144 18145 27168
rect 17825 26080 17833 26144
rect 17897 26080 17913 26144
rect 17977 26080 17993 26144
rect 18057 26080 18073 26144
rect 18137 26080 18145 26144
rect 17825 25056 18145 26080
rect 17825 24992 17833 25056
rect 17897 24992 17913 25056
rect 17977 24992 17993 25056
rect 18057 24992 18073 25056
rect 18137 24992 18145 25056
rect 17825 23968 18145 24992
rect 17825 23904 17833 23968
rect 17897 23904 17913 23968
rect 17977 23904 17993 23968
rect 18057 23904 18073 23968
rect 18137 23904 18145 23968
rect 17825 22880 18145 23904
rect 17825 22816 17833 22880
rect 17897 22816 17913 22880
rect 17977 22816 17993 22880
rect 18057 22816 18073 22880
rect 18137 22816 18145 22880
rect 17825 21792 18145 22816
rect 17825 21728 17833 21792
rect 17897 21728 17913 21792
rect 17977 21728 17993 21792
rect 18057 21728 18073 21792
rect 18137 21728 18145 21792
rect 17825 20704 18145 21728
rect 17825 20640 17833 20704
rect 17897 20640 17913 20704
rect 17977 20640 17993 20704
rect 18057 20640 18073 20704
rect 18137 20640 18145 20704
rect 17825 19616 18145 20640
rect 17825 19552 17833 19616
rect 17897 19552 17913 19616
rect 17977 19552 17993 19616
rect 18057 19552 18073 19616
rect 18137 19552 18145 19616
rect 17825 18528 18145 19552
rect 17825 18464 17833 18528
rect 17897 18464 17913 18528
rect 17977 18464 17993 18528
rect 18057 18464 18073 18528
rect 18137 18464 18145 18528
rect 17825 17440 18145 18464
rect 17825 17376 17833 17440
rect 17897 17376 17913 17440
rect 17977 17376 17993 17440
rect 18057 17376 18073 17440
rect 18137 17376 18145 17440
rect 17825 16352 18145 17376
rect 17825 16288 17833 16352
rect 17897 16288 17913 16352
rect 17977 16288 17993 16352
rect 18057 16288 18073 16352
rect 18137 16288 18145 16352
rect 17825 15264 18145 16288
rect 17825 15200 17833 15264
rect 17897 15200 17913 15264
rect 17977 15200 17993 15264
rect 18057 15200 18073 15264
rect 18137 15200 18145 15264
rect 17825 14176 18145 15200
rect 17825 14112 17833 14176
rect 17897 14112 17913 14176
rect 17977 14112 17993 14176
rect 18057 14112 18073 14176
rect 18137 14112 18145 14176
rect 17825 13088 18145 14112
rect 17825 13024 17833 13088
rect 17897 13024 17913 13088
rect 17977 13024 17993 13088
rect 18057 13024 18073 13088
rect 18137 13024 18145 13088
rect 17825 12000 18145 13024
rect 17825 11936 17833 12000
rect 17897 11936 17913 12000
rect 17977 11936 17993 12000
rect 18057 11936 18073 12000
rect 18137 11936 18145 12000
rect 17825 10912 18145 11936
rect 17825 10848 17833 10912
rect 17897 10848 17913 10912
rect 17977 10848 17993 10912
rect 18057 10848 18073 10912
rect 18137 10848 18145 10912
rect 17825 9824 18145 10848
rect 17825 9760 17833 9824
rect 17897 9760 17913 9824
rect 17977 9760 17993 9824
rect 18057 9760 18073 9824
rect 18137 9760 18145 9824
rect 17825 8736 18145 9760
rect 17825 8672 17833 8736
rect 17897 8672 17913 8736
rect 17977 8672 17993 8736
rect 18057 8672 18073 8736
rect 18137 8672 18145 8736
rect 17825 7648 18145 8672
rect 17825 7584 17833 7648
rect 17897 7584 17913 7648
rect 17977 7584 17993 7648
rect 18057 7584 18073 7648
rect 18137 7584 18145 7648
rect 17825 6560 18145 7584
rect 17825 6496 17833 6560
rect 17897 6496 17913 6560
rect 17977 6496 17993 6560
rect 18057 6496 18073 6560
rect 18137 6496 18145 6560
rect 17825 5472 18145 6496
rect 17825 5408 17833 5472
rect 17897 5408 17913 5472
rect 17977 5408 17993 5472
rect 18057 5408 18073 5472
rect 18137 5408 18145 5472
rect 17825 4384 18145 5408
rect 17825 4320 17833 4384
rect 17897 4320 17913 4384
rect 17977 4320 17993 4384
rect 18057 4320 18073 4384
rect 18137 4320 18145 4384
rect 17825 3296 18145 4320
rect 17825 3232 17833 3296
rect 17897 3232 17913 3296
rect 17977 3232 17993 3296
rect 18057 3232 18073 3296
rect 18137 3232 18145 3296
rect 17825 2208 18145 3232
rect 17825 2144 17833 2208
rect 17897 2144 17913 2208
rect 17977 2144 17993 2208
rect 18057 2144 18073 2208
rect 18137 2144 18145 2208
rect 17825 2128 18145 2144
rect 22046 39744 22366 39760
rect 22046 39680 22054 39744
rect 22118 39680 22134 39744
rect 22198 39680 22214 39744
rect 22278 39680 22294 39744
rect 22358 39680 22366 39744
rect 22046 38656 22366 39680
rect 22046 38592 22054 38656
rect 22118 38592 22134 38656
rect 22198 38592 22214 38656
rect 22278 38592 22294 38656
rect 22358 38592 22366 38656
rect 22046 37568 22366 38592
rect 22046 37504 22054 37568
rect 22118 37504 22134 37568
rect 22198 37504 22214 37568
rect 22278 37504 22294 37568
rect 22358 37504 22366 37568
rect 22046 36480 22366 37504
rect 26266 39200 26586 39760
rect 26266 39136 26274 39200
rect 26338 39136 26354 39200
rect 26418 39136 26434 39200
rect 26498 39136 26514 39200
rect 26578 39136 26586 39200
rect 26266 38112 26586 39136
rect 26266 38048 26274 38112
rect 26338 38048 26354 38112
rect 26418 38048 26434 38112
rect 26498 38048 26514 38112
rect 26578 38048 26586 38112
rect 24715 37092 24781 37093
rect 24715 37028 24716 37092
rect 24780 37028 24781 37092
rect 24715 37027 24781 37028
rect 22046 36416 22054 36480
rect 22118 36416 22134 36480
rect 22198 36416 22214 36480
rect 22278 36416 22294 36480
rect 22358 36416 22366 36480
rect 22046 35392 22366 36416
rect 22046 35328 22054 35392
rect 22118 35328 22134 35392
rect 22198 35328 22214 35392
rect 22278 35328 22294 35392
rect 22358 35328 22366 35392
rect 22046 34304 22366 35328
rect 23427 34644 23493 34645
rect 23427 34580 23428 34644
rect 23492 34580 23493 34644
rect 23427 34579 23493 34580
rect 22046 34240 22054 34304
rect 22118 34240 22134 34304
rect 22198 34240 22214 34304
rect 22278 34240 22294 34304
rect 22358 34240 22366 34304
rect 22046 33216 22366 34240
rect 22046 33152 22054 33216
rect 22118 33152 22134 33216
rect 22198 33152 22214 33216
rect 22278 33152 22294 33216
rect 22358 33152 22366 33216
rect 22046 32128 22366 33152
rect 22046 32064 22054 32128
rect 22118 32064 22134 32128
rect 22198 32064 22214 32128
rect 22278 32064 22294 32128
rect 22358 32064 22366 32128
rect 22046 31040 22366 32064
rect 22046 30976 22054 31040
rect 22118 30976 22134 31040
rect 22198 30976 22214 31040
rect 22278 30976 22294 31040
rect 22358 30976 22366 31040
rect 22046 29952 22366 30976
rect 22046 29888 22054 29952
rect 22118 29888 22134 29952
rect 22198 29888 22214 29952
rect 22278 29888 22294 29952
rect 22358 29888 22366 29952
rect 22046 28864 22366 29888
rect 22046 28800 22054 28864
rect 22118 28800 22134 28864
rect 22198 28800 22214 28864
rect 22278 28800 22294 28864
rect 22358 28800 22366 28864
rect 22046 27776 22366 28800
rect 23430 28661 23490 34579
rect 23427 28660 23493 28661
rect 23427 28596 23428 28660
rect 23492 28596 23493 28660
rect 23427 28595 23493 28596
rect 22046 27712 22054 27776
rect 22118 27712 22134 27776
rect 22198 27712 22214 27776
rect 22278 27712 22294 27776
rect 22358 27712 22366 27776
rect 22046 26688 22366 27712
rect 22046 26624 22054 26688
rect 22118 26624 22134 26688
rect 22198 26624 22214 26688
rect 22278 26624 22294 26688
rect 22358 26624 22366 26688
rect 22046 25600 22366 26624
rect 22046 25536 22054 25600
rect 22118 25536 22134 25600
rect 22198 25536 22214 25600
rect 22278 25536 22294 25600
rect 22358 25536 22366 25600
rect 22046 24512 22366 25536
rect 22046 24448 22054 24512
rect 22118 24448 22134 24512
rect 22198 24448 22214 24512
rect 22278 24448 22294 24512
rect 22358 24448 22366 24512
rect 22046 23424 22366 24448
rect 22046 23360 22054 23424
rect 22118 23360 22134 23424
rect 22198 23360 22214 23424
rect 22278 23360 22294 23424
rect 22358 23360 22366 23424
rect 22046 22336 22366 23360
rect 22046 22272 22054 22336
rect 22118 22272 22134 22336
rect 22198 22272 22214 22336
rect 22278 22272 22294 22336
rect 22358 22272 22366 22336
rect 22046 21248 22366 22272
rect 22046 21184 22054 21248
rect 22118 21184 22134 21248
rect 22198 21184 22214 21248
rect 22278 21184 22294 21248
rect 22358 21184 22366 21248
rect 22046 20160 22366 21184
rect 22046 20096 22054 20160
rect 22118 20096 22134 20160
rect 22198 20096 22214 20160
rect 22278 20096 22294 20160
rect 22358 20096 22366 20160
rect 22046 19072 22366 20096
rect 22046 19008 22054 19072
rect 22118 19008 22134 19072
rect 22198 19008 22214 19072
rect 22278 19008 22294 19072
rect 22358 19008 22366 19072
rect 22046 17984 22366 19008
rect 24531 18596 24597 18597
rect 24531 18532 24532 18596
rect 24596 18532 24597 18596
rect 24531 18531 24597 18532
rect 22046 17920 22054 17984
rect 22118 17920 22134 17984
rect 22198 17920 22214 17984
rect 22278 17920 22294 17984
rect 22358 17920 22366 17984
rect 22046 16896 22366 17920
rect 22046 16832 22054 16896
rect 22118 16832 22134 16896
rect 22198 16832 22214 16896
rect 22278 16832 22294 16896
rect 22358 16832 22366 16896
rect 22046 15808 22366 16832
rect 24534 16557 24594 18531
rect 24531 16556 24597 16557
rect 24531 16492 24532 16556
rect 24596 16492 24597 16556
rect 24531 16491 24597 16492
rect 22046 15744 22054 15808
rect 22118 15744 22134 15808
rect 22198 15744 22214 15808
rect 22278 15744 22294 15808
rect 22358 15744 22366 15808
rect 22046 14720 22366 15744
rect 24718 15061 24778 37027
rect 26266 37024 26586 38048
rect 30487 39744 30807 39760
rect 30487 39680 30495 39744
rect 30559 39680 30575 39744
rect 30639 39680 30655 39744
rect 30719 39680 30735 39744
rect 30799 39680 30807 39744
rect 30487 38656 30807 39680
rect 30971 39404 31037 39405
rect 30971 39340 30972 39404
rect 31036 39340 31037 39404
rect 30971 39339 31037 39340
rect 30487 38592 30495 38656
rect 30559 38592 30575 38656
rect 30639 38592 30655 38656
rect 30719 38592 30735 38656
rect 30799 38592 30807 38656
rect 28763 37636 28829 37637
rect 28763 37572 28764 37636
rect 28828 37572 28829 37636
rect 28763 37571 28829 37572
rect 26266 36960 26274 37024
rect 26338 36960 26354 37024
rect 26418 36960 26434 37024
rect 26498 36960 26514 37024
rect 26578 36960 26586 37024
rect 26266 35936 26586 36960
rect 27659 36004 27725 36005
rect 27659 35940 27660 36004
rect 27724 35940 27725 36004
rect 27659 35939 27725 35940
rect 26266 35872 26274 35936
rect 26338 35872 26354 35936
rect 26418 35872 26434 35936
rect 26498 35872 26514 35936
rect 26578 35872 26586 35936
rect 26266 34848 26586 35872
rect 26266 34784 26274 34848
rect 26338 34784 26354 34848
rect 26418 34784 26434 34848
rect 26498 34784 26514 34848
rect 26578 34784 26586 34848
rect 26266 33760 26586 34784
rect 26266 33696 26274 33760
rect 26338 33696 26354 33760
rect 26418 33696 26434 33760
rect 26498 33696 26514 33760
rect 26578 33696 26586 33760
rect 26266 32672 26586 33696
rect 26266 32608 26274 32672
rect 26338 32608 26354 32672
rect 26418 32608 26434 32672
rect 26498 32608 26514 32672
rect 26578 32608 26586 32672
rect 26266 31584 26586 32608
rect 26266 31520 26274 31584
rect 26338 31520 26354 31584
rect 26418 31520 26434 31584
rect 26498 31520 26514 31584
rect 26578 31520 26586 31584
rect 26266 30496 26586 31520
rect 26266 30432 26274 30496
rect 26338 30432 26354 30496
rect 26418 30432 26434 30496
rect 26498 30432 26514 30496
rect 26578 30432 26586 30496
rect 26266 29408 26586 30432
rect 27662 29885 27722 35939
rect 28766 33557 28826 37571
rect 30487 37568 30807 38592
rect 30487 37504 30495 37568
rect 30559 37504 30575 37568
rect 30639 37504 30655 37568
rect 30719 37504 30735 37568
rect 30799 37504 30807 37568
rect 28947 37500 29013 37501
rect 28947 37436 28948 37500
rect 29012 37436 29013 37500
rect 28947 37435 29013 37436
rect 29315 37500 29381 37501
rect 29315 37436 29316 37500
rect 29380 37436 29381 37500
rect 29315 37435 29381 37436
rect 28950 35189 29010 37435
rect 29131 36548 29197 36549
rect 29131 36484 29132 36548
rect 29196 36484 29197 36548
rect 29131 36483 29197 36484
rect 29134 35869 29194 36483
rect 29131 35868 29197 35869
rect 29131 35804 29132 35868
rect 29196 35804 29197 35868
rect 29131 35803 29197 35804
rect 28947 35188 29013 35189
rect 28947 35124 28948 35188
rect 29012 35124 29013 35188
rect 28947 35123 29013 35124
rect 28763 33556 28829 33557
rect 28763 33492 28764 33556
rect 28828 33492 28829 33556
rect 28763 33491 28829 33492
rect 27659 29884 27725 29885
rect 27659 29820 27660 29884
rect 27724 29820 27725 29884
rect 27659 29819 27725 29820
rect 26266 29344 26274 29408
rect 26338 29344 26354 29408
rect 26418 29344 26434 29408
rect 26498 29344 26514 29408
rect 26578 29344 26586 29408
rect 26266 28320 26586 29344
rect 29318 29010 29378 37435
rect 29499 36548 29565 36549
rect 29499 36484 29500 36548
rect 29564 36484 29565 36548
rect 29499 36483 29565 36484
rect 29502 31109 29562 36483
rect 30487 36480 30807 37504
rect 30974 37093 31034 39339
rect 34707 39200 35027 39760
rect 34707 39136 34715 39200
rect 34779 39136 34795 39200
rect 34859 39136 34875 39200
rect 34939 39136 34955 39200
rect 35019 39136 35027 39200
rect 34707 38112 35027 39136
rect 34707 38048 34715 38112
rect 34779 38048 34795 38112
rect 34859 38048 34875 38112
rect 34939 38048 34955 38112
rect 35019 38048 35027 38112
rect 31523 37228 31589 37229
rect 31523 37164 31524 37228
rect 31588 37164 31589 37228
rect 31523 37163 31589 37164
rect 30971 37092 31037 37093
rect 30971 37028 30972 37092
rect 31036 37028 31037 37092
rect 30971 37027 31037 37028
rect 30487 36416 30495 36480
rect 30559 36416 30575 36480
rect 30639 36416 30655 36480
rect 30719 36416 30735 36480
rect 30799 36416 30807 36480
rect 30235 36412 30301 36413
rect 30235 36348 30236 36412
rect 30300 36348 30301 36412
rect 30235 36347 30301 36348
rect 29499 31108 29565 31109
rect 29499 31044 29500 31108
rect 29564 31044 29565 31108
rect 29499 31043 29565 31044
rect 30238 29613 30298 36347
rect 30487 35392 30807 36416
rect 31155 36412 31221 36413
rect 31155 36348 31156 36412
rect 31220 36348 31221 36412
rect 31155 36347 31221 36348
rect 30487 35328 30495 35392
rect 30559 35328 30575 35392
rect 30639 35328 30655 35392
rect 30719 35328 30735 35392
rect 30799 35328 30807 35392
rect 30487 34304 30807 35328
rect 30487 34240 30495 34304
rect 30559 34240 30575 34304
rect 30639 34240 30655 34304
rect 30719 34240 30735 34304
rect 30799 34240 30807 34304
rect 30487 33216 30807 34240
rect 30487 33152 30495 33216
rect 30559 33152 30575 33216
rect 30639 33152 30655 33216
rect 30719 33152 30735 33216
rect 30799 33152 30807 33216
rect 30487 32128 30807 33152
rect 31158 32605 31218 36347
rect 31526 33693 31586 37163
rect 34707 37024 35027 38048
rect 34707 36960 34715 37024
rect 34779 36960 34795 37024
rect 34859 36960 34875 37024
rect 34939 36960 34955 37024
rect 35019 36960 35027 37024
rect 34707 35936 35027 36960
rect 34707 35872 34715 35936
rect 34779 35872 34795 35936
rect 34859 35872 34875 35936
rect 34939 35872 34955 35936
rect 35019 35872 35027 35936
rect 32259 35460 32325 35461
rect 32259 35396 32260 35460
rect 32324 35396 32325 35460
rect 32259 35395 32325 35396
rect 31523 33692 31589 33693
rect 31523 33628 31524 33692
rect 31588 33628 31589 33692
rect 31523 33627 31589 33628
rect 31155 32604 31221 32605
rect 31155 32540 31156 32604
rect 31220 32540 31221 32604
rect 31155 32539 31221 32540
rect 30487 32064 30495 32128
rect 30559 32064 30575 32128
rect 30639 32064 30655 32128
rect 30719 32064 30735 32128
rect 30799 32064 30807 32128
rect 30487 31040 30807 32064
rect 30487 30976 30495 31040
rect 30559 30976 30575 31040
rect 30639 30976 30655 31040
rect 30719 30976 30735 31040
rect 30799 30976 30807 31040
rect 30487 29952 30807 30976
rect 30487 29888 30495 29952
rect 30559 29888 30575 29952
rect 30639 29888 30655 29952
rect 30719 29888 30735 29952
rect 30799 29888 30807 29952
rect 30235 29612 30301 29613
rect 30235 29548 30236 29612
rect 30300 29548 30301 29612
rect 30235 29547 30301 29548
rect 26266 28256 26274 28320
rect 26338 28256 26354 28320
rect 26418 28256 26434 28320
rect 26498 28256 26514 28320
rect 26578 28256 26586 28320
rect 26266 27232 26586 28256
rect 29134 28950 29378 29010
rect 29134 28117 29194 28950
rect 30487 28864 30807 29888
rect 32262 29205 32322 35395
rect 34707 34848 35027 35872
rect 34707 34784 34715 34848
rect 34779 34784 34795 34848
rect 34859 34784 34875 34848
rect 34939 34784 34955 34848
rect 35019 34784 35027 34848
rect 34707 33760 35027 34784
rect 34707 33696 34715 33760
rect 34779 33696 34795 33760
rect 34859 33696 34875 33760
rect 34939 33696 34955 33760
rect 35019 33696 35027 33760
rect 34707 32672 35027 33696
rect 34707 32608 34715 32672
rect 34779 32608 34795 32672
rect 34859 32608 34875 32672
rect 34939 32608 34955 32672
rect 35019 32608 35027 32672
rect 34707 31584 35027 32608
rect 34707 31520 34715 31584
rect 34779 31520 34795 31584
rect 34859 31520 34875 31584
rect 34939 31520 34955 31584
rect 35019 31520 35027 31584
rect 34707 30496 35027 31520
rect 34707 30432 34715 30496
rect 34779 30432 34795 30496
rect 34859 30432 34875 30496
rect 34939 30432 34955 30496
rect 35019 30432 35027 30496
rect 34707 29408 35027 30432
rect 34707 29344 34715 29408
rect 34779 29344 34795 29408
rect 34859 29344 34875 29408
rect 34939 29344 34955 29408
rect 35019 29344 35027 29408
rect 32259 29204 32325 29205
rect 32259 29140 32260 29204
rect 32324 29140 32325 29204
rect 32259 29139 32325 29140
rect 30487 28800 30495 28864
rect 30559 28800 30575 28864
rect 30639 28800 30655 28864
rect 30719 28800 30735 28864
rect 30799 28800 30807 28864
rect 29131 28116 29197 28117
rect 29131 28052 29132 28116
rect 29196 28052 29197 28116
rect 29131 28051 29197 28052
rect 26266 27168 26274 27232
rect 26338 27168 26354 27232
rect 26418 27168 26434 27232
rect 26498 27168 26514 27232
rect 26578 27168 26586 27232
rect 26266 26144 26586 27168
rect 26266 26080 26274 26144
rect 26338 26080 26354 26144
rect 26418 26080 26434 26144
rect 26498 26080 26514 26144
rect 26578 26080 26586 26144
rect 26266 25056 26586 26080
rect 26266 24992 26274 25056
rect 26338 24992 26354 25056
rect 26418 24992 26434 25056
rect 26498 24992 26514 25056
rect 26578 24992 26586 25056
rect 26266 23968 26586 24992
rect 26266 23904 26274 23968
rect 26338 23904 26354 23968
rect 26418 23904 26434 23968
rect 26498 23904 26514 23968
rect 26578 23904 26586 23968
rect 26266 22880 26586 23904
rect 30487 27776 30807 28800
rect 30487 27712 30495 27776
rect 30559 27712 30575 27776
rect 30639 27712 30655 27776
rect 30719 27712 30735 27776
rect 30799 27712 30807 27776
rect 30487 26688 30807 27712
rect 34707 28320 35027 29344
rect 34707 28256 34715 28320
rect 34779 28256 34795 28320
rect 34859 28256 34875 28320
rect 34939 28256 34955 28320
rect 35019 28256 35027 28320
rect 32075 27572 32141 27573
rect 32075 27508 32076 27572
rect 32140 27508 32141 27572
rect 32075 27507 32141 27508
rect 30487 26624 30495 26688
rect 30559 26624 30575 26688
rect 30639 26624 30655 26688
rect 30719 26624 30735 26688
rect 30799 26624 30807 26688
rect 30487 25600 30807 26624
rect 30487 25536 30495 25600
rect 30559 25536 30575 25600
rect 30639 25536 30655 25600
rect 30719 25536 30735 25600
rect 30799 25536 30807 25600
rect 30487 24512 30807 25536
rect 31523 24988 31589 24989
rect 31523 24924 31524 24988
rect 31588 24924 31589 24988
rect 31523 24923 31589 24924
rect 31339 24716 31405 24717
rect 31339 24652 31340 24716
rect 31404 24652 31405 24716
rect 31339 24651 31405 24652
rect 30487 24448 30495 24512
rect 30559 24448 30575 24512
rect 30639 24448 30655 24512
rect 30719 24448 30735 24512
rect 30799 24448 30807 24512
rect 29499 23628 29565 23629
rect 29499 23564 29500 23628
rect 29564 23564 29565 23628
rect 29499 23563 29565 23564
rect 26739 23492 26805 23493
rect 26739 23428 26740 23492
rect 26804 23428 26805 23492
rect 26739 23427 26805 23428
rect 26266 22816 26274 22880
rect 26338 22816 26354 22880
rect 26418 22816 26434 22880
rect 26498 22816 26514 22880
rect 26578 22816 26586 22880
rect 26266 21792 26586 22816
rect 26266 21728 26274 21792
rect 26338 21728 26354 21792
rect 26418 21728 26434 21792
rect 26498 21728 26514 21792
rect 26578 21728 26586 21792
rect 25635 20772 25701 20773
rect 25635 20708 25636 20772
rect 25700 20708 25701 20772
rect 25635 20707 25701 20708
rect 25638 15333 25698 20707
rect 26266 20704 26586 21728
rect 26266 20640 26274 20704
rect 26338 20640 26354 20704
rect 26418 20640 26434 20704
rect 26498 20640 26514 20704
rect 26578 20640 26586 20704
rect 26266 19616 26586 20640
rect 26266 19552 26274 19616
rect 26338 19552 26354 19616
rect 26418 19552 26434 19616
rect 26498 19552 26514 19616
rect 26578 19552 26586 19616
rect 26266 18528 26586 19552
rect 26266 18464 26274 18528
rect 26338 18464 26354 18528
rect 26418 18464 26434 18528
rect 26498 18464 26514 18528
rect 26578 18464 26586 18528
rect 26266 17440 26586 18464
rect 26266 17376 26274 17440
rect 26338 17376 26354 17440
rect 26418 17376 26434 17440
rect 26498 17376 26514 17440
rect 26578 17376 26586 17440
rect 26266 16352 26586 17376
rect 26266 16288 26274 16352
rect 26338 16288 26354 16352
rect 26418 16288 26434 16352
rect 26498 16288 26514 16352
rect 26578 16288 26586 16352
rect 25635 15332 25701 15333
rect 25635 15268 25636 15332
rect 25700 15268 25701 15332
rect 25635 15267 25701 15268
rect 26266 15264 26586 16288
rect 26266 15200 26274 15264
rect 26338 15200 26354 15264
rect 26418 15200 26434 15264
rect 26498 15200 26514 15264
rect 26578 15200 26586 15264
rect 24715 15060 24781 15061
rect 24715 14996 24716 15060
rect 24780 14996 24781 15060
rect 24715 14995 24781 14996
rect 22046 14656 22054 14720
rect 22118 14656 22134 14720
rect 22198 14656 22214 14720
rect 22278 14656 22294 14720
rect 22358 14656 22366 14720
rect 22046 13632 22366 14656
rect 22046 13568 22054 13632
rect 22118 13568 22134 13632
rect 22198 13568 22214 13632
rect 22278 13568 22294 13632
rect 22358 13568 22366 13632
rect 22046 12544 22366 13568
rect 22046 12480 22054 12544
rect 22118 12480 22134 12544
rect 22198 12480 22214 12544
rect 22278 12480 22294 12544
rect 22358 12480 22366 12544
rect 22046 11456 22366 12480
rect 22046 11392 22054 11456
rect 22118 11392 22134 11456
rect 22198 11392 22214 11456
rect 22278 11392 22294 11456
rect 22358 11392 22366 11456
rect 22046 10368 22366 11392
rect 22046 10304 22054 10368
rect 22118 10304 22134 10368
rect 22198 10304 22214 10368
rect 22278 10304 22294 10368
rect 22358 10304 22366 10368
rect 22046 9280 22366 10304
rect 22046 9216 22054 9280
rect 22118 9216 22134 9280
rect 22198 9216 22214 9280
rect 22278 9216 22294 9280
rect 22358 9216 22366 9280
rect 22046 8192 22366 9216
rect 22046 8128 22054 8192
rect 22118 8128 22134 8192
rect 22198 8128 22214 8192
rect 22278 8128 22294 8192
rect 22358 8128 22366 8192
rect 22046 7104 22366 8128
rect 22046 7040 22054 7104
rect 22118 7040 22134 7104
rect 22198 7040 22214 7104
rect 22278 7040 22294 7104
rect 22358 7040 22366 7104
rect 22046 6016 22366 7040
rect 22046 5952 22054 6016
rect 22118 5952 22134 6016
rect 22198 5952 22214 6016
rect 22278 5952 22294 6016
rect 22358 5952 22366 6016
rect 22046 4928 22366 5952
rect 22046 4864 22054 4928
rect 22118 4864 22134 4928
rect 22198 4864 22214 4928
rect 22278 4864 22294 4928
rect 22358 4864 22366 4928
rect 22046 3840 22366 4864
rect 22046 3776 22054 3840
rect 22118 3776 22134 3840
rect 22198 3776 22214 3840
rect 22278 3776 22294 3840
rect 22358 3776 22366 3840
rect 22046 2752 22366 3776
rect 22046 2688 22054 2752
rect 22118 2688 22134 2752
rect 22198 2688 22214 2752
rect 22278 2688 22294 2752
rect 22358 2688 22366 2752
rect 22046 2128 22366 2688
rect 26266 14176 26586 15200
rect 26266 14112 26274 14176
rect 26338 14112 26354 14176
rect 26418 14112 26434 14176
rect 26498 14112 26514 14176
rect 26578 14112 26586 14176
rect 26266 13088 26586 14112
rect 26742 13973 26802 23427
rect 29131 21860 29197 21861
rect 29131 21796 29132 21860
rect 29196 21796 29197 21860
rect 29131 21795 29197 21796
rect 27659 18732 27725 18733
rect 27659 18668 27660 18732
rect 27724 18668 27725 18732
rect 27659 18667 27725 18668
rect 27662 15061 27722 18667
rect 27659 15060 27725 15061
rect 27659 14996 27660 15060
rect 27724 14996 27725 15060
rect 27659 14995 27725 14996
rect 26739 13972 26805 13973
rect 26739 13908 26740 13972
rect 26804 13908 26805 13972
rect 26739 13907 26805 13908
rect 29134 13429 29194 21795
rect 29502 15197 29562 23563
rect 30487 23424 30807 24448
rect 30487 23360 30495 23424
rect 30559 23360 30575 23424
rect 30639 23360 30655 23424
rect 30719 23360 30735 23424
rect 30799 23360 30807 23424
rect 30487 22336 30807 23360
rect 30487 22272 30495 22336
rect 30559 22272 30575 22336
rect 30639 22272 30655 22336
rect 30719 22272 30735 22336
rect 30799 22272 30807 22336
rect 29683 22268 29749 22269
rect 29683 22204 29684 22268
rect 29748 22204 29749 22268
rect 29683 22203 29749 22204
rect 29686 16557 29746 22203
rect 30487 21248 30807 22272
rect 30487 21184 30495 21248
rect 30559 21184 30575 21248
rect 30639 21184 30655 21248
rect 30719 21184 30735 21248
rect 30799 21184 30807 21248
rect 30487 20160 30807 21184
rect 30971 20772 31037 20773
rect 30971 20708 30972 20772
rect 31036 20708 31037 20772
rect 30971 20707 31037 20708
rect 31155 20772 31221 20773
rect 31155 20708 31156 20772
rect 31220 20708 31221 20772
rect 31155 20707 31221 20708
rect 30487 20096 30495 20160
rect 30559 20096 30575 20160
rect 30639 20096 30655 20160
rect 30719 20096 30735 20160
rect 30799 20096 30807 20160
rect 30487 19072 30807 20096
rect 30487 19008 30495 19072
rect 30559 19008 30575 19072
rect 30639 19008 30655 19072
rect 30719 19008 30735 19072
rect 30799 19008 30807 19072
rect 30487 17984 30807 19008
rect 30487 17920 30495 17984
rect 30559 17920 30575 17984
rect 30639 17920 30655 17984
rect 30719 17920 30735 17984
rect 30799 17920 30807 17984
rect 30487 16896 30807 17920
rect 30487 16832 30495 16896
rect 30559 16832 30575 16896
rect 30639 16832 30655 16896
rect 30719 16832 30735 16896
rect 30799 16832 30807 16896
rect 29683 16556 29749 16557
rect 29683 16492 29684 16556
rect 29748 16492 29749 16556
rect 29683 16491 29749 16492
rect 30487 15808 30807 16832
rect 30974 16285 31034 20707
rect 31158 16829 31218 20707
rect 31342 16829 31402 24651
rect 31155 16828 31221 16829
rect 31155 16764 31156 16828
rect 31220 16764 31221 16828
rect 31155 16763 31221 16764
rect 31339 16828 31405 16829
rect 31339 16764 31340 16828
rect 31404 16764 31405 16828
rect 31339 16763 31405 16764
rect 31526 16285 31586 24923
rect 31891 23764 31957 23765
rect 31891 23700 31892 23764
rect 31956 23700 31957 23764
rect 31891 23699 31957 23700
rect 30971 16284 31037 16285
rect 30971 16220 30972 16284
rect 31036 16220 31037 16284
rect 30971 16219 31037 16220
rect 31523 16284 31589 16285
rect 31523 16220 31524 16284
rect 31588 16220 31589 16284
rect 31523 16219 31589 16220
rect 30487 15744 30495 15808
rect 30559 15744 30575 15808
rect 30639 15744 30655 15808
rect 30719 15744 30735 15808
rect 30799 15744 30807 15808
rect 29499 15196 29565 15197
rect 29499 15132 29500 15196
rect 29564 15132 29565 15196
rect 29499 15131 29565 15132
rect 30487 14720 30807 15744
rect 30487 14656 30495 14720
rect 30559 14656 30575 14720
rect 30639 14656 30655 14720
rect 30719 14656 30735 14720
rect 30799 14656 30807 14720
rect 30487 13632 30807 14656
rect 30487 13568 30495 13632
rect 30559 13568 30575 13632
rect 30639 13568 30655 13632
rect 30719 13568 30735 13632
rect 30799 13568 30807 13632
rect 29131 13428 29197 13429
rect 29131 13364 29132 13428
rect 29196 13364 29197 13428
rect 29131 13363 29197 13364
rect 26266 13024 26274 13088
rect 26338 13024 26354 13088
rect 26418 13024 26434 13088
rect 26498 13024 26514 13088
rect 26578 13024 26586 13088
rect 26266 12000 26586 13024
rect 26266 11936 26274 12000
rect 26338 11936 26354 12000
rect 26418 11936 26434 12000
rect 26498 11936 26514 12000
rect 26578 11936 26586 12000
rect 26266 10912 26586 11936
rect 26266 10848 26274 10912
rect 26338 10848 26354 10912
rect 26418 10848 26434 10912
rect 26498 10848 26514 10912
rect 26578 10848 26586 10912
rect 26266 9824 26586 10848
rect 26266 9760 26274 9824
rect 26338 9760 26354 9824
rect 26418 9760 26434 9824
rect 26498 9760 26514 9824
rect 26578 9760 26586 9824
rect 26266 8736 26586 9760
rect 26266 8672 26274 8736
rect 26338 8672 26354 8736
rect 26418 8672 26434 8736
rect 26498 8672 26514 8736
rect 26578 8672 26586 8736
rect 26266 7648 26586 8672
rect 26266 7584 26274 7648
rect 26338 7584 26354 7648
rect 26418 7584 26434 7648
rect 26498 7584 26514 7648
rect 26578 7584 26586 7648
rect 26266 6560 26586 7584
rect 26266 6496 26274 6560
rect 26338 6496 26354 6560
rect 26418 6496 26434 6560
rect 26498 6496 26514 6560
rect 26578 6496 26586 6560
rect 26266 5472 26586 6496
rect 26266 5408 26274 5472
rect 26338 5408 26354 5472
rect 26418 5408 26434 5472
rect 26498 5408 26514 5472
rect 26578 5408 26586 5472
rect 26266 4384 26586 5408
rect 26266 4320 26274 4384
rect 26338 4320 26354 4384
rect 26418 4320 26434 4384
rect 26498 4320 26514 4384
rect 26578 4320 26586 4384
rect 26266 3296 26586 4320
rect 26266 3232 26274 3296
rect 26338 3232 26354 3296
rect 26418 3232 26434 3296
rect 26498 3232 26514 3296
rect 26578 3232 26586 3296
rect 26266 2208 26586 3232
rect 26266 2144 26274 2208
rect 26338 2144 26354 2208
rect 26418 2144 26434 2208
rect 26498 2144 26514 2208
rect 26578 2144 26586 2208
rect 26266 2128 26586 2144
rect 30487 12544 30807 13568
rect 31894 13565 31954 23699
rect 32078 16693 32138 27507
rect 34707 27232 35027 28256
rect 34707 27168 34715 27232
rect 34779 27168 34795 27232
rect 34859 27168 34875 27232
rect 34939 27168 34955 27232
rect 35019 27168 35027 27232
rect 34707 26144 35027 27168
rect 34707 26080 34715 26144
rect 34779 26080 34795 26144
rect 34859 26080 34875 26144
rect 34939 26080 34955 26144
rect 35019 26080 35027 26144
rect 34707 25056 35027 26080
rect 34707 24992 34715 25056
rect 34779 24992 34795 25056
rect 34859 24992 34875 25056
rect 34939 24992 34955 25056
rect 35019 24992 35027 25056
rect 32811 24716 32877 24717
rect 32811 24652 32812 24716
rect 32876 24652 32877 24716
rect 32811 24651 32877 24652
rect 32259 20908 32325 20909
rect 32259 20844 32260 20908
rect 32324 20844 32325 20908
rect 32259 20843 32325 20844
rect 32262 19005 32322 20843
rect 32259 19004 32325 19005
rect 32259 18940 32260 19004
rect 32324 18940 32325 19004
rect 32259 18939 32325 18940
rect 32814 18053 32874 24651
rect 34707 23968 35027 24992
rect 34707 23904 34715 23968
rect 34779 23904 34795 23968
rect 34859 23904 34875 23968
rect 34939 23904 34955 23968
rect 35019 23904 35027 23968
rect 33731 23900 33797 23901
rect 33731 23836 33732 23900
rect 33796 23836 33797 23900
rect 33731 23835 33797 23836
rect 32811 18052 32877 18053
rect 32811 17988 32812 18052
rect 32876 17988 32877 18052
rect 32811 17987 32877 17988
rect 32075 16692 32141 16693
rect 32075 16628 32076 16692
rect 32140 16628 32141 16692
rect 32075 16627 32141 16628
rect 33734 13565 33794 23835
rect 33915 23492 33981 23493
rect 33915 23428 33916 23492
rect 33980 23428 33981 23492
rect 33915 23427 33981 23428
rect 33918 15061 33978 23427
rect 34707 22880 35027 23904
rect 34707 22816 34715 22880
rect 34779 22816 34795 22880
rect 34859 22816 34875 22880
rect 34939 22816 34955 22880
rect 35019 22816 35027 22880
rect 34099 22676 34165 22677
rect 34099 22612 34100 22676
rect 34164 22612 34165 22676
rect 34099 22611 34165 22612
rect 33915 15060 33981 15061
rect 33915 14996 33916 15060
rect 33980 14996 33981 15060
rect 33915 14995 33981 14996
rect 31891 13564 31957 13565
rect 31891 13500 31892 13564
rect 31956 13500 31957 13564
rect 31891 13499 31957 13500
rect 33731 13564 33797 13565
rect 33731 13500 33732 13564
rect 33796 13500 33797 13564
rect 33731 13499 33797 13500
rect 30487 12480 30495 12544
rect 30559 12480 30575 12544
rect 30639 12480 30655 12544
rect 30719 12480 30735 12544
rect 30799 12480 30807 12544
rect 30487 11456 30807 12480
rect 34102 11797 34162 22611
rect 34707 21792 35027 22816
rect 34707 21728 34715 21792
rect 34779 21728 34795 21792
rect 34859 21728 34875 21792
rect 34939 21728 34955 21792
rect 35019 21728 35027 21792
rect 34707 20704 35027 21728
rect 34707 20640 34715 20704
rect 34779 20640 34795 20704
rect 34859 20640 34875 20704
rect 34939 20640 34955 20704
rect 35019 20640 35027 20704
rect 34707 19616 35027 20640
rect 34707 19552 34715 19616
rect 34779 19552 34795 19616
rect 34859 19552 34875 19616
rect 34939 19552 34955 19616
rect 35019 19552 35027 19616
rect 34707 18528 35027 19552
rect 34707 18464 34715 18528
rect 34779 18464 34795 18528
rect 34859 18464 34875 18528
rect 34939 18464 34955 18528
rect 35019 18464 35027 18528
rect 34707 17440 35027 18464
rect 34707 17376 34715 17440
rect 34779 17376 34795 17440
rect 34859 17376 34875 17440
rect 34939 17376 34955 17440
rect 35019 17376 35027 17440
rect 34707 16352 35027 17376
rect 34707 16288 34715 16352
rect 34779 16288 34795 16352
rect 34859 16288 34875 16352
rect 34939 16288 34955 16352
rect 35019 16288 35027 16352
rect 34707 15264 35027 16288
rect 34707 15200 34715 15264
rect 34779 15200 34795 15264
rect 34859 15200 34875 15264
rect 34939 15200 34955 15264
rect 35019 15200 35027 15264
rect 34707 14176 35027 15200
rect 34707 14112 34715 14176
rect 34779 14112 34795 14176
rect 34859 14112 34875 14176
rect 34939 14112 34955 14176
rect 35019 14112 35027 14176
rect 34707 13088 35027 14112
rect 34707 13024 34715 13088
rect 34779 13024 34795 13088
rect 34859 13024 34875 13088
rect 34939 13024 34955 13088
rect 35019 13024 35027 13088
rect 34707 12000 35027 13024
rect 34707 11936 34715 12000
rect 34779 11936 34795 12000
rect 34859 11936 34875 12000
rect 34939 11936 34955 12000
rect 35019 11936 35027 12000
rect 34099 11796 34165 11797
rect 34099 11732 34100 11796
rect 34164 11732 34165 11796
rect 34099 11731 34165 11732
rect 30487 11392 30495 11456
rect 30559 11392 30575 11456
rect 30639 11392 30655 11456
rect 30719 11392 30735 11456
rect 30799 11392 30807 11456
rect 30487 10368 30807 11392
rect 30487 10304 30495 10368
rect 30559 10304 30575 10368
rect 30639 10304 30655 10368
rect 30719 10304 30735 10368
rect 30799 10304 30807 10368
rect 30487 9280 30807 10304
rect 30487 9216 30495 9280
rect 30559 9216 30575 9280
rect 30639 9216 30655 9280
rect 30719 9216 30735 9280
rect 30799 9216 30807 9280
rect 30487 8192 30807 9216
rect 30487 8128 30495 8192
rect 30559 8128 30575 8192
rect 30639 8128 30655 8192
rect 30719 8128 30735 8192
rect 30799 8128 30807 8192
rect 30487 7104 30807 8128
rect 30487 7040 30495 7104
rect 30559 7040 30575 7104
rect 30639 7040 30655 7104
rect 30719 7040 30735 7104
rect 30799 7040 30807 7104
rect 30487 6016 30807 7040
rect 30487 5952 30495 6016
rect 30559 5952 30575 6016
rect 30639 5952 30655 6016
rect 30719 5952 30735 6016
rect 30799 5952 30807 6016
rect 30487 4928 30807 5952
rect 30487 4864 30495 4928
rect 30559 4864 30575 4928
rect 30639 4864 30655 4928
rect 30719 4864 30735 4928
rect 30799 4864 30807 4928
rect 30487 3840 30807 4864
rect 30487 3776 30495 3840
rect 30559 3776 30575 3840
rect 30639 3776 30655 3840
rect 30719 3776 30735 3840
rect 30799 3776 30807 3840
rect 30487 2752 30807 3776
rect 30487 2688 30495 2752
rect 30559 2688 30575 2752
rect 30639 2688 30655 2752
rect 30719 2688 30735 2752
rect 30799 2688 30807 2752
rect 30487 2128 30807 2688
rect 34707 10912 35027 11936
rect 34707 10848 34715 10912
rect 34779 10848 34795 10912
rect 34859 10848 34875 10912
rect 34939 10848 34955 10912
rect 35019 10848 35027 10912
rect 34707 9824 35027 10848
rect 34707 9760 34715 9824
rect 34779 9760 34795 9824
rect 34859 9760 34875 9824
rect 34939 9760 34955 9824
rect 35019 9760 35027 9824
rect 34707 8736 35027 9760
rect 34707 8672 34715 8736
rect 34779 8672 34795 8736
rect 34859 8672 34875 8736
rect 34939 8672 34955 8736
rect 35019 8672 35027 8736
rect 34707 7648 35027 8672
rect 34707 7584 34715 7648
rect 34779 7584 34795 7648
rect 34859 7584 34875 7648
rect 34939 7584 34955 7648
rect 35019 7584 35027 7648
rect 34707 6560 35027 7584
rect 34707 6496 34715 6560
rect 34779 6496 34795 6560
rect 34859 6496 34875 6560
rect 34939 6496 34955 6560
rect 35019 6496 35027 6560
rect 34707 5472 35027 6496
rect 34707 5408 34715 5472
rect 34779 5408 34795 5472
rect 34859 5408 34875 5472
rect 34939 5408 34955 5472
rect 35019 5408 35027 5472
rect 34707 4384 35027 5408
rect 34707 4320 34715 4384
rect 34779 4320 34795 4384
rect 34859 4320 34875 4384
rect 34939 4320 34955 4384
rect 35019 4320 35027 4384
rect 34707 3296 35027 4320
rect 34707 3232 34715 3296
rect 34779 3232 34795 3296
rect 34859 3232 34875 3296
rect 34939 3232 34955 3296
rect 35019 3232 35027 3296
rect 34707 2208 35027 3232
rect 34707 2144 34715 2208
rect 34779 2144 34795 2208
rect 34859 2144 34875 2208
rect 34939 2144 34955 2208
rect 35019 2144 35027 2208
rect 34707 2128 35027 2144
use sky130_fd_sc_hd__diode_2  ANTENNA_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 32568 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1666464484
transform 1 0 31464 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1666464484
transform 1 0 17112 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1666464484
transform 1 0 31280 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1666464484
transform 1 0 13156 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1666464484
transform 1 0 20884 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26
timestamp 1666464484
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1666464484
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1666464484
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80
timestamp 1666464484
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1666464484
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_108
timestamp 1666464484
transform 1 0 11040 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1666464484
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1666464484
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_153
timestamp 1666464484
transform 1 0 15180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_157 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 15548 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_161 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 15916 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1666464484
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_169
timestamp 1666464484
transform 1 0 16652 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_175 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 17204 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_183
timestamp 1666464484
transform 1 0 17940 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_188
timestamp 1666464484
transform 1 0 18400 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1666464484
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_202
timestamp 1666464484
transform 1 0 19688 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_217
timestamp 1666464484
transform 1 0 21068 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1666464484
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1666464484
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1666464484
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1666464484
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1666464484
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1666464484
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1666464484
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_281
timestamp 1666464484
transform 1 0 26956 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_292
timestamp 1666464484
transform 1 0 27968 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_299
timestamp 1666464484
transform 1 0 28612 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_306
timestamp 1666464484
transform 1 0 29256 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_309
timestamp 1666464484
transform 1 0 29532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_334
timestamp 1666464484
transform 1 0 31832 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1666464484
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_360
timestamp 1666464484
transform 1 0 34224 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3
timestamp 1666464484
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_7
timestamp 1666464484
transform 1 0 1748 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_29
timestamp 1666464484
transform 1 0 3772 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1666464484
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_57
timestamp 1666464484
transform 1 0 6348 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_63
timestamp 1666464484
transform 1 0 6900 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_85
timestamp 1666464484
transform 1 0 8924 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1666464484
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1666464484
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_125
timestamp 1666464484
transform 1 0 12604 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_134
timestamp 1666464484
transform 1 0 13432 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_142
timestamp 1666464484
transform 1 0 14168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_164
timestamp 1666464484
transform 1 0 16192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1666464484
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_192
timestamp 1666464484
transform 1 0 18768 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_198
timestamp 1666464484
transform 1 0 19320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_220
timestamp 1666464484
transform 1 0 21344 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp 1666464484
transform 1 0 21804 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_230
timestamp 1666464484
transform 1 0 22264 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_242
timestamp 1666464484
transform 1 0 23368 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_246
timestamp 1666464484
transform 1 0 23736 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_268
timestamp 1666464484
transform 1 0 25760 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_281
timestamp 1666464484
transform 1 0 26956 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_292
timestamp 1666464484
transform 1 0 27968 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_299
timestamp 1666464484
transform 1 0 28612 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_306
timestamp 1666464484
transform 1 0 29256 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_331
timestamp 1666464484
transform 1 0 31556 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1666464484
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_337
timestamp 1666464484
transform 1 0 32108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_360
timestamp 1666464484
transform 1 0 34224 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1666464484
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1666464484
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1666464484
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_34
timestamp 1666464484
transform 1 0 4232 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_41
timestamp 1666464484
transform 1 0 4876 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_48
timestamp 1666464484
transform 1 0 5520 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_73
timestamp 1666464484
transform 1 0 7820 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_80
timestamp 1666464484
transform 1 0 8464 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_85
timestamp 1666464484
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_90
timestamp 1666464484
transform 1 0 9384 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_94
timestamp 1666464484
transform 1 0 9752 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_98
timestamp 1666464484
transform 1 0 10120 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_105
timestamp 1666464484
transform 1 0 10764 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_117
timestamp 1666464484
transform 1 0 11868 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_125
timestamp 1666464484
transform 1 0 12604 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_131
timestamp 1666464484
transform 1 0 13156 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1666464484
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_141
timestamp 1666464484
transform 1 0 14076 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_147
timestamp 1666464484
transform 1 0 14628 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_155
timestamp 1666464484
transform 1 0 15364 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_178
timestamp 1666464484
transform 1 0 17480 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_190
timestamp 1666464484
transform 1 0 18584 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1666464484
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_202
timestamp 1666464484
transform 1 0 19688 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_209
timestamp 1666464484
transform 1 0 20332 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_234
timestamp 1666464484
transform 1 0 22632 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_246
timestamp 1666464484
transform 1 0 23736 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1666464484
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1666464484
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_258
timestamp 1666464484
transform 1 0 24840 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_270
timestamp 1666464484
transform 1 0 25944 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_282
timestamp 1666464484
transform 1 0 27048 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_288
timestamp 1666464484
transform 1 0 27600 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_292
timestamp 1666464484
transform 1 0 27968 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_299
timestamp 1666464484
transform 1 0 28612 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_306
timestamp 1666464484
transform 1 0 29256 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_309
timestamp 1666464484
transform 1 0 29532 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_314
timestamp 1666464484
transform 1 0 29992 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_321
timestamp 1666464484
transform 1 0 30636 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_346
timestamp 1666464484
transform 1 0 32936 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_353
timestamp 1666464484
transform 1 0 33580 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_360
timestamp 1666464484
transform 1 0 34224 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 1666464484
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_7
timestamp 1666464484
transform 1 0 1748 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_11
timestamp 1666464484
transform 1 0 2116 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_15
timestamp 1666464484
transform 1 0 2484 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_37
timestamp 1666464484
transform 1 0 4508 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_41
timestamp 1666464484
transform 1 0 4876 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_45
timestamp 1666464484
transform 1 0 5244 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_52
timestamp 1666464484
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1666464484
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_62
timestamp 1666464484
transform 1 0 6808 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_69
timestamp 1666464484
transform 1 0 7452 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_3_78
timestamp 1666464484
transform 1 0 8280 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_86
timestamp 1666464484
transform 1 0 9016 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_90
timestamp 1666464484
transform 1 0 9384 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_102
timestamp 1666464484
transform 1 0 10488 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1666464484
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1666464484
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_125
timestamp 1666464484
transform 1 0 12604 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_129
timestamp 1666464484
transform 1 0 12972 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_151
timestamp 1666464484
transform 1 0 14996 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_3_160
timestamp 1666464484
transform 1 0 15824 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_169
timestamp 1666464484
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_174
timestamp 1666464484
transform 1 0 17112 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_186
timestamp 1666464484
transform 1 0 18216 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_198
timestamp 1666464484
transform 1 0 19320 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_222
timestamp 1666464484
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1666464484
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1666464484
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1666464484
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1666464484
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1666464484
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1666464484
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1666464484
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_293
timestamp 1666464484
transform 1 0 28060 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_302
timestamp 1666464484
transform 1 0 28888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_309
timestamp 1666464484
transform 1 0 29532 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_334
timestamp 1666464484
transform 1 0 31832 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_337
timestamp 1666464484
transform 1 0 32108 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_362
timestamp 1666464484
transform 1 0 34408 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1666464484
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_26
timestamp 1666464484
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1666464484
transform 1 0 3772 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_52
timestamp 1666464484
transform 1 0 5888 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_59
timestamp 1666464484
transform 1 0 6532 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_66
timestamp 1666464484
transform 1 0 7176 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_73
timestamp 1666464484
transform 1 0 7820 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_80
timestamp 1666464484
transform 1 0 8464 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1666464484
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1666464484
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1666464484
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1666464484
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1666464484
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1666464484
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1666464484
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1666464484
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1666464484
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1666464484
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1666464484
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1666464484
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_197
timestamp 1666464484
transform 1 0 19228 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_208
timestamp 1666464484
transform 1 0 20240 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_220
timestamp 1666464484
transform 1 0 21344 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_232
timestamp 1666464484
transform 1 0 22448 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_244
timestamp 1666464484
transform 1 0 23552 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1666464484
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1666464484
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1666464484
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1666464484
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_301
timestamp 1666464484
transform 1 0 28796 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_306
timestamp 1666464484
transform 1 0 29256 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_309
timestamp 1666464484
transform 1 0 29532 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_315
timestamp 1666464484
transform 1 0 30084 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_337
timestamp 1666464484
transform 1 0 32108 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_362
timestamp 1666464484
transform 1 0 34408 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1666464484
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_28
timestamp 1666464484
transform 1 0 3680 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_53
timestamp 1666464484
transform 1 0 5980 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_57
timestamp 1666464484
transform 1 0 6348 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_62
timestamp 1666464484
transform 1 0 6808 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1666464484
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1666464484
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1666464484
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1666464484
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1666464484
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1666464484
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1666464484
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1666464484
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1666464484
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1666464484
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1666464484
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1666464484
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1666464484
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1666464484
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1666464484
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1666464484
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1666464484
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1666464484
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1666464484
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1666464484
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1666464484
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1666464484
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1666464484
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1666464484
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1666464484
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_305
timestamp 1666464484
transform 1 0 29164 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_316
timestamp 1666464484
transform 1 0 30176 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_324
timestamp 1666464484
transform 1 0 30912 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_328
timestamp 1666464484
transform 1 0 31280 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_337
timestamp 1666464484
transform 1 0 32108 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_362
timestamp 1666464484
transform 1 0 34408 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1666464484
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_26
timestamp 1666464484
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1666464484
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_34
timestamp 1666464484
transform 1 0 4232 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_41
timestamp 1666464484
transform 1 0 4876 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_48
timestamp 1666464484
transform 1 0 5520 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_55
timestamp 1666464484
transform 1 0 6164 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_62
timestamp 1666464484
transform 1 0 6808 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_69
timestamp 1666464484
transform 1 0 7452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_81
timestamp 1666464484
transform 1 0 8556 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1666464484
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1666464484
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1666464484
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1666464484
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1666464484
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1666464484
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1666464484
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1666464484
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1666464484
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1666464484
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1666464484
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1666464484
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1666464484
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1666464484
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1666464484
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1666464484
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1666464484
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1666464484
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1666464484
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1666464484
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1666464484
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1666464484
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1666464484
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1666464484
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_309
timestamp 1666464484
transform 1 0 29532 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_317
timestamp 1666464484
transform 1 0 30268 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_323
timestamp 1666464484
transform 1 0 30820 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_330
timestamp 1666464484
transform 1 0 31464 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_337
timestamp 1666464484
transform 1 0 32108 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_362
timestamp 1666464484
transform 1 0 34408 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3
timestamp 1666464484
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_28
timestamp 1666464484
transform 1 0 3680 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_35
timestamp 1666464484
transform 1 0 4324 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_42
timestamp 1666464484
transform 1 0 4968 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_49
timestamp 1666464484
transform 1 0 5612 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1666464484
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1666464484
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1666464484
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1666464484
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1666464484
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1666464484
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1666464484
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1666464484
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1666464484
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1666464484
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1666464484
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1666464484
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1666464484
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1666464484
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1666464484
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1666464484
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1666464484
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1666464484
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1666464484
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1666464484
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1666464484
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1666464484
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1666464484
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1666464484
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1666464484
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1666464484
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1666464484
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1666464484
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1666464484
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_329
timestamp 1666464484
transform 1 0 31372 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_334
timestamp 1666464484
transform 1 0 31832 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_337
timestamp 1666464484
transform 1 0 32108 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_362
timestamp 1666464484
transform 1 0 34408 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3
timestamp 1666464484
transform 1 0 1380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_9
timestamp 1666464484
transform 1 0 1932 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_13
timestamp 1666464484
transform 1 0 2300 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_20
timestamp 1666464484
transform 1 0 2944 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1666464484
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_34
timestamp 1666464484
transform 1 0 4232 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_41
timestamp 1666464484
transform 1 0 4876 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_48
timestamp 1666464484
transform 1 0 5520 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_60
timestamp 1666464484
transform 1 0 6624 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_72
timestamp 1666464484
transform 1 0 7728 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_85
timestamp 1666464484
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_99
timestamp 1666464484
transform 1 0 10212 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_111
timestamp 1666464484
transform 1 0 11316 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_123
timestamp 1666464484
transform 1 0 12420 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_135
timestamp 1666464484
transform 1 0 13524 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1666464484
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1666464484
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1666464484
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1666464484
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1666464484
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1666464484
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1666464484
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1666464484
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1666464484
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1666464484
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1666464484
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1666464484
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1666464484
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1666464484
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1666464484
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1666464484
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1666464484
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1666464484
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1666464484
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1666464484
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1666464484
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_333
timestamp 1666464484
transform 1 0 31740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_337
timestamp 1666464484
transform 1 0 32108 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_362
timestamp 1666464484
transform 1 0 34408 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3
timestamp 1666464484
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_28
timestamp 1666464484
transform 1 0 3680 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_35
timestamp 1666464484
transform 1 0 4324 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_47
timestamp 1666464484
transform 1 0 5428 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1666464484
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1666464484
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1666464484
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1666464484
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1666464484
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1666464484
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1666464484
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1666464484
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1666464484
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1666464484
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1666464484
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1666464484
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1666464484
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1666464484
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1666464484
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1666464484
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1666464484
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1666464484
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1666464484
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1666464484
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1666464484
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1666464484
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1666464484
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1666464484
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1666464484
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1666464484
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1666464484
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1666464484
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1666464484
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1666464484
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1666464484
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_337
timestamp 1666464484
transform 1 0 32108 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_345
timestamp 1666464484
transform 1 0 32844 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_351
timestamp 1666464484
transform 1 0 33396 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_358
timestamp 1666464484
transform 1 0 34040 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_3
timestamp 1666464484
transform 1 0 1380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_7
timestamp 1666464484
transform 1 0 1748 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_11
timestamp 1666464484
transform 1 0 2116 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_18
timestamp 1666464484
transform 1 0 2760 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_25
timestamp 1666464484
transform 1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1666464484
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1666464484
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1666464484
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1666464484
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1666464484
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1666464484
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1666464484
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1666464484
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1666464484
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1666464484
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1666464484
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1666464484
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1666464484
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1666464484
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1666464484
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1666464484
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1666464484
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1666464484
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1666464484
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1666464484
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1666464484
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1666464484
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1666464484
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1666464484
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1666464484
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1666464484
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1666464484
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1666464484
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1666464484
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1666464484
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1666464484
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1666464484
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1666464484
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_345
timestamp 1666464484
transform 1 0 32844 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_351
timestamp 1666464484
transform 1 0 33396 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_358
timestamp 1666464484
transform 1 0 34040 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1666464484
transform 1 0 1380 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_28
timestamp 1666464484
transform 1 0 3680 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_40
timestamp 1666464484
transform 1 0 4784 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_52
timestamp 1666464484
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1666464484
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1666464484
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1666464484
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1666464484
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1666464484
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1666464484
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1666464484
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1666464484
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1666464484
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1666464484
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1666464484
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1666464484
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1666464484
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1666464484
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1666464484
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1666464484
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1666464484
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1666464484
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1666464484
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1666464484
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1666464484
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1666464484
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1666464484
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1666464484
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1666464484
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1666464484
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1666464484
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1666464484
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1666464484
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1666464484
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_337
timestamp 1666464484
transform 1 0 32108 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_362
timestamp 1666464484
transform 1 0 34408 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1666464484
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1666464484
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1666464484
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1666464484
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1666464484
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1666464484
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1666464484
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1666464484
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1666464484
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1666464484
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1666464484
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1666464484
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1666464484
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1666464484
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1666464484
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1666464484
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1666464484
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1666464484
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1666464484
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1666464484
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1666464484
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1666464484
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1666464484
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1666464484
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1666464484
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1666464484
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1666464484
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1666464484
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1666464484
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1666464484
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1666464484
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1666464484
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1666464484
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1666464484
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1666464484
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_345
timestamp 1666464484
transform 1 0 32844 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_353
timestamp 1666464484
transform 1 0 33580 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_358
timestamp 1666464484
transform 1 0 34040 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1666464484
transform 1 0 1380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_7
timestamp 1666464484
transform 1 0 1748 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_11
timestamp 1666464484
transform 1 0 2116 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_18
timestamp 1666464484
transform 1 0 2760 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_30
timestamp 1666464484
transform 1 0 3864 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_42
timestamp 1666464484
transform 1 0 4968 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1666464484
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1666464484
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1666464484
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1666464484
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1666464484
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1666464484
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1666464484
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1666464484
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1666464484
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1666464484
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1666464484
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1666464484
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1666464484
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1666464484
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1666464484
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1666464484
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1666464484
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1666464484
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1666464484
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1666464484
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1666464484
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1666464484
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1666464484
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1666464484
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1666464484
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1666464484
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1666464484
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1666464484
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1666464484
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1666464484
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1666464484
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1666464484
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1666464484
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_361
timestamp 1666464484
transform 1 0 34316 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_14_3
timestamp 1666464484
transform 1 0 1380 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_12
timestamp 1666464484
transform 1 0 2208 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_24
timestamp 1666464484
transform 1 0 3312 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1666464484
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1666464484
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1666464484
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1666464484
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1666464484
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1666464484
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1666464484
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1666464484
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1666464484
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1666464484
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1666464484
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1666464484
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1666464484
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1666464484
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1666464484
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1666464484
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1666464484
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1666464484
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1666464484
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1666464484
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1666464484
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1666464484
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1666464484
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1666464484
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1666464484
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1666464484
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1666464484
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1666464484
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1666464484
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1666464484
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1666464484
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1666464484
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1666464484
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1666464484
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_357
timestamp 1666464484
transform 1 0 33948 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_362
timestamp 1666464484
transform 1 0 34408 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_3
timestamp 1666464484
transform 1 0 1380 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_28
timestamp 1666464484
transform 1 0 3680 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_40
timestamp 1666464484
transform 1 0 4784 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_52
timestamp 1666464484
transform 1 0 5888 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1666464484
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1666464484
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1666464484
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1666464484
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1666464484
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1666464484
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1666464484
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1666464484
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1666464484
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1666464484
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1666464484
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1666464484
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1666464484
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1666464484
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1666464484
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1666464484
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1666464484
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1666464484
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1666464484
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1666464484
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1666464484
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1666464484
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1666464484
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1666464484
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1666464484
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1666464484
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_305
timestamp 1666464484
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1666464484
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1666464484
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1666464484
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_337
timestamp 1666464484
transform 1 0 32108 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_345
timestamp 1666464484
transform 1 0 32844 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_351
timestamp 1666464484
transform 1 0 33396 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_358
timestamp 1666464484
transform 1 0 34040 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_3
timestamp 1666464484
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_7
timestamp 1666464484
transform 1 0 1748 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_11
timestamp 1666464484
transform 1 0 2116 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_18
timestamp 1666464484
transform 1 0 2760 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1666464484
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1666464484
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1666464484
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1666464484
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1666464484
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1666464484
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1666464484
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1666464484
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1666464484
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1666464484
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1666464484
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1666464484
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1666464484
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1666464484
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1666464484
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1666464484
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1666464484
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1666464484
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1666464484
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1666464484
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1666464484
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_221
timestamp 1666464484
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_233
timestamp 1666464484
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1666464484
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1666464484
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1666464484
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1666464484
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1666464484
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1666464484
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1666464484
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1666464484
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1666464484
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1666464484
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_333
timestamp 1666464484
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_345
timestamp 1666464484
transform 1 0 32844 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_351
timestamp 1666464484
transform 1 0 33396 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_358
timestamp 1666464484
transform 1 0 34040 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_3
timestamp 1666464484
transform 1 0 1380 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_28
timestamp 1666464484
transform 1 0 3680 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_40
timestamp 1666464484
transform 1 0 4784 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_52
timestamp 1666464484
transform 1 0 5888 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1666464484
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1666464484
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1666464484
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1666464484
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1666464484
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1666464484
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1666464484
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1666464484
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1666464484
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1666464484
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1666464484
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1666464484
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1666464484
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1666464484
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1666464484
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1666464484
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1666464484
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1666464484
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1666464484
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1666464484
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1666464484
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1666464484
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1666464484
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1666464484
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1666464484
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1666464484
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1666464484
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1666464484
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1666464484
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1666464484
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_337
timestamp 1666464484
transform 1 0 32108 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_344
timestamp 1666464484
transform 1 0 32752 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_351
timestamp 1666464484
transform 1 0 33396 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_358
timestamp 1666464484
transform 1 0 34040 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_18_3
timestamp 1666464484
transform 1 0 1380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_9
timestamp 1666464484
transform 1 0 1932 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_13
timestamp 1666464484
transform 1 0 2300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_25
timestamp 1666464484
transform 1 0 3404 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1666464484
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1666464484
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1666464484
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1666464484
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1666464484
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1666464484
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1666464484
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1666464484
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1666464484
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1666464484
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1666464484
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1666464484
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1666464484
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1666464484
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1666464484
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1666464484
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1666464484
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1666464484
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1666464484
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1666464484
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1666464484
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_233
timestamp 1666464484
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1666464484
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1666464484
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1666464484
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1666464484
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1666464484
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_289
timestamp 1666464484
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1666464484
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1666464484
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1666464484
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_321
timestamp 1666464484
transform 1 0 30636 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_330
timestamp 1666464484
transform 1 0 31464 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_337
timestamp 1666464484
transform 1 0 32108 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_362
timestamp 1666464484
transform 1 0 34408 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_3
timestamp 1666464484
transform 1 0 1380 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_9
timestamp 1666464484
transform 1 0 1932 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_13
timestamp 1666464484
transform 1 0 2300 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_25
timestamp 1666464484
transform 1 0 3404 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_37
timestamp 1666464484
transform 1 0 4508 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_49
timestamp 1666464484
transform 1 0 5612 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1666464484
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1666464484
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1666464484
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1666464484
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1666464484
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1666464484
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1666464484
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1666464484
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1666464484
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1666464484
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1666464484
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1666464484
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1666464484
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1666464484
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1666464484
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1666464484
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1666464484
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1666464484
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1666464484
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1666464484
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1666464484
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1666464484
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_261
timestamp 1666464484
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1666464484
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1666464484
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1666464484
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1666464484
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1666464484
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_317
timestamp 1666464484
transform 1 0 30268 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_325
timestamp 1666464484
transform 1 0 31004 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_330
timestamp 1666464484
transform 1 0 31464 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_337
timestamp 1666464484
transform 1 0 32108 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_362
timestamp 1666464484
transform 1 0 34408 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_3
timestamp 1666464484
transform 1 0 1380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_7
timestamp 1666464484
transform 1 0 1748 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_11
timestamp 1666464484
transform 1 0 2116 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_18
timestamp 1666464484
transform 1 0 2760 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1666464484
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1666464484
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1666464484
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1666464484
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1666464484
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1666464484
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1666464484
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1666464484
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1666464484
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1666464484
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1666464484
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1666464484
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1666464484
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1666464484
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1666464484
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1666464484
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1666464484
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1666464484
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1666464484
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1666464484
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1666464484
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_221
timestamp 1666464484
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_233
timestamp 1666464484
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1666464484
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1666464484
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1666464484
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 1666464484
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_277
timestamp 1666464484
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_289
timestamp 1666464484
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1666464484
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1666464484
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1666464484
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_321
timestamp 1666464484
transform 1 0 30636 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_325
timestamp 1666464484
transform 1 0 31004 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_329
timestamp 1666464484
transform 1 0 31372 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_336
timestamp 1666464484
transform 1 0 32016 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_343
timestamp 1666464484
transform 1 0 32660 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_351
timestamp 1666464484
transform 1 0 33396 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_356
timestamp 1666464484
transform 1 0 33856 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_3
timestamp 1666464484
transform 1 0 1380 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_28
timestamp 1666464484
transform 1 0 3680 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_40
timestamp 1666464484
transform 1 0 4784 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_52
timestamp 1666464484
transform 1 0 5888 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1666464484
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1666464484
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1666464484
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1666464484
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1666464484
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1666464484
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1666464484
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1666464484
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1666464484
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1666464484
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1666464484
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1666464484
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1666464484
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1666464484
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1666464484
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1666464484
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1666464484
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1666464484
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1666464484
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_237
timestamp 1666464484
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_249
timestamp 1666464484
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_261
timestamp 1666464484
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1666464484
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1666464484
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1666464484
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1666464484
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_305
timestamp 1666464484
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_320
timestamp 1666464484
transform 1 0 30544 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_327
timestamp 1666464484
transform 1 0 31188 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_334
timestamp 1666464484
transform 1 0 31832 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_337
timestamp 1666464484
transform 1 0 32108 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_362
timestamp 1666464484
transform 1 0 34408 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1666464484
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1666464484
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1666464484
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1666464484
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1666464484
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1666464484
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1666464484
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1666464484
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1666464484
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1666464484
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1666464484
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1666464484
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1666464484
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1666464484
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1666464484
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1666464484
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1666464484
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1666464484
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1666464484
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1666464484
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1666464484
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1666464484
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1666464484
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_233
timestamp 1666464484
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1666464484
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1666464484
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_253
timestamp 1666464484
transform 1 0 24380 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_22_264
timestamp 1666464484
transform 1 0 25392 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_273
timestamp 1666464484
transform 1 0 26220 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_280
timestamp 1666464484
transform 1 0 26864 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_292
timestamp 1666464484
transform 1 0 27968 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_304
timestamp 1666464484
transform 1 0 29072 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_309
timestamp 1666464484
transform 1 0 29532 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_320
timestamp 1666464484
transform 1 0 30544 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_327
timestamp 1666464484
transform 1 0 31188 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_334
timestamp 1666464484
transform 1 0 31832 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_340
timestamp 1666464484
transform 1 0 32384 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_362
timestamp 1666464484
transform 1 0 34408 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_3
timestamp 1666464484
transform 1 0 1380 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_14
timestamp 1666464484
transform 1 0 2392 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_21
timestamp 1666464484
transform 1 0 3036 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_33
timestamp 1666464484
transform 1 0 4140 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_45
timestamp 1666464484
transform 1 0 5244 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_53
timestamp 1666464484
transform 1 0 5980 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1666464484
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1666464484
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1666464484
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1666464484
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1666464484
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1666464484
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1666464484
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1666464484
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1666464484
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1666464484
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1666464484
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1666464484
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1666464484
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1666464484
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1666464484
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1666464484
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1666464484
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1666464484
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1666464484
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_237
timestamp 1666464484
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_249
timestamp 1666464484
transform 1 0 24012 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_260
timestamp 1666464484
transform 1 0 25024 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_267
timestamp 1666464484
transform 1 0 25668 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_274
timestamp 1666464484
transform 1 0 26312 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_281
timestamp 1666464484
transform 1 0 26956 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_286
timestamp 1666464484
transform 1 0 27416 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_295
timestamp 1666464484
transform 1 0 28244 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_302
timestamp 1666464484
transform 1 0 28888 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_309
timestamp 1666464484
transform 1 0 29532 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_316
timestamp 1666464484
transform 1 0 30176 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_323
timestamp 1666464484
transform 1 0 30820 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_330
timestamp 1666464484
transform 1 0 31464 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_337
timestamp 1666464484
transform 1 0 32108 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_342
timestamp 1666464484
transform 1 0 32568 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_349
timestamp 1666464484
transform 1 0 33212 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_356
timestamp 1666464484
transform 1 0 33856 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1666464484
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp 1666464484
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1666464484
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1666464484
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1666464484
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1666464484
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1666464484
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1666464484
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1666464484
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1666464484
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1666464484
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1666464484
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1666464484
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1666464484
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1666464484
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1666464484
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1666464484
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1666464484
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1666464484
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1666464484
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1666464484
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1666464484
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_221
timestamp 1666464484
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_233
timestamp 1666464484
transform 1 0 22540 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_237
timestamp 1666464484
transform 1 0 22908 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_241
timestamp 1666464484
transform 1 0 23276 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 1666464484
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_253
timestamp 1666464484
transform 1 0 24380 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_264
timestamp 1666464484
transform 1 0 25392 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_271
timestamp 1666464484
transform 1 0 26036 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_281
timestamp 1666464484
transform 1 0 26956 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_288
timestamp 1666464484
transform 1 0 27600 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_294
timestamp 1666464484
transform 1 0 28152 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1666464484
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1666464484
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_309
timestamp 1666464484
transform 1 0 29532 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_314
timestamp 1666464484
transform 1 0 29992 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_320
timestamp 1666464484
transform 1 0 30544 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_324
timestamp 1666464484
transform 1 0 30912 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_331
timestamp 1666464484
transform 1 0 31556 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_338
timestamp 1666464484
transform 1 0 32200 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_345
timestamp 1666464484
transform 1 0 32844 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_353
timestamp 1666464484
transform 1 0 33580 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_358
timestamp 1666464484
transform 1 0 34040 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_3
timestamp 1666464484
transform 1 0 1380 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_7
timestamp 1666464484
transform 1 0 1748 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_11
timestamp 1666464484
transform 1 0 2116 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_23
timestamp 1666464484
transform 1 0 3220 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_35
timestamp 1666464484
transform 1 0 4324 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_47
timestamp 1666464484
transform 1 0 5428 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1666464484
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1666464484
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1666464484
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1666464484
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1666464484
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1666464484
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1666464484
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1666464484
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1666464484
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1666464484
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1666464484
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1666464484
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1666464484
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1666464484
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1666464484
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1666464484
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1666464484
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1666464484
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1666464484
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_225
timestamp 1666464484
transform 1 0 21804 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_232
timestamp 1666464484
transform 1 0 22448 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_236
timestamp 1666464484
transform 1 0 22816 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_240
timestamp 1666464484
transform 1 0 23184 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_244
timestamp 1666464484
transform 1 0 23552 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_249
timestamp 1666464484
transform 1 0 24012 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_256
timestamp 1666464484
transform 1 0 24656 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_262
timestamp 1666464484
transform 1 0 25208 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_267
timestamp 1666464484
transform 1 0 25668 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_275
timestamp 1666464484
transform 1 0 26404 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1666464484
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_281
timestamp 1666464484
transform 1 0 26956 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_290
timestamp 1666464484
transform 1 0 27784 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_301
timestamp 1666464484
transform 1 0 28796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_308
timestamp 1666464484
transform 1 0 29440 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_315
timestamp 1666464484
transform 1 0 30084 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_322
timestamp 1666464484
transform 1 0 30728 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_328
timestamp 1666464484
transform 1 0 31280 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_332
timestamp 1666464484
transform 1 0 31648 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_337
timestamp 1666464484
transform 1 0 32108 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_342
timestamp 1666464484
transform 1 0 32568 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_349
timestamp 1666464484
transform 1 0 33212 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_353
timestamp 1666464484
transform 1 0 33580 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_357
timestamp 1666464484
transform 1 0 33948 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_363
timestamp 1666464484
transform 1 0 34500 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_3
timestamp 1666464484
transform 1 0 1380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_7
timestamp 1666464484
transform 1 0 1748 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_11
timestamp 1666464484
transform 1 0 2116 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_18
timestamp 1666464484
transform 1 0 2760 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 1666464484
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1666464484
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1666464484
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1666464484
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1666464484
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1666464484
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1666464484
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1666464484
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1666464484
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1666464484
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1666464484
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1666464484
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1666464484
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1666464484
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1666464484
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1666464484
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1666464484
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1666464484
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1666464484
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1666464484
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_209
timestamp 1666464484
transform 1 0 20332 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_26_216
timestamp 1666464484
transform 1 0 20976 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_222
timestamp 1666464484
transform 1 0 21528 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_226
timestamp 1666464484
transform 1 0 21896 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_234
timestamp 1666464484
transform 1 0 22632 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_241
timestamp 1666464484
transform 1 0 23276 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_245
timestamp 1666464484
transform 1 0 23644 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp 1666464484
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1666464484
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_259
timestamp 1666464484
transform 1 0 24932 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_267
timestamp 1666464484
transform 1 0 25668 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_271
timestamp 1666464484
transform 1 0 26036 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_277
timestamp 1666464484
transform 1 0 26588 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_291
timestamp 1666464484
transform 1 0 27876 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_302
timestamp 1666464484
transform 1 0 28888 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_309
timestamp 1666464484
transform 1 0 29532 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_315
timestamp 1666464484
transform 1 0 30084 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_321
timestamp 1666464484
transform 1 0 30636 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_325
timestamp 1666464484
transform 1 0 31004 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_26_334
timestamp 1666464484
transform 1 0 31832 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_340
timestamp 1666464484
transform 1 0 32384 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_362
timestamp 1666464484
transform 1 0 34408 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1666464484
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_28
timestamp 1666464484
transform 1 0 3680 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_40
timestamp 1666464484
transform 1 0 4784 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_52
timestamp 1666464484
transform 1 0 5888 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1666464484
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1666464484
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1666464484
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1666464484
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1666464484
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1666464484
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1666464484
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1666464484
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1666464484
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1666464484
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1666464484
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1666464484
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1666464484
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1666464484
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_193
timestamp 1666464484
transform 1 0 18860 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_200
timestamp 1666464484
transform 1 0 19504 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1666464484
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_225
timestamp 1666464484
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_232
timestamp 1666464484
transform 1 0 22448 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_252
timestamp 1666464484
transform 1 0 24288 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_263
timestamp 1666464484
transform 1 0 25300 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_271
timestamp 1666464484
transform 1 0 26036 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_278
timestamp 1666464484
transform 1 0 26680 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_281
timestamp 1666464484
transform 1 0 26956 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_299
timestamp 1666464484
transform 1 0 28612 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_310
timestamp 1666464484
transform 1 0 29624 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_318
timestamp 1666464484
transform 1 0 30360 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_326
timestamp 1666464484
transform 1 0 31096 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_334
timestamp 1666464484
transform 1 0 31832 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_337
timestamp 1666464484
transform 1 0 32108 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_362
timestamp 1666464484
transform 1 0 34408 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_3
timestamp 1666464484
transform 1 0 1380 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_9
timestamp 1666464484
transform 1 0 1932 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_13
timestamp 1666464484
transform 1 0 2300 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_25
timestamp 1666464484
transform 1 0 3404 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1666464484
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1666464484
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1666464484
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1666464484
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1666464484
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1666464484
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1666464484
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1666464484
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1666464484
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1666464484
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1666464484
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1666464484
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1666464484
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1666464484
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1666464484
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1666464484
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1666464484
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1666464484
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1666464484
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_215
timestamp 1666464484
transform 1 0 20884 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_221
timestamp 1666464484
transform 1 0 21436 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_238
timestamp 1666464484
transform 1 0 23000 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_242
timestamp 1666464484
transform 1 0 23368 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_249
timestamp 1666464484
transform 1 0 24012 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1666464484
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_271
timestamp 1666464484
transform 1 0 26036 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_291
timestamp 1666464484
transform 1 0 27876 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_295
timestamp 1666464484
transform 1 0 28244 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_304
timestamp 1666464484
transform 1 0 29072 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_309
timestamp 1666464484
transform 1 0 29532 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_328
timestamp 1666464484
transform 1 0 31280 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_336
timestamp 1666464484
transform 1 0 32016 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_340
timestamp 1666464484
transform 1 0 32384 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_362
timestamp 1666464484
transform 1 0 34408 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1666464484
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_28
timestamp 1666464484
transform 1 0 3680 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_40
timestamp 1666464484
transform 1 0 4784 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_52
timestamp 1666464484
transform 1 0 5888 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1666464484
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1666464484
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1666464484
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1666464484
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1666464484
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1666464484
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1666464484
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1666464484
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1666464484
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1666464484
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1666464484
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1666464484
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1666464484
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_178
timestamp 1666464484
transform 1 0 17480 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_186
timestamp 1666464484
transform 1 0 18216 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_204
timestamp 1666464484
transform 1 0 19872 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_214
timestamp 1666464484
transform 1 0 20792 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_222
timestamp 1666464484
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1666464484
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_243
timestamp 1666464484
transform 1 0 23460 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_263
timestamp 1666464484
transform 1 0 25300 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_272
timestamp 1666464484
transform 1 0 26128 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_281
timestamp 1666464484
transform 1 0 26956 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_293
timestamp 1666464484
transform 1 0 28060 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_313
timestamp 1666464484
transform 1 0 29900 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_321
timestamp 1666464484
transform 1 0 30636 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_329
timestamp 1666464484
transform 1 0 31372 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_334
timestamp 1666464484
transform 1 0 31832 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_337
timestamp 1666464484
transform 1 0 32108 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_343
timestamp 1666464484
transform 1 0 32660 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_351
timestamp 1666464484
transform 1 0 33396 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_359
timestamp 1666464484
transform 1 0 34132 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_363
timestamp 1666464484
transform 1 0 34500 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_3
timestamp 1666464484
transform 1 0 1380 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_7
timestamp 1666464484
transform 1 0 1748 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_11
timestamp 1666464484
transform 1 0 2116 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_18
timestamp 1666464484
transform 1 0 2760 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_26
timestamp 1666464484
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1666464484
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1666464484
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1666464484
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1666464484
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1666464484
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1666464484
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1666464484
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1666464484
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1666464484
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1666464484
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1666464484
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1666464484
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1666464484
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1666464484
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_165
timestamp 1666464484
transform 1 0 16284 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_173
timestamp 1666464484
transform 1 0 17020 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_182
timestamp 1666464484
transform 1 0 17848 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1666464484
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_197
timestamp 1666464484
transform 1 0 19228 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_201
timestamp 1666464484
transform 1 0 19596 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_218
timestamp 1666464484
transform 1 0 21160 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_227
timestamp 1666464484
transform 1 0 21988 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_236
timestamp 1666464484
transform 1 0 22816 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_244
timestamp 1666464484
transform 1 0 23552 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1666464484
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1666464484
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_261
timestamp 1666464484
transform 1 0 25116 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_267
timestamp 1666464484
transform 1 0 25668 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_274
timestamp 1666464484
transform 1 0 26312 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_287
timestamp 1666464484
transform 1 0 27508 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_298
timestamp 1666464484
transform 1 0 28520 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_306
timestamp 1666464484
transform 1 0 29256 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_309
timestamp 1666464484
transform 1 0 29532 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_317
timestamp 1666464484
transform 1 0 30268 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_325
timestamp 1666464484
transform 1 0 31004 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_342
timestamp 1666464484
transform 1 0 32568 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_350
timestamp 1666464484
transform 1 0 33304 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_358
timestamp 1666464484
transform 1 0 34040 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1666464484
transform 1 0 1380 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_28
timestamp 1666464484
transform 1 0 3680 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_40
timestamp 1666464484
transform 1 0 4784 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_52
timestamp 1666464484
transform 1 0 5888 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1666464484
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1666464484
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1666464484
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1666464484
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1666464484
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1666464484
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1666464484
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1666464484
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1666464484
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_149
timestamp 1666464484
transform 1 0 14812 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_153
timestamp 1666464484
transform 1 0 15180 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_157
timestamp 1666464484
transform 1 0 15548 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1666464484
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1666464484
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_178
timestamp 1666464484
transform 1 0 17480 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_186
timestamp 1666464484
transform 1 0 18216 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_192
timestamp 1666464484
transform 1 0 18768 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_199
timestamp 1666464484
transform 1 0 19412 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_206
timestamp 1666464484
transform 1 0 20056 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_216
timestamp 1666464484
transform 1 0 20976 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1666464484
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_233
timestamp 1666464484
transform 1 0 22540 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_243
timestamp 1666464484
transform 1 0 23460 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_252
timestamp 1666464484
transform 1 0 24288 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_258
timestamp 1666464484
transform 1 0 24840 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_264
timestamp 1666464484
transform 1 0 25392 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_268
timestamp 1666464484
transform 1 0 25760 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_276
timestamp 1666464484
transform 1 0 26496 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_281
timestamp 1666464484
transform 1 0 26956 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_290
timestamp 1666464484
transform 1 0 27784 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_296
timestamp 1666464484
transform 1 0 28336 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_305
timestamp 1666464484
transform 1 0 29164 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_313
timestamp 1666464484
transform 1 0 29900 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_317
timestamp 1666464484
transform 1 0 30268 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_334
timestamp 1666464484
transform 1 0 31832 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_337
timestamp 1666464484
transform 1 0 32108 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_362
timestamp 1666464484
transform 1 0 34408 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_3
timestamp 1666464484
transform 1 0 1380 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_9
timestamp 1666464484
transform 1 0 1932 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_13
timestamp 1666464484
transform 1 0 2300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_25
timestamp 1666464484
transform 1 0 3404 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1666464484
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1666464484
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1666464484
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1666464484
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1666464484
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1666464484
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1666464484
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1666464484
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1666464484
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1666464484
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1666464484
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1666464484
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1666464484
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_153
timestamp 1666464484
transform 1 0 15180 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_161
timestamp 1666464484
transform 1 0 15916 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_165
timestamp 1666464484
transform 1 0 16284 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_175
timestamp 1666464484
transform 1 0 17204 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_179
timestamp 1666464484
transform 1 0 17572 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_183
timestamp 1666464484
transform 1 0 17940 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_193
timestamp 1666464484
transform 1 0 18860 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_197
timestamp 1666464484
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_215
timestamp 1666464484
transform 1 0 20884 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_226
timestamp 1666464484
transform 1 0 21896 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_230
timestamp 1666464484
transform 1 0 22264 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_247
timestamp 1666464484
transform 1 0 23828 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1666464484
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 1666464484
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_271
timestamp 1666464484
transform 1 0 26036 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_275
timestamp 1666464484
transform 1 0 26404 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_284
timestamp 1666464484
transform 1 0 27232 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_288
timestamp 1666464484
transform 1 0 27600 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_297
timestamp 1666464484
transform 1 0 28428 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_306
timestamp 1666464484
transform 1 0 29256 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_309
timestamp 1666464484
transform 1 0 29532 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_327
timestamp 1666464484
transform 1 0 31188 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_336
timestamp 1666464484
transform 1 0 32016 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_340
timestamp 1666464484
transform 1 0 32384 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_362
timestamp 1666464484
transform 1 0 34408 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1666464484
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1666464484
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1666464484
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1666464484
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1666464484
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1666464484
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1666464484
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1666464484
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1666464484
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1666464484
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1666464484
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1666464484
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1666464484
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1666464484
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1666464484
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1666464484
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_161
timestamp 1666464484
transform 1 0 15916 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_165
timestamp 1666464484
transform 1 0 16284 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_169
timestamp 1666464484
transform 1 0 16652 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_173
timestamp 1666464484
transform 1 0 17020 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_180
timestamp 1666464484
transform 1 0 17664 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_189
timestamp 1666464484
transform 1 0 18492 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_197
timestamp 1666464484
transform 1 0 19228 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_215
timestamp 1666464484
transform 1 0 20884 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1666464484
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1666464484
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_243
timestamp 1666464484
transform 1 0 23460 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_253
timestamp 1666464484
transform 1 0 24380 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_267
timestamp 1666464484
transform 1 0 25668 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_278
timestamp 1666464484
transform 1 0 26680 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_281
timestamp 1666464484
transform 1 0 26956 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_299
timestamp 1666464484
transform 1 0 28612 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_310
timestamp 1666464484
transform 1 0 29624 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_321
timestamp 1666464484
transform 1 0 30636 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_331
timestamp 1666464484
transform 1 0 31556 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1666464484
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_337
timestamp 1666464484
transform 1 0 32108 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_355
timestamp 1666464484
transform 1 0 33764 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_362
timestamp 1666464484
transform 1 0 34408 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1666464484
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1666464484
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1666464484
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1666464484
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1666464484
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1666464484
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1666464484
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1666464484
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1666464484
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1666464484
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1666464484
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1666464484
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1666464484
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1666464484
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1666464484
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1666464484
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_153
timestamp 1666464484
transform 1 0 15180 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_161
timestamp 1666464484
transform 1 0 15916 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_170
timestamp 1666464484
transform 1 0 16744 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_182
timestamp 1666464484
transform 1 0 17848 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1666464484
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1666464484
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_202
timestamp 1666464484
transform 1 0 19688 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_210
timestamp 1666464484
transform 1 0 20424 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_234
timestamp 1666464484
transform 1 0 22632 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_242
timestamp 1666464484
transform 1 0 23368 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1666464484
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_253
timestamp 1666464484
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_261
timestamp 1666464484
transform 1 0 25116 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_269
timestamp 1666464484
transform 1 0 25852 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_291
timestamp 1666464484
transform 1 0 27876 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_304
timestamp 1666464484
transform 1 0 29072 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_309
timestamp 1666464484
transform 1 0 29532 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_316
timestamp 1666464484
transform 1 0 30176 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_325
timestamp 1666464484
transform 1 0 31004 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_331
timestamp 1666464484
transform 1 0 31556 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_337
timestamp 1666464484
transform 1 0 32108 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_362
timestamp 1666464484
transform 1 0 34408 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1666464484
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1666464484
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1666464484
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1666464484
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1666464484
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1666464484
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1666464484
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1666464484
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1666464484
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1666464484
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1666464484
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1666464484
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1666464484
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1666464484
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1666464484
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_149
timestamp 1666464484
transform 1 0 14812 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_155
timestamp 1666464484
transform 1 0 15364 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1666464484
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_169
timestamp 1666464484
transform 1 0 16652 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_173
timestamp 1666464484
transform 1 0 17020 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_182
timestamp 1666464484
transform 1 0 17848 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_190
timestamp 1666464484
transform 1 0 18584 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_207
timestamp 1666464484
transform 1 0 20148 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_35_222
timestamp 1666464484
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1666464484
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_234
timestamp 1666464484
transform 1 0 22632 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_242
timestamp 1666464484
transform 1 0 23368 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_259
timestamp 1666464484
transform 1 0 24932 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_267
timestamp 1666464484
transform 1 0 25668 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_278
timestamp 1666464484
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_281
timestamp 1666464484
transform 1 0 26956 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_285
timestamp 1666464484
transform 1 0 27324 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_302
timestamp 1666464484
transform 1 0 28888 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_311
timestamp 1666464484
transform 1 0 29716 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_322
timestamp 1666464484
transform 1 0 30728 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_331
timestamp 1666464484
transform 1 0 31556 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1666464484
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_337
timestamp 1666464484
transform 1 0 32108 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_361
timestamp 1666464484
transform 1 0 34316 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1666464484
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1666464484
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1666464484
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1666464484
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1666464484
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1666464484
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1666464484
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1666464484
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1666464484
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1666464484
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1666464484
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1666464484
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1666464484
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1666464484
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1666464484
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1666464484
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_153
timestamp 1666464484
transform 1 0 15180 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_168
timestamp 1666464484
transform 1 0 16560 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_172
timestamp 1666464484
transform 1 0 16928 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_180
timestamp 1666464484
transform 1 0 17664 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_194
timestamp 1666464484
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_197
timestamp 1666464484
transform 1 0 19228 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_205
timestamp 1666464484
transform 1 0 19964 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_216
timestamp 1666464484
transform 1 0 20976 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_222
timestamp 1666464484
transform 1 0 21528 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_231
timestamp 1666464484
transform 1 0 22356 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_242
timestamp 1666464484
transform 1 0 23368 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1666464484
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1666464484
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_261
timestamp 1666464484
transform 1 0 25116 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_269
timestamp 1666464484
transform 1 0 25852 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_278
timestamp 1666464484
transform 1 0 26680 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_284
timestamp 1666464484
transform 1 0 27232 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_293
timestamp 1666464484
transform 1 0 28060 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_304
timestamp 1666464484
transform 1 0 29072 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_309
timestamp 1666464484
transform 1 0 29532 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_327
timestamp 1666464484
transform 1 0 31188 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_337
timestamp 1666464484
transform 1 0 32108 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_343
timestamp 1666464484
transform 1 0 32660 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_360
timestamp 1666464484
transform 1 0 34224 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1666464484
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1666464484
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1666464484
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1666464484
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1666464484
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1666464484
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1666464484
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1666464484
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1666464484
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1666464484
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1666464484
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1666464484
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1666464484
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1666464484
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1666464484
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1666464484
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1666464484
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1666464484
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_169
timestamp 1666464484
transform 1 0 16652 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_179
timestamp 1666464484
transform 1 0 17572 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_187
timestamp 1666464484
transform 1 0 18308 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_204
timestamp 1666464484
transform 1 0 19872 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_219
timestamp 1666464484
transform 1 0 21252 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1666464484
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_225
timestamp 1666464484
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_243
timestamp 1666464484
transform 1 0 23460 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_263
timestamp 1666464484
transform 1 0 25300 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_271
timestamp 1666464484
transform 1 0 26036 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_278
timestamp 1666464484
transform 1 0 26680 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_281
timestamp 1666464484
transform 1 0 26956 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_287
timestamp 1666464484
transform 1 0 27508 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_296
timestamp 1666464484
transform 1 0 28336 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_306
timestamp 1666464484
transform 1 0 29256 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_37_330
timestamp 1666464484
transform 1 0 31464 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_37_337
timestamp 1666464484
transform 1 0 32108 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_355
timestamp 1666464484
transform 1 0 33764 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_362
timestamp 1666464484
transform 1 0 34408 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1666464484
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1666464484
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1666464484
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1666464484
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1666464484
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1666464484
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1666464484
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1666464484
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1666464484
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1666464484
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1666464484
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1666464484
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1666464484
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1666464484
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1666464484
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1666464484
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1666464484
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_165
timestamp 1666464484
transform 1 0 16284 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_171
timestamp 1666464484
transform 1 0 16836 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_183
timestamp 1666464484
transform 1 0 17940 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_189
timestamp 1666464484
transform 1 0 18492 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_194
timestamp 1666464484
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1666464484
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_205
timestamp 1666464484
transform 1 0 19964 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_213
timestamp 1666464484
transform 1 0 20700 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_234
timestamp 1666464484
transform 1 0 22632 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_244
timestamp 1666464484
transform 1 0 23552 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1666464484
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_261
timestamp 1666464484
transform 1 0 25116 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_281
timestamp 1666464484
transform 1 0 26956 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_291
timestamp 1666464484
transform 1 0 27876 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_38_306
timestamp 1666464484
transform 1 0 29256 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_309
timestamp 1666464484
transform 1 0 29532 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_326
timestamp 1666464484
transform 1 0 31096 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_330
timestamp 1666464484
transform 1 0 31464 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_337
timestamp 1666464484
transform 1 0 32108 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_362
timestamp 1666464484
transform 1 0 34408 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1666464484
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1666464484
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1666464484
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1666464484
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1666464484
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1666464484
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1666464484
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1666464484
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1666464484
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1666464484
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1666464484
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1666464484
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1666464484
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1666464484
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1666464484
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_149
timestamp 1666464484
transform 1 0 14812 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_157
timestamp 1666464484
transform 1 0 15548 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_166
timestamp 1666464484
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_169
timestamp 1666464484
transform 1 0 16652 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_178
timestamp 1666464484
transform 1 0 17480 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_191
timestamp 1666464484
transform 1 0 18676 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_211
timestamp 1666464484
transform 1 0 20516 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_222
timestamp 1666464484
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 1666464484
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_233
timestamp 1666464484
transform 1 0 22540 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_240
timestamp 1666464484
transform 1 0 23184 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_260
timestamp 1666464484
transform 1 0 25024 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_272
timestamp 1666464484
transform 1 0 26128 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_281
timestamp 1666464484
transform 1 0 26956 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_290
timestamp 1666464484
transform 1 0 27784 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_298
timestamp 1666464484
transform 1 0 28520 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_319
timestamp 1666464484
transform 1 0 30452 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1666464484
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1666464484
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_337
timestamp 1666464484
transform 1 0 32108 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_362
timestamp 1666464484
transform 1 0 34408 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1666464484
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1666464484
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1666464484
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1666464484
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1666464484
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1666464484
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1666464484
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1666464484
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1666464484
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1666464484
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1666464484
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1666464484
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1666464484
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1666464484
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1666464484
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1666464484
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_153
timestamp 1666464484
transform 1 0 15180 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_160
timestamp 1666464484
transform 1 0 15824 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_171
timestamp 1666464484
transform 1 0 16836 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_181
timestamp 1666464484
transform 1 0 17756 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_185
timestamp 1666464484
transform 1 0 18124 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_194
timestamp 1666464484
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1666464484
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_215
timestamp 1666464484
transform 1 0 20884 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_223
timestamp 1666464484
transform 1 0 21620 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_230
timestamp 1666464484
transform 1 0 22264 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_240
timestamp 1666464484
transform 1 0 23184 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_249
timestamp 1666464484
transform 1 0 24012 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_40_253
timestamp 1666464484
transform 1 0 24380 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_263
timestamp 1666464484
transform 1 0 25300 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_273
timestamp 1666464484
transform 1 0 26220 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_40_286
timestamp 1666464484
transform 1 0 27416 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1666464484
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1666464484
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_309
timestamp 1666464484
transform 1 0 29532 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_317
timestamp 1666464484
transform 1 0 30268 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_327
timestamp 1666464484
transform 1 0 31188 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_337
timestamp 1666464484
transform 1 0 32108 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_362
timestamp 1666464484
transform 1 0 34408 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_3
timestamp 1666464484
transform 1 0 1380 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_9
timestamp 1666464484
transform 1 0 1932 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_13
timestamp 1666464484
transform 1 0 2300 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_25
timestamp 1666464484
transform 1 0 3404 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_37
timestamp 1666464484
transform 1 0 4508 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_49
timestamp 1666464484
transform 1 0 5612 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1666464484
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1666464484
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1666464484
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1666464484
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1666464484
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1666464484
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1666464484
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1666464484
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1666464484
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1666464484
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1666464484
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_161
timestamp 1666464484
transform 1 0 15916 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_166
timestamp 1666464484
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_169
timestamp 1666464484
transform 1 0 16652 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_182
timestamp 1666464484
transform 1 0 17848 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_189
timestamp 1666464484
transform 1 0 18492 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_196
timestamp 1666464484
transform 1 0 19136 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_203
timestamp 1666464484
transform 1 0 19780 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_213
timestamp 1666464484
transform 1 0 20700 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_222
timestamp 1666464484
transform 1 0 21528 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_225
timestamp 1666464484
transform 1 0 21804 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_231
timestamp 1666464484
transform 1 0 22356 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_248
timestamp 1666464484
transform 1 0 23920 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_268
timestamp 1666464484
transform 1 0 25760 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_278
timestamp 1666464484
transform 1 0 26680 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_281
timestamp 1666464484
transform 1 0 26956 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_293
timestamp 1666464484
transform 1 0 28060 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_313
timestamp 1666464484
transform 1 0 29900 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_322
timestamp 1666464484
transform 1 0 30728 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_41_333
timestamp 1666464484
transform 1 0 31740 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_337
timestamp 1666464484
transform 1 0 32108 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_346
timestamp 1666464484
transform 1 0 32936 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_357
timestamp 1666464484
transform 1 0 33948 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_363
timestamp 1666464484
transform 1 0 34500 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_3
timestamp 1666464484
transform 1 0 1380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_26
timestamp 1666464484
transform 1 0 3496 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1666464484
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1666464484
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1666464484
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1666464484
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1666464484
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1666464484
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1666464484
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1666464484
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1666464484
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1666464484
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1666464484
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1666464484
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1666464484
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_153
timestamp 1666464484
transform 1 0 15180 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_157
timestamp 1666464484
transform 1 0 15548 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_164
timestamp 1666464484
transform 1 0 16192 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_171
timestamp 1666464484
transform 1 0 16836 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_180
timestamp 1666464484
transform 1 0 17664 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_184
timestamp 1666464484
transform 1 0 18032 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_192
timestamp 1666464484
transform 1 0 18768 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_197
timestamp 1666464484
transform 1 0 19228 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_207
timestamp 1666464484
transform 1 0 20148 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_213
timestamp 1666464484
transform 1 0 20700 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_230
timestamp 1666464484
transform 1 0 22264 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_243
timestamp 1666464484
transform 1 0 23460 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_250
timestamp 1666464484
transform 1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_253
timestamp 1666464484
transform 1 0 24380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_261
timestamp 1666464484
transform 1 0 25116 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_276
timestamp 1666464484
transform 1 0 26496 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_287
timestamp 1666464484
transform 1 0 27508 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_297
timestamp 1666464484
transform 1 0 28428 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_306
timestamp 1666464484
transform 1 0 29256 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_309
timestamp 1666464484
transform 1 0 29532 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_324
timestamp 1666464484
transform 1 0 30912 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_337
timestamp 1666464484
transform 1 0 32108 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_362
timestamp 1666464484
transform 1 0 34408 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_3
timestamp 1666464484
transform 1 0 1380 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_7
timestamp 1666464484
transform 1 0 1748 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_11
timestamp 1666464484
transform 1 0 2116 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_23
timestamp 1666464484
transform 1 0 3220 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_35
timestamp 1666464484
transform 1 0 4324 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_47
timestamp 1666464484
transform 1 0 5428 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1666464484
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1666464484
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1666464484
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1666464484
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1666464484
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1666464484
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1666464484
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1666464484
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1666464484
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1666464484
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_149
timestamp 1666464484
transform 1 0 14812 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_155
timestamp 1666464484
transform 1 0 15364 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_159
timestamp 1666464484
transform 1 0 15732 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_166
timestamp 1666464484
transform 1 0 16376 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_169
timestamp 1666464484
transform 1 0 16652 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_175
timestamp 1666464484
transform 1 0 17204 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_184
timestamp 1666464484
transform 1 0 18032 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_194
timestamp 1666464484
transform 1 0 18952 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_214
timestamp 1666464484
transform 1 0 20792 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_222
timestamp 1666464484
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_225
timestamp 1666464484
transform 1 0 21804 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_230
timestamp 1666464484
transform 1 0 22264 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_250
timestamp 1666464484
transform 1 0 24104 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_270
timestamp 1666464484
transform 1 0 25944 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_278
timestamp 1666464484
transform 1 0 26680 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_281
timestamp 1666464484
transform 1 0 26956 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_295
timestamp 1666464484
transform 1 0 28244 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_315
timestamp 1666464484
transform 1 0 30084 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_323
timestamp 1666464484
transform 1 0 30820 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_333
timestamp 1666464484
transform 1 0 31740 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_337
timestamp 1666464484
transform 1 0 32108 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_362
timestamp 1666464484
transform 1 0 34408 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1666464484
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1666464484
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1666464484
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1666464484
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1666464484
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1666464484
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1666464484
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1666464484
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1666464484
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1666464484
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1666464484
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1666464484
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1666464484
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1666464484
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1666464484
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1666464484
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1666464484
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_165
timestamp 1666464484
transform 1 0 16284 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_174
timestamp 1666464484
transform 1 0 17112 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_187
timestamp 1666464484
transform 1 0 18308 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_194
timestamp 1666464484
transform 1 0 18952 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_197
timestamp 1666464484
transform 1 0 19228 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_202
timestamp 1666464484
transform 1 0 19688 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_206
timestamp 1666464484
transform 1 0 20056 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_210
timestamp 1666464484
transform 1 0 20424 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_234
timestamp 1666464484
transform 1 0 22632 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_246
timestamp 1666464484
transform 1 0 23736 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_44_253
timestamp 1666464484
transform 1 0 24380 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_262
timestamp 1666464484
transform 1 0 25208 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_274
timestamp 1666464484
transform 1 0 26312 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_282
timestamp 1666464484
transform 1 0 27048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_299
timestamp 1666464484
transform 1 0 28612 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_306
timestamp 1666464484
transform 1 0 29256 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_309
timestamp 1666464484
transform 1 0 29532 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_44_321
timestamp 1666464484
transform 1 0 30636 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_329
timestamp 1666464484
transform 1 0 31372 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_338
timestamp 1666464484
transform 1 0 32200 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_360
timestamp 1666464484
transform 1 0 34224 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1666464484
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1666464484
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1666464484
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1666464484
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1666464484
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1666464484
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_57
timestamp 1666464484
transform 1 0 6348 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_62
timestamp 1666464484
transform 1 0 6808 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_74
timestamp 1666464484
transform 1 0 7912 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_82
timestamp 1666464484
transform 1 0 8648 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_86
timestamp 1666464484
transform 1 0 9016 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_98
timestamp 1666464484
transform 1 0 10120 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_110
timestamp 1666464484
transform 1 0 11224 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1666464484
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1666464484
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1666464484
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1666464484
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_161
timestamp 1666464484
transform 1 0 15916 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_166
timestamp 1666464484
transform 1 0 16376 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_169
timestamp 1666464484
transform 1 0 16652 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_174
timestamp 1666464484
transform 1 0 17112 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_185
timestamp 1666464484
transform 1 0 18124 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_194
timestamp 1666464484
transform 1 0 18952 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_198
timestamp 1666464484
transform 1 0 19320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_215
timestamp 1666464484
transform 1 0 20884 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_222
timestamp 1666464484
transform 1 0 21528 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_225
timestamp 1666464484
transform 1 0 21804 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_243
timestamp 1666464484
transform 1 0 23460 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_247
timestamp 1666464484
transform 1 0 23828 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_254
timestamp 1666464484
transform 1 0 24472 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_278
timestamp 1666464484
transform 1 0 26680 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_281
timestamp 1666464484
transform 1 0 26956 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_303
timestamp 1666464484
transform 1 0 28980 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_315
timestamp 1666464484
transform 1 0 30084 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_323
timestamp 1666464484
transform 1 0 30820 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_334
timestamp 1666464484
transform 1 0 31832 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_337
timestamp 1666464484
transform 1 0 32108 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_346
timestamp 1666464484
transform 1 0 32936 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_356
timestamp 1666464484
transform 1 0 33856 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1666464484
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1666464484
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1666464484
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1666464484
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1666464484
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_53
timestamp 1666464484
transform 1 0 5980 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_57
timestamp 1666464484
transform 1 0 6348 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_79
timestamp 1666464484
transform 1 0 8372 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1666464484
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1666464484
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1666464484
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1666464484
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1666464484
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1666464484
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1666464484
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1666464484
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_153
timestamp 1666464484
transform 1 0 15180 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_159
timestamp 1666464484
transform 1 0 15732 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_163
timestamp 1666464484
transform 1 0 16100 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_173
timestamp 1666464484
transform 1 0 17020 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_185
timestamp 1666464484
transform 1 0 18124 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_194
timestamp 1666464484
transform 1 0 18952 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_197
timestamp 1666464484
transform 1 0 19228 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_215
timestamp 1666464484
transform 1 0 20884 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_235
timestamp 1666464484
transform 1 0 22724 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_246
timestamp 1666464484
transform 1 0 23736 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_46_253
timestamp 1666464484
transform 1 0 24380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_259
timestamp 1666464484
transform 1 0 24932 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_271
timestamp 1666464484
transform 1 0 26036 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_281
timestamp 1666464484
transform 1 0 26956 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_289
timestamp 1666464484
transform 1 0 27692 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_296
timestamp 1666464484
transform 1 0 28336 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_306
timestamp 1666464484
transform 1 0 29256 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_309
timestamp 1666464484
transform 1 0 29532 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_318
timestamp 1666464484
transform 1 0 30360 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_326
timestamp 1666464484
transform 1 0 31096 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_334
timestamp 1666464484
transform 1 0 31832 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_340
timestamp 1666464484
transform 1 0 32384 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_344
timestamp 1666464484
transform 1 0 32752 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_362
timestamp 1666464484
transform 1 0 34408 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1666464484
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1666464484
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1666464484
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1666464484
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1666464484
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1666464484
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1666464484
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1666464484
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1666464484
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1666464484
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1666464484
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1666464484
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1666464484
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1666464484
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1666464484
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_149
timestamp 1666464484
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_161
timestamp 1666464484
transform 1 0 15916 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_166
timestamp 1666464484
transform 1 0 16376 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_47_169
timestamp 1666464484
transform 1 0 16652 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_175
timestamp 1666464484
transform 1 0 17204 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_185
timestamp 1666464484
transform 1 0 18124 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_205
timestamp 1666464484
transform 1 0 19964 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_213
timestamp 1666464484
transform 1 0 20700 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_222
timestamp 1666464484
transform 1 0 21528 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_47_225
timestamp 1666464484
transform 1 0 21804 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_244
timestamp 1666464484
transform 1 0 23552 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_251
timestamp 1666464484
transform 1 0 24196 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_271
timestamp 1666464484
transform 1 0 26036 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_278
timestamp 1666464484
transform 1 0 26680 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_281
timestamp 1666464484
transform 1 0 26956 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_47_288
timestamp 1666464484
transform 1 0 27600 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_294
timestamp 1666464484
transform 1 0 28152 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_302
timestamp 1666464484
transform 1 0 28888 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_315
timestamp 1666464484
transform 1 0 30084 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_323
timestamp 1666464484
transform 1 0 30820 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_334
timestamp 1666464484
transform 1 0 31832 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_337
timestamp 1666464484
transform 1 0 32108 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_362
timestamp 1666464484
transform 1 0 34408 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1666464484
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1666464484
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1666464484
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1666464484
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1666464484
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1666464484
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1666464484
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1666464484
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1666464484
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1666464484
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1666464484
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1666464484
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1666464484
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1666464484
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1666464484
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1666464484
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_153
timestamp 1666464484
transform 1 0 15180 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_161
timestamp 1666464484
transform 1 0 15916 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_166
timestamp 1666464484
transform 1 0 16376 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_173
timestamp 1666464484
transform 1 0 17020 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_180
timestamp 1666464484
transform 1 0 17664 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1666464484
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1666464484
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_197
timestamp 1666464484
transform 1 0 19228 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_204
timestamp 1666464484
transform 1 0 19872 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_212
timestamp 1666464484
transform 1 0 20608 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_234
timestamp 1666464484
transform 1 0 22632 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_243
timestamp 1666464484
transform 1 0 23460 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_250
timestamp 1666464484
transform 1 0 24104 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_253
timestamp 1666464484
transform 1 0 24380 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_271
timestamp 1666464484
transform 1 0 26036 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_291
timestamp 1666464484
transform 1 0 27876 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_306
timestamp 1666464484
transform 1 0 29256 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_309
timestamp 1666464484
transform 1 0 29532 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_327
timestamp 1666464484
transform 1 0 31188 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_335
timestamp 1666464484
transform 1 0 31924 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_347
timestamp 1666464484
transform 1 0 33028 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_358
timestamp 1666464484
transform 1 0 34040 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1666464484
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1666464484
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1666464484
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1666464484
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1666464484
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1666464484
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1666464484
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1666464484
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1666464484
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1666464484
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1666464484
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1666464484
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1666464484
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1666464484
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1666464484
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1666464484
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1666464484
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1666464484
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_169
timestamp 1666464484
transform 1 0 16652 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_175
timestamp 1666464484
transform 1 0 17204 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_192
timestamp 1666464484
transform 1 0 18768 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_212
timestamp 1666464484
transform 1 0 20608 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_222
timestamp 1666464484
transform 1 0 21528 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_225
timestamp 1666464484
transform 1 0 21804 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_232
timestamp 1666464484
transform 1 0 22448 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_49_256
timestamp 1666464484
transform 1 0 24656 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_268
timestamp 1666464484
transform 1 0 25760 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_278
timestamp 1666464484
transform 1 0 26680 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_281
timestamp 1666464484
transform 1 0 26956 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_285
timestamp 1666464484
transform 1 0 27324 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_295
timestamp 1666464484
transform 1 0 28244 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_319
timestamp 1666464484
transform 1 0 30452 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_325
timestamp 1666464484
transform 1 0 31004 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_334
timestamp 1666464484
transform 1 0 31832 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_337
timestamp 1666464484
transform 1 0 32108 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_345
timestamp 1666464484
transform 1 0 32844 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_349
timestamp 1666464484
transform 1 0 33212 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_356
timestamp 1666464484
transform 1 0 33856 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1666464484
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1666464484
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1666464484
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1666464484
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1666464484
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1666464484
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1666464484
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1666464484
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1666464484
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1666464484
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1666464484
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1666464484
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1666464484
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1666464484
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1666464484
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1666464484
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_153
timestamp 1666464484
transform 1 0 15180 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_161
timestamp 1666464484
transform 1 0 15916 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_167
timestamp 1666464484
transform 1 0 16468 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_172
timestamp 1666464484
transform 1 0 16928 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_176
timestamp 1666464484
transform 1 0 17296 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_182
timestamp 1666464484
transform 1 0 17848 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_194
timestamp 1666464484
transform 1 0 18952 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_197
timestamp 1666464484
transform 1 0 19228 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_210
timestamp 1666464484
transform 1 0 20424 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_230
timestamp 1666464484
transform 1 0 22264 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_239
timestamp 1666464484
transform 1 0 23092 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_248
timestamp 1666464484
transform 1 0 23920 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_253
timestamp 1666464484
transform 1 0 24380 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_263
timestamp 1666464484
transform 1 0 25300 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_274
timestamp 1666464484
transform 1 0 26312 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_50_290
timestamp 1666464484
transform 1 0 27784 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_298
timestamp 1666464484
transform 1 0 28520 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_306
timestamp 1666464484
transform 1 0 29256 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_309
timestamp 1666464484
transform 1 0 29532 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_318
timestamp 1666464484
transform 1 0 30360 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_325
timestamp 1666464484
transform 1 0 31004 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_345
timestamp 1666464484
transform 1 0 32844 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_355
timestamp 1666464484
transform 1 0 33764 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_362
timestamp 1666464484
transform 1 0 34408 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1666464484
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1666464484
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1666464484
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1666464484
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1666464484
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1666464484
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1666464484
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1666464484
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1666464484
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1666464484
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1666464484
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1666464484
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1666464484
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1666464484
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1666464484
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_149
timestamp 1666464484
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1666464484
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1666464484
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_169
timestamp 1666464484
transform 1 0 16652 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_177
timestamp 1666464484
transform 1 0 17388 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_181
timestamp 1666464484
transform 1 0 17756 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_201
timestamp 1666464484
transform 1 0 19596 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_51_221
timestamp 1666464484
transform 1 0 21436 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_51_225
timestamp 1666464484
transform 1 0 21804 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_243
timestamp 1666464484
transform 1 0 23460 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_252
timestamp 1666464484
transform 1 0 24288 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_256
timestamp 1666464484
transform 1 0 24656 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1666464484
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1666464484
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_281
timestamp 1666464484
transform 1 0 26956 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_51_303
timestamp 1666464484
transform 1 0 28980 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_309
timestamp 1666464484
transform 1 0 29532 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_317
timestamp 1666464484
transform 1 0 30268 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_328
timestamp 1666464484
transform 1 0 31280 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_337
timestamp 1666464484
transform 1 0 32108 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_342
timestamp 1666464484
transform 1 0 32568 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_362
timestamp 1666464484
transform 1 0 34408 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_3
timestamp 1666464484
transform 1 0 1380 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_9
timestamp 1666464484
transform 1 0 1932 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_13
timestamp 1666464484
transform 1 0 2300 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_25
timestamp 1666464484
transform 1 0 3404 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1666464484
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1666464484
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1666464484
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1666464484
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1666464484
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1666464484
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1666464484
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1666464484
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1666464484
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1666464484
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1666464484
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1666464484
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1666464484
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1666464484
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_165
timestamp 1666464484
transform 1 0 16284 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_176
timestamp 1666464484
transform 1 0 17296 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_185
timestamp 1666464484
transform 1 0 18124 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_194
timestamp 1666464484
transform 1 0 18952 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_197
timestamp 1666464484
transform 1 0 19228 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_204
timestamp 1666464484
transform 1 0 19872 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_208
timestamp 1666464484
transform 1 0 20240 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_225
timestamp 1666464484
transform 1 0 21804 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_235
timestamp 1666464484
transform 1 0 22724 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_250
timestamp 1666464484
transform 1 0 24104 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_253
timestamp 1666464484
transform 1 0 24380 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_260
timestamp 1666464484
transform 1 0 25024 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_268
timestamp 1666464484
transform 1 0 25760 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_291
timestamp 1666464484
transform 1 0 27876 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1666464484
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1666464484
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_309
timestamp 1666464484
transform 1 0 29532 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_318
timestamp 1666464484
transform 1 0 30360 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_329
timestamp 1666464484
transform 1 0 31372 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_335
timestamp 1666464484
transform 1 0 31924 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_352
timestamp 1666464484
transform 1 0 33488 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_52_361
timestamp 1666464484
transform 1 0 34316 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_3
timestamp 1666464484
transform 1 0 1380 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_28
timestamp 1666464484
transform 1 0 3680 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_40
timestamp 1666464484
transform 1 0 4784 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_52
timestamp 1666464484
transform 1 0 5888 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1666464484
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1666464484
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1666464484
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1666464484
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1666464484
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1666464484
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1666464484
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1666464484
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1666464484
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1666464484
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1666464484
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1666464484
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_169
timestamp 1666464484
transform 1 0 16652 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_176
timestamp 1666464484
transform 1 0 17296 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_183
timestamp 1666464484
transform 1 0 17940 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_203
timestamp 1666464484
transform 1 0 19780 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_211
timestamp 1666464484
transform 1 0 20516 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_220
timestamp 1666464484
transform 1 0 21344 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_53_225
timestamp 1666464484
transform 1 0 21804 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_244
timestamp 1666464484
transform 1 0 23552 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_251
timestamp 1666464484
transform 1 0 24196 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_271
timestamp 1666464484
transform 1 0 26036 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_278
timestamp 1666464484
transform 1 0 26680 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_281
timestamp 1666464484
transform 1 0 26956 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_299
timestamp 1666464484
transform 1 0 28612 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_323
timestamp 1666464484
transform 1 0 30820 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_334
timestamp 1666464484
transform 1 0 31832 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_337
timestamp 1666464484
transform 1 0 32108 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_362
timestamp 1666464484
transform 1 0 34408 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_3
timestamp 1666464484
transform 1 0 1380 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_7
timestamp 1666464484
transform 1 0 1748 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_11
timestamp 1666464484
transform 1 0 2116 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_23
timestamp 1666464484
transform 1 0 3220 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1666464484
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1666464484
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1666464484
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1666464484
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1666464484
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1666464484
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1666464484
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1666464484
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1666464484
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1666464484
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1666464484
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1666464484
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1666464484
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1666464484
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1666464484
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1666464484
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_180
timestamp 1666464484
transform 1 0 17664 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1666464484
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1666464484
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_197
timestamp 1666464484
transform 1 0 19228 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_54_208
timestamp 1666464484
transform 1 0 20240 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_214
timestamp 1666464484
transform 1 0 20792 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_231
timestamp 1666464484
transform 1 0 22356 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_241
timestamp 1666464484
transform 1 0 23276 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_250
timestamp 1666464484
transform 1 0 24104 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_253
timestamp 1666464484
transform 1 0 24380 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_261
timestamp 1666464484
transform 1 0 25116 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_270
timestamp 1666464484
transform 1 0 25944 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_276
timestamp 1666464484
transform 1 0 26496 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_293
timestamp 1666464484
transform 1 0 28060 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_297
timestamp 1666464484
transform 1 0 28428 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_304
timestamp 1666464484
transform 1 0 29072 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_309
timestamp 1666464484
transform 1 0 29532 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_316
timestamp 1666464484
transform 1 0 30176 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_328
timestamp 1666464484
transform 1 0 31280 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_336
timestamp 1666464484
transform 1 0 32016 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_356
timestamp 1666464484
transform 1 0 33856 0 1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1666464484
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1666464484
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1666464484
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1666464484
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1666464484
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1666464484
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1666464484
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1666464484
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1666464484
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1666464484
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1666464484
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1666464484
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1666464484
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1666464484
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1666464484
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1666464484
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1666464484
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1666464484
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1666464484
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_181
timestamp 1666464484
transform 1 0 17756 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_201
timestamp 1666464484
transform 1 0 19596 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_212
timestamp 1666464484
transform 1 0 20608 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_55_221
timestamp 1666464484
transform 1 0 21436 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_225
timestamp 1666464484
transform 1 0 21804 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_230
timestamp 1666464484
transform 1 0 22264 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_250
timestamp 1666464484
transform 1 0 24104 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_259
timestamp 1666464484
transform 1 0 24932 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_265
timestamp 1666464484
transform 1 0 25484 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_274
timestamp 1666464484
transform 1 0 26312 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_55_281
timestamp 1666464484
transform 1 0 26956 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_290
timestamp 1666464484
transform 1 0 27784 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_300
timestamp 1666464484
transform 1 0 28704 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_309
timestamp 1666464484
transform 1 0 29532 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_318
timestamp 1666464484
transform 1 0 30360 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_326
timestamp 1666464484
transform 1 0 31096 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_334
timestamp 1666464484
transform 1 0 31832 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_337
timestamp 1666464484
transform 1 0 32108 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_362
timestamp 1666464484
transform 1 0 34408 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_3
timestamp 1666464484
transform 1 0 1380 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_8
timestamp 1666464484
transform 1 0 1840 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_20
timestamp 1666464484
transform 1 0 2944 0 1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1666464484
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1666464484
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1666464484
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1666464484
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1666464484
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1666464484
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1666464484
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1666464484
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1666464484
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1666464484
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1666464484
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1666464484
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1666464484
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1666464484
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1666464484
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1666464484
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_189
timestamp 1666464484
transform 1 0 18492 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_194
timestamp 1666464484
transform 1 0 18952 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_56_197
timestamp 1666464484
transform 1 0 19228 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_216
timestamp 1666464484
transform 1 0 20976 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_225
timestamp 1666464484
transform 1 0 21804 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_233
timestamp 1666464484
transform 1 0 22540 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_240
timestamp 1666464484
transform 1 0 23184 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_250
timestamp 1666464484
transform 1 0 24104 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_56_253
timestamp 1666464484
transform 1 0 24380 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_261
timestamp 1666464484
transform 1 0 25116 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_281
timestamp 1666464484
transform 1 0 26956 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_289
timestamp 1666464484
transform 1 0 27692 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_306
timestamp 1666464484
transform 1 0 29256 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_309
timestamp 1666464484
transform 1 0 29532 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_316
timestamp 1666464484
transform 1 0 30176 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_320
timestamp 1666464484
transform 1 0 30544 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_328
timestamp 1666464484
transform 1 0 31280 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_332
timestamp 1666464484
transform 1 0 31648 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_350
timestamp 1666464484
transform 1 0 33304 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_359
timestamp 1666464484
transform 1 0 34132 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1666464484
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_3
timestamp 1666464484
transform 1 0 1380 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_9
timestamp 1666464484
transform 1 0 1932 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_13
timestamp 1666464484
transform 1 0 2300 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_20
timestamp 1666464484
transform 1 0 2944 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_32
timestamp 1666464484
transform 1 0 4048 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_44
timestamp 1666464484
transform 1 0 5152 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1666464484
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1666464484
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1666464484
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1666464484
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1666464484
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1666464484
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1666464484
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1666464484
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1666464484
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1666464484
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1666464484
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1666464484
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1666464484
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_181
timestamp 1666464484
transform 1 0 17756 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_201
timestamp 1666464484
transform 1 0 19596 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_214
timestamp 1666464484
transform 1 0 20792 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_222
timestamp 1666464484
transform 1 0 21528 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_225
timestamp 1666464484
transform 1 0 21804 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_243
timestamp 1666464484
transform 1 0 23460 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_250
timestamp 1666464484
transform 1 0 24104 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_270
timestamp 1666464484
transform 1 0 25944 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_278
timestamp 1666464484
transform 1 0 26680 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_281
timestamp 1666464484
transform 1 0 26956 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_286
timestamp 1666464484
transform 1 0 27416 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_306
timestamp 1666464484
transform 1 0 29256 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_312
timestamp 1666464484
transform 1 0 29808 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1666464484
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1666464484
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_337
timestamp 1666464484
transform 1 0 32108 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_362
timestamp 1666464484
transform 1 0 34408 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_3
timestamp 1666464484
transform 1 0 1380 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_10
timestamp 1666464484
transform 1 0 2024 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_23
timestamp 1666464484
transform 1 0 3220 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1666464484
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1666464484
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1666464484
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1666464484
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1666464484
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1666464484
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1666464484
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1666464484
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1666464484
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1666464484
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1666464484
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1666464484
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1666464484
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1666464484
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1666464484
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1666464484
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_177
timestamp 1666464484
transform 1 0 17388 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_186
timestamp 1666464484
transform 1 0 18216 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_190
timestamp 1666464484
transform 1 0 18584 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_194
timestamp 1666464484
transform 1 0 18952 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_58_197
timestamp 1666464484
transform 1 0 19228 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_203
timestamp 1666464484
transform 1 0 19780 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_211
timestamp 1666464484
transform 1 0 20516 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_231
timestamp 1666464484
transform 1 0 22356 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_235
timestamp 1666464484
transform 1 0 22724 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_243
timestamp 1666464484
transform 1 0 23460 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_250
timestamp 1666464484
transform 1 0 24104 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_253
timestamp 1666464484
transform 1 0 24380 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_271
timestamp 1666464484
transform 1 0 26036 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_291
timestamp 1666464484
transform 1 0 27876 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_302
timestamp 1666464484
transform 1 0 28888 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_58_309
timestamp 1666464484
transform 1 0 29532 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_327
timestamp 1666464484
transform 1 0 31188 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_337
timestamp 1666464484
transform 1 0 32108 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_362
timestamp 1666464484
transform 1 0 34408 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_3
timestamp 1666464484
transform 1 0 1380 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_28
timestamp 1666464484
transform 1 0 3680 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_40
timestamp 1666464484
transform 1 0 4784 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_52
timestamp 1666464484
transform 1 0 5888 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1666464484
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1666464484
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1666464484
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1666464484
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1666464484
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1666464484
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1666464484
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1666464484
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1666464484
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1666464484
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1666464484
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1666464484
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_169
timestamp 1666464484
transform 1 0 16652 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_193
timestamp 1666464484
transform 1 0 18860 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_213
timestamp 1666464484
transform 1 0 20700 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_222
timestamp 1666464484
transform 1 0 21528 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_225
timestamp 1666464484
transform 1 0 21804 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_243
timestamp 1666464484
transform 1 0 23460 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_263
timestamp 1666464484
transform 1 0 25300 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_272
timestamp 1666464484
transform 1 0 26128 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_281
timestamp 1666464484
transform 1 0 26956 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_299
timestamp 1666464484
transform 1 0 28612 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_303
timestamp 1666464484
transform 1 0 28980 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_309
timestamp 1666464484
transform 1 0 29532 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_315
timestamp 1666464484
transform 1 0 30084 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_332
timestamp 1666464484
transform 1 0 31648 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_337
timestamp 1666464484
transform 1 0 32108 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_362
timestamp 1666464484
transform 1 0 34408 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_3
timestamp 1666464484
transform 1 0 1380 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_26
timestamp 1666464484
transform 1 0 3496 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_29
timestamp 1666464484
transform 1 0 3772 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_43
timestamp 1666464484
transform 1 0 5060 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_55
timestamp 1666464484
transform 1 0 6164 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_67
timestamp 1666464484
transform 1 0 7268 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_79
timestamp 1666464484
transform 1 0 8372 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1666464484
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1666464484
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1666464484
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1666464484
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1666464484
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1666464484
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1666464484
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1666464484
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1666464484
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_165
timestamp 1666464484
transform 1 0 16284 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_173
timestamp 1666464484
transform 1 0 17020 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_181
timestamp 1666464484
transform 1 0 17756 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_190
timestamp 1666464484
transform 1 0 18584 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_60_197
timestamp 1666464484
transform 1 0 19228 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_204
timestamp 1666464484
transform 1 0 19872 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_215
timestamp 1666464484
transform 1 0 20884 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_224
timestamp 1666464484
transform 1 0 21712 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_233
timestamp 1666464484
transform 1 0 22540 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_243
timestamp 1666464484
transform 1 0 23460 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_250
timestamp 1666464484
transform 1 0 24104 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_253
timestamp 1666464484
transform 1 0 24380 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_271
timestamp 1666464484
transform 1 0 26036 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_280
timestamp 1666464484
transform 1 0 26864 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_304
timestamp 1666464484
transform 1 0 29072 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_309
timestamp 1666464484
transform 1 0 29532 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_316
timestamp 1666464484
transform 1 0 30176 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_320
timestamp 1666464484
transform 1 0 30544 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_337
timestamp 1666464484
transform 1 0 32108 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_362
timestamp 1666464484
transform 1 0 34408 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_3
timestamp 1666464484
transform 1 0 1380 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_17
timestamp 1666464484
transform 1 0 2668 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_33
timestamp 1666464484
transform 1 0 4140 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_49
timestamp 1666464484
transform 1 0 5612 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1666464484
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1666464484
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1666464484
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1666464484
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1666464484
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1666464484
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1666464484
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1666464484
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1666464484
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1666464484
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1666464484
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1666464484
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1666464484
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_169
timestamp 1666464484
transform 1 0 16652 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_177
timestamp 1666464484
transform 1 0 17388 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_181
timestamp 1666464484
transform 1 0 17756 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_201
timestamp 1666464484
transform 1 0 19596 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_208
timestamp 1666464484
transform 1 0 20240 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_219
timestamp 1666464484
transform 1 0 21252 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1666464484
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_61_225
timestamp 1666464484
transform 1 0 21804 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_61_233
timestamp 1666464484
transform 1 0 22540 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_241
timestamp 1666464484
transform 1 0 23276 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_258
timestamp 1666464484
transform 1 0 24840 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_267
timestamp 1666464484
transform 1 0 25668 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_276
timestamp 1666464484
transform 1 0 26496 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_281
timestamp 1666464484
transform 1 0 26956 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_288
timestamp 1666464484
transform 1 0 27600 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_297
timestamp 1666464484
transform 1 0 28428 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_301
timestamp 1666464484
transform 1 0 28796 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_307
timestamp 1666464484
transform 1 0 29348 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_316
timestamp 1666464484
transform 1 0 30176 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_325
timestamp 1666464484
transform 1 0 31004 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_334
timestamp 1666464484
transform 1 0 31832 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_61_337
timestamp 1666464484
transform 1 0 32108 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_345
timestamp 1666464484
transform 1 0 32844 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_354
timestamp 1666464484
transform 1 0 33672 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_362
timestamp 1666464484
transform 1 0 34408 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_3
timestamp 1666464484
transform 1 0 1380 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_10
timestamp 1666464484
transform 1 0 2024 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_26
timestamp 1666464484
transform 1 0 3496 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_29
timestamp 1666464484
transform 1 0 3772 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_43
timestamp 1666464484
transform 1 0 5060 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_59
timestamp 1666464484
transform 1 0 6532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_71
timestamp 1666464484
transform 1 0 7636 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1666464484
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1666464484
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1666464484
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1666464484
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1666464484
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1666464484
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1666464484
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1666464484
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1666464484
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1666464484
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_177
timestamp 1666464484
transform 1 0 17388 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_185
timestamp 1666464484
transform 1 0 18124 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1666464484
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1666464484
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_197
timestamp 1666464484
transform 1 0 19228 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_206
timestamp 1666464484
transform 1 0 20056 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_213
timestamp 1666464484
transform 1 0 20700 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_220
timestamp 1666464484
transform 1 0 21344 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_227
timestamp 1666464484
transform 1 0 21988 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_238
timestamp 1666464484
transform 1 0 23000 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_247
timestamp 1666464484
transform 1 0 23828 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1666464484
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_253
timestamp 1666464484
transform 1 0 24380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_62_258
timestamp 1666464484
transform 1 0 24840 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_266
timestamp 1666464484
transform 1 0 25576 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_272
timestamp 1666464484
transform 1 0 26128 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_281
timestamp 1666464484
transform 1 0 26956 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_290
timestamp 1666464484
transform 1 0 27784 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_297
timestamp 1666464484
transform 1 0 28428 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_301
timestamp 1666464484
transform 1 0 28796 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_306
timestamp 1666464484
transform 1 0 29256 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_62_309
timestamp 1666464484
transform 1 0 29532 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_317
timestamp 1666464484
transform 1 0 30268 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_326
timestamp 1666464484
transform 1 0 31096 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_335
timestamp 1666464484
transform 1 0 31924 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_62_362
timestamp 1666464484
transform 1 0 34408 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_3
timestamp 1666464484
transform 1 0 1380 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_28
timestamp 1666464484
transform 1 0 3680 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_44
timestamp 1666464484
transform 1 0 5152 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1666464484
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1666464484
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_57
timestamp 1666464484
transform 1 0 6348 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_62
timestamp 1666464484
transform 1 0 6808 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1666464484
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1666464484
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1666464484
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1666464484
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1666464484
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1666464484
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1666464484
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1666464484
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1666464484
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1666464484
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1666464484
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_169
timestamp 1666464484
transform 1 0 16652 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_180
timestamp 1666464484
transform 1 0 17664 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_187
timestamp 1666464484
transform 1 0 18308 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_194
timestamp 1666464484
transform 1 0 18952 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_201
timestamp 1666464484
transform 1 0 19596 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_208
timestamp 1666464484
transform 1 0 20240 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_213
timestamp 1666464484
transform 1 0 20700 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_217
timestamp 1666464484
transform 1 0 21068 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_222
timestamp 1666464484
transform 1 0 21528 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_225
timestamp 1666464484
transform 1 0 21804 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_232
timestamp 1666464484
transform 1 0 22448 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_241
timestamp 1666464484
transform 1 0 23276 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_248
timestamp 1666464484
transform 1 0 23920 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_255
timestamp 1666464484
transform 1 0 24564 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_262
timestamp 1666464484
transform 1 0 25208 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_266
timestamp 1666464484
transform 1 0 25576 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_270
timestamp 1666464484
transform 1 0 25944 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_278
timestamp 1666464484
transform 1 0 26680 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_281
timestamp 1666464484
transform 1 0 26956 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_286
timestamp 1666464484
transform 1 0 27416 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_293
timestamp 1666464484
transform 1 0 28060 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_300
timestamp 1666464484
transform 1 0 28704 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_307
timestamp 1666464484
transform 1 0 29348 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_319
timestamp 1666464484
transform 1 0 30452 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_328
timestamp 1666464484
transform 1 0 31280 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_337
timestamp 1666464484
transform 1 0 32108 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_362
timestamp 1666464484
transform 1 0 34408 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_3
timestamp 1666464484
transform 1 0 1380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_26
timestamp 1666464484
transform 1 0 3496 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_29
timestamp 1666464484
transform 1 0 3772 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_43
timestamp 1666464484
transform 1 0 5060 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_50
timestamp 1666464484
transform 1 0 5704 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_57
timestamp 1666464484
transform 1 0 6348 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_64
timestamp 1666464484
transform 1 0 6992 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_71
timestamp 1666464484
transform 1 0 7636 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_78
timestamp 1666464484
transform 1 0 8280 0 1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1666464484
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1666464484
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_109
timestamp 1666464484
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_121
timestamp 1666464484
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1666464484
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1666464484
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1666464484
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_153
timestamp 1666464484
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_165
timestamp 1666464484
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_180
timestamp 1666464484
transform 1 0 17664 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_187
timestamp 1666464484
transform 1 0 18308 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_194
timestamp 1666464484
transform 1 0 18952 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_197
timestamp 1666464484
transform 1 0 19228 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_208
timestamp 1666464484
transform 1 0 20240 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_215
timestamp 1666464484
transform 1 0 20884 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_222
timestamp 1666464484
transform 1 0 21528 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_229
timestamp 1666464484
transform 1 0 22172 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_236
timestamp 1666464484
transform 1 0 22816 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_243
timestamp 1666464484
transform 1 0 23460 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_250
timestamp 1666464484
transform 1 0 24104 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_64_253
timestamp 1666464484
transform 1 0 24380 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_259
timestamp 1666464484
transform 1 0 24932 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_266
timestamp 1666464484
transform 1 0 25576 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_277
timestamp 1666464484
transform 1 0 26588 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_281
timestamp 1666464484
transform 1 0 26956 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_285
timestamp 1666464484
transform 1 0 27324 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_291
timestamp 1666464484
transform 1 0 27876 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_295
timestamp 1666464484
transform 1 0 28244 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_306
timestamp 1666464484
transform 1 0 29256 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_309
timestamp 1666464484
transform 1 0 29532 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_319
timestamp 1666464484
transform 1 0 30452 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_328
timestamp 1666464484
transform 1 0 31280 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_337
timestamp 1666464484
transform 1 0 32108 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_362
timestamp 1666464484
transform 1 0 34408 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_65_3
timestamp 1666464484
transform 1 0 1380 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_17
timestamp 1666464484
transform 1 0 2668 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_42
timestamp 1666464484
transform 1 0 4968 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_46
timestamp 1666464484
transform 1 0 5336 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_65_50
timestamp 1666464484
transform 1 0 5704 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_65_57
timestamp 1666464484
transform 1 0 6348 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_65_68
timestamp 1666464484
transform 1 0 7360 0 -1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_65_95
timestamp 1666464484
transform 1 0 9844 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_107
timestamp 1666464484
transform 1 0 10948 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1666464484
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_113
timestamp 1666464484
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_125
timestamp 1666464484
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_137
timestamp 1666464484
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_149
timestamp 1666464484
transform 1 0 14812 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_155
timestamp 1666464484
transform 1 0 15364 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_159
timestamp 1666464484
transform 1 0 15732 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_166
timestamp 1666464484
transform 1 0 16376 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_65_169
timestamp 1666464484
transform 1 0 16652 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_175
timestamp 1666464484
transform 1 0 17204 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_182
timestamp 1666464484
transform 1 0 17848 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_190
timestamp 1666464484
transform 1 0 18584 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_195
timestamp 1666464484
transform 1 0 19044 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_202
timestamp 1666464484
transform 1 0 19688 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_209
timestamp 1666464484
transform 1 0 20332 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_217
timestamp 1666464484
transform 1 0 21068 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_222
timestamp 1666464484
transform 1 0 21528 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_65_225
timestamp 1666464484
transform 1 0 21804 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_231
timestamp 1666464484
transform 1 0 22356 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_235
timestamp 1666464484
transform 1 0 22724 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_242
timestamp 1666464484
transform 1 0 23368 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_249
timestamp 1666464484
transform 1 0 24012 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_256
timestamp 1666464484
transform 1 0 24656 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_263
timestamp 1666464484
transform 1 0 25300 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_269
timestamp 1666464484
transform 1 0 25852 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_65_273
timestamp 1666464484
transform 1 0 26220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1666464484
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_281
timestamp 1666464484
transform 1 0 26956 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_286
timestamp 1666464484
transform 1 0 27416 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_293
timestamp 1666464484
transform 1 0 28060 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_297
timestamp 1666464484
transform 1 0 28428 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_319
timestamp 1666464484
transform 1 0 30452 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_327
timestamp 1666464484
transform 1 0 31188 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_334
timestamp 1666464484
transform 1 0 31832 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_337
timestamp 1666464484
transform 1 0 32108 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_362
timestamp 1666464484
transform 1 0 34408 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_3
timestamp 1666464484
transform 1 0 1380 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_26
timestamp 1666464484
transform 1 0 3496 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_29
timestamp 1666464484
transform 1 0 3772 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_34
timestamp 1666464484
transform 1 0 4232 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_41
timestamp 1666464484
transform 1 0 4876 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_66_50
timestamp 1666464484
transform 1 0 5704 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_57
timestamp 1666464484
transform 1 0 6348 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_82
timestamp 1666464484
transform 1 0 8648 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_85
timestamp 1666464484
transform 1 0 8924 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_90
timestamp 1666464484
transform 1 0 9384 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_97
timestamp 1666464484
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_109
timestamp 1666464484
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_121
timestamp 1666464484
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1666464484
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1666464484
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_141
timestamp 1666464484
transform 1 0 14076 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_66_146
timestamp 1666464484
transform 1 0 14536 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_66_155
timestamp 1666464484
transform 1 0 15364 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_162
timestamp 1666464484
transform 1 0 16008 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_187
timestamp 1666464484
transform 1 0 18308 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_194
timestamp 1666464484
transform 1 0 18952 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_66_197
timestamp 1666464484
transform 1 0 19228 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_66_226
timestamp 1666464484
transform 1 0 21896 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_233
timestamp 1666464484
transform 1 0 22540 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_239
timestamp 1666464484
transform 1 0 23092 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_243
timestamp 1666464484
transform 1 0 23460 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_250
timestamp 1666464484
transform 1 0 24104 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_66_253
timestamp 1666464484
transform 1 0 24380 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_66_280
timestamp 1666464484
transform 1 0 26864 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_287
timestamp 1666464484
transform 1 0 27508 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_291
timestamp 1666464484
transform 1 0 27876 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_295
timestamp 1666464484
transform 1 0 28244 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_302
timestamp 1666464484
transform 1 0 28888 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_66_309
timestamp 1666464484
transform 1 0 29532 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_66_333
timestamp 1666464484
transform 1 0 31740 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_362
timestamp 1666464484
transform 1 0 34408 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_3
timestamp 1666464484
transform 1 0 1380 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_28
timestamp 1666464484
transform 1 0 3680 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_32
timestamp 1666464484
transform 1 0 4048 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_54
timestamp 1666464484
transform 1 0 6072 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_67_57
timestamp 1666464484
transform 1 0 6348 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_67_68
timestamp 1666464484
transform 1 0 7360 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_75
timestamp 1666464484
transform 1 0 8004 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_100
timestamp 1666464484
transform 1 0 10304 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_107
timestamp 1666464484
transform 1 0 10948 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1666464484
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_113
timestamp 1666464484
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_125
timestamp 1666464484
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_137
timestamp 1666464484
transform 1 0 13708 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_141
timestamp 1666464484
transform 1 0 14076 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_166
timestamp 1666464484
transform 1 0 16376 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_169
timestamp 1666464484
transform 1 0 16652 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_192
timestamp 1666464484
transform 1 0 18768 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1666464484
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1666464484
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_225
timestamp 1666464484
transform 1 0 21804 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_248
timestamp 1666464484
transform 1 0 23920 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_252
timestamp 1666464484
transform 1 0 24288 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_67_274
timestamp 1666464484
transform 1 0 26312 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_67_281
timestamp 1666464484
transform 1 0 26956 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_304
timestamp 1666464484
transform 1 0 29072 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_329
timestamp 1666464484
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1666464484
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_67_337
timestamp 1666464484
transform 1 0 32108 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_67_361
timestamp 1666464484
transform 1 0 34316 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_68_3
timestamp 1666464484
transform 1 0 1380 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_26
timestamp 1666464484
transform 1 0 3496 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_29
timestamp 1666464484
transform 1 0 3772 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_68_34
timestamp 1666464484
transform 1 0 4232 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_42
timestamp 1666464484
transform 1 0 4968 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_47
timestamp 1666464484
transform 1 0 5428 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_54
timestamp 1666464484
transform 1 0 6072 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_57
timestamp 1666464484
transform 1 0 6348 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_80
timestamp 1666464484
transform 1 0 8464 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_85
timestamp 1666464484
transform 1 0 8924 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_90
timestamp 1666464484
transform 1 0 9384 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_97
timestamp 1666464484
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_109
timestamp 1666464484
transform 1 0 11132 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_113
timestamp 1666464484
transform 1 0 11500 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_125
timestamp 1666464484
transform 1 0 12604 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_68_133
timestamp 1666464484
transform 1 0 13340 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_138
timestamp 1666464484
transform 1 0 13800 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_141
timestamp 1666464484
transform 1 0 14076 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_164
timestamp 1666464484
transform 1 0 16192 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_169
timestamp 1666464484
transform 1 0 16652 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_174
timestamp 1666464484
transform 1 0 17112 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_178
timestamp 1666464484
transform 1 0 17480 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_182
timestamp 1666464484
transform 1 0 17848 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_190
timestamp 1666464484
transform 1 0 18584 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_194
timestamp 1666464484
transform 1 0 18952 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_197
timestamp 1666464484
transform 1 0 19228 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_202
timestamp 1666464484
transform 1 0 19688 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_209
timestamp 1666464484
transform 1 0 20332 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_217
timestamp 1666464484
transform 1 0 21068 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_222
timestamp 1666464484
transform 1 0 21528 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_225
timestamp 1666464484
transform 1 0 21804 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_232
timestamp 1666464484
transform 1 0 22448 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_68_243
timestamp 1666464484
transform 1 0 23460 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_250
timestamp 1666464484
transform 1 0 24104 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_253
timestamp 1666464484
transform 1 0 24380 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_258
timestamp 1666464484
transform 1 0 24840 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_265
timestamp 1666464484
transform 1 0 25484 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_272
timestamp 1666464484
transform 1 0 26128 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_68_281
timestamp 1666464484
transform 1 0 26956 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_68_287
timestamp 1666464484
transform 1 0 27508 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_294
timestamp 1666464484
transform 1 0 28152 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_301
timestamp 1666464484
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1666464484
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_309
timestamp 1666464484
transform 1 0 29532 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_314
timestamp 1666464484
transform 1 0 29992 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_321
timestamp 1666464484
transform 1 0 30636 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_328
timestamp 1666464484
transform 1 0 31280 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_68_337
timestamp 1666464484
transform 1 0 32108 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_362
timestamp 1666464484
transform 1 0 34408 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1666464484
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1666464484
transform -1 0 34868 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1666464484
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1666464484
transform -1 0 34868 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1666464484
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1666464484
transform -1 0 34868 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1666464484
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1666464484
transform -1 0 34868 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1666464484
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1666464484
transform -1 0 34868 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1666464484
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1666464484
transform -1 0 34868 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1666464484
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1666464484
transform -1 0 34868 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1666464484
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1666464484
transform -1 0 34868 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1666464484
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1666464484
transform -1 0 34868 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1666464484
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1666464484
transform -1 0 34868 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1666464484
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1666464484
transform -1 0 34868 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1666464484
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1666464484
transform -1 0 34868 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1666464484
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1666464484
transform -1 0 34868 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1666464484
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1666464484
transform -1 0 34868 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1666464484
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1666464484
transform -1 0 34868 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1666464484
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1666464484
transform -1 0 34868 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1666464484
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1666464484
transform -1 0 34868 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1666464484
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1666464484
transform -1 0 34868 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1666464484
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1666464484
transform -1 0 34868 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1666464484
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1666464484
transform -1 0 34868 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1666464484
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1666464484
transform -1 0 34868 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1666464484
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1666464484
transform -1 0 34868 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1666464484
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1666464484
transform -1 0 34868 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1666464484
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1666464484
transform -1 0 34868 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1666464484
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1666464484
transform -1 0 34868 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1666464484
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1666464484
transform -1 0 34868 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1666464484
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1666464484
transform -1 0 34868 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1666464484
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1666464484
transform -1 0 34868 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1666464484
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1666464484
transform -1 0 34868 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1666464484
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1666464484
transform -1 0 34868 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1666464484
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1666464484
transform -1 0 34868 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1666464484
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1666464484
transform -1 0 34868 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1666464484
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1666464484
transform -1 0 34868 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1666464484
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1666464484
transform -1 0 34868 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1666464484
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1666464484
transform -1 0 34868 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1666464484
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1666464484
transform -1 0 34868 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1666464484
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1666464484
transform -1 0 34868 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1666464484
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1666464484
transform -1 0 34868 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1666464484
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1666464484
transform -1 0 34868 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1666464484
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1666464484
transform -1 0 34868 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1666464484
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1666464484
transform -1 0 34868 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1666464484
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1666464484
transform -1 0 34868 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1666464484
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1666464484
transform -1 0 34868 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1666464484
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1666464484
transform -1 0 34868 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1666464484
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1666464484
transform -1 0 34868 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1666464484
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1666464484
transform -1 0 34868 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1666464484
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1666464484
transform -1 0 34868 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1666464484
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1666464484
transform -1 0 34868 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1666464484
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1666464484
transform -1 0 34868 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1666464484
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1666464484
transform -1 0 34868 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1666464484
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1666464484
transform -1 0 34868 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1666464484
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1666464484
transform -1 0 34868 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1666464484
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1666464484
transform -1 0 34868 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1666464484
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1666464484
transform -1 0 34868 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1666464484
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1666464484
transform -1 0 34868 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1666464484
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1666464484
transform -1 0 34868 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1666464484
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1666464484
transform -1 0 34868 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1666464484
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1666464484
transform -1 0 34868 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1666464484
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1666464484
transform -1 0 34868 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1666464484
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1666464484
transform -1 0 34868 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1666464484
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1666464484
transform -1 0 34868 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1666464484
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1666464484
transform -1 0 34868 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1666464484
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1666464484
transform -1 0 34868 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1666464484
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1666464484
transform -1 0 34868 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1666464484
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1666464484
transform -1 0 34868 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1666464484
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1666464484
transform -1 0 34868 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1666464484
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1666464484
transform -1 0 34868 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1666464484
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1666464484
transform -1 0 34868 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1666464484
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1666464484
transform -1 0 34868 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1666464484
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1666464484
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1666464484
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1666464484
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1666464484
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1666464484
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1666464484
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1666464484
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1666464484
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1666464484
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1666464484
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1666464484
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1666464484
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1666464484
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1666464484
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1666464484
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1666464484
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1666464484
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1666464484
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1666464484
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1666464484
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1666464484
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1666464484
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1666464484
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1666464484
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1666464484
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1666464484
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1666464484
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1666464484
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1666464484
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1666464484
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1666464484
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1666464484
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1666464484
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1666464484
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1666464484
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1666464484
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1666464484
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1666464484
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1666464484
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1666464484
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1666464484
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1666464484
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1666464484
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1666464484
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1666464484
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1666464484
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1666464484
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1666464484
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1666464484
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1666464484
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1666464484
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1666464484
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1666464484
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1666464484
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1666464484
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1666464484
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1666464484
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1666464484
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1666464484
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1666464484
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1666464484
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1666464484
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1666464484
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1666464484
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1666464484
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1666464484
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1666464484
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1666464484
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1666464484
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1666464484
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1666464484
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1666464484
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1666464484
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1666464484
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1666464484
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1666464484
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1666464484
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1666464484
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1666464484
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1666464484
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1666464484
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1666464484
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1666464484
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1666464484
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1666464484
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1666464484
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1666464484
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1666464484
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1666464484
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1666464484
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1666464484
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1666464484
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1666464484
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1666464484
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1666464484
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1666464484
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1666464484
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1666464484
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1666464484
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1666464484
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1666464484
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1666464484
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1666464484
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1666464484
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1666464484
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1666464484
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1666464484
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1666464484
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1666464484
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1666464484
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1666464484
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1666464484
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1666464484
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1666464484
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1666464484
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1666464484
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1666464484
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1666464484
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1666464484
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1666464484
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1666464484
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1666464484
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1666464484
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1666464484
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1666464484
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1666464484
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1666464484
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1666464484
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1666464484
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1666464484
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1666464484
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1666464484
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1666464484
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1666464484
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1666464484
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1666464484
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1666464484
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1666464484
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1666464484
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1666464484
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1666464484
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1666464484
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1666464484
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1666464484
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1666464484
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1666464484
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1666464484
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1666464484
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1666464484
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1666464484
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1666464484
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1666464484
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1666464484
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1666464484
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1666464484
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1666464484
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1666464484
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1666464484
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1666464484
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1666464484
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1666464484
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1666464484
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1666464484
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1666464484
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1666464484
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1666464484
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1666464484
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1666464484
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1666464484
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1666464484
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1666464484
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1666464484
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1666464484
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1666464484
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1666464484
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1666464484
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1666464484
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1666464484
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1666464484
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1666464484
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1666464484
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1666464484
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1666464484
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1666464484
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1666464484
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1666464484
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1666464484
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1666464484
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1666464484
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1666464484
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1666464484
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1666464484
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1666464484
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1666464484
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1666464484
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1666464484
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1666464484
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1666464484
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1666464484
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1666464484
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1666464484
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1666464484
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1666464484
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1666464484
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1666464484
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1666464484
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1666464484
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1666464484
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1666464484
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1666464484
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1666464484
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1666464484
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1666464484
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1666464484
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1666464484
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1666464484
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1666464484
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1666464484
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1666464484
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1666464484
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1666464484
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1666464484
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1666464484
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1666464484
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1666464484
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1666464484
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1666464484
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1666464484
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1666464484
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1666464484
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1666464484
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1666464484
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1666464484
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1666464484
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1666464484
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1666464484
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1666464484
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1666464484
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1666464484
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1666464484
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1666464484
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1666464484
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1666464484
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1666464484
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1666464484
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1666464484
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1666464484
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1666464484
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1666464484
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1666464484
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1666464484
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1666464484
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1666464484
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1666464484
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1666464484
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1666464484
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1666464484
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1666464484
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1666464484
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1666464484
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1666464484
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1666464484
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1666464484
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1666464484
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1666464484
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1666464484
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1666464484
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1666464484
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1666464484
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1666464484
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1666464484
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1666464484
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1666464484
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1666464484
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1666464484
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1666464484
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1666464484
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1666464484
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1666464484
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1666464484
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1666464484
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1666464484
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1666464484
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1666464484
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1666464484
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1666464484
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1666464484
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1666464484
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1666464484
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1666464484
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1666464484
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1666464484
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1666464484
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1666464484
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1666464484
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1666464484
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1666464484
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1666464484
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1666464484
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1666464484
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1666464484
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1666464484
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1666464484
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1666464484
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1666464484
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1666464484
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1666464484
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1666464484
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1666464484
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1666464484
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1666464484
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1666464484
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1666464484
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1666464484
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1666464484
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1666464484
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1666464484
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1666464484
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1666464484
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1666464484
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1666464484
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1666464484
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1666464484
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1666464484
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1666464484
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1666464484
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1666464484
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1666464484
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1666464484
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1666464484
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1666464484
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1666464484
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1666464484
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1666464484
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1666464484
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1666464484
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1666464484
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1666464484
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1666464484
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1666464484
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1666464484
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1666464484
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1666464484
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1666464484
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1666464484
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1666464484
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1666464484
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1666464484
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1666464484
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1666464484
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1666464484
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1666464484
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1666464484
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1666464484
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1666464484
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1666464484
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1666464484
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1666464484
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1666464484
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1666464484
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1666464484
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1666464484
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1666464484
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1666464484
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1666464484
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1666464484
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1666464484
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1666464484
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1666464484
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1666464484
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1666464484
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1666464484
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1666464484
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1666464484
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1666464484
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1666464484
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1666464484
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1666464484
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1666464484
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1666464484
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1666464484
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1666464484
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1666464484
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1666464484
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1666464484
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1666464484
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1666464484
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1666464484
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1666464484
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1666464484
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1666464484
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1666464484
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1666464484
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1666464484
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1666464484
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1666464484
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1666464484
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1666464484
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1666464484
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1666464484
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1666464484
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1666464484
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1666464484
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1666464484
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1666464484
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1666464484
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1666464484
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1666464484
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1666464484
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1666464484
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1666464484
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1666464484
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1666464484
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1666464484
transform 1 0 6256 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1666464484
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1666464484
transform 1 0 11408 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1666464484
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1666464484
transform 1 0 16560 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1666464484
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1666464484
transform 1 0 21712 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1666464484
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1666464484
transform 1 0 26864 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1666464484
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1666464484
transform 1 0 32016 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_8  _0668_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1656 0 -1 38080
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_8  _0669_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1564 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  _0670_
timestamp 1666464484
transform 1 0 2392 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0671_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 6532 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0672_
timestamp 1666464484
transform 1 0 2024 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0673_
timestamp 1666464484
transform 1 0 15640 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0674_
timestamp 1666464484
transform 1 0 2024 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0675_
timestamp 1666464484
transform 1 0 22540 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0676_
timestamp 1666464484
transform 1 0 19320 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0677_
timestamp 1666464484
transform 1 0 31188 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0678_
timestamp 1666464484
transform 1 0 6532 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0679_
timestamp 1666464484
transform 1 0 16928 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0680_
timestamp 1666464484
transform 1 0 31556 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0681_
timestamp 1666464484
transform 1 0 9108 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0682_
timestamp 1666464484
transform 1 0 21252 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0683_
timestamp 1666464484
transform 1 0 7544 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0684_
timestamp 1666464484
transform 1 0 7360 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0685_
timestamp 1666464484
transform 1 0 17572 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0686_
timestamp 1666464484
transform 1 0 7176 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0687_
timestamp 1666464484
transform 1 0 31096 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0688_
timestamp 1666464484
transform 1 0 27968 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0689_
timestamp 1666464484
transform 1 0 7176 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0690_
timestamp 1666464484
transform 1 0 30268 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0691_
timestamp 1666464484
transform 1 0 2484 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0692_
timestamp 1666464484
transform 1 0 4048 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0693_
timestamp 1666464484
transform 1 0 33120 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0694_
timestamp 1666464484
transform 1 0 5244 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0695_
timestamp 1666464484
transform 1 0 3956 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0696_
timestamp 1666464484
transform 1 0 30912 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0697_
timestamp 1666464484
transform 1 0 27692 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0698_
timestamp 1666464484
transform 1 0 9108 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0699_
timestamp 1666464484
transform 1 0 5612 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0700_
timestamp 1666464484
transform 1 0 20056 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0701_
timestamp 1666464484
transform 1 0 33120 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0702_
timestamp 1666464484
transform 1 0 20608 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0703_
timestamp 1666464484
transform 1 0 3956 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0704_
timestamp 1666464484
transform 1 0 22172 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0705_
timestamp 1666464484
transform 1 0 4968 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0706_
timestamp 1666464484
transform 1 0 1748 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0707_
timestamp 1666464484
transform 1 0 15272 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0708_
timestamp 1666464484
transform 1 0 14260 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0709_
timestamp 1666464484
transform 1 0 21252 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0710_
timestamp 1666464484
transform 1 0 3956 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0711_
timestamp 1666464484
transform 1 0 4600 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0712_
timestamp 1666464484
transform 1 0 28980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0713_
timestamp 1666464484
transform 1 0 29256 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0714_
timestamp 1666464484
transform 1 0 4508 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0715_
timestamp 1666464484
transform 1 0 27048 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0716_
timestamp 1666464484
transform 1 0 2024 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0717_
timestamp 1666464484
transform 1 0 6532 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0718_
timestamp 1666464484
transform 1 0 14352 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0719_
timestamp 1666464484
transform 1 0 31740 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0720_
timestamp 1666464484
transform 1 0 23828 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0721_
timestamp 1666464484
transform 1 0 28336 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0722_
timestamp 1666464484
transform 1 0 2024 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0723_
timestamp 1666464484
transform 1 0 28520 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0724_
timestamp 1666464484
transform 1 0 2024 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0725_
timestamp 1666464484
transform 1 0 3956 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0726_
timestamp 1666464484
transform 1 0 23828 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0727_
timestamp 1666464484
transform 1 0 31188 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0728_
timestamp 1666464484
transform 1 0 33948 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0729_
timestamp 1666464484
transform 1 0 13156 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0730_
timestamp 1666464484
transform 1 0 4600 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0731_
timestamp 1666464484
transform 1 0 27140 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0732_
timestamp 1666464484
transform 1 0 1932 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0733_
timestamp 1666464484
transform 1 0 6532 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0734_
timestamp 1666464484
transform 1 0 5520 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0735_
timestamp 1666464484
transform 1 0 25024 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0736_
timestamp 1666464484
transform 1 0 3956 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0737_
timestamp 1666464484
transform 1 0 33764 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0738_
timestamp 1666464484
transform 1 0 25300 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0739_
timestamp 1666464484
transform 1 0 23736 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0740_
timestamp 1666464484
transform 1 0 9108 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0741_
timestamp 1666464484
transform 1 0 22448 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0742_
timestamp 1666464484
transform 1 0 28980 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0743_
timestamp 1666464484
transform 1 0 18676 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0744_
timestamp 1666464484
transform 1 0 19412 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0745_
timestamp 1666464484
transform 1 0 8004 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0746_
timestamp 1666464484
transform 1 0 6900 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0747_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2392 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0748_
timestamp 1666464484
transform 1 0 2024 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0749_
timestamp 1666464484
transform 1 0 5428 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0750_
timestamp 1666464484
transform 1 0 17480 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0751_
timestamp 1666464484
transform 1 0 29900 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0752_
timestamp 1666464484
transform 1 0 33764 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0753_
timestamp 1666464484
transform 1 0 2024 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0754_
timestamp 1666464484
transform 1 0 30912 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0755_
timestamp 1666464484
transform 1 0 2668 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0756_
timestamp 1666464484
transform 1 0 7084 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0757_
timestamp 1666464484
transform 1 0 31556 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0758_
timestamp 1666464484
transform 1 0 3036 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0759_
timestamp 1666464484
transform 1 0 10488 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0760_
timestamp 1666464484
transform 1 0 24564 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0761_
timestamp 1666464484
transform 1 0 7084 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0762_
timestamp 1666464484
transform 1 0 32292 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0763_
timestamp 1666464484
transform 1 0 3956 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0764_
timestamp 1666464484
transform 1 0 4692 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0765_
timestamp 1666464484
transform 1 0 15088 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0766_
timestamp 1666464484
transform 1 0 16836 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0767_
timestamp 1666464484
transform 1 0 28336 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0768_
timestamp 1666464484
transform 1 0 27692 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0769_
timestamp 1666464484
transform 1 0 5428 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0770_
timestamp 1666464484
transform 1 0 23092 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0771_
timestamp 1666464484
transform 1 0 2116 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0772_
timestamp 1666464484
transform 1 0 21988 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0773_
timestamp 1666464484
transform 1 0 31832 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0774_
timestamp 1666464484
transform 1 0 24656 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0775_
timestamp 1666464484
transform 1 0 18676 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0776_
timestamp 1666464484
transform 1 0 28336 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0777_
timestamp 1666464484
transform 1 0 17388 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0778_
timestamp 1666464484
transform 1 0 6532 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0779_
timestamp 1666464484
transform 1 0 28980 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0780_
timestamp 1666464484
transform 1 0 2024 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0781_
timestamp 1666464484
transform 1 0 29900 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0782_
timestamp 1666464484
transform 1 0 5428 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0783_
timestamp 1666464484
transform 1 0 2484 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0784_
timestamp 1666464484
transform 1 0 2484 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0785_
timestamp 1666464484
transform 1 0 2760 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0786_
timestamp 1666464484
transform 1 0 19964 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0787_
timestamp 1666464484
transform 1 0 24380 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0788_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 24564 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0789_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 26312 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _0790_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 27324 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0791_
timestamp 1666464484
transform 1 0 27968 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0792_
timestamp 1666464484
transform 1 0 27140 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0793_
timestamp 1666464484
transform 1 0 27324 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0794_
timestamp 1666464484
transform 1 0 25116 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0795_
timestamp 1666464484
transform 1 0 24748 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0796_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 25852 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0797_
timestamp 1666464484
transform 1 0 25944 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0798_
timestamp 1666464484
transform 1 0 26036 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0799_
timestamp 1666464484
transform 1 0 26036 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0800_
timestamp 1666464484
transform 1 0 19412 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0801_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 25392 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0802_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28888 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0803_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 26036 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0804_
timestamp 1666464484
transform 1 0 26036 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0805_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 25116 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0806_
timestamp 1666464484
transform 1 0 27140 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0807_
timestamp 1666464484
transform 1 0 25760 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _0808_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 26680 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0809_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 27324 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0810_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28612 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0811_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 33580 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0812_
timestamp 1666464484
transform 1 0 21988 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0813_
timestamp 1666464484
transform 1 0 23828 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0814_
timestamp 1666464484
transform 1 0 23000 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0815_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 21988 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0816_
timestamp 1666464484
transform 1 0 19780 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0817_
timestamp 1666464484
transform 1 0 24380 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0818_
timestamp 1666464484
transform 1 0 21252 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0819_
timestamp 1666464484
transform 1 0 17664 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0820_
timestamp 1666464484
transform 1 0 21252 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0821_
timestamp 1666464484
transform 1 0 20332 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0822_
timestamp 1666464484
transform 1 0 20148 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0823_
timestamp 1666464484
transform 1 0 22908 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0824_
timestamp 1666464484
transform 1 0 20332 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0825_
timestamp 1666464484
transform 1 0 20608 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0826_
timestamp 1666464484
transform 1 0 21988 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0827_
timestamp 1666464484
transform 1 0 23000 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0828_
timestamp 1666464484
transform 1 0 22724 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _0829_
timestamp 1666464484
transform 1 0 23828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _0830_
timestamp 1666464484
transform 1 0 20700 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0831_
timestamp 1666464484
transform 1 0 21620 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0832_
timestamp 1666464484
transform 1 0 21804 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0833_
timestamp 1666464484
transform 1 0 8740 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0834_
timestamp 1666464484
transform 1 0 30636 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0835_
timestamp 1666464484
transform 1 0 32292 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0836_
timestamp 1666464484
transform 1 0 31372 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0837_
timestamp 1666464484
transform 1 0 33764 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0838_
timestamp 1666464484
transform 1 0 32936 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0839_
timestamp 1666464484
transform 1 0 32936 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0840_
timestamp 1666464484
transform 1 0 31556 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0841_
timestamp 1666464484
transform 1 0 31924 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0842_
timestamp 1666464484
transform 1 0 31280 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0843_
timestamp 1666464484
transform 1 0 31096 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0844_
timestamp 1666464484
transform 1 0 15916 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0845_
timestamp 1666464484
transform 1 0 30452 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0846_
timestamp 1666464484
transform 1 0 32016 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0847_
timestamp 1666464484
transform 1 0 30268 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0848_
timestamp 1666464484
transform 1 0 32292 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0849_
timestamp 1666464484
transform 1 0 31556 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0850_
timestamp 1666464484
transform 1 0 33304 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0851_
timestamp 1666464484
transform 1 0 33304 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _0852_
timestamp 1666464484
transform 1 0 31280 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0853_
timestamp 1666464484
transform 1 0 31004 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0854_
timestamp 1666464484
transform 1 0 30268 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0855_
timestamp 1666464484
transform 1 0 16100 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0856_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 24564 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0857_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 25116 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0858_
timestamp 1666464484
transform 1 0 24564 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0859_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 20056 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0860_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 23552 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0861_
timestamp 1666464484
transform 1 0 23736 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0862_
timestamp 1666464484
transform 1 0 24932 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0863_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 24564 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0864_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 25668 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _0865_
timestamp 1666464484
transform 1 0 23552 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0866_
timestamp 1666464484
transform 1 0 23736 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0867_
timestamp 1666464484
transform 1 0 23828 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0868_
timestamp 1666464484
transform 1 0 23644 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0869_
timestamp 1666464484
transform 1 0 23460 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0870_
timestamp 1666464484
transform 1 0 25300 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0871_
timestamp 1666464484
transform 1 0 24840 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0872_
timestamp 1666464484
transform 1 0 25300 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0873_
timestamp 1666464484
transform 1 0 26128 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0874_
timestamp 1666464484
transform 1 0 26036 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0875_
timestamp 1666464484
transform 1 0 26588 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0876_
timestamp 1666464484
transform 1 0 26588 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0877_
timestamp 1666464484
transform 1 0 26128 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0878_
timestamp 1666464484
transform 1 0 19228 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0879_
timestamp 1666464484
transform 1 0 21160 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0880_
timestamp 1666464484
transform 1 0 20240 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0881_
timestamp 1666464484
transform 1 0 20608 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0882_
timestamp 1666464484
transform 1 0 21528 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0883_
timestamp 1666464484
transform 1 0 20608 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0884_
timestamp 1666464484
transform 1 0 21988 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0885_
timestamp 1666464484
transform 1 0 22080 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0886_
timestamp 1666464484
transform 1 0 21620 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0887_
timestamp 1666464484
transform 1 0 22356 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0888_
timestamp 1666464484
transform 1 0 22264 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0889_
timestamp 1666464484
transform 1 0 23000 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0890_
timestamp 1666464484
transform 1 0 23828 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0891_
timestamp 1666464484
transform 1 0 25760 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0892_
timestamp 1666464484
transform 1 0 22908 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0893_
timestamp 1666464484
transform 1 0 19504 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0894_
timestamp 1666464484
transform 1 0 23736 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0895_
timestamp 1666464484
transform 1 0 22908 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0896_
timestamp 1666464484
transform 1 0 25668 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0897_
timestamp 1666464484
transform 1 0 24564 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0898_
timestamp 1666464484
transform 1 0 30636 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0899_
timestamp 1666464484
transform 1 0 21160 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0900_
timestamp 1666464484
transform 1 0 31556 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0901_
timestamp 1666464484
transform 1 0 32292 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0902_
timestamp 1666464484
transform 1 0 31648 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0903_
timestamp 1666464484
transform 1 0 33028 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0904_
timestamp 1666464484
transform 1 0 30544 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0905_
timestamp 1666464484
transform 1 0 33764 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0906_
timestamp 1666464484
transform 1 0 32568 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0907_
timestamp 1666464484
transform 1 0 31648 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0908_
timestamp 1666464484
transform 1 0 31004 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0909_
timestamp 1666464484
transform 1 0 31464 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0910_
timestamp 1666464484
transform 1 0 31556 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0911_
timestamp 1666464484
transform 1 0 33672 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0912_
timestamp 1666464484
transform 1 0 31096 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0913_
timestamp 1666464484
transform 1 0 30268 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0914_
timestamp 1666464484
transform 1 0 33672 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0915_
timestamp 1666464484
transform 1 0 31464 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0916_
timestamp 1666464484
transform 1 0 30820 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0917_
timestamp 1666464484
transform 1 0 27140 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0918_
timestamp 1666464484
transform 1 0 23920 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0919_
timestamp 1666464484
transform 1 0 24656 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0920_
timestamp 1666464484
transform 1 0 26404 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0921_
timestamp 1666464484
transform 1 0 28796 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0922_
timestamp 1666464484
transform 1 0 26404 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _0923_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 25576 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0924_
timestamp 1666464484
transform 1 0 29532 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0925_
timestamp 1666464484
transform 1 0 25300 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0926_
timestamp 1666464484
transform 1 0 24564 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _0927_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 25300 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0928_
timestamp 1666464484
transform 1 0 26128 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0929_
timestamp 1666464484
transform 1 0 27324 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0930_
timestamp 1666464484
transform 1 0 34132 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _0931_
timestamp 1666464484
transform 1 0 25668 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0932_
timestamp 1666464484
transform 1 0 28980 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0933_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 24656 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0934_
timestamp 1666464484
transform 1 0 26404 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0935_
timestamp 1666464484
transform 1 0 24564 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0936_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 25392 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0937_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 26864 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0938_
timestamp 1666464484
transform 1 0 25668 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0939_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 26772 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0940_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 30268 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0941_
timestamp 1666464484
transform 1 0 34132 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _0942_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 27600 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _0943_
timestamp 1666464484
transform 1 0 27324 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0944_
timestamp 1666464484
transform 1 0 30728 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0945_
timestamp 1666464484
transform 1 0 27140 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0946_
timestamp 1666464484
transform 1 0 29256 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0947_
timestamp 1666464484
transform 1 0 28704 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0948_
timestamp 1666464484
transform 1 0 31556 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0949_
timestamp 1666464484
transform 1 0 22724 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _0950_
timestamp 1666464484
transform 1 0 28428 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0951_
timestamp 1666464484
transform 1 0 29716 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0952_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28152 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0953_
timestamp 1666464484
transform 1 0 27876 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0954_
timestamp 1666464484
transform 1 0 28796 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0955_
timestamp 1666464484
transform 1 0 29164 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _0956_
timestamp 1666464484
transform 1 0 27692 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _0957_
timestamp 1666464484
transform 1 0 26496 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _0958_
timestamp 1666464484
transform 1 0 28428 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _0959_
timestamp 1666464484
transform 1 0 28428 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0960_
timestamp 1666464484
transform 1 0 29992 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0961_
timestamp 1666464484
transform 1 0 29992 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0962_
timestamp 1666464484
transform 1 0 32936 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0963_
timestamp 1666464484
transform 1 0 28612 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0964_
timestamp 1666464484
transform 1 0 27324 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0965_
timestamp 1666464484
transform 1 0 29716 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0966_
timestamp 1666464484
transform 1 0 29716 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0967_
timestamp 1666464484
transform 1 0 28980 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0968_
timestamp 1666464484
transform 1 0 28152 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0969_
timestamp 1666464484
transform 1 0 29808 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0970_
timestamp 1666464484
transform 1 0 28336 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0971_
timestamp 1666464484
transform 1 0 28244 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0972_
timestamp 1666464484
transform 1 0 28244 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0973_
timestamp 1666464484
transform 1 0 28980 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0974_
timestamp 1666464484
transform 1 0 30728 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0975_
timestamp 1666464484
transform 1 0 29716 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0976_
timestamp 1666464484
transform 1 0 20976 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0977_
timestamp 1666464484
transform 1 0 18032 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0978_
timestamp 1666464484
transform 1 0 16928 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0979_
timestamp 1666464484
transform 1 0 24656 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0980_
timestamp 1666464484
transform 1 0 15824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0981_
timestamp 1666464484
transform 1 0 17572 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0982_
timestamp 1666464484
transform 1 0 16468 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0983_
timestamp 1666464484
transform 1 0 18492 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0984_
timestamp 1666464484
transform 1 0 16836 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _0985_
timestamp 1666464484
transform 1 0 17296 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0986_
timestamp 1666464484
transform 1 0 18400 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0987_
timestamp 1666464484
transform 1 0 18584 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0988_
timestamp 1666464484
transform 1 0 19412 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _0989_
timestamp 1666464484
transform 1 0 17388 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0990_
timestamp 1666464484
transform 1 0 16560 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0991_
timestamp 1666464484
transform 1 0 16008 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0992_
timestamp 1666464484
transform 1 0 16560 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _0993_
timestamp 1666464484
transform 1 0 17480 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0994_
timestamp 1666464484
transform 1 0 18676 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0995_
timestamp 1666464484
transform 1 0 18124 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0996_
timestamp 1666464484
transform 1 0 18860 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0997_
timestamp 1666464484
transform 1 0 19412 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0998_
timestamp 1666464484
transform 1 0 17480 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0999_
timestamp 1666464484
transform 1 0 18400 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1000_
timestamp 1666464484
transform 1 0 16192 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1001_
timestamp 1666464484
transform 1 0 17204 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1002_
timestamp 1666464484
transform 1 0 15548 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1003_
timestamp 1666464484
transform 1 0 17204 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1004_
timestamp 1666464484
transform 1 0 18216 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1005_
timestamp 1666464484
transform 1 0 16560 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1006_
timestamp 1666464484
transform 1 0 15732 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1007_
timestamp 1666464484
transform 1 0 17388 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1008_
timestamp 1666464484
transform 1 0 17204 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1009_
timestamp 1666464484
transform 1 0 18216 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1010_
timestamp 1666464484
transform 1 0 17848 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1011_
timestamp 1666464484
transform 1 0 17020 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1012_
timestamp 1666464484
transform 1 0 16836 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1013_
timestamp 1666464484
transform 1 0 15916 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1014_
timestamp 1666464484
transform 1 0 18032 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1015_
timestamp 1666464484
transform 1 0 15088 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1016_
timestamp 1666464484
transform 1 0 17112 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1017_
timestamp 1666464484
transform 1 0 18216 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1018_
timestamp 1666464484
transform 1 0 16100 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1019_
timestamp 1666464484
transform 1 0 17112 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1020_
timestamp 1666464484
transform 1 0 17020 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1021_
timestamp 1666464484
transform 1 0 19136 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _1022_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 18400 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1023_
timestamp 1666464484
transform 1 0 15272 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1024_
timestamp 1666464484
transform 1 0 15916 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1025_
timestamp 1666464484
transform 1 0 16008 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1026_
timestamp 1666464484
transform 1 0 17112 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1027_
timestamp 1666464484
transform 1 0 15732 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1028_
timestamp 1666464484
transform 1 0 16836 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1029_
timestamp 1666464484
transform 1 0 17572 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1030_
timestamp 1666464484
transform 1 0 18216 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1031_
timestamp 1666464484
transform 1 0 16652 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1032_
timestamp 1666464484
transform 1 0 16376 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1033_
timestamp 1666464484
transform 1 0 16836 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1034_
timestamp 1666464484
transform 1 0 16008 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _1035_
timestamp 1666464484
transform 1 0 18308 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1036_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 20332 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1037_
timestamp 1666464484
transform 1 0 29716 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1038_
timestamp 1666464484
transform 1 0 27140 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1039_
timestamp 1666464484
transform 1 0 20148 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1040_
timestamp 1666464484
transform 1 0 18676 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1041_
timestamp 1666464484
transform 1 0 26128 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1042_
timestamp 1666464484
transform 1 0 25208 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1043_
timestamp 1666464484
transform 1 0 33856 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1044_
timestamp 1666464484
transform 1 0 28152 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1045_
timestamp 1666464484
transform 1 0 29716 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_2  _1046_
timestamp 1666464484
transform 1 0 30084 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1047_
timestamp 1666464484
transform 1 0 31556 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1048_
timestamp 1666464484
transform 1 0 27508 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1049_
timestamp 1666464484
transform 1 0 30452 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__and4b_1  _1050_
timestamp 1666464484
transform 1 0 27048 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1051_
timestamp 1666464484
transform 1 0 28244 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1052_
timestamp 1666464484
transform 1 0 28520 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1053_
timestamp 1666464484
transform 1 0 16100 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1054_
timestamp 1666464484
transform 1 0 27416 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1055_
timestamp 1666464484
transform 1 0 16100 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1056_
timestamp 1666464484
transform 1 0 31648 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1057_
timestamp 1666464484
transform 1 0 32292 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1058_
timestamp 1666464484
transform 1 0 27876 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1059_
timestamp 1666464484
transform 1 0 27508 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1060_
timestamp 1666464484
transform 1 0 28612 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1061_
timestamp 1666464484
transform 1 0 27784 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1062_
timestamp 1666464484
transform 1 0 28244 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1063_
timestamp 1666464484
transform 1 0 29716 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1064_
timestamp 1666464484
transform 1 0 29072 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1065_
timestamp 1666464484
transform 1 0 28704 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1066_
timestamp 1666464484
transform 1 0 29348 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1067_
timestamp 1666464484
transform 1 0 29716 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1068_
timestamp 1666464484
transform 1 0 29624 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1069_
timestamp 1666464484
transform 1 0 31648 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1070_
timestamp 1666464484
transform 1 0 28612 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1071_
timestamp 1666464484
transform 1 0 29256 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1072_
timestamp 1666464484
transform 1 0 30084 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1073_
timestamp 1666464484
transform 1 0 29716 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1074_
timestamp 1666464484
transform 1 0 31188 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1075_
timestamp 1666464484
transform 1 0 33672 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1076_
timestamp 1666464484
transform 1 0 34132 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1077_
timestamp 1666464484
transform 1 0 33304 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1078_
timestamp 1666464484
transform 1 0 31096 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1079_
timestamp 1666464484
transform 1 0 32292 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1080_
timestamp 1666464484
transform 1 0 32292 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1081_
timestamp 1666464484
transform 1 0 33396 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1082_
timestamp 1666464484
transform 1 0 28888 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1083_
timestamp 1666464484
transform 1 0 17480 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1084_
timestamp 1666464484
transform 1 0 27232 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1085_
timestamp 1666464484
transform 1 0 32384 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1086_
timestamp 1666464484
transform 1 0 19780 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1087_
timestamp 1666464484
transform 1 0 33212 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1088_
timestamp 1666464484
transform 1 0 31188 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1089_
timestamp 1666464484
transform 1 0 30636 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1090_
timestamp 1666464484
transform 1 0 33212 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1091_
timestamp 1666464484
transform 1 0 31096 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1092_
timestamp 1666464484
transform 1 0 32292 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1093_
timestamp 1666464484
transform 1 0 30728 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1094_
timestamp 1666464484
transform 1 0 29716 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1095_
timestamp 1666464484
transform 1 0 30084 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1096_
timestamp 1666464484
transform 1 0 34040 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1097_
timestamp 1666464484
transform 1 0 18492 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1098_
timestamp 1666464484
transform 1 0 19412 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1099_
timestamp 1666464484
transform 1 0 22632 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1100_
timestamp 1666464484
transform 1 0 26404 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1101_
timestamp 1666464484
transform 1 0 23828 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1102_
timestamp 1666464484
transform 1 0 16744 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1103_
timestamp 1666464484
transform 1 0 21988 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1104_
timestamp 1666464484
transform 1 0 23920 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1105_
timestamp 1666464484
transform 1 0 21068 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1106_
timestamp 1666464484
transform 1 0 21988 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1107_
timestamp 1666464484
transform 1 0 21068 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1108_
timestamp 1666464484
transform 1 0 21252 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1109_
timestamp 1666464484
transform 1 0 23552 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1110_
timestamp 1666464484
transform 1 0 23828 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1111_
timestamp 1666464484
transform 1 0 21068 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1112_
timestamp 1666464484
transform 1 0 19504 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1113_
timestamp 1666464484
transform 1 0 29072 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1114_
timestamp 1666464484
transform 1 0 27784 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1115_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 22816 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1116_
timestamp 1666464484
transform 1 0 23092 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1117_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 23920 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1118_
timestamp 1666464484
transform 1 0 22632 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1119_
timestamp 1666464484
transform 1 0 23000 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1120_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 23000 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1121_
timestamp 1666464484
transform 1 0 30820 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1122_
timestamp 1666464484
transform 1 0 28612 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1123_
timestamp 1666464484
transform 1 0 29716 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1124_
timestamp 1666464484
transform 1 0 27140 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1125_
timestamp 1666464484
transform 1 0 29900 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1126_
timestamp 1666464484
transform 1 0 23828 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1127_
timestamp 1666464484
transform 1 0 25484 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1128_
timestamp 1666464484
transform 1 0 16100 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1129_
timestamp 1666464484
transform 1 0 26312 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1130_
timestamp 1666464484
transform 1 0 24472 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1131_
timestamp 1666464484
transform 1 0 30728 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1132_
timestamp 1666464484
transform 1 0 24564 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1133_
timestamp 1666464484
transform 1 0 17480 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1134_
timestamp 1666464484
transform 1 0 22724 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1135_
timestamp 1666464484
transform 1 0 23828 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1136_
timestamp 1666464484
transform 1 0 25668 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1137_
timestamp 1666464484
transform 1 0 23828 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1138_
timestamp 1666464484
transform 1 0 23460 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1139_
timestamp 1666464484
transform 1 0 29072 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1140_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 25208 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1141_
timestamp 1666464484
transform 1 0 24564 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1142_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 25668 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1143_
timestamp 1666464484
transform 1 0 24564 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1144_
timestamp 1666464484
transform 1 0 17296 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1145_
timestamp 1666464484
transform 1 0 17940 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1146_
timestamp 1666464484
transform 1 0 19780 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1147_
timestamp 1666464484
transform 1 0 17664 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1148_
timestamp 1666464484
transform 1 0 18032 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1149_
timestamp 1666464484
transform 1 0 17388 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1150_
timestamp 1666464484
transform 1 0 17664 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1151_
timestamp 1666464484
transform 1 0 17020 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1152_
timestamp 1666464484
transform 1 0 19412 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1153_
timestamp 1666464484
transform 1 0 16652 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1154_
timestamp 1666464484
transform 1 0 23460 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1155_
timestamp 1666464484
transform 1 0 17388 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1156_
timestamp 1666464484
transform 1 0 23644 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1157_
timestamp 1666464484
transform 1 0 21988 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1158_
timestamp 1666464484
transform 1 0 20976 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1159_
timestamp 1666464484
transform 1 0 17020 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1160_
timestamp 1666464484
transform 1 0 20700 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1161_
timestamp 1666464484
transform 1 0 18492 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1162_
timestamp 1666464484
transform 1 0 19412 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1163_
timestamp 1666464484
transform 1 0 22172 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1164_
timestamp 1666464484
transform 1 0 19780 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1165_
timestamp 1666464484
transform 1 0 18216 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1166_
timestamp 1666464484
transform 1 0 18124 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1167_
timestamp 1666464484
transform 1 0 18216 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1168_
timestamp 1666464484
transform 1 0 21160 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1169_
timestamp 1666464484
transform 1 0 19412 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1170_
timestamp 1666464484
transform 1 0 18676 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1171_
timestamp 1666464484
transform 1 0 21068 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1172_
timestamp 1666464484
transform 1 0 19964 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1173_
timestamp 1666464484
transform 1 0 20792 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1174_
timestamp 1666464484
transform 1 0 21068 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1175_
timestamp 1666464484
transform 1 0 21344 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1176_
timestamp 1666464484
transform 1 0 21712 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1177_
timestamp 1666464484
transform 1 0 22080 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1178_
timestamp 1666464484
transform 1 0 22172 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1179_
timestamp 1666464484
transform 1 0 22540 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1180_
timestamp 1666464484
transform 1 0 23644 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1181_
timestamp 1666464484
transform 1 0 22080 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1182_
timestamp 1666464484
transform 1 0 24288 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1183_
timestamp 1666464484
transform 1 0 22816 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1184_
timestamp 1666464484
transform 1 0 20240 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1185_
timestamp 1666464484
transform 1 0 22908 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1186_
timestamp 1666464484
transform 1 0 21252 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _1187_
timestamp 1666464484
transform 1 0 20148 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1188_
timestamp 1666464484
transform 1 0 19872 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1189_
timestamp 1666464484
transform 1 0 23368 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1190_
timestamp 1666464484
transform 1 0 24564 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1191_
timestamp 1666464484
transform 1 0 26404 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1192_
timestamp 1666464484
transform 1 0 25668 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1193_
timestamp 1666464484
transform 1 0 27324 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1194_
timestamp 1666464484
transform 1 0 25944 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1195_
timestamp 1666464484
transform 1 0 26036 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1196_
timestamp 1666464484
transform 1 0 24932 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1197_
timestamp 1666464484
transform 1 0 25668 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1198_
timestamp 1666464484
transform 1 0 26312 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1199_
timestamp 1666464484
transform 1 0 26312 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1200_
timestamp 1666464484
transform 1 0 27968 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1201_
timestamp 1666464484
transform 1 0 27968 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1202_
timestamp 1666464484
transform 1 0 28888 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1203_
timestamp 1666464484
transform 1 0 28980 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1204_
timestamp 1666464484
transform 1 0 29716 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1205_
timestamp 1666464484
transform 1 0 28428 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1206_
timestamp 1666464484
transform 1 0 28244 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1207_
timestamp 1666464484
transform 1 0 26496 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1208_
timestamp 1666464484
transform 1 0 27140 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1209_
timestamp 1666464484
transform 1 0 28152 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1210_
timestamp 1666464484
transform 1 0 27140 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1211_
timestamp 1666464484
transform 1 0 25576 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1212_
timestamp 1666464484
transform 1 0 31372 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1213_
timestamp 1666464484
transform 1 0 16928 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1214_
timestamp 1666464484
transform 1 0 29716 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1215_
timestamp 1666464484
transform 1 0 20424 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1216_
timestamp 1666464484
transform 1 0 31372 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1217_
timestamp 1666464484
transform 1 0 18032 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1218_
timestamp 1666464484
transform 1 0 30820 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1219_
timestamp 1666464484
transform 1 0 13524 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1220_
timestamp 1666464484
transform 1 0 31648 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1221_
timestamp 1666464484
transform 1 0 17388 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1222_
timestamp 1666464484
transform 1 0 31464 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1223_
timestamp 1666464484
transform 1 0 30360 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1224_
timestamp 1666464484
transform 1 0 29808 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1225_
timestamp 1666464484
transform 1 0 31004 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1226_
timestamp 1666464484
transform 1 0 30636 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1227_
timestamp 1666464484
transform 1 0 18676 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1228_
timestamp 1666464484
transform 1 0 30636 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1229_
timestamp 1666464484
transform 1 0 31188 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1230_
timestamp 1666464484
transform 1 0 31280 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1231_
timestamp 1666464484
transform 1 0 31556 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1232_
timestamp 1666464484
transform 1 0 30544 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1233_
timestamp 1666464484
transform 1 0 30544 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1234_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 23828 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1235_
timestamp 1666464484
transform 1 0 23460 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1236_
timestamp 1666464484
transform 1 0 24564 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1237_
timestamp 1666464484
transform 1 0 23828 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1238_
timestamp 1666464484
transform 1 0 22816 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1239_
timestamp 1666464484
transform 1 0 24564 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1240_
timestamp 1666464484
transform 1 0 26404 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1241_
timestamp 1666464484
transform 1 0 27140 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1242_
timestamp 1666464484
transform 1 0 19412 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1243_
timestamp 1666464484
transform 1 0 19688 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1244_
timestamp 1666464484
transform 1 0 20056 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1245_
timestamp 1666464484
transform 1 0 21528 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1246_
timestamp 1666464484
transform 1 0 21988 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1247_
timestamp 1666464484
transform 1 0 22356 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1248_
timestamp 1666464484
transform 1 0 21988 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1249_
timestamp 1666464484
transform 1 0 21988 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1250_
timestamp 1666464484
transform 1 0 31096 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1251_
timestamp 1666464484
transform 1 0 32752 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1252_
timestamp 1666464484
transform 1 0 32292 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1253_
timestamp 1666464484
transform 1 0 32844 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1254_
timestamp 1666464484
transform 1 0 30360 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1255_
timestamp 1666464484
transform 1 0 32292 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1256_
timestamp 1666464484
transform 1 0 29624 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1257_
timestamp 1666464484
transform 1 0 29992 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1258_
timestamp 1666464484
transform 1 0 24472 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1259_
timestamp 1666464484
transform 1 0 23552 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1260_
timestamp 1666464484
transform 1 0 25484 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1261_
timestamp 1666464484
transform 1 0 27416 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1262_
timestamp 1666464484
transform 1 0 29716 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1263_
timestamp 1666464484
transform 1 0 27140 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1264_
timestamp 1666464484
transform 1 0 29716 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1265_
timestamp 1666464484
transform 1 0 28428 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1266_
timestamp 1666464484
transform 1 0 29808 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1267_
timestamp 1666464484
transform 1 0 18492 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1268_
timestamp 1666464484
transform 1 0 25208 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1269_
timestamp 1666464484
transform 1 0 18400 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1270_
timestamp 1666464484
transform 1 0 19320 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1271_
timestamp 1666464484
transform 1 0 19412 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1272_
timestamp 1666464484
transform 1 0 19044 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1273_
timestamp 1666464484
transform 1 0 19412 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1274_
timestamp 1666464484
transform 1 0 18676 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1275_
timestamp 1666464484
transform 1 0 18400 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1276_
timestamp 1666464484
transform 1 0 19412 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1277_
timestamp 1666464484
transform 1 0 26404 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1278_
timestamp 1666464484
transform 1 0 19412 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1279_
timestamp 1666464484
transform 1 0 28428 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1280_
timestamp 1666464484
transform 1 0 27140 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1281_
timestamp 1666464484
transform 1 0 28612 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1282_
timestamp 1666464484
transform 1 0 29716 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1283_
timestamp 1666464484
transform 1 0 32752 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1284_
timestamp 1666464484
transform 1 0 32936 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1285_
timestamp 1666464484
transform 1 0 31372 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1286_
timestamp 1666464484
transform 1 0 29348 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1287_
timestamp 1666464484
transform 1 0 19412 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1288_
timestamp 1666464484
transform 1 0 20792 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1289_
timestamp 1666464484
transform 1 0 22080 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1290_
timestamp 1666464484
transform 1 0 21988 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1291_
timestamp 1666464484
transform 1 0 21252 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1292_
timestamp 1666464484
transform 1 0 20792 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1293_
timestamp 1666464484
transform 1 0 22448 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1294_
timestamp 1666464484
transform 1 0 24288 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1295_
timestamp 1666464484
transform 1 0 27140 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1296_
timestamp 1666464484
transform 1 0 22632 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1297_
timestamp 1666464484
transform 1 0 27508 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1298_
timestamp 1666464484
transform 1 0 24748 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1299_
timestamp 1666464484
transform 1 0 24564 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1300_
timestamp 1666464484
transform 1 0 24564 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1301_
timestamp 1666464484
transform 1 0 23184 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1302_
timestamp 1666464484
transform 1 0 21988 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1303_
timestamp 1666464484
transform 1 0 22080 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1304_
timestamp 1666464484
transform 1 0 22632 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1305_
timestamp 1666464484
transform 1 0 24564 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1306_
timestamp 1666464484
transform 1 0 18124 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1307_
timestamp 1666464484
transform 1 0 18308 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1308_
timestamp 1666464484
transform 1 0 18124 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1309_
timestamp 1666464484
transform 1 0 18124 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1310_
timestamp 1666464484
transform 1 0 19136 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1311_
timestamp 1666464484
transform 1 0 19964 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1312_
timestamp 1666464484
transform 1 0 20332 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1313_
timestamp 1666464484
transform 1 0 20884 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1314_
timestamp 1666464484
transform 1 0 17296 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1315_
timestamp 1666464484
transform 1 0 18124 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1316_
timestamp 1666464484
transform 1 0 17388 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1317_
timestamp 1666464484
transform 1 0 19228 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1318_
timestamp 1666464484
transform 1 0 20884 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1319_
timestamp 1666464484
transform 1 0 21988 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1320_
timestamp 1666464484
transform 1 0 21988 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1321_
timestamp 1666464484
transform 1 0 23828 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1322_
timestamp 1666464484
transform 1 0 23368 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1323_
timestamp 1666464484
transform 1 0 19504 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1324_
timestamp 1666464484
transform 1 0 24564 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1325_
timestamp 1666464484
transform 1 0 24472 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1326_
timestamp 1666464484
transform 1 0 26404 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1327_
timestamp 1666464484
transform 1 0 24564 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1328_
timestamp 1666464484
transform 1 0 27140 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1329_
timestamp 1666464484
transform 1 0 27600 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1330_
timestamp 1666464484
transform 1 0 27784 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1331_
timestamp 1666464484
transform 1 0 27784 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1332_
timestamp 1666464484
transform 1 0 25484 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1333_
timestamp 1666464484
transform 1 0 32936 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1334_
timestamp 1666464484
transform 1 0 32016 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1335_
timestamp 1666464484
transform 1 0 32384 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1336_
timestamp 1666464484
transform 1 0 31832 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1337_
timestamp 1666464484
transform 1 0 30636 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1338_
timestamp 1666464484
transform 1 0 30176 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1339_
timestamp 1666464484
transform 1 0 29716 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1340_
timestamp 1666464484
transform 1 0 29900 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1341_
timestamp 1666464484
transform 1 0 26588 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1447__9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 5244 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1447_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 5888 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1448_
timestamp 1666464484
transform 1 0 1564 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1448__10
timestamp 1666464484
transform 1 0 2668 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1449__11
timestamp 1666464484
transform 1 0 15548 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1449_
timestamp 1666464484
transform 1 0 15548 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1450__12
timestamp 1666464484
transform 1 0 3128 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1450_
timestamp 1666464484
transform 1 0 1748 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1451__13
timestamp 1666464484
transform 1 0 30544 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1451_
timestamp 1666464484
transform 1 0 32476 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1452__14
timestamp 1666464484
transform 1 0 4048 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1452_
timestamp 1666464484
transform 1 0 1564 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1453_
timestamp 1666464484
transform 1 0 32476 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1453__15
timestamp 1666464484
transform 1 0 30544 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1454__16
timestamp 1666464484
transform 1 0 7176 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1454_
timestamp 1666464484
transform 1 0 6532 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1455__17
timestamp 1666464484
transform 1 0 27876 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1455_
timestamp 1666464484
transform 1 0 32476 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1456__18
timestamp 1666464484
transform 1 0 23184 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1456_
timestamp 1666464484
transform 1 0 32476 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1457_
timestamp 1666464484
transform 1 0 32476 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1457__19
timestamp 1666464484
transform 1 0 33120 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1458__20
timestamp 1666464484
transform 1 0 16836 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1458_
timestamp 1666464484
transform 1 0 16836 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1459_
timestamp 1666464484
transform 1 0 32476 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1459__21
timestamp 1666464484
transform 1 0 19964 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1460__22
timestamp 1666464484
transform 1 0 9752 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1460_
timestamp 1666464484
transform 1 0 1564 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1461_
timestamp 1666464484
transform 1 0 16836 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1461__23
timestamp 1666464484
transform 1 0 17572 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1462__24
timestamp 1666464484
transform 1 0 5244 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1462_
timestamp 1666464484
transform 1 0 4048 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1463_
timestamp 1666464484
transform 1 0 32476 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1463__25
timestamp 1666464484
transform 1 0 32476 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1464__26
timestamp 1666464484
transform 1 0 27784 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1464_
timestamp 1666464484
transform 1 0 32476 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1465__27
timestamp 1666464484
transform 1 0 9752 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1465_
timestamp 1666464484
transform 1 0 1564 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1466_
timestamp 1666464484
transform 1 0 32476 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1466__28
timestamp 1666464484
transform 1 0 33764 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1467_
timestamp 1666464484
transform 1 0 1748 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1467__29
timestamp 1666464484
transform 1 0 1840 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1468__30
timestamp 1666464484
transform 1 0 21896 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1468_
timestamp 1666464484
transform 1 0 32476 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1469__31
timestamp 1666464484
transform 1 0 20056 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1469_
timestamp 1666464484
transform 1 0 19964 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1470__32
timestamp 1666464484
transform 1 0 9108 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1470_
timestamp 1666464484
transform 1 0 9108 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1471_
timestamp 1666464484
transform 1 0 32476 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1471__33
timestamp 1666464484
transform 1 0 33120 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1472__34
timestamp 1666464484
transform 1 0 6256 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1472_
timestamp 1666464484
transform 1 0 2576 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1473__35
timestamp 1666464484
transform 1 0 33764 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1473_
timestamp 1666464484
transform 1 0 32476 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1474__36
timestamp 1666464484
transform 1 0 4600 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1474_
timestamp 1666464484
transform 1 0 1564 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1475_
timestamp 1666464484
transform 1 0 30176 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1475__37
timestamp 1666464484
transform 1 0 28980 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1476__38
timestamp 1666464484
transform 1 0 3956 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1476_
timestamp 1666464484
transform 1 0 4140 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1477_
timestamp 1666464484
transform 1 0 32476 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1477__39
timestamp 1666464484
transform 1 0 31188 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1478_
timestamp 1666464484
transform 1 0 32476 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1478__40
timestamp 1666464484
transform 1 0 20424 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1479_
timestamp 1666464484
transform 1 0 29808 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1479__41
timestamp 1666464484
transform 1 0 23828 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1480__42
timestamp 1666464484
transform 1 0 22264 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1480_
timestamp 1666464484
transform 1 0 21988 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1481__43
timestamp 1666464484
transform 1 0 4600 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1481_
timestamp 1666464484
transform 1 0 4140 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1482__44
timestamp 1666464484
transform 1 0 1748 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1482_
timestamp 1666464484
transform 1 0 1748 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1483_
timestamp 1666464484
transform 1 0 32476 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1483__45
timestamp 1666464484
transform 1 0 15456 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1484_
timestamp 1666464484
transform 1 0 14260 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1484__46
timestamp 1666464484
transform 1 0 13800 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1485_
timestamp 1666464484
transform 1 0 32476 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1485__47
timestamp 1666464484
transform 1 0 19412 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1486__48
timestamp 1666464484
transform 1 0 1840 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1486_
timestamp 1666464484
transform 1 0 1564 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1487__49
timestamp 1666464484
transform 1 0 13524 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1487_
timestamp 1666464484
transform 1 0 14260 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1488_
timestamp 1666464484
transform 1 0 1748 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1488__50
timestamp 1666464484
transform 1 0 1840 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1489_
timestamp 1666464484
transform 1 0 32476 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1489__51
timestamp 1666464484
transform 1 0 33580 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1490__52
timestamp 1666464484
transform 1 0 8188 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1490_
timestamp 1666464484
transform 1 0 1564 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1491__53
timestamp 1666464484
transform 1 0 4048 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1491_
timestamp 1666464484
transform 1 0 1564 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1492__54
timestamp 1666464484
transform 1 0 30360 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1492_
timestamp 1666464484
transform 1 0 29900 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1493_
timestamp 1666464484
transform 1 0 32476 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1494_
timestamp 1666464484
transform 1 0 6440 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1495_
timestamp 1666464484
transform 1 0 32476 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1496__55
timestamp 1666464484
transform 1 0 23184 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1496_
timestamp 1666464484
transform 1 0 32384 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1497_
timestamp 1666464484
transform 1 0 29900 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1497__56
timestamp 1666464484
transform 1 0 27692 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1498__57
timestamp 1666464484
transform 1 0 2484 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1498_
timestamp 1666464484
transform 1 0 1748 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1499_
timestamp 1666464484
transform 1 0 29440 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1499__58
timestamp 1666464484
transform 1 0 18768 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1500__59
timestamp 1666464484
transform 1 0 1840 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1500_
timestamp 1666464484
transform 1 0 1748 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1501__60
timestamp 1666464484
transform 1 0 24564 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1501_
timestamp 1666464484
transform 1 0 23828 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1502_
timestamp 1666464484
transform 1 0 32476 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1502__61
timestamp 1666464484
transform 1 0 32384 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1503_
timestamp 1666464484
transform 1 0 20700 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1503__62
timestamp 1666464484
transform 1 0 20792 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1504__63
timestamp 1666464484
transform 1 0 25852 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1504_
timestamp 1666464484
transform 1 0 24932 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1505__64
timestamp 1666464484
transform 1 0 5888 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1505_
timestamp 1666464484
transform 1 0 1564 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1506_
timestamp 1666464484
transform 1 0 27140 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1506__65
timestamp 1666464484
transform 1 0 19964 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1507_
timestamp 1666464484
transform 1 0 13064 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1507__66
timestamp 1666464484
transform 1 0 12880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1508__67
timestamp 1666464484
transform 1 0 31832 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1508_
timestamp 1666464484
transform 1 0 32476 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1509_
timestamp 1666464484
transform 1 0 1748 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1509__68
timestamp 1666464484
transform 1 0 1840 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1510__69
timestamp 1666464484
transform 1 0 2484 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1510_
timestamp 1666464484
transform 1 0 1748 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1511__70
timestamp 1666464484
transform 1 0 5428 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1511_
timestamp 1666464484
transform 1 0 1748 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1512__71
timestamp 1666464484
transform 1 0 33764 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1512_
timestamp 1666464484
transform 1 0 32476 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1513__72
timestamp 1666464484
transform 1 0 23828 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1513_
timestamp 1666464484
transform 1 0 32476 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1514__73
timestamp 1666464484
transform 1 0 23184 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1514_
timestamp 1666464484
transform 1 0 32476 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1515__74
timestamp 1666464484
transform 1 0 7728 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1515_
timestamp 1666464484
transform 1 0 8372 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1516_
timestamp 1666464484
transform 1 0 32476 0 -1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1516__75
timestamp 1666464484
transform 1 0 21252 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1517_
timestamp 1666464484
transform 1 0 19596 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1517__76
timestamp 1666464484
transform 1 0 20056 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1518__77
timestamp 1666464484
transform 1 0 29716 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1518_
timestamp 1666464484
transform 1 0 29624 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1519__78
timestamp 1666464484
transform 1 0 27232 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1519_
timestamp 1666464484
transform 1 0 28520 0 -1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1520__79
timestamp 1666464484
transform 1 0 19412 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1520_
timestamp 1666464484
transform 1 0 19412 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1521__80
timestamp 1666464484
transform 1 0 31188 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1521_
timestamp 1666464484
transform 1 0 32476 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1522__81
timestamp 1666464484
transform 1 0 1840 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1522_
timestamp 1666464484
transform 1 0 1564 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1523_
timestamp 1666464484
transform 1 0 32476 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1523__82
timestamp 1666464484
transform 1 0 31556 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1524__83
timestamp 1666464484
transform 1 0 5796 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1524_
timestamp 1666464484
transform 1 0 6532 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1525__84
timestamp 1666464484
transform 1 0 5336 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1525_
timestamp 1666464484
transform 1 0 1840 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1526__85
timestamp 1666464484
transform 1 0 8188 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1526_
timestamp 1666464484
transform 1 0 6992 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1527_
timestamp 1666464484
transform 1 0 1748 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1527__86
timestamp 1666464484
transform 1 0 2484 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1528__87
timestamp 1666464484
transform 1 0 16100 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1528_
timestamp 1666464484
transform 1 0 32476 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1529_
timestamp 1666464484
transform 1 0 32476 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1529__88
timestamp 1666464484
transform 1 0 30268 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1530_
timestamp 1666464484
transform 1 0 32476 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1530__89
timestamp 1666464484
transform 1 0 31832 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1531__90
timestamp 1666464484
transform 1 0 3956 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1531_
timestamp 1666464484
transform 1 0 1748 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1532__91
timestamp 1666464484
transform 1 0 6072 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1532_
timestamp 1666464484
transform 1 0 6716 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1533__92
timestamp 1666464484
transform 1 0 33120 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1533_
timestamp 1666464484
transform 1 0 32476 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1534__93
timestamp 1666464484
transform 1 0 9844 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1534_
timestamp 1666464484
transform 1 0 9292 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1535__94
timestamp 1666464484
transform 1 0 25208 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1535_
timestamp 1666464484
transform 1 0 24380 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1536__95
timestamp 1666464484
transform 1 0 9108 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1536_
timestamp 1666464484
transform 1 0 7912 0 -1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1537_
timestamp 1666464484
transform 1 0 32476 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1537__96
timestamp 1666464484
transform 1 0 33764 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1538_
timestamp 1666464484
transform 1 0 3036 0 -1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1538__97
timestamp 1666464484
transform 1 0 6072 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1539_
timestamp 1666464484
transform 1 0 3956 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1539__98
timestamp 1666464484
transform 1 0 7176 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1540_
timestamp 1666464484
transform 1 0 14444 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1540__99
timestamp 1666464484
transform 1 0 15456 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1541__100
timestamp 1666464484
transform 1 0 15732 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1541_
timestamp 1666464484
transform 1 0 16376 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1542_
timestamp 1666464484
transform 1 0 32476 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1542__101
timestamp 1666464484
transform 1 0 28612 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1543__102
timestamp 1666464484
transform 1 0 23000 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1543_
timestamp 1666464484
transform 1 0 32476 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1544__103
timestamp 1666464484
transform 1 0 19412 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1544_
timestamp 1666464484
transform 1 0 19136 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1545__104
timestamp 1666464484
transform 1 0 29256 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1545_
timestamp 1666464484
transform 1 0 32292 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1546__105
timestamp 1666464484
transform 1 0 18032 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1546_
timestamp 1666464484
transform 1 0 32476 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1547_
timestamp 1666464484
transform 1 0 1748 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1547__106
timestamp 1666464484
transform 1 0 8004 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1548__107
timestamp 1666464484
transform 1 0 33304 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1548_
timestamp 1666464484
transform 1 0 32292 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1549_
timestamp 1666464484
transform 1 0 1748 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1549__108
timestamp 1666464484
transform 1 0 1840 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1550__109
timestamp 1666464484
transform 1 0 31004 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1550_
timestamp 1666464484
transform 1 0 31004 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1551__110
timestamp 1666464484
transform 1 0 5152 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1551_
timestamp 1666464484
transform 1 0 4140 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1552_
timestamp 1666464484
transform 1 0 1748 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1552__111
timestamp 1666464484
transform 1 0 1840 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1553__112
timestamp 1666464484
transform 1 0 1840 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1553_
timestamp 1666464484
transform 1 0 1564 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1554_
timestamp 1666464484
transform 1 0 1564 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1554__113
timestamp 1666464484
transform 1 0 1840 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 27140 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_wb_clk_i
timestamp 1666464484
transform 1 0 20792 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_wb_clk_i
timestamp 1666464484
transform 1 0 20792 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_wb_clk_i
timestamp 1666464484
transform 1 0 26036 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_wb_clk_i
timestamp 1666464484
transform 1 0 28612 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_wb_clk_i
timestamp 1666464484
transform 1 0 20792 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_wb_clk_i
timestamp 1666464484
transform 1 0 20792 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_wb_clk_i
timestamp 1666464484
transform 1 0 28612 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_wb_clk_i
timestamp 1666464484
transform 1 0 26036 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1666464484
transform 1 0 1564 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1666464484
transform 1 0 18676 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1666464484
transform 1 0 10672 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1666464484
transform 1 0 21252 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1666464484
transform 1 0 18124 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1666464484
transform 1 0 16192 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1666464484
transform 1 0 6716 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input8
timestamp 1666464484
transform 1 0 34040 0 1 9792
box -38 -48 406 592
<< labels >>
flabel metal3 s 200 35988 800 36228 0 FreeSans 960 0 0 0 active
port 0 nsew signal input
flabel metal2 s 11582 200 11694 800 0 FreeSans 448 90 0 0 io_in[0]
port 1 nsew signal input
flabel metal2 s 18666 41200 18778 41800 0 FreeSans 448 90 0 0 io_in[10]
port 2 nsew signal input
flabel metal3 s 200 38708 800 38948 0 FreeSans 960 0 0 0 io_in[11]
port 3 nsew signal input
flabel metal3 s 35200 35988 35800 36228 0 FreeSans 960 0 0 0 io_in[12]
port 4 nsew signal input
flabel metal2 s 18022 200 18134 800 0 FreeSans 448 90 0 0 io_in[13]
port 5 nsew signal input
flabel metal2 s 11582 41200 11694 41800 0 FreeSans 448 90 0 0 io_in[14]
port 6 nsew signal input
flabel metal3 s 35200 37348 35800 37588 0 FreeSans 960 0 0 0 io_in[15]
port 7 nsew signal input
flabel metal3 s 35200 6068 35800 6308 0 FreeSans 960 0 0 0 io_in[16]
port 8 nsew signal input
flabel metal2 s 5142 41200 5254 41800 0 FreeSans 448 90 0 0 io_in[17]
port 9 nsew signal input
flabel metal2 s 6430 41200 6542 41800 0 FreeSans 448 90 0 0 io_in[18]
port 10 nsew signal input
flabel metal2 s 33478 200 33590 800 0 FreeSans 448 90 0 0 io_in[19]
port 11 nsew signal input
flabel metal3 s 200 12188 800 12428 0 FreeSans 960 0 0 0 io_in[1]
port 12 nsew signal input
flabel metal3 s 200 22388 800 22628 0 FreeSans 960 0 0 0 io_in[20]
port 13 nsew signal input
flabel metal3 s 200 14908 800 15148 0 FreeSans 960 0 0 0 io_in[21]
port 14 nsew signal input
flabel metal3 s 35200 15588 35800 15828 0 FreeSans 960 0 0 0 io_in[22]
port 15 nsew signal input
flabel metal2 s 4498 41200 4610 41800 0 FreeSans 448 90 0 0 io_in[23]
port 16 nsew signal input
flabel metal2 s 1922 41200 2034 41800 0 FreeSans 448 90 0 0 io_in[24]
port 17 nsew signal input
flabel metal2 s 28970 200 29082 800 0 FreeSans 448 90 0 0 io_in[25]
port 18 nsew signal input
flabel metal2 s 28326 200 28438 800 0 FreeSans 448 90 0 0 io_in[26]
port 19 nsew signal input
flabel metal3 s 35200 11508 35800 11748 0 FreeSans 960 0 0 0 io_in[27]
port 20 nsew signal input
flabel metal2 s 25750 200 25862 800 0 FreeSans 448 90 0 0 io_in[28]
port 21 nsew signal input
flabel metal2 s 35410 41200 35522 41800 0 FreeSans 448 90 0 0 io_in[29]
port 22 nsew signal input
flabel metal2 s 12870 200 12982 800 0 FreeSans 448 90 0 0 io_in[2]
port 23 nsew signal input
flabel metal3 s 35200 18308 35800 18548 0 FreeSans 960 0 0 0 io_in[30]
port 24 nsew signal input
flabel metal3 s 200 34628 800 34868 0 FreeSans 960 0 0 0 io_in[31]
port 25 nsew signal input
flabel metal2 s 23818 200 23930 800 0 FreeSans 448 90 0 0 io_in[32]
port 26 nsew signal input
flabel metal3 s 200 20348 800 20588 0 FreeSans 960 0 0 0 io_in[33]
port 27 nsew signal input
flabel metal2 s 26394 41200 26506 41800 0 FreeSans 448 90 0 0 io_in[34]
port 28 nsew signal input
flabel metal2 s 30902 41200 31014 41800 0 FreeSans 448 90 0 0 io_in[35]
port 29 nsew signal input
flabel metal3 s 35200 27148 35800 27388 0 FreeSans 960 0 0 0 io_in[36]
port 30 nsew signal input
flabel metal2 s 31546 41200 31658 41800 0 FreeSans 448 90 0 0 io_in[37]
port 31 nsew signal input
flabel metal2 s 19310 41200 19422 41800 0 FreeSans 448 90 0 0 io_in[3]
port 32 nsew signal input
flabel metal3 s 35200 26468 35800 26708 0 FreeSans 960 0 0 0 io_in[4]
port 33 nsew signal input
flabel metal3 s 35200 40068 35800 40308 0 FreeSans 960 0 0 0 io_in[5]
port 34 nsew signal input
flabel metal3 s 200 23748 800 23988 0 FreeSans 960 0 0 0 io_in[6]
port 35 nsew signal input
flabel metal3 s 200 16268 800 16508 0 FreeSans 960 0 0 0 io_in[7]
port 36 nsew signal input
flabel metal3 s 35200 29188 35800 29428 0 FreeSans 960 0 0 0 io_in[8]
port 37 nsew signal input
flabel metal2 s 3210 41200 3322 41800 0 FreeSans 448 90 0 0 io_in[9]
port 38 nsew signal input
flabel metal2 s 20598 200 20710 800 0 FreeSans 448 90 0 0 io_oeb[0]
port 39 nsew signal tristate
flabel metal3 s 200 13548 800 13788 0 FreeSans 960 0 0 0 io_oeb[10]
port 40 nsew signal tristate
flabel metal3 s 35200 25108 35800 25348 0 FreeSans 960 0 0 0 io_oeb[11]
port 41 nsew signal tristate
flabel metal3 s 35200 14228 35800 14468 0 FreeSans 960 0 0 0 io_oeb[12]
port 42 nsew signal tristate
flabel metal3 s 35200 13548 35800 13788 0 FreeSans 960 0 0 0 io_oeb[13]
port 43 nsew signal tristate
flabel metal3 s 200 3348 800 3588 0 FreeSans 960 0 0 0 io_oeb[14]
port 44 nsew signal tristate
flabel metal2 s 7718 41200 7830 41800 0 FreeSans 448 90 0 0 io_oeb[15]
port 45 nsew signal tristate
flabel metal3 s 35200 4708 35800 4948 0 FreeSans 960 0 0 0 io_oeb[16]
port 46 nsew signal tristate
flabel metal2 s 10294 200 10406 800 0 FreeSans 448 90 0 0 io_oeb[17]
port 47 nsew signal tristate
flabel metal2 s 25106 41200 25218 41800 0 FreeSans 448 90 0 0 io_oeb[18]
port 48 nsew signal tristate
flabel metal2 s 8362 41200 8474 41800 0 FreeSans 448 90 0 0 io_oeb[19]
port 49 nsew signal tristate
flabel metal2 s 30258 200 30370 800 0 FreeSans 448 90 0 0 io_oeb[1]
port 50 nsew signal tristate
flabel metal3 s 35200 19668 35800 19908 0 FreeSans 960 0 0 0 io_oeb[20]
port 51 nsew signal tristate
flabel metal3 s 200 40748 800 40988 0 FreeSans 960 0 0 0 io_oeb[21]
port 52 nsew signal tristate
flabel metal2 s 3854 200 3966 800 0 FreeSans 448 90 0 0 io_oeb[22]
port 53 nsew signal tristate
flabel metal2 s 16090 41200 16202 41800 0 FreeSans 448 90 0 0 io_oeb[23]
port 54 nsew signal tristate
flabel metal2 s 17378 41200 17490 41800 0 FreeSans 448 90 0 0 io_oeb[24]
port 55 nsew signal tristate
flabel metal3 s 35200 628 35800 868 0 FreeSans 960 0 0 0 io_oeb[25]
port 56 nsew signal tristate
flabel metal3 s 35200 33268 35800 33508 0 FreeSans 960 0 0 0 io_oeb[26]
port 57 nsew signal tristate
flabel metal2 s 19954 41200 20066 41800 0 FreeSans 448 90 0 0 io_oeb[27]
port 58 nsew signal tristate
flabel metal2 s 32834 200 32946 800 0 FreeSans 448 90 0 0 io_oeb[28]
port 59 nsew signal tristate
flabel metal3 s 35200 27828 35800 28068 0 FreeSans 960 0 0 0 io_oeb[29]
port 60 nsew signal tristate
flabel metal2 s 28970 41200 29082 41800 0 FreeSans 448 90 0 0 io_oeb[2]
port 61 nsew signal tristate
flabel metal3 s 200 41428 800 41668 0 FreeSans 960 0 0 0 io_oeb[30]
port 62 nsew signal tristate
flabel metal2 s 32190 200 32302 800 0 FreeSans 448 90 0 0 io_oeb[31]
port 63 nsew signal tristate
flabel metal3 s 200 18988 800 19228 0 FreeSans 960 0 0 0 io_oeb[32]
port 64 nsew signal tristate
flabel metal3 s 35200 1988 35800 2228 0 FreeSans 960 0 0 0 io_oeb[33]
port 65 nsew signal tristate
flabel metal2 s 5786 41200 5898 41800 0 FreeSans 448 90 0 0 io_oeb[34]
port 66 nsew signal tristate
flabel metal3 s 200 16948 800 17188 0 FreeSans 960 0 0 0 io_oeb[35]
port 67 nsew signal tristate
flabel metal3 s 200 8788 800 9028 0 FreeSans 960 0 0 0 io_oeb[36]
port 68 nsew signal tristate
flabel metal3 s 200 14228 800 14468 0 FreeSans 960 0 0 0 io_oeb[37]
port 69 nsew signal tristate
flabel metal2 s 19954 200 20066 800 0 FreeSans 448 90 0 0 io_oeb[3]
port 70 nsew signal tristate
flabel metal3 s 35200 3348 35800 3588 0 FreeSans 960 0 0 0 io_oeb[4]
port 71 nsew signal tristate
flabel metal3 s 200 25108 800 25348 0 FreeSans 960 0 0 0 io_oeb[5]
port 72 nsew signal tristate
flabel metal3 s 35200 16948 35800 17188 0 FreeSans 960 0 0 0 io_oeb[6]
port 73 nsew signal tristate
flabel metal2 s 7074 41200 7186 41800 0 FreeSans 448 90 0 0 io_oeb[7]
port 74 nsew signal tristate
flabel metal2 s 3210 200 3322 800 0 FreeSans 448 90 0 0 io_oeb[8]
port 75 nsew signal tristate
flabel metal2 s 8362 200 8474 800 0 FreeSans 448 90 0 0 io_oeb[9]
port 76 nsew signal tristate
flabel metal3 s 35200 39388 35800 39628 0 FreeSans 960 0 0 0 io_out[0]
port 77 nsew signal tristate
flabel metal3 s 35200 24428 35800 24668 0 FreeSans 960 0 0 0 io_out[10]
port 78 nsew signal tristate
flabel metal3 s 200 1988 800 2228 0 FreeSans 960 0 0 0 io_out[11]
port 79 nsew signal tristate
flabel metal3 s 200 5388 800 5628 0 FreeSans 960 0 0 0 io_out[12]
port 80 nsew signal tristate
flabel metal2 s 30902 200 31014 800 0 FreeSans 448 90 0 0 io_out[13]
port 81 nsew signal tristate
flabel metal3 s 35200 33948 35800 34188 0 FreeSans 960 0 0 0 io_out[14]
port 82 nsew signal tristate
flabel metal3 s 200 31908 800 32148 0 FreeSans 960 0 0 0 io_out[15]
port 83 nsew signal tristate
flabel metal3 s 35200 23748 35800 23988 0 FreeSans 960 0 0 0 io_out[16]
port 84 nsew signal tristate
flabel metal2 s 32834 41200 32946 41800 0 FreeSans 448 90 0 0 io_out[17]
port 85 nsew signal tristate
flabel metal3 s 35200 -52 35800 188 0 FreeSans 960 0 0 0 io_out[18]
port 86 nsew signal tristate
flabel metal3 s 200 18308 800 18548 0 FreeSans 960 0 0 0 io_out[19]
port 87 nsew signal tristate
flabel metal2 s 22530 41200 22642 41800 0 FreeSans 448 90 0 0 io_out[1]
port 88 nsew signal tristate
flabel metal2 s 28326 41200 28438 41800 0 FreeSans 448 90 0 0 io_out[20]
port 89 nsew signal tristate
flabel metal3 s 200 31228 800 31468 0 FreeSans 960 0 0 0 io_out[21]
port 90 nsew signal tristate
flabel metal2 s 24462 200 24574 800 0 FreeSans 448 90 0 0 io_out[22]
port 91 nsew signal tristate
flabel metal3 s 35200 20348 35800 20588 0 FreeSans 960 0 0 0 io_out[23]
port 92 nsew signal tristate
flabel metal2 s 21242 200 21354 800 0 FreeSans 448 90 0 0 io_out[24]
port 93 nsew signal tristate
flabel metal2 s 25750 41200 25862 41800 0 FreeSans 448 90 0 0 io_out[25]
port 94 nsew signal tristate
flabel metal3 s 200 4028 800 4268 0 FreeSans 960 0 0 0 io_out[26]
port 95 nsew signal tristate
flabel metal2 s 27038 41200 27150 41800 0 FreeSans 448 90 0 0 io_out[27]
port 96 nsew signal tristate
flabel metal2 s 13514 200 13626 800 0 FreeSans 448 90 0 0 io_out[28]
port 97 nsew signal tristate
flabel metal3 s 35200 4028 35800 4268 0 FreeSans 960 0 0 0 io_out[29]
port 98 nsew signal tristate
flabel metal2 s 5142 200 5254 800 0 FreeSans 448 90 0 0 io_out[2]
port 99 nsew signal tristate
flabel metal3 s 200 4708 800 4948 0 FreeSans 960 0 0 0 io_out[30]
port 100 nsew signal tristate
flabel metal3 s 200 10828 800 11068 0 FreeSans 960 0 0 0 io_out[31]
port 101 nsew signal tristate
flabel metal3 s 200 36668 800 36908 0 FreeSans 960 0 0 0 io_out[32]
port 102 nsew signal tristate
flabel metal3 s 35200 8788 35800 9028 0 FreeSans 960 0 0 0 io_out[33]
port 103 nsew signal tristate
flabel metal3 s 35200 34628 35800 34868 0 FreeSans 960 0 0 0 io_out[34]
port 104 nsew signal tristate
flabel metal3 s 35200 32588 35800 32828 0 FreeSans 960 0 0 0 io_out[35]
port 105 nsew signal tristate
flabel metal2 s 9006 41200 9118 41800 0 FreeSans 448 90 0 0 io_out[36]
port 106 nsew signal tristate
flabel metal3 s 35200 38028 35800 38268 0 FreeSans 960 0 0 0 io_out[37]
port 107 nsew signal tristate
flabel metal3 s 200 33948 800 34188 0 FreeSans 960 0 0 0 io_out[3]
port 108 nsew signal tristate
flabel metal3 s 35200 25788 35800 26028 0 FreeSans 960 0 0 0 io_out[4]
port 109 nsew signal tristate
flabel metal2 s 14802 41200 14914 41800 0 FreeSans 448 90 0 0 io_out[5]
port 110 nsew signal tristate
flabel metal2 s 34122 41200 34234 41800 0 FreeSans 448 90 0 0 io_out[6]
port 111 nsew signal tristate
flabel metal3 s 200 15588 800 15828 0 FreeSans 960 0 0 0 io_out[7]
port 112 nsew signal tristate
flabel metal2 s 14802 200 14914 800 0 FreeSans 448 90 0 0 io_out[8]
port 113 nsew signal tristate
flabel metal3 s 200 11508 800 11748 0 FreeSans 960 0 0 0 io_out[9]
port 114 nsew signal tristate
flabel metal3 s 35200 9468 35800 9708 0 FreeSans 960 0 0 0 la1_data_in[0]
port 115 nsew signal input
flabel metal2 s 16734 200 16846 800 0 FreeSans 448 90 0 0 la1_data_in[10]
port 116 nsew signal input
flabel metal3 s 35200 7428 35800 7668 0 FreeSans 960 0 0 0 la1_data_in[11]
port 117 nsew signal input
flabel metal3 s 200 29188 800 29428 0 FreeSans 960 0 0 0 la1_data_in[12]
port 118 nsew signal input
flabel metal2 s 26394 200 26506 800 0 FreeSans 448 90 0 0 la1_data_in[13]
port 119 nsew signal input
flabel metal3 s 200 10148 800 10388 0 FreeSans 960 0 0 0 la1_data_in[14]
port 120 nsew signal input
flabel metal2 s 9650 41200 9762 41800 0 FreeSans 448 90 0 0 la1_data_in[15]
port 121 nsew signal input
flabel metal2 s 21242 41200 21354 41800 0 FreeSans 448 90 0 0 la1_data_in[16]
port 122 nsew signal input
flabel metal2 s 15446 41200 15558 41800 0 FreeSans 448 90 0 0 la1_data_in[17]
port 123 nsew signal input
flabel metal2 s 34122 200 34234 800 0 FreeSans 448 90 0 0 la1_data_in[18]
port 124 nsew signal input
flabel metal2 s 10938 41200 11050 41800 0 FreeSans 448 90 0 0 la1_data_in[19]
port 125 nsew signal input
flabel metal2 s 15446 200 15558 800 0 FreeSans 448 90 0 0 la1_data_in[1]
port 126 nsew signal input
flabel metal3 s 200 28508 800 28748 0 FreeSans 960 0 0 0 la1_data_in[20]
port 127 nsew signal input
flabel metal2 s 34766 41200 34878 41800 0 FreeSans 448 90 0 0 la1_data_in[21]
port 128 nsew signal input
flabel metal3 s 35200 10148 35800 10388 0 FreeSans 960 0 0 0 la1_data_in[22]
port 129 nsew signal input
flabel metal3 s 200 628 800 868 0 FreeSans 960 0 0 0 la1_data_in[23]
port 130 nsew signal input
flabel metal2 s 10938 200 11050 800 0 FreeSans 448 90 0 0 la1_data_in[24]
port 131 nsew signal input
flabel metal3 s 200 29868 800 30108 0 FreeSans 960 0 0 0 la1_data_in[25]
port 132 nsew signal input
flabel metal3 s 35200 5388 35800 5628 0 FreeSans 960 0 0 0 la1_data_in[26]
port 133 nsew signal input
flabel metal2 s 22530 200 22642 800 0 FreeSans 448 90 0 0 la1_data_in[27]
port 134 nsew signal input
flabel metal3 s 200 25788 800 26028 0 FreeSans 960 0 0 0 la1_data_in[28]
port 135 nsew signal input
flabel metal3 s 200 39388 800 39628 0 FreeSans 960 0 0 0 la1_data_in[29]
port 136 nsew signal input
flabel metal2 s 9006 200 9118 800 0 FreeSans 448 90 0 0 la1_data_in[2]
port 137 nsew signal input
flabel metal2 s 1278 200 1390 800 0 FreeSans 448 90 0 0 la1_data_in[30]
port 138 nsew signal input
flabel metal2 s 29614 200 29726 800 0 FreeSans 448 90 0 0 la1_data_in[31]
port 139 nsew signal input
flabel metal3 s 200 24428 800 24668 0 FreeSans 960 0 0 0 la1_data_in[3]
port 140 nsew signal input
flabel metal2 s 30258 41200 30370 41800 0 FreeSans 448 90 0 0 la1_data_in[4]
port 141 nsew signal input
flabel metal3 s 35200 22388 35800 22628 0 FreeSans 960 0 0 0 la1_data_in[5]
port 142 nsew signal input
flabel metal2 s 12226 41200 12338 41800 0 FreeSans 448 90 0 0 la1_data_in[6]
port 143 nsew signal input
flabel metal3 s 200 17628 800 17868 0 FreeSans 960 0 0 0 la1_data_in[7]
port 144 nsew signal input
flabel metal2 s 12870 41200 12982 41800 0 FreeSans 448 90 0 0 la1_data_in[8]
port 145 nsew signal input
flabel metal3 s 200 27148 800 27388 0 FreeSans 960 0 0 0 la1_data_in[9]
port 146 nsew signal input
flabel metal2 s 6430 200 6542 800 0 FreeSans 448 90 0 0 la1_data_out[0]
port 147 nsew signal tristate
flabel metal3 s 35200 12188 35800 12428 0 FreeSans 960 0 0 0 la1_data_out[10]
port 148 nsew signal tristate
flabel metal2 s 17378 200 17490 800 0 FreeSans 448 90 0 0 la1_data_out[11]
port 149 nsew signal tristate
flabel metal3 s 35200 38708 35800 38948 0 FreeSans 960 0 0 0 la1_data_out[12]
port 150 nsew signal tristate
flabel metal2 s 634 41200 746 41800 0 FreeSans 448 90 0 0 la1_data_out[13]
port 151 nsew signal tristate
flabel metal2 s 18022 41200 18134 41800 0 FreeSans 448 90 0 0 la1_data_out[14]
port 152 nsew signal tristate
flabel metal3 s 200 1308 800 1548 0 FreeSans 960 0 0 0 la1_data_out[15]
port 153 nsew signal tristate
flabel metal3 s 35200 16268 35800 16508 0 FreeSans 960 0 0 0 la1_data_out[16]
port 154 nsew signal tristate
flabel metal3 s 35200 31228 35800 31468 0 FreeSans 960 0 0 0 la1_data_out[17]
port 155 nsew signal tristate
flabel metal2 s 1278 41200 1390 41800 0 FreeSans 448 90 0 0 la1_data_out[18]
port 156 nsew signal tristate
flabel metal3 s 35200 23068 35800 23308 0 FreeSans 960 0 0 0 la1_data_out[19]
port 157 nsew signal tristate
flabel metal3 s 200 35308 800 35548 0 FreeSans 960 0 0 0 la1_data_out[1]
port 158 nsew signal tristate
flabel metal3 s 200 8108 800 8348 0 FreeSans 960 0 0 0 la1_data_out[20]
port 159 nsew signal tristate
flabel metal3 s 35200 36668 35800 36908 0 FreeSans 960 0 0 0 la1_data_out[21]
port 160 nsew signal tristate
flabel metal2 s 20598 41200 20710 41800 0 FreeSans 448 90 0 0 la1_data_out[22]
port 161 nsew signal tristate
flabel metal2 s 9650 200 9762 800 0 FreeSans 448 90 0 0 la1_data_out[23]
port 162 nsew signal tristate
flabel metal3 s 35200 17628 35800 17868 0 FreeSans 960 0 0 0 la1_data_out[24]
port 163 nsew signal tristate
flabel metal3 s 200 2668 800 2908 0 FreeSans 960 0 0 0 la1_data_out[25]
port 164 nsew signal tristate
flabel metal3 s 35200 6748 35800 6988 0 FreeSans 960 0 0 0 la1_data_out[26]
port 165 nsew signal tristate
flabel metal3 s 200 37348 800 37588 0 FreeSans 960 0 0 0 la1_data_out[27]
port 166 nsew signal tristate
flabel metal2 s 34766 200 34878 800 0 FreeSans 448 90 0 0 la1_data_out[28]
port 167 nsew signal tristate
flabel metal2 s 4498 200 4610 800 0 FreeSans 448 90 0 0 la1_data_out[29]
port 168 nsew signal tristate
flabel metal2 s 16090 200 16202 800 0 FreeSans 448 90 0 0 la1_data_out[2]
port 169 nsew signal tristate
flabel metal3 s 35200 12868 35800 13108 0 FreeSans 960 0 0 0 la1_data_out[30]
port 170 nsew signal tristate
flabel metal3 s 35200 40748 35800 40988 0 FreeSans 960 0 0 0 la1_data_out[31]
port 171 nsew signal tristate
flabel metal3 s 200 7428 800 7668 0 FreeSans 960 0 0 0 la1_data_out[3]
port 172 nsew signal tristate
flabel metal2 s 35410 200 35522 800 0 FreeSans 448 90 0 0 la1_data_out[4]
port 173 nsew signal tristate
flabel metal2 s 2566 200 2678 800 0 FreeSans 448 90 0 0 la1_data_out[5]
port 174 nsew signal tristate
flabel metal3 s 35200 18988 35800 19228 0 FreeSans 960 0 0 0 la1_data_out[6]
port 175 nsew signal tristate
flabel metal2 s 634 200 746 800 0 FreeSans 448 90 0 0 la1_data_out[7]
port 176 nsew signal tristate
flabel metal3 s 35200 31908 35800 32148 0 FreeSans 960 0 0 0 la1_data_out[8]
port 177 nsew signal tristate
flabel metal2 s 33478 41200 33590 41800 0 FreeSans 448 90 0 0 la1_data_out[9]
port 178 nsew signal tristate
flabel metal3 s 35200 2668 35800 2908 0 FreeSans 960 0 0 0 la1_oenb[0]
port 179 nsew signal input
flabel metal2 s 32190 41200 32302 41800 0 FreeSans 448 90 0 0 la1_oenb[10]
port 180 nsew signal input
flabel metal3 s 200 21708 800 21948 0 FreeSans 960 0 0 0 la1_oenb[11]
port 181 nsew signal input
flabel metal3 s 200 23068 800 23308 0 FreeSans 960 0 0 0 la1_oenb[12]
port 182 nsew signal input
flabel metal2 s 23174 200 23286 800 0 FreeSans 448 90 0 0 la1_oenb[13]
port 183 nsew signal input
flabel metal2 s -10 200 102 800 0 FreeSans 448 90 0 0 la1_oenb[14]
port 184 nsew signal input
flabel metal2 s 27682 200 27794 800 0 FreeSans 448 90 0 0 la1_oenb[15]
port 185 nsew signal input
flabel metal3 s 200 27828 800 28068 0 FreeSans 960 0 0 0 la1_oenb[16]
port 186 nsew signal input
flabel metal2 s -10 41200 102 41800 0 FreeSans 448 90 0 0 la1_oenb[17]
port 187 nsew signal input
flabel metal2 s 14158 41200 14270 41800 0 FreeSans 448 90 0 0 la1_oenb[18]
port 188 nsew signal input
flabel metal3 s 200 21028 800 21268 0 FreeSans 960 0 0 0 la1_oenb[19]
port 189 nsew signal input
flabel metal2 s 7074 200 7186 800 0 FreeSans 448 90 0 0 la1_oenb[1]
port 190 nsew signal input
flabel metal2 s 1922 200 2034 800 0 FreeSans 448 90 0 0 la1_oenb[20]
port 191 nsew signal input
flabel metal2 s 21886 41200 21998 41800 0 FreeSans 448 90 0 0 la1_oenb[21]
port 192 nsew signal input
flabel metal2 s 13514 41200 13626 41800 0 FreeSans 448 90 0 0 la1_oenb[22]
port 193 nsew signal input
flabel metal2 s 19310 200 19422 800 0 FreeSans 448 90 0 0 la1_oenb[23]
port 194 nsew signal input
flabel metal2 s 27682 41200 27794 41800 0 FreeSans 448 90 0 0 la1_oenb[24]
port 195 nsew signal input
flabel metal3 s 35200 10828 35800 11068 0 FreeSans 960 0 0 0 la1_oenb[25]
port 196 nsew signal input
flabel metal3 s 200 30548 800 30788 0 FreeSans 960 0 0 0 la1_oenb[26]
port 197 nsew signal input
flabel metal3 s 35200 30548 35800 30788 0 FreeSans 960 0 0 0 la1_oenb[27]
port 198 nsew signal input
flabel metal2 s 7718 200 7830 800 0 FreeSans 448 90 0 0 la1_oenb[28]
port 199 nsew signal input
flabel metal2 s 14158 200 14270 800 0 FreeSans 448 90 0 0 la1_oenb[29]
port 200 nsew signal input
flabel metal3 s 200 6748 800 6988 0 FreeSans 960 0 0 0 la1_oenb[2]
port 201 nsew signal input
flabel metal3 s 35200 29868 35800 30108 0 FreeSans 960 0 0 0 la1_oenb[30]
port 202 nsew signal input
flabel metal2 s 21886 200 21998 800 0 FreeSans 448 90 0 0 la1_oenb[31]
port 203 nsew signal input
flabel metal2 s 24462 41200 24574 41800 0 FreeSans 448 90 0 0 la1_oenb[3]
port 204 nsew signal input
flabel metal2 s 23818 41200 23930 41800 0 FreeSans 448 90 0 0 la1_oenb[4]
port 205 nsew signal input
flabel metal3 s 200 38028 800 38268 0 FreeSans 960 0 0 0 la1_oenb[5]
port 206 nsew signal input
flabel metal2 s 2566 41200 2678 41800 0 FreeSans 448 90 0 0 la1_oenb[6]
port 207 nsew signal input
flabel metal2 s 27038 200 27150 800 0 FreeSans 448 90 0 0 la1_oenb[7]
port 208 nsew signal input
flabel metal3 s 200 9468 800 9708 0 FreeSans 960 0 0 0 la1_oenb[8]
port 209 nsew signal input
flabel metal3 s 200 32588 800 32828 0 FreeSans 960 0 0 0 la1_oenb[9]
port 210 nsew signal input
flabel metal4 s 5164 2128 5484 39760 0 FreeSans 1920 90 0 0 vccd1
port 211 nsew power bidirectional
flabel metal4 s 13605 2128 13925 39760 0 FreeSans 1920 90 0 0 vccd1
port 211 nsew power bidirectional
flabel metal4 s 22046 2128 22366 39760 0 FreeSans 1920 90 0 0 vccd1
port 211 nsew power bidirectional
flabel metal4 s 30487 2128 30807 39760 0 FreeSans 1920 90 0 0 vccd1
port 211 nsew power bidirectional
flabel metal4 s 9384 2128 9704 39760 0 FreeSans 1920 90 0 0 vssd1
port 212 nsew ground bidirectional
flabel metal4 s 17825 2128 18145 39760 0 FreeSans 1920 90 0 0 vssd1
port 212 nsew ground bidirectional
flabel metal4 s 26266 2128 26586 39760 0 FreeSans 1920 90 0 0 vssd1
port 212 nsew ground bidirectional
flabel metal4 s 34707 2128 35027 39760 0 FreeSans 1920 90 0 0 vssd1
port 212 nsew ground bidirectional
flabel metal3 s 35200 21028 35800 21268 0 FreeSans 960 0 0 0 wb_clk_i
port 213 nsew signal input
rlabel metal1 17986 39712 17986 39712 0 vccd1
rlabel via1 18065 39168 18065 39168 0 vssd1
rlabel metal1 24656 15674 24656 15674 0 _0000_
rlabel metal2 23598 21318 23598 21318 0 _0001_
rlabel metal2 24794 18224 24794 18224 0 _0002_
rlabel metal1 23920 15674 23920 15674 0 _0003_
rlabel metal1 23317 17238 23317 17238 0 _0004_
rlabel metal1 25111 17578 25111 17578 0 _0005_
rlabel metal1 26680 14586 26680 14586 0 _0006_
rlabel metal1 26802 17238 26802 17238 0 _0007_
rlabel metal2 19366 17442 19366 17442 0 _0008_
rlabel metal2 20286 18530 20286 18530 0 _0009_
rlabel metal2 20654 16966 20654 16966 0 _0010_
rlabel metal2 21666 17170 21666 17170 0 _0011_
rlabel metal1 22954 15674 22954 15674 0 _0012_
rlabel metal2 22954 19618 22954 19618 0 _0013_
rlabel metal1 22908 16218 22908 16218 0 _0014_
rlabel metal1 23455 22678 23455 22678 0 _0015_
rlabel metal1 30774 15674 30774 15674 0 _0016_
rlabel metal1 32322 21930 32322 21930 0 _0017_
rlabel metal1 33028 18394 33028 18394 0 _0018_
rlabel metal1 32890 15674 32890 15674 0 _0019_
rlabel metal1 30861 19346 30861 19346 0 _0020_
rlabel metal2 33718 19686 33718 19686 0 _0021_
rlabel metal1 34178 16218 34178 16218 0 _0022_
rlabel metal1 30585 22678 30585 22678 0 _0023_
rlabel metal1 23782 26418 23782 26418 0 _0024_
rlabel metal1 24518 22202 24518 22202 0 _0025_
rlabel metal1 25606 23018 25606 23018 0 _0026_
rlabel metal1 27538 21590 27538 21590 0 _0027_
rlabel metal1 29614 21998 29614 21998 0 _0028_
rlabel metal1 26910 20026 26910 20026 0 _0029_
rlabel metal2 30866 19346 30866 19346 0 _0030_
rlabel metal2 28382 18054 28382 18054 0 _0031_
rlabel metal1 29930 17578 29930 17578 0 _0032_
rlabel metal1 18712 28050 18712 28050 0 _0033_
rlabel metal1 21390 26792 21390 26792 0 _0034_
rlabel metal1 19085 22610 19085 22610 0 _0035_
rlabel metal2 19458 25670 19458 25670 0 _0036_
rlabel metal1 18982 24106 18982 24106 0 _0037_
rlabel metal1 18982 23766 18982 23766 0 _0038_
rlabel metal1 19534 20502 19534 20502 0 _0039_
rlabel via1 18993 21522 18993 21522 0 _0040_
rlabel metal1 18620 18258 18620 18258 0 _0041_
rlabel metal1 19258 19754 19258 19754 0 _0042_
rlabel metal1 26956 33286 26956 33286 0 _0043_
rlabel metal1 19688 33082 19688 33082 0 _0044_
rlabel metal1 29435 24786 29435 24786 0 _0045_
rlabel metal2 27554 26112 27554 26112 0 _0046_
rlabel metal1 29159 25874 29159 25874 0 _0047_
rlabel metal2 30038 28288 30038 28288 0 _0048_
rlabel metal2 32430 26588 32430 26588 0 _0049_
rlabel metal1 20930 27030 20930 27030 0 _0050_
rlabel metal2 31142 29376 31142 29376 0 _0051_
rlabel metal1 33902 35462 33902 35462 0 _0052_
rlabel metal2 19504 26486 19504 26486 0 _0053_
rlabel metal1 26680 27914 26680 27914 0 _0054_
rlabel metal2 16790 28288 16790 28288 0 _0055_
rlabel metal1 22949 26962 22949 26962 0 _0056_
rlabel via1 22034 25755 22034 25755 0 _0057_
rlabel metal1 21201 25194 21201 25194 0 _0058_
rlabel via1 22765 24786 22765 24786 0 _0059_
rlabel metal1 20815 24650 20815 24650 0 _0060_
rlabel metal1 27262 31382 27262 31382 0 _0061_
rlabel metal1 22995 25942 22995 25942 0 _0062_
rlabel metal1 28520 38182 28520 38182 0 _0063_
rlabel metal3 26266 36108 26266 36108 0 _0064_
rlabel metal1 24380 34918 24380 34918 0 _0065_
rlabel metal1 18722 28730 18722 28730 0 _0066_
rlabel metal2 30774 29376 30774 29376 0 _0067_
rlabel via2 19642 30277 19642 30277 0 _0068_
rlabel metal1 23690 33286 23690 33286 0 _0069_
rlabel metal1 23409 32470 23409 32470 0 _0070_
rlabel via1 24881 28526 24881 28526 0 _0071_
rlabel via1 18441 33490 18441 33490 0 _0072_
rlabel via1 18625 31314 18625 31314 0 _0073_
rlabel metal2 17434 32232 17434 32232 0 _0074_
rlabel metal1 18712 30294 18712 30294 0 _0075_
rlabel metal1 19120 29206 19120 29206 0 _0076_
rlabel metal1 18124 28662 18124 28662 0 _0077_
rlabel metal1 21758 32198 21758 32198 0 _0078_
rlabel metal1 18952 31450 18952 31450 0 _0079_
rlabel via1 17613 29138 17613 29138 0 _0080_
rlabel metal1 18338 35734 18338 35734 0 _0081_
rlabel metal2 18722 34374 18722 34374 0 _0082_
rlabel metal1 19775 34646 19775 34646 0 _0083_
rlabel viali 21201 33966 21201 33966 0 _0084_
rlabel metal2 22494 34782 22494 34782 0 _0085_
rlabel metal1 22443 34578 22443 34578 0 _0086_
rlabel metal1 23904 34646 23904 34646 0 _0087_
rlabel metal1 24007 35734 24007 35734 0 _0088_
rlabel via1 19821 32878 19821 32878 0 _0089_
rlabel metal1 24784 33966 24784 33966 0 _0090_
rlabel metal1 25249 33558 25249 33558 0 _0091_
rlabel metal1 26342 33898 26342 33898 0 _0092_
rlabel via1 24881 35054 24881 35054 0 _0093_
rlabel metal1 27216 34646 27216 34646 0 _0094_
rlabel metal1 27963 34986 27963 34986 0 _0095_
rlabel metal2 29302 34051 29302 34051 0 _0096_
rlabel metal1 28285 32810 28285 32810 0 _0097_
rlabel metal2 25622 32674 25622 32674 0 _0098_
rlabel metal2 21206 35785 21206 35785 0 _0099_
rlabel metal2 20654 32640 20654 32640 0 _0100_
rlabel metal1 19918 33388 19918 33388 0 _0101_
rlabel via2 20654 32963 20654 32963 0 _0102_
rlabel metal1 20102 35564 20102 35564 0 _0103_
rlabel metal2 30498 35258 30498 35258 0 _0104_
rlabel metal1 31004 39270 31004 39270 0 _0105_
rlabel metal2 19090 35360 19090 35360 0 _0106_
rlabel metal1 30406 31790 30406 31790 0 _0107_
rlabel metal1 3496 37230 3496 37230 0 _0108_
rlabel metal1 2024 19822 2024 19822 0 _0109_
rlabel metal1 2208 6766 2208 6766 0 _0110_
rlabel metal1 2530 7888 2530 7888 0 _0111_
rlabel metal1 5198 5678 5198 5678 0 _0112_
rlabel metal1 4186 5678 4186 5678 0 _0113_
rlabel metal1 2116 17646 2116 17646 0 _0114_
rlabel metal1 6532 5202 6532 5202 0 _0115_
rlabel metal2 5060 5508 5060 5508 0 _0116_
rlabel metal2 2070 21794 2070 21794 0 _0117_
rlabel metal1 4324 6290 4324 6290 0 _0118_
rlabel metal1 6302 36040 6302 36040 0 _0119_
rlabel metal2 29992 32878 29992 32878 0 _0120_
rlabel metal1 28888 21930 28888 21930 0 _0121_
rlabel metal1 29210 18734 29210 18734 0 _0122_
rlabel metal2 28106 16694 28106 16694 0 _0123_
rlabel metal1 27462 18326 27462 18326 0 _0124_
rlabel viali 27566 19346 27566 19346 0 _0125_
rlabel metal1 26128 19278 26128 19278 0 _0126_
rlabel metal1 25484 19346 25484 19346 0 _0127_
rlabel metal2 26174 18938 26174 18938 0 _0128_
rlabel metal1 26772 14518 26772 14518 0 _0129_
rlabel metal1 26266 21488 26266 21488 0 _0130_
rlabel metal1 25806 20570 25806 20570 0 _0131_
rlabel metal2 19550 19737 19550 19737 0 _0132_
rlabel metal2 25622 15215 25622 15215 0 _0133_
rlabel metal1 28796 18938 28796 18938 0 _0134_
rlabel metal1 25714 20434 25714 20434 0 _0135_
rlabel metal1 25346 20400 25346 20400 0 _0136_
rlabel metal1 26450 18734 26450 18734 0 _0137_
rlabel metal1 25990 18700 25990 18700 0 _0138_
rlabel metal1 26726 18768 26726 18768 0 _0139_
rlabel metal2 27370 18428 27370 18428 0 _0140_
rlabel metal2 28014 20128 28014 20128 0 _0141_
rlabel metal2 33810 13345 33810 13345 0 _0142_
rlabel metal1 21528 24378 21528 24378 0 _0143_
rlabel metal1 23092 22066 23092 22066 0 _0144_
rlabel metal1 21942 21896 21942 21896 0 _0145_
rlabel metal1 20930 21454 20930 21454 0 _0146_
rlabel metal1 22080 19958 22080 19958 0 _0147_
rlabel metal2 21482 19652 21482 19652 0 _0148_
rlabel metal2 22586 20978 22586 20978 0 _0149_
rlabel metal1 20976 22066 20976 22066 0 _0150_
rlabel metal1 20562 21964 20562 21964 0 _0151_
rlabel metal2 20378 22542 20378 22542 0 _0152_
rlabel metal1 20378 24752 20378 24752 0 _0153_
rlabel metal1 21459 22678 21459 22678 0 _0154_
rlabel metal2 20654 23596 20654 23596 0 _0155_
rlabel metal2 23506 22916 23506 22916 0 _0156_
rlabel metal1 22908 21658 22908 21658 0 _0157_
rlabel metal1 22908 22950 22908 22950 0 _0158_
rlabel via2 21022 21539 21022 21539 0 _0159_
rlabel metal1 20746 21420 20746 21420 0 _0160_
rlabel metal2 21482 21828 21482 21828 0 _0161_
rlabel metal1 22356 21862 22356 21862 0 _0162_
rlabel metal2 8970 25398 8970 25398 0 _0163_
rlabel metal2 32246 25772 32246 25772 0 _0164_
rlabel via2 32430 16235 32430 16235 0 _0165_
rlabel metal2 31510 16507 31510 16507 0 _0166_
rlabel metal1 33994 15674 33994 15674 0 _0167_
rlabel metal1 33304 16218 33304 16218 0 _0168_
rlabel metal2 33074 16575 33074 16575 0 _0169_
rlabel metal2 33718 26758 33718 26758 0 _0170_
rlabel metal2 32062 18877 32062 18877 0 _0171_
rlabel metal1 31510 15674 31510 15674 0 _0172_
rlabel metal1 31142 24140 31142 24140 0 _0173_
rlabel metal2 32062 27489 32062 27489 0 _0174_
rlabel metal1 30728 16218 30728 16218 0 _0175_
rlabel metal1 30222 25262 30222 25262 0 _0176_
rlabel metal2 32062 24633 32062 24633 0 _0177_
rlabel metal1 31832 24174 31832 24174 0 _0178_
rlabel metal2 33074 25636 33074 25636 0 _0179_
rlabel metal1 33718 24650 33718 24650 0 _0180_
rlabel metal1 31234 25262 31234 25262 0 _0181_
rlabel metal2 31050 25670 31050 25670 0 _0182_
rlabel metal1 31112 21590 31112 21590 0 _0183_
rlabel metal1 16376 37842 16376 37842 0 _0184_
rlabel metal1 18906 19822 18906 19822 0 _0185_
rlabel metal1 20056 20842 20056 20842 0 _0186_
rlabel metal1 23782 20978 23782 20978 0 _0187_
rlabel metal1 24242 16694 24242 16694 0 _0188_
rlabel metal1 25622 18258 25622 18258 0 _0189_
rlabel metal1 25592 17238 25592 17238 0 _0190_
rlabel metal2 31878 17918 31878 17918 0 _0191_
rlabel metal2 23874 15946 23874 15946 0 _0192_
rlabel metal2 23690 16796 23690 16796 0 _0193_
rlabel metal2 25438 16252 25438 16252 0 _0194_
rlabel metal1 25300 16082 25300 16082 0 _0195_
rlabel metal2 26910 14926 26910 14926 0 _0196_
rlabel metal2 26634 15130 26634 15130 0 _0197_
rlabel metal1 26588 17170 26588 17170 0 _0198_
rlabel metal1 20470 18190 20470 18190 0 _0199_
rlabel metal2 20746 17918 20746 17918 0 _0200_
rlabel metal1 21574 16524 21574 16524 0 _0201_
rlabel metal2 21850 16762 21850 16762 0 _0202_
rlabel metal1 21666 16592 21666 16592 0 _0203_
rlabel metal2 19734 21488 19734 21488 0 _0204_
rlabel metal2 23046 15946 23046 15946 0 _0205_
rlabel metal2 24242 17442 24242 17442 0 _0206_
rlabel metal1 24472 15606 24472 15606 0 _0207_
rlabel metal2 20562 18955 20562 18955 0 _0208_
rlabel metal1 22954 16116 22954 16116 0 _0209_
rlabel metal1 25530 22474 25530 22474 0 _0210_
rlabel metal2 32430 24072 32430 24072 0 _0211_
rlabel metal1 32752 18122 32752 18122 0 _0212_
rlabel metal1 33212 18258 33212 18258 0 _0213_
rlabel metal1 31832 17170 31832 17170 0 _0214_
rlabel metal1 32614 15504 32614 15504 0 _0215_
rlabel metal1 31464 17850 31464 17850 0 _0216_
rlabel metal2 32706 17918 32706 17918 0 _0217_
rlabel metal1 32154 19686 32154 19686 0 _0218_
rlabel metal1 31326 21318 31326 21318 0 _0219_
rlabel metal1 31970 18156 31970 18156 0 _0220_
rlabel metal1 31280 23698 31280 23698 0 _0221_
rlabel metal1 27324 28186 27324 28186 0 _0222_
rlabel metal1 25714 26418 25714 26418 0 _0223_
rlabel metal2 26174 26928 26174 26928 0 _0224_
rlabel metal2 26082 25330 26082 25330 0 _0225_
rlabel metal1 26404 26350 26404 26350 0 _0226_
rlabel metal1 29762 17102 29762 17102 0 _0227_
rlabel metal1 26910 19856 26910 19856 0 _0228_
rlabel metal1 25070 21386 25070 21386 0 _0229_
rlabel metal1 26358 24820 26358 24820 0 _0230_
rlabel metal2 27094 24412 27094 24412 0 _0231_
rlabel metal1 34178 22678 34178 22678 0 _0232_
rlabel metal2 34270 24786 34270 24786 0 _0233_
rlabel metal1 26496 25330 26496 25330 0 _0234_
rlabel metal2 24978 24735 24978 24735 0 _0235_
rlabel metal1 26450 22644 26450 22644 0 _0236_
rlabel metal2 26634 23188 26634 23188 0 _0237_
rlabel metal2 27922 18666 27922 18666 0 _0238_
rlabel metal1 26542 24174 26542 24174 0 _0239_
rlabel metal1 26657 24038 26657 24038 0 _0240_
rlabel metal1 30268 24786 30268 24786 0 _0241_
rlabel metal1 28014 22508 28014 22508 0 _0242_
rlabel metal1 29624 21318 29624 21318 0 _0243_
rlabel metal1 28060 22406 28060 22406 0 _0244_
rlabel metal2 29992 16422 29992 16422 0 _0245_
rlabel metal1 29164 21522 29164 21522 0 _0246_
rlabel metal2 29670 21760 29670 21760 0 _0247_
rlabel metal3 30475 16524 30475 16524 0 _0248_
rlabel metal3 30038 16660 30038 16660 0 _0249_
rlabel metal1 20194 33830 20194 33830 0 _0250_
rlabel metal1 29210 24174 29210 24174 0 _0251_
rlabel metal1 28980 19754 28980 19754 0 _0252_
rlabel metal2 28842 19278 28842 19278 0 _0253_
rlabel metal1 28658 19890 28658 19890 0 _0254_
rlabel metal1 28888 19346 28888 19346 0 _0255_
rlabel metal1 27002 19788 27002 19788 0 _0256_
rlabel metal1 29118 20434 29118 20434 0 _0257_
rlabel metal1 29624 19482 29624 19482 0 _0258_
rlabel metal2 31970 20162 31970 20162 0 _0259_
rlabel metal2 30314 17952 30314 17952 0 _0260_
rlabel metal1 29302 15062 29302 15062 0 _0261_
rlabel metal2 28474 15674 28474 15674 0 _0262_
rlabel metal1 29256 15334 29256 15334 0 _0263_
rlabel metal1 29624 18938 29624 18938 0 _0264_
rlabel metal1 28566 16014 28566 16014 0 _0265_
rlabel metal1 28750 15980 28750 15980 0 _0266_
rlabel metal1 29440 16218 29440 16218 0 _0267_
rlabel metal1 28750 15674 28750 15674 0 _0268_
rlabel metal2 28842 16932 28842 16932 0 _0269_
rlabel metal2 30038 16796 30038 16796 0 _0270_
rlabel metal1 30084 16490 30084 16490 0 _0271_
rlabel metal1 17434 35020 17434 35020 0 _0272_
rlabel metal2 17158 28254 17158 28254 0 _0273_
rlabel metal1 18032 32742 18032 32742 0 _0274_
rlabel metal1 17802 26928 17802 26928 0 _0275_
rlabel metal1 17802 26316 17802 26316 0 _0276_
rlabel metal2 17894 26588 17894 26588 0 _0277_
rlabel metal2 17066 26554 17066 26554 0 _0278_
rlabel metal1 17664 20774 17664 20774 0 _0279_
rlabel metal2 19090 24990 19090 24990 0 _0280_
rlabel metal1 19642 23120 19642 23120 0 _0281_
rlabel metal1 17986 26996 17986 26996 0 _0282_
rlabel metal2 16054 25534 16054 25534 0 _0283_
rlabel metal1 16652 18802 16652 18802 0 _0284_
rlabel metal1 17756 25466 17756 25466 0 _0285_
rlabel metal1 18492 26350 18492 26350 0 _0286_
rlabel metal2 18446 25772 18446 25772 0 _0287_
rlabel metal2 18906 24956 18906 24956 0 _0288_
rlabel metal1 19458 24854 19458 24854 0 _0289_
rlabel metal1 18906 25908 18906 25908 0 _0290_
rlabel metal2 17434 25466 17434 25466 0 _0291_
rlabel metal1 16836 24378 16836 24378 0 _0292_
rlabel metal2 17618 24140 17618 24140 0 _0293_
rlabel metal1 17710 24140 17710 24140 0 _0294_
rlabel metal1 18170 23290 18170 23290 0 _0295_
rlabel metal1 17158 24038 17158 24038 0 _0296_
rlabel metal1 17480 24174 17480 24174 0 _0297_
rlabel metal1 18078 23732 18078 23732 0 _0298_
rlabel metal2 17250 24582 17250 24582 0 _0299_
rlabel metal1 18262 23698 18262 23698 0 _0300_
rlabel metal1 17204 22746 17204 22746 0 _0301_
rlabel metal2 16146 20978 16146 20978 0 _0302_
rlabel metal2 16054 21454 16054 21454 0 _0303_
rlabel metal1 18354 20570 18354 20570 0 _0304_
rlabel metal1 16238 21658 16238 21658 0 _0305_
rlabel metal1 18743 20978 18743 20978 0 _0306_
rlabel metal2 16698 21556 16698 21556 0 _0307_
rlabel metal1 17572 21658 17572 21658 0 _0308_
rlabel metal1 18032 22134 18032 22134 0 _0309_
rlabel metal1 18952 19210 18952 19210 0 _0310_
rlabel metal1 15824 19414 15824 19414 0 _0311_
rlabel metal1 16192 19482 16192 19482 0 _0312_
rlabel metal2 17066 20026 17066 20026 0 _0313_
rlabel metal1 17020 20570 17020 20570 0 _0314_
rlabel metal1 17158 19856 17158 19856 0 _0315_
rlabel metal2 17434 18564 17434 18564 0 _0316_
rlabel metal1 18722 18836 18722 18836 0 _0317_
rlabel metal1 16882 19346 16882 19346 0 _0318_
rlabel metal2 16974 19108 16974 19108 0 _0319_
rlabel metal1 17894 19210 17894 19210 0 _0320_
rlabel metal1 18216 19822 18216 19822 0 _0321_
rlabel metal1 21298 24820 21298 24820 0 _0322_
rlabel metal2 30130 32946 30130 32946 0 _0323_
rlabel metal1 19734 32538 19734 32538 0 _0324_
rlabel metal1 27968 29138 27968 29138 0 _0325_
rlabel metal1 28934 29070 28934 29070 0 _0326_
rlabel viali 29946 29614 29946 29614 0 _0327_
rlabel metal1 28796 30702 28796 30702 0 _0328_
rlabel metal1 29854 36754 29854 36754 0 _0329_
rlabel metal3 30107 36380 30107 36380 0 _0330_
rlabel metal1 27922 25909 27922 25909 0 _0331_
rlabel metal1 27968 24718 27968 24718 0 _0332_
rlabel metal2 29118 29818 29118 29818 0 _0333_
rlabel metal2 28566 29937 28566 29937 0 _0334_
rlabel metal1 32338 28594 32338 28594 0 _0335_
rlabel metal2 16330 27404 16330 27404 0 _0336_
rlabel metal2 16974 26724 16974 26724 0 _0337_
rlabel metal2 16146 26622 16146 26622 0 _0338_
rlabel metal1 32016 23290 32016 23290 0 _0339_
rlabel metal2 28382 25364 28382 25364 0 _0340_
rlabel metal1 27968 25466 27968 25466 0 _0341_
rlabel metal2 28290 28458 28290 28458 0 _0342_
rlabel metal1 30038 20910 30038 20910 0 _0343_
rlabel metal1 29808 20910 29808 20910 0 _0344_
rlabel metal1 29808 21114 29808 21114 0 _0345_
rlabel metal1 28934 28492 28934 28492 0 _0346_
rlabel metal1 29854 26996 29854 26996 0 _0347_
rlabel metal1 31142 39610 31142 39610 0 _0348_
rlabel metal1 28842 28628 28842 28628 0 _0349_
rlabel metal1 29486 28083 29486 28083 0 _0350_
rlabel viali 29575 28050 29575 28050 0 _0351_
rlabel metal1 30176 26554 30176 26554 0 _0352_
rlabel metal2 31602 27676 31602 27676 0 _0353_
rlabel metal1 33764 32810 33764 32810 0 _0354_
rlabel metal1 33856 29274 33856 29274 0 _0355_
rlabel metal2 33810 28798 33810 28798 0 _0356_
rlabel metal1 32292 27030 32292 27030 0 _0357_
rlabel metal2 32890 27710 32890 27710 0 _0358_
rlabel metal1 33258 28594 33258 28594 0 _0359_
rlabel metal2 17894 29665 17894 29665 0 _0360_
rlabel metal2 19642 29937 19642 29937 0 _0361_
rlabel metal1 26266 39610 26266 39610 0 _0362_
rlabel metal2 19826 35853 19826 35853 0 _0363_
rlabel metal2 20010 31212 20010 31212 0 _0364_
rlabel metal1 32062 27982 32062 27982 0 _0365_
rlabel metal1 31096 28186 31096 28186 0 _0366_
rlabel via1 31507 29139 31507 29139 0 _0367_
rlabel metal1 31648 29138 31648 29138 0 _0368_
rlabel metal1 32246 29138 32246 29138 0 _0369_
rlabel viali 30033 30770 30033 30770 0 _0370_
rlabel metal1 33948 35598 33948 35598 0 _0371_
rlabel metal2 34086 36584 34086 36584 0 _0372_
rlabel metal1 19504 26350 19504 26350 0 _0373_
rlabel metal1 26404 28050 26404 28050 0 _0374_
rlabel metal1 20194 29104 20194 29104 0 _0375_
rlabel metal2 24150 28628 24150 28628 0 _0376_
rlabel metal2 22402 26860 22402 26860 0 _0377_
rlabel metal2 21482 25874 21482 25874 0 _0378_
rlabel metal1 24012 24378 24012 24378 0 _0379_
rlabel metal1 21114 23562 21114 23562 0 _0380_
rlabel metal1 29394 34714 29394 34714 0 _0381_
rlabel metal1 23368 25466 23368 25466 0 _0382_
rlabel metal2 23230 26860 23230 26860 0 _0383_
rlabel metal2 24426 27642 24426 27642 0 _0384_
rlabel metal2 23138 26418 23138 26418 0 _0385_
rlabel via1 23519 26350 23519 26350 0 _0386_
rlabel metal2 31234 37502 31234 37502 0 _0387_
rlabel metal1 29992 32742 29992 32742 0 _0388_
rlabel metal1 30268 32538 30268 32538 0 _0389_
rlabel metal1 17434 32538 17434 32538 0 _0390_
rlabel metal2 19090 29546 19090 29546 0 _0391_
rlabel metal1 26450 32198 26450 32198 0 _0392_
rlabel metal1 18262 30192 18262 30192 0 _0393_
rlabel metal1 23598 33082 23598 33082 0 _0394_
rlabel metal1 24150 33966 24150 33966 0 _0395_
rlabel metal1 29264 32470 29264 32470 0 _0396_
rlabel metal2 29440 31212 29440 31212 0 _0397_
rlabel metal2 26036 33422 26036 33422 0 _0398_
rlabel metal2 25070 30668 25070 30668 0 _0399_
rlabel metal1 25415 29546 25415 29546 0 _0400_
rlabel metal1 18262 33966 18262 33966 0 _0401_
rlabel metal2 17618 31654 17618 31654 0 _0402_
rlabel metal1 17618 31824 17618 31824 0 _0403_
rlabel metal1 17250 30736 17250 30736 0 _0404_
rlabel metal1 19596 28594 19596 28594 0 _0405_
rlabel metal2 21850 29376 21850 29376 0 _0406_
rlabel metal1 24012 31994 24012 31994 0 _0407_
rlabel metal1 21068 32198 21068 32198 0 _0408_
rlabel metal1 19336 30634 19336 30634 0 _0409_
rlabel metal2 18446 30226 18446 30226 0 _0410_
rlabel metal1 19964 29750 19964 29750 0 _0411_
rlabel metal2 20194 30158 20194 30158 0 _0412_
rlabel via2 19274 29563 19274 29563 0 _0413_
rlabel metal1 18492 35258 18492 35258 0 _0414_
rlabel metal1 25898 36176 25898 36176 0 _0415_
rlabel metal1 19366 33966 19366 33966 0 _0416_
rlabel metal1 21114 34714 21114 34714 0 _0417_
rlabel metal1 21252 35802 21252 35802 0 _0418_
rlabel metal1 21850 33082 21850 33082 0 _0419_
rlabel metal1 22448 35802 22448 35802 0 _0420_
rlabel metal2 22954 36550 22954 36550 0 _0421_
rlabel metal1 22448 35258 22448 35258 0 _0422_
rlabel metal1 20838 33932 20838 33932 0 _0423_
rlabel metal1 20102 34068 20102 34068 0 _0424_
rlabel metal1 21298 35088 21298 35088 0 _0425_
rlabel metal1 21114 33422 21114 33422 0 _0426_
rlabel metal1 20286 33626 20286 33626 0 _0427_
rlabel metal1 24288 36142 24288 36142 0 _0428_
rlabel metal1 26358 35258 26358 35258 0 _0429_
rlabel metal1 27646 36346 27646 36346 0 _0430_
rlabel metal1 25806 35802 25806 35802 0 _0431_
rlabel metal2 26082 36788 26082 36788 0 _0432_
rlabel metal1 28198 35700 28198 35700 0 _0433_
rlabel metal1 28290 35802 28290 35802 0 _0434_
rlabel metal1 29256 35802 29256 35802 0 _0435_
rlabel metal1 30084 35802 30084 35802 0 _0436_
rlabel metal1 28152 34170 28152 34170 0 _0437_
rlabel metal1 25806 32436 25806 32436 0 _0438_
rlabel metal1 27508 32402 27508 32402 0 _0439_
rlabel metal1 28106 32266 28106 32266 0 _0440_
rlabel metal1 26657 32402 26657 32402 0 _0441_
rlabel metal1 18722 34680 18722 34680 0 _0442_
rlabel metal1 30130 35224 30130 35224 0 _0443_
rlabel metal2 18262 37468 18262 37468 0 _0444_
rlabel via2 13754 39389 13754 39389 0 _0445_
rlabel via2 17618 36771 17618 36771 0 _0446_
rlabel metal1 31832 36346 31832 36346 0 _0447_
rlabel metal1 30360 39338 30360 39338 0 _0448_
rlabel via2 18906 37213 18906 37213 0 _0449_
rlabel metal1 30866 31824 30866 31824 0 _0450_
rlabel metal2 31786 31722 31786 31722 0 _0451_
rlabel metal2 31786 33235 31786 33235 0 _0452_
rlabel metal1 32016 33830 32016 33830 0 _0453_
rlabel via1 31063 31722 31063 31722 0 _0454_
rlabel metal2 6118 3740 6118 3740 0 _0455_
rlabel metal2 2162 34306 2162 34306 0 _0456_
rlabel metal2 15778 3026 15778 3026 0 _0457_
rlabel metal1 2070 6970 2070 6970 0 _0458_
rlabel metal2 32706 3604 32706 3604 0 _0459_
rlabel metal2 5842 3400 5842 3400 0 _0460_
rlabel metal1 32706 19448 32706 19448 0 _0461_
rlabel metal2 6762 4012 6762 4012 0 _0462_
rlabel metal1 21850 34136 21850 34136 0 _0463_
rlabel metal2 30038 37247 30038 37247 0 _0464_
rlabel metal1 32016 12138 32016 12138 0 _0465_
rlabel metal2 17066 2788 17066 2788 0 _0466_
rlabel metal1 27048 39474 27048 39474 0 _0467_
rlabel metal1 5658 38216 5658 38216 0 _0468_
rlabel metal2 17066 39134 17066 39134 0 _0469_
rlabel metal1 5796 5270 5796 5270 0 _0470_
rlabel metal2 32706 16218 32706 16218 0 _0471_
rlabel metal1 32292 31382 32292 31382 0 _0472_
rlabel metal1 5474 39372 5474 39372 0 _0473_
rlabel metal2 32706 21879 32706 21879 0 _0474_
rlabel metal2 2622 8228 2622 8228 0 _0475_
rlabel via2 25346 37893 25346 37893 0 _0476_
rlabel metal2 20194 38114 20194 38114 0 _0477_
rlabel via1 9338 2363 9338 2363 0 _0478_
rlabel metal2 31050 16150 31050 16150 0 _0479_
rlabel metal1 3496 4046 3496 4046 0 _0480_
rlabel metal1 32982 6834 32982 6834 0 _0481_
rlabel metal1 2944 37162 2944 37162 0 _0482_
rlabel metal1 29348 2618 29348 2618 0 _0483_
rlabel metal1 5060 2346 5060 2346 0 _0484_
rlabel metal1 33212 11322 33212 11322 0 _0485_
rlabel metal2 20746 36992 20746 36992 0 _0486_
rlabel metal2 24518 38080 24518 38080 0 _0487_
rlabel metal2 22218 39134 22218 39134 0 _0488_
rlabel metal2 4370 3502 4370 3502 0 _0489_
rlabel metal1 1932 34170 1932 34170 0 _0490_
rlabel metal1 16422 25126 16422 25126 0 _0491_
rlabel metal1 14444 38522 14444 38522 0 _0492_
rlabel metal2 21390 37859 21390 37859 0 _0493_
rlabel metal1 2024 15130 2024 15130 0 _0494_
rlabel metal2 14490 3230 14490 3230 0 _0495_
rlabel metal2 1978 11934 1978 11934 0 _0496_
rlabel via2 32706 23613 32706 23613 0 _0497_
rlabel metal1 2392 3434 2392 3434 0 _0498_
rlabel metal1 2944 5746 2944 5746 0 _0499_
rlabel metal1 29624 2346 29624 2346 0 _0500_
rlabel metal2 32338 35241 32338 35241 0 _0501_
rlabel metal2 6670 27234 6670 27234 0 _0502_
rlabel via2 31878 13515 31878 13515 0 _0503_
rlabel metal2 32614 39406 32614 39406 0 _0504_
rlabel metal1 29302 3706 29302 3706 0 _0505_
rlabel metal1 2070 17850 2070 17850 0 _0506_
rlabel metal2 29670 39134 29670 39134 0 _0507_
rlabel metal2 2162 31076 2162 31076 0 _0508_
rlabel metal2 24058 3230 24058 3230 0 _0509_
rlabel metal1 31786 20808 31786 20808 0 _0510_
rlabel metal2 22126 3298 22126 3298 0 _0511_
rlabel metal2 25162 38080 25162 38080 0 _0512_
rlabel metal1 1840 4658 1840 4658 0 _0513_
rlabel metal1 27324 37706 27324 37706 0 _0514_
rlabel metal2 13294 3604 13294 3604 0 _0515_
rlabel metal1 33396 5270 33396 5270 0 _0516_
rlabel metal1 1978 5304 1978 5304 0 _0517_
rlabel metal2 2070 10404 2070 10404 0 _0518_
rlabel metal1 3818 36822 3818 36822 0 _0519_
rlabel metal2 33902 8228 33902 8228 0 _0520_
rlabel metal1 32223 34646 32223 34646 0 _0521_
rlabel metal1 32223 35122 32223 35122 0 _0522_
rlabel metal1 8924 38522 8924 38522 0 _0523_
rlabel metal2 30130 37672 30130 37672 0 _0524_
rlabel metal2 19826 4318 19826 4318 0 _0525_
rlabel metal1 29486 3094 29486 3094 0 _0526_
rlabel metal1 20930 36720 20930 36720 0 _0527_
rlabel metal1 19596 2618 19596 2618 0 _0528_
rlabel metal2 32706 5644 32706 5644 0 _0529_
rlabel metal1 1978 24922 1978 24922 0 _0530_
rlabel metal1 32706 17272 32706 17272 0 _0531_
rlabel metal1 6164 38522 6164 38522 0 _0532_
rlabel metal1 2070 3128 2070 3128 0 _0533_
rlabel metal2 7222 3502 7222 3502 0 _0534_
rlabel metal1 2070 12954 2070 12954 0 _0535_
rlabel metal2 17618 35037 17618 35037 0 _0536_
rlabel metal1 33304 10778 33304 10778 0 _0537_
rlabel metal1 31878 13974 31878 13974 0 _0538_
rlabel metal2 1978 6494 1978 6494 0 _0539_
rlabel metal2 7222 38114 7222 38114 0 _0540_
rlabel metal1 32200 6358 32200 6358 0 _0541_
rlabel metal1 9660 3094 9660 3094 0 _0542_
rlabel metal2 24610 39134 24610 39134 0 _0543_
rlabel metal2 8142 38318 8142 38318 0 _0544_
rlabel metal1 32614 15130 32614 15130 0 _0545_
rlabel metal2 3266 38590 3266 38590 0 _0546_
rlabel metal1 4508 4658 4508 4658 0 _0547_
rlabel metal2 15226 38692 15226 38692 0 _0548_
rlabel metal2 16606 38828 16606 38828 0 _0549_
rlabel metal1 32430 5610 32430 5610 0 _0550_
rlabel metal2 28566 34017 28566 34017 0 _0551_
rlabel metal1 19090 38522 19090 38522 0 _0552_
rlabel metal2 30222 2584 30222 2584 0 _0553_
rlabel metal1 18078 31654 18078 31654 0 _0554_
rlabel metal1 5888 36686 5888 36686 0 _0555_
rlabel metal2 32522 3230 32522 3230 0 _0556_
rlabel metal2 1978 19550 1978 19550 0 _0557_
rlabel metal1 31142 3434 31142 3434 0 _0558_
rlabel metal2 5566 38420 5566 38420 0 _0559_
rlabel metal2 2622 16932 2622 16932 0 _0560_
rlabel metal1 2208 9010 2208 9010 0 _0561_
rlabel metal2 1794 14620 1794 14620 0 _0562_
rlabel metal3 1786 36108 1786 36108 0 active
rlabel metal1 20884 20910 20884 20910 0 clknet_0_wb_clk_i
rlabel metal2 19458 20876 19458 20876 0 clknet_3_0__leaf_wb_clk_i
rlabel metal1 21988 20434 21988 20434 0 clknet_3_1__leaf_wb_clk_i
rlabel metal1 32844 21522 32844 21522 0 clknet_3_2__leaf_wb_clk_i
rlabel metal2 32338 24480 32338 24480 0 clknet_3_3__leaf_wb_clk_i
rlabel metal1 22034 30090 22034 30090 0 clknet_3_4__leaf_wb_clk_i
rlabel metal1 18216 33490 18216 33490 0 clknet_3_5__leaf_wb_clk_i
rlabel metal1 32982 27540 32982 27540 0 clknet_3_6__leaf_wb_clk_i
rlabel metal1 28336 32878 28336 32878 0 clknet_3_7__leaf_wb_clk_i
rlabel metal1 18814 39406 18814 39406 0 io_in[10]
rlabel metal3 2108 38828 2108 38828 0 io_in[11]
rlabel metal1 21482 36720 21482 36720 0 io_in[12]
rlabel metal2 18078 1095 18078 1095 0 io_in[13]
rlabel metal1 16422 29716 16422 29716 0 io_in[8]
rlabel metal1 6854 37264 6854 37264 0 io_in[9]
rlabel metal2 20654 2404 20654 2404 0 io_oeb[0]
rlabel metal3 1740 13668 1740 13668 0 io_oeb[10]
rlabel metal3 34784 25228 34784 25228 0 io_oeb[11]
rlabel metal3 34784 14348 34784 14348 0 io_oeb[12]
rlabel metal3 34784 13668 34784 13668 0 io_oeb[13]
rlabel metal3 1786 3468 1786 3468 0 io_oeb[14]
rlabel metal2 7774 39824 7774 39824 0 io_oeb[15]
rlabel metal2 34362 5525 34362 5525 0 io_oeb[16]
rlabel metal2 10350 1860 10350 1860 0 io_oeb[17]
rlabel metal2 25162 40062 25162 40062 0 io_oeb[18]
rlabel metal1 9430 37842 9430 37842 0 io_oeb[19]
rlabel metal2 30314 1860 30314 1860 0 io_oeb[1]
rlabel metal3 34784 19788 34784 19788 0 io_oeb[20]
rlabel metal1 3496 37774 3496 37774 0 io_oeb[21]
rlabel metal2 3910 1826 3910 1826 0 io_oeb[22]
rlabel metal2 16146 40062 16146 40062 0 io_oeb[23]
rlabel metal2 17434 39824 17434 39824 0 io_oeb[24]
rlabel metal1 34500 5610 34500 5610 0 io_oeb[25]
rlabel metal3 34784 33388 34784 33388 0 io_oeb[26]
rlabel metal2 20010 40062 20010 40062 0 io_oeb[27]
rlabel metal2 32890 1622 32890 1622 0 io_oeb[28]
rlabel metal3 34784 27948 34784 27948 0 io_oeb[29]
rlabel metal2 29026 39518 29026 39518 0 io_oeb[2]
rlabel metal2 2806 40205 2806 40205 0 io_oeb[30]
rlabel metal2 32246 1826 32246 1826 0 io_oeb[31]
rlabel metal3 1464 19108 1464 19108 0 io_oeb[32]
rlabel metal2 35926 2771 35926 2771 0 io_oeb[33]
rlabel metal2 5842 40062 5842 40062 0 io_oeb[34]
rlabel metal3 1740 17068 1740 17068 0 io_oeb[35]
rlabel metal3 1740 8908 1740 8908 0 io_oeb[36]
rlabel metal3 1740 14348 1740 14348 0 io_oeb[37]
rlabel metal2 20010 1860 20010 1860 0 io_oeb[3]
rlabel metal3 34784 3468 34784 3468 0 io_oeb[4]
rlabel metal3 1740 25228 1740 25228 0 io_oeb[5]
rlabel metal3 34784 17068 34784 17068 0 io_oeb[6]
rlabel metal2 7130 40368 7130 40368 0 io_oeb[7]
rlabel metal2 3266 1860 3266 1860 0 io_oeb[8]
rlabel metal2 8418 1860 8418 1860 0 io_oeb[9]
rlabel metal2 32246 38913 32246 38913 0 io_out[0]
rlabel metal3 34830 24548 34830 24548 0 io_out[10]
rlabel metal3 1740 2108 1740 2108 0 io_out[11]
rlabel metal3 2062 5508 2062 5508 0 io_out[12]
rlabel metal2 30958 1622 30958 1622 0 io_out[13]
rlabel metal3 34830 34068 34830 34068 0 io_out[14]
rlabel metal3 2108 32028 2108 32028 0 io_out[15]
rlabel metal2 34362 23919 34362 23919 0 io_out[16]
rlabel metal2 32890 40062 32890 40062 0 io_out[17]
rlabel metal1 31832 4046 31832 4046 0 io_out[18]
rlabel metal2 2806 18309 2806 18309 0 io_out[19]
rlabel metal2 22586 40062 22586 40062 0 io_out[1]
rlabel metal1 29946 38828 29946 38828 0 io_out[20]
rlabel metal3 1740 31348 1740 31348 0 io_out[21]
rlabel metal2 24518 1860 24518 1860 0 io_out[22]
rlabel metal3 34784 20468 34784 20468 0 io_out[23]
rlabel metal2 21298 2166 21298 2166 0 io_out[24]
rlabel metal1 26358 38420 26358 38420 0 io_out[25]
rlabel metal3 1740 4148 1740 4148 0 io_out[26]
rlabel metal1 27600 38862 27600 38862 0 io_out[27]
rlabel metal2 13570 1503 13570 1503 0 io_out[28]
rlabel metal2 33074 4641 33074 4641 0 io_out[29]
rlabel metal2 5198 1231 5198 1231 0 io_out[2]
rlabel metal3 1740 4828 1740 4828 0 io_out[30]
rlabel metal2 2806 10761 2806 10761 0 io_out[31]
rlabel metal3 1740 36788 1740 36788 0 io_out[32]
rlabel metal3 34784 8908 34784 8908 0 io_out[33]
rlabel metal3 35198 34748 35198 34748 0 io_out[34]
rlabel metal1 34500 34986 34500 34986 0 io_out[35]
rlabel metal2 9062 40062 9062 40062 0 io_out[36]
rlabel metal3 35198 38148 35198 38148 0 io_out[37]
rlabel metal3 1740 34068 1740 34068 0 io_out[3]
rlabel metal3 34784 25908 34784 25908 0 io_out[4]
rlabel metal2 14858 40368 14858 40368 0 io_out[5]
rlabel metal2 34178 39824 34178 39824 0 io_out[6]
rlabel metal2 2806 15623 2806 15623 0 io_out[7]
rlabel metal2 14858 1860 14858 1860 0 io_out[8]
rlabel metal3 1740 11628 1740 11628 0 io_out[9]
rlabel metal2 34086 9809 34086 9809 0 la1_data_in[0]
rlabel metal2 6486 2166 6486 2166 0 la1_data_out[0]
rlabel metal3 34784 12308 34784 12308 0 la1_data_out[10]
rlabel metal2 17434 1860 17434 1860 0 la1_data_out[11]
rlabel metal3 34784 38828 34784 38828 0 la1_data_out[12]
rlabel metal1 2070 38250 2070 38250 0 la1_data_out[13]
rlabel metal2 18078 40657 18078 40657 0 la1_data_out[14]
rlabel metal3 2384 1428 2384 1428 0 la1_data_out[15]
rlabel metal1 34776 16490 34776 16490 0 la1_data_out[16]
rlabel metal3 34784 31348 34784 31348 0 la1_data_out[17]
rlabel metal1 2392 39338 2392 39338 0 la1_data_out[18]
rlabel metal3 34784 23188 34784 23188 0 la1_data_out[19]
rlabel metal2 2806 35275 2806 35275 0 la1_data_out[1]
rlabel metal3 1740 8228 1740 8228 0 la1_data_out[20]
rlabel metal3 34784 36788 34784 36788 0 la1_data_out[21]
rlabel metal1 20700 38386 20700 38386 0 la1_data_out[22]
rlabel metal2 9706 1027 9706 1027 0 la1_data_out[23]
rlabel metal3 34784 17748 34784 17748 0 la1_data_out[24]
rlabel metal3 2338 2788 2338 2788 0 la1_data_out[25]
rlabel metal3 34784 6868 34784 6868 0 la1_data_out[26]
rlabel metal2 2070 37383 2070 37383 0 la1_data_out[27]
rlabel metal1 32062 4488 32062 4488 0 la1_data_out[28]
rlabel metal2 4554 1622 4554 1622 0 la1_data_out[29]
rlabel metal2 16146 2166 16146 2166 0 la1_data_out[2]
rlabel metal3 35198 12988 35198 12988 0 la1_data_out[30]
rlabel metal3 34140 40868 34140 40868 0 la1_data_out[31]
rlabel metal2 2806 7429 2806 7429 0 la1_data_out[3]
rlabel metal2 35466 2404 35466 2404 0 la1_data_out[4]
rlabel metal2 2622 1622 2622 1622 0 la1_data_out[5]
rlabel metal3 34784 19108 34784 19108 0 la1_data_out[6]
rlabel metal2 690 1792 690 1792 0 la1_data_out[7]
rlabel metal3 34784 32028 34784 32028 0 la1_data_out[8]
rlabel metal2 33534 38974 33534 38974 0 la1_data_out[9]
rlabel metal1 1656 33082 1656 33082 0 net1
rlabel metal2 2898 34204 2898 34204 0 net10
rlabel metal1 16192 38318 16192 38318 0 net100
rlabel metal2 28842 4930 28842 4930 0 net101
rlabel metal2 23506 34952 23506 34952 0 net102
rlabel metal2 19182 39168 19182 39168 0 net103
rlabel metal2 31694 3196 31694 3196 0 net104
rlabel metal1 18722 37298 18722 37298 0 net105
rlabel metal2 4002 38080 4002 38080 0 net106
rlabel metal1 32936 2958 32936 2958 0 net107
rlabel metal1 1932 18938 1932 18938 0 net108
rlabel metal1 31142 3570 31142 3570 0 net109
rlabel metal2 15594 3740 15594 3740 0 net11
rlabel metal2 4186 39168 4186 39168 0 net110
rlabel metal1 1932 16762 1932 16762 0 net111
rlabel metal2 1610 9180 1610 9180 0 net112
rlabel metal1 1840 13430 1840 13430 0 net113
rlabel metal2 1794 7582 1794 7582 0 net12
rlabel metal2 31326 4896 31326 4896 0 net13
rlabel metal1 2944 2550 2944 2550 0 net14
rlabel metal2 32154 17136 32154 17136 0 net15
rlabel metal1 6578 2516 6578 2516 0 net16
rlabel metal1 32522 32436 32522 32436 0 net17
rlabel metal2 25714 37383 25714 37383 0 net18
rlabel metal2 33350 11458 33350 11458 0 net19
rlabel metal2 18354 37162 18354 37162 0 net2
rlabel metal2 16882 3468 16882 3468 0 net20
rlabel metal1 20286 37434 20286 37434 0 net21
rlabel metal1 1610 38420 1610 38420 0 net22
rlabel metal1 17756 37842 17756 37842 0 net23
rlabel metal1 4508 5134 4508 5134 0 net24
rlabel metal1 32798 11730 32798 11730 0 net25
rlabel metal1 32154 37740 32154 37740 0 net26
rlabel metal1 1610 39508 1610 39508 0 net27
rlabel via2 33994 11747 33994 11747 0 net28
rlabel metal1 1932 8058 1932 8058 0 net29
rlabel metal2 16698 36924 16698 36924 0 net3
rlabel metal2 22494 36805 22494 36805 0 net30
rlabel metal1 20148 38386 20148 38386 0 net31
rlabel metal1 9246 2482 9246 2482 0 net32
rlabel metal1 33304 11730 33304 11730 0 net33
rlabel metal1 2622 4012 2622 4012 0 net34
rlabel metal1 33258 6698 33258 6698 0 net35
rlabel metal1 1610 37162 1610 37162 0 net36
rlabel metal1 29716 4590 29716 4590 0 net37
rlabel metal2 4186 2992 4186 2992 0 net38
rlabel metal1 31970 12750 31970 12750 0 net39
rlabel metal1 26542 36652 26542 36652 0 net4
rlabel via2 20654 36669 20654 36669 0 net40
rlabel metal2 29394 38454 29394 38454 0 net41
rlabel metal1 22448 38522 22448 38522 0 net42
rlabel metal1 4508 2958 4508 2958 0 net43
rlabel metal1 1886 36142 1886 36142 0 net44
rlabel metal1 15686 25942 15686 25942 0 net45
rlabel metal2 14030 39168 14030 39168 0 net46
rlabel metal1 32522 38284 32522 38284 0 net47
rlabel metal2 1610 15708 1610 15708 0 net48
rlabel metal2 14306 3264 14306 3264 0 net49
rlabel metal1 18630 2618 18630 2618 0 net5
rlabel metal2 2070 11492 2070 11492 0 net50
rlabel via2 33810 15011 33810 15011 0 net51
rlabel metal1 1610 3604 1610 3604 0 net52
rlabel metal2 1610 5916 1610 5916 0 net53
rlabel metal1 30176 2482 30176 2482 0 net54
rlabel metal1 32085 38930 32085 38930 0 net55
rlabel metal2 27922 3876 27922 3876 0 net56
rlabel metal2 1794 18496 1794 18496 0 net57
rlabel metal2 18998 38726 18998 38726 0 net58
rlabel metal2 1794 31552 1794 31552 0 net59
rlabel metal2 16238 31688 16238 31688 0 net6
rlabel metal1 23874 3094 23874 3094 0 net60
rlabel metal2 32614 17204 32614 17204 0 net61
rlabel metal1 20884 2618 20884 2618 0 net62
rlabel metal1 25530 38386 25530 38386 0 net63
rlabel metal1 1610 4692 1610 4692 0 net64
rlabel metal1 20378 36754 20378 36754 0 net65
rlabel metal2 13110 3876 13110 3876 0 net66
rlabel metal1 32292 5202 32292 5202 0 net67
rlabel metal1 1932 4114 1932 4114 0 net68
rlabel metal2 1794 10880 1794 10880 0 net69
rlabel metal1 6762 37128 6762 37128 0 net7
rlabel metal1 1794 36822 1794 36822 0 net70
rlabel metal2 32522 8704 32522 8704 0 net71
rlabel metal2 32522 34867 32522 34867 0 net72
rlabel metal1 23506 37230 23506 37230 0 net73
rlabel metal1 8188 38862 8188 38862 0 net74
rlabel metal2 21482 37468 21482 37468 0 net75
rlabel metal2 20286 3876 20286 3876 0 net76
rlabel metal2 29670 3264 29670 3264 0 net77
rlabel metal1 28014 37842 28014 37842 0 net78
rlabel metal2 19458 3264 19458 3264 0 net79
rlabel metal2 34270 12818 34270 12818 0 net8
rlabel metal1 32200 4658 32200 4658 0 net80
rlabel metal2 1610 25500 1610 25500 0 net81
rlabel metal1 32154 14586 32154 14586 0 net82
rlabel metal1 6302 39406 6302 39406 0 net83
rlabel metal1 2484 2958 2484 2958 0 net84
rlabel metal2 7038 3230 7038 3230 0 net85
rlabel metal1 2254 13498 2254 13498 0 net86
rlabel via2 29027 25381 29027 25381 0 net87
rlabel metal1 31510 14450 31510 14450 0 net88
rlabel metal1 32292 12410 32292 12410 0 net89
rlabel metal1 5704 3502 5704 3502 0 net9
rlabel metal2 1794 6494 1794 6494 0 net90
rlabel metal1 6532 38318 6532 38318 0 net91
rlabel metal1 32936 6222 32936 6222 0 net92
rlabel metal1 9706 2958 9706 2958 0 net93
rlabel metal2 24426 39134 24426 39134 0 net94
rlabel metal1 8648 37774 8648 37774 0 net95
rlabel metal1 33718 11322 33718 11322 0 net96
rlabel metal1 4692 37434 4692 37434 0 net97
rlabel metal2 5566 4284 5566 4284 0 net98
rlabel metal2 15686 38318 15686 38318 0 net99
rlabel metal1 32338 30056 32338 30056 0 rgb_mixer0.debounce0_a.button_hist\[0\]
rlabel metal1 31602 32436 31602 32436 0 rgb_mixer0.debounce0_a.button_hist\[1\]
rlabel metal2 31326 32521 31326 32521 0 rgb_mixer0.debounce0_a.button_hist\[2\]
rlabel metal2 31510 34850 31510 34850 0 rgb_mixer0.debounce0_a.button_hist\[3\]
rlabel metal1 31694 34136 31694 34136 0 rgb_mixer0.debounce0_a.button_hist\[4\]
rlabel metal1 31464 34714 31464 34714 0 rgb_mixer0.debounce0_a.button_hist\[5\]
rlabel metal2 31142 35190 31142 35190 0 rgb_mixer0.debounce0_a.button_hist\[6\]
rlabel metal2 31326 33830 31326 33830 0 rgb_mixer0.debounce0_a.button_hist\[7\]
rlabel metal1 29256 34510 29256 34510 0 rgb_mixer0.debounce0_a.debounced
rlabel metal2 26542 35258 26542 35258 0 rgb_mixer0.debounce0_b.button_hist\[0\]
rlabel metal1 27048 35598 27048 35598 0 rgb_mixer0.debounce0_b.button_hist\[1\]
rlabel metal1 27646 33830 27646 33830 0 rgb_mixer0.debounce0_b.button_hist\[2\]
rlabel metal1 25944 34918 25944 34918 0 rgb_mixer0.debounce0_b.button_hist\[3\]
rlabel metal2 28566 35156 28566 35156 0 rgb_mixer0.debounce0_b.button_hist\[4\]
rlabel metal2 28290 33150 28290 33150 0 rgb_mixer0.debounce0_b.button_hist\[5\]
rlabel metal2 29210 34442 29210 34442 0 rgb_mixer0.debounce0_b.button_hist\[6\]
rlabel metal1 28474 32334 28474 32334 0 rgb_mixer0.debounce0_b.button_hist\[7\]
rlabel metal2 26450 29104 26450 29104 0 rgb_mixer0.debounce0_b.debounced
rlabel metal2 20470 34204 20470 34204 0 rgb_mixer0.debounce1_a.button_hist\[0\]
rlabel metal2 20286 34850 20286 34850 0 rgb_mixer0.debounce1_a.button_hist\[1\]
rlabel metal2 20654 34816 20654 34816 0 rgb_mixer0.debounce1_a.button_hist\[2\]
rlabel metal1 21482 32844 21482 32844 0 rgb_mixer0.debounce1_a.button_hist\[3\]
rlabel metal2 22954 35428 22954 35428 0 rgb_mixer0.debounce1_a.button_hist\[4\]
rlabel metal1 23046 34714 23046 34714 0 rgb_mixer0.debounce1_a.button_hist\[5\]
rlabel metal1 23363 33830 23363 33830 0 rgb_mixer0.debounce1_a.button_hist\[6\]
rlabel metal2 23138 34680 23138 34680 0 rgb_mixer0.debounce1_a.button_hist\[7\]
rlabel metal1 19918 32334 19918 32334 0 rgb_mixer0.debounce1_a.debounced
rlabel metal1 19688 31858 19688 31858 0 rgb_mixer0.debounce1_b.button_hist\[0\]
rlabel metal2 18538 31178 18538 31178 0 rgb_mixer0.debounce1_b.button_hist\[1\]
rlabel metal1 19458 32198 19458 32198 0 rgb_mixer0.debounce1_b.button_hist\[2\]
rlabel metal2 19550 29274 19550 29274 0 rgb_mixer0.debounce1_b.button_hist\[3\]
rlabel metal1 20746 31314 20746 31314 0 rgb_mixer0.debounce1_b.button_hist\[4\]
rlabel metal2 21390 30770 21390 30770 0 rgb_mixer0.debounce1_b.button_hist\[5\]
rlabel metal1 21436 30906 21436 30906 0 rgb_mixer0.debounce1_b.button_hist\[6\]
rlabel metal1 22448 31654 22448 31654 0 rgb_mixer0.debounce1_b.button_hist\[7\]
rlabel metal1 19817 29648 19817 29648 0 rgb_mixer0.debounce1_b.debounced
rlabel metal1 29486 32878 29486 32878 0 rgb_mixer0.debounce2_a.button_hist\[0\]
rlabel metal3 25484 31892 25484 31892 0 rgb_mixer0.debounce2_a.button_hist\[1\]
rlabel metal2 25530 31926 25530 31926 0 rgb_mixer0.debounce2_a.button_hist\[2\]
rlabel metal1 24610 32436 24610 32436 0 rgb_mixer0.debounce2_a.button_hist\[3\]
rlabel metal1 24564 31994 24564 31994 0 rgb_mixer0.debounce2_a.button_hist\[4\]
rlabel metal1 23414 30838 23414 30838 0 rgb_mixer0.debounce2_a.button_hist\[5\]
rlabel metal1 25070 34578 25070 34578 0 rgb_mixer0.debounce2_a.button_hist\[6\]
rlabel metal2 24702 32028 24702 32028 0 rgb_mixer0.debounce2_a.button_hist\[7\]
rlabel metal1 25116 32810 25116 32810 0 rgb_mixer0.debounce2_a.debounced
rlabel metal1 21459 27302 21459 27302 0 rgb_mixer0.debounce2_b.button_hist\[0\]
rlabel metal1 23184 27302 23184 27302 0 rgb_mixer0.debounce2_b.button_hist\[1\]
rlabel metal1 23552 28186 23552 28186 0 rgb_mixer0.debounce2_b.button_hist\[2\]
rlabel metal1 21206 28084 21206 28084 0 rgb_mixer0.debounce2_b.button_hist\[3\]
rlabel metal2 22862 26316 22862 26316 0 rgb_mixer0.debounce2_b.button_hist\[4\]
rlabel metal1 22632 25126 22632 25126 0 rgb_mixer0.debounce2_b.button_hist\[5\]
rlabel metal2 22678 23868 22678 23868 0 rgb_mixer0.debounce2_b.button_hist\[6\]
rlabel metal1 23092 25262 23092 25262 0 rgb_mixer0.debounce2_b.button_hist\[7\]
rlabel metal1 24702 26486 24702 26486 0 rgb_mixer0.debounce2_b.debounced
rlabel metal1 15962 25330 15962 25330 0 rgb_mixer0.enc0\[0\]
rlabel metal2 17066 27846 17066 27846 0 rgb_mixer0.enc0\[1\]
rlabel metal1 29900 39406 29900 39406 0 rgb_mixer0.enc0\[2\]
rlabel metal1 31878 26316 31878 26316 0 rgb_mixer0.enc0\[3\]
rlabel metal1 33718 26214 33718 26214 0 rgb_mixer0.enc0\[4\]
rlabel metal1 32890 26962 32890 26962 0 rgb_mixer0.enc0\[5\]
rlabel metal2 31970 26741 31970 26741 0 rgb_mixer0.enc0\[6\]
rlabel metal2 31418 25126 31418 25126 0 rgb_mixer0.enc0\[7\]
rlabel metal2 18814 26146 18814 26146 0 rgb_mixer0.enc1\[0\]
rlabel metal1 17434 26350 17434 26350 0 rgb_mixer0.enc1\[1\]
rlabel metal1 21160 21998 21160 21998 0 rgb_mixer0.enc1\[2\]
rlabel metal2 17526 23052 17526 23052 0 rgb_mixer0.enc1\[3\]
rlabel metal1 16146 21964 16146 21964 0 rgb_mixer0.enc1\[4\]
rlabel metal2 19366 19516 19366 19516 0 rgb_mixer0.enc1\[5\]
rlabel metal1 21252 21522 21252 21522 0 rgb_mixer0.enc1\[6\]
rlabel metal1 21114 19958 21114 19958 0 rgb_mixer0.enc1\[7\]
rlabel metal1 19918 20842 19918 20842 0 rgb_mixer0.enc2\[0\]
rlabel metal1 28934 22712 28934 22712 0 rgb_mixer0.enc2\[1\]
rlabel metal1 27876 21318 27876 21318 0 rgb_mixer0.enc2\[2\]
rlabel metal2 26358 20128 26358 20128 0 rgb_mixer0.enc2\[3\]
rlabel metal1 28796 19278 28796 19278 0 rgb_mixer0.enc2\[4\]
rlabel metal2 30222 19244 30222 19244 0 rgb_mixer0.enc2\[5\]
rlabel metal1 27462 16116 27462 16116 0 rgb_mixer0.enc2\[6\]
rlabel metal2 28474 16898 28474 16898 0 rgb_mixer0.enc2\[7\]
rlabel metal2 34086 30906 34086 30906 0 rgb_mixer0.encoder0.old_a
rlabel metal3 27991 35972 27991 35972 0 rgb_mixer0.encoder0.old_b
rlabel metal1 18722 27030 18722 27030 0 rgb_mixer0.encoder1.old_a
rlabel metal2 18538 27404 18538 27404 0 rgb_mixer0.encoder1.old_b
rlabel metal1 26864 26758 26864 26758 0 rgb_mixer0.encoder2.old_a
rlabel metal1 26818 31314 26818 31314 0 rgb_mixer0.encoder2.old_b
rlabel via1 31886 20774 31886 20774 0 rgb_mixer0.pwm0.count\[0\]
rlabel metal2 32430 20876 32430 20876 0 rgb_mixer0.pwm0.count\[1\]
rlabel metal1 31694 20876 31694 20876 0 rgb_mixer0.pwm0.count\[2\]
rlabel metal1 33718 18258 33718 18258 0 rgb_mixer0.pwm0.count\[3\]
rlabel metal1 32430 17510 32430 17510 0 rgb_mixer0.pwm0.count\[4\]
rlabel metal2 33810 16218 33810 16218 0 rgb_mixer0.pwm0.count\[5\]
rlabel metal1 30268 18258 30268 18258 0 rgb_mixer0.pwm0.count\[6\]
rlabel metal2 30820 19890 30820 19890 0 rgb_mixer0.pwm0.count\[7\]
rlabel metal2 22034 34034 22034 34034 0 rgb_mixer0.pwm0.out
rlabel metal1 20976 18190 20976 18190 0 rgb_mixer0.pwm1.count\[0\]
rlabel metal2 20838 19890 20838 19890 0 rgb_mixer0.pwm1.count\[1\]
rlabel metal2 20700 19346 20700 19346 0 rgb_mixer0.pwm1.count\[2\]
rlabel metal2 22126 15980 22126 15980 0 rgb_mixer0.pwm1.count\[3\]
rlabel metal1 21022 19380 21022 19380 0 rgb_mixer0.pwm1.count\[4\]
rlabel metal1 20792 22202 20792 22202 0 rgb_mixer0.pwm1.count\[5\]
rlabel metal1 20010 21930 20010 21930 0 rgb_mixer0.pwm1.count\[6\]
rlabel metal1 25162 23086 25162 23086 0 rgb_mixer0.pwm1.count\[7\]
rlabel metal1 8234 27098 8234 27098 0 rgb_mixer0.pwm1.out
rlabel metal2 20378 19822 20378 19822 0 rgb_mixer0.pwm2.count\[0\]
rlabel metal1 20286 20944 20286 20944 0 rgb_mixer0.pwm2.count\[1\]
rlabel metal2 25990 17034 25990 17034 0 rgb_mixer0.pwm2.count\[2\]
rlabel metal1 25254 18156 25254 18156 0 rgb_mixer0.pwm2.count\[3\]
rlabel metal2 25530 15470 25530 15470 0 rgb_mixer0.pwm2.count\[4\]
rlabel metal1 25530 16490 25530 16490 0 rgb_mixer0.pwm2.count\[5\]
rlabel metal2 26174 17034 26174 17034 0 rgb_mixer0.pwm2.count\[6\]
rlabel metal1 27600 16558 27600 16558 0 rgb_mixer0.pwm2.count\[7\]
rlabel via2 33626 13515 33626 13515 0 rgb_mixer0.pwm2.out
rlabel metal2 33074 21403 33074 21403 0 wb_clk_i
<< properties >>
string FIXED_BBOX 0 0 36000 42000
<< end >>
