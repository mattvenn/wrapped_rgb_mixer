VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_rgb_mixer
  CLASS BLOCK ;
  FOREIGN wrapped_rgb_mixer ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 300.000 ;
  PIN active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 296.000 26.130 300.000 ;
    END
  END active
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 0.720 300.000 1.320 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 79.600 300.000 80.200 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 87.080 300.000 87.680 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 95.240 300.000 95.840 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 102.720 300.000 103.320 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 110.880 300.000 111.480 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 119.040 300.000 119.640 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 126.520 300.000 127.120 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 134.680 300.000 135.280 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 142.160 300.000 142.760 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 150.320 300.000 150.920 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 8.200 300.000 8.800 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 158.480 300.000 159.080 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 165.960 300.000 166.560 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 174.120 300.000 174.720 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 181.600 300.000 182.200 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 189.760 300.000 190.360 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 197.920 300.000 198.520 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 205.400 300.000 206.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 213.560 300.000 214.160 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 221.040 300.000 221.640 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 229.200 300.000 229.800 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 16.360 300.000 16.960 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 237.360 300.000 237.960 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 244.840 300.000 245.440 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 253.000 300.000 253.600 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 260.480 300.000 261.080 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 268.640 300.000 269.240 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 276.800 300.000 277.400 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 284.280 300.000 284.880 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 292.440 300.000 293.040 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 23.840 300.000 24.440 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 32.000 300.000 32.600 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 40.160 300.000 40.760 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 47.640 300.000 48.240 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 55.800 300.000 56.400 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 63.280 300.000 63.880 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 71.440 300.000 72.040 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 5.480 300.000 6.080 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 84.360 300.000 84.960 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 92.520 300.000 93.120 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 100.680 300.000 101.280 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 108.160 300.000 108.760 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 116.320 300.000 116.920 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 123.800 300.000 124.400 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 131.960 300.000 132.560 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 140.120 300.000 140.720 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 147.600 300.000 148.200 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 155.760 300.000 156.360 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 13.640 300.000 14.240 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 163.240 300.000 163.840 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 171.400 300.000 172.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 179.560 300.000 180.160 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 187.040 300.000 187.640 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 195.200 300.000 195.800 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 202.680 300.000 203.280 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 210.840 300.000 211.440 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 219.000 300.000 219.600 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 226.480 300.000 227.080 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 234.640 300.000 235.240 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 21.120 300.000 21.720 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 242.120 300.000 242.720 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 250.280 300.000 250.880 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 258.440 300.000 259.040 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 265.920 300.000 266.520 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 274.080 300.000 274.680 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 281.560 300.000 282.160 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 289.720 300.000 290.320 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 297.880 300.000 298.480 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 29.280 300.000 29.880 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 37.440 300.000 38.040 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 44.920 300.000 45.520 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 53.080 300.000 53.680 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 60.560 300.000 61.160 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 68.720 300.000 69.320 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 76.880 300.000 77.480 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 2.760 300.000 3.360 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 81.640 300.000 82.240 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 89.800 300.000 90.400 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 97.960 300.000 98.560 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 105.440 300.000 106.040 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 113.600 300.000 114.200 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 121.080 300.000 121.680 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 129.240 300.000 129.840 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 137.400 300.000 138.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 144.880 300.000 145.480 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 153.040 300.000 153.640 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 10.920 300.000 11.520 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 160.520 300.000 161.120 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 168.680 300.000 169.280 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 176.840 300.000 177.440 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 184.320 300.000 184.920 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 192.480 300.000 193.080 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 200.640 300.000 201.240 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 208.120 300.000 208.720 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 216.280 300.000 216.880 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 223.760 300.000 224.360 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 231.920 300.000 232.520 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 19.080 300.000 19.680 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 240.080 300.000 240.680 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 247.560 300.000 248.160 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 255.720 300.000 256.320 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 263.200 300.000 263.800 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 271.360 300.000 271.960 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 279.520 300.000 280.120 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 287.000 300.000 287.600 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 295.160 300.000 295.760 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 26.560 300.000 27.160 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 34.720 300.000 35.320 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 42.200 300.000 42.800 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 50.360 300.000 50.960 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 58.520 300.000 59.120 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 66.000 300.000 66.600 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 74.160 300.000 74.760 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 0.000 54.190 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 0.000 58.790 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.110 0.000 63.390 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 0.000 72.590 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 0.000 82.250 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.570 0.000 86.850 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 0.000 91.450 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 0.000 96.050 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.370 0.000 100.650 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.430 0.000 105.710 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.030 0.000 110.310 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.630 0.000 114.910 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.830 0.000 124.110 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 0.000 133.770 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 0.000 138.370 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 0.000 147.570 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 0.000 25.670 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 0.000 30.730 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.350 0.000 152.630 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.810 0.000 199.090 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.870 0.000 204.150 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.470 0.000 208.750 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.070 0.000 213.350 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.670 0.000 217.950 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.330 0.000 227.610 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.530 0.000 236.810 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.130 0.000 241.410 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.950 0.000 157.230 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.730 0.000 246.010 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.330 0.000 250.610 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 0.000 255.670 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.990 0.000 260.270 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.590 0.000 264.870 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.190 0.000 269.470 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 0.000 274.070 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.850 0.000 279.130 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 0.000 283.730 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.050 0.000 288.330 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.550 0.000 161.830 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.650 0.000 292.930 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.250 0.000 297.530 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.150 0.000 166.430 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.350 0.000 175.630 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 0.000 185.290 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.610 0.000 189.890 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.210 0.000 194.490 4.000 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.680 4.000 152.280 ;
    END
  END la_oen[0]
  PIN la_oen[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 4.000 199.200 ;
    END
  END la_oen[10]
  PIN la_oen[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 203.360 4.000 203.960 ;
    END
  END la_oen[11]
  PIN la_oen[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.120 4.000 208.720 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.880 4.000 213.480 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.960 4.000 217.560 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.720 4.000 222.320 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 226.480 4.000 227.080 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.000 4.000 236.600 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.760 4.000 241.360 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 245.520 4.000 246.120 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.280 4.000 250.880 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.040 4.000 255.640 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.120 4.000 259.720 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 263.880 4.000 264.480 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.640 4.000 269.240 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 273.400 4.000 274.000 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.160 4.000 278.760 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.920 4.000 283.520 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.680 4.000 288.280 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.200 4.000 161.800 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.200 4.000 297.800 ;
    END
  END la_oen[31]
  PIN la_oen[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.960 4.000 166.560 ;
    END
  END la_oen[3]
  PIN la_oen[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.720 4.000 171.320 ;
    END
  END la_oen[4]
  PIN la_oen[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.800 4.000 175.400 ;
    END
  END la_oen[5]
  PIN la_oen[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.560 4.000 180.160 ;
    END
  END la_oen[6]
  PIN la_oen[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 184.320 4.000 184.920 ;
    END
  END la_oen[7]
  PIN la_oen[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.080 4.000 189.680 ;
    END
  END la_oen[8]
  PIN la_oen[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END la_oen[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 296.000 2.210 300.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 296.000 5.890 300.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.710 296.000 21.990 300.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 296.000 45.910 300.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 296.000 85.930 300.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 296.000 90.070 300.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 296.000 93.750 300.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 296.000 97.890 300.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.750 296.000 102.030 300.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 296.000 106.170 300.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 296.000 109.850 300.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.710 296.000 113.990 300.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 296.000 118.130 300.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.530 296.000 121.810 300.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 296.000 50.050 300.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 296.000 125.950 300.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 296.000 130.090 300.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 296.000 133.770 300.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.630 296.000 137.910 300.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 296.000 142.050 300.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.450 296.000 145.730 300.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 296.000 149.870 300.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.730 296.000 154.010 300.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 296.000 158.150 300.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.550 296.000 161.830 300.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 296.000 54.190 300.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 296.000 165.970 300.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.830 296.000 170.110 300.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 296.000 57.870 300.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 296.000 62.010 300.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 296.000 66.150 300.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 296.000 69.830 300.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 296.000 73.970 300.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 296.000 78.110 300.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.510 296.000 81.790 300.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 296.000 14.170 300.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.510 296.000 173.790 300.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.530 296.000 213.810 300.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.670 296.000 217.950 300.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.810 296.000 222.090 300.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 296.000 225.770 300.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.630 296.000 229.910 300.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.770 296.000 234.050 300.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.450 296.000 237.730 300.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 296.000 241.870 300.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.730 296.000 246.010 300.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.410 296.000 249.690 300.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.650 296.000 177.930 300.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.550 296.000 253.830 300.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 296.000 257.970 300.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.830 296.000 262.110 300.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.510 296.000 265.790 300.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.650 296.000 269.930 300.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 296.000 274.070 300.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.470 296.000 277.750 300.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.610 296.000 281.890 300.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.750 296.000 286.030 300.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.430 296.000 289.710 300.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.790 296.000 182.070 300.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.570 296.000 293.850 300.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.710 296.000 297.990 300.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.470 296.000 185.750 300.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.610 296.000 189.890 300.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.750 296.000 194.030 300.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.430 296.000 197.710 300.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.570 296.000 201.850 300.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 296.000 205.990 300.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 296.000 210.130 300.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.080 4.000 2.680 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.320 4.000 48.920 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 4.000 53.680 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 4.000 63.200 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 67.360 4.000 67.960 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 4.000 72.720 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.880 4.000 77.480 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 86.400 4.000 87.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 90.480 4.000 91.080 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.160 4.000 6.760 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 4.000 100.600 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 4.000 105.360 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 109.520 4.000 110.120 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.280 4.000 114.880 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.800 4.000 124.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 128.560 4.000 129.160 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.160 4.000 142.760 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.920 4.000 147.520 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.680 4.000 16.280 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.200 4.000 25.800 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 4.000 30.560 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.720 4.000 35.320 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 296.000 29.810 300.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 296.000 33.950 300.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 296.000 38.090 300.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.490 296.000 41.770 300.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 296.000 10.030 300.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 296.000 17.850 300.000 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 288.560 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 288.560 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 288.560 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 288.560 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 177.940 10.880 179.540 288.320 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.880 25.940 288.320 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 254.740 10.880 256.340 288.320 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 101.140 10.880 102.740 288.320 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 181.240 10.880 182.840 288.320 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 27.640 10.880 29.240 288.320 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 258.040 10.880 259.640 288.320 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 104.440 10.880 106.040 288.320 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 184.540 10.880 186.140 288.320 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 30.940 10.880 32.540 288.320 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 261.340 10.880 262.940 288.320 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 107.740 10.880 109.340 288.320 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 294.400 288.405 ;
      LAYER met1 ;
        RECT 1.910 4.120 298.010 288.560 ;
      LAYER met2 ;
        RECT 2.490 295.720 5.330 298.365 ;
        RECT 6.170 295.720 9.470 298.365 ;
        RECT 10.310 295.720 13.610 298.365 ;
        RECT 14.450 295.720 17.290 298.365 ;
        RECT 18.130 295.720 21.430 298.365 ;
        RECT 22.270 295.720 25.570 298.365 ;
        RECT 26.410 295.720 29.250 298.365 ;
        RECT 30.090 295.720 33.390 298.365 ;
        RECT 34.230 295.720 37.530 298.365 ;
        RECT 38.370 295.720 41.210 298.365 ;
        RECT 42.050 295.720 45.350 298.365 ;
        RECT 46.190 295.720 49.490 298.365 ;
        RECT 50.330 295.720 53.630 298.365 ;
        RECT 54.470 295.720 57.310 298.365 ;
        RECT 58.150 295.720 61.450 298.365 ;
        RECT 62.290 295.720 65.590 298.365 ;
        RECT 66.430 295.720 69.270 298.365 ;
        RECT 70.110 295.720 73.410 298.365 ;
        RECT 74.250 295.720 77.550 298.365 ;
        RECT 78.390 295.720 81.230 298.365 ;
        RECT 82.070 295.720 85.370 298.365 ;
        RECT 86.210 295.720 89.510 298.365 ;
        RECT 90.350 295.720 93.190 298.365 ;
        RECT 94.030 295.720 97.330 298.365 ;
        RECT 98.170 295.720 101.470 298.365 ;
        RECT 102.310 295.720 105.610 298.365 ;
        RECT 106.450 295.720 109.290 298.365 ;
        RECT 110.130 295.720 113.430 298.365 ;
        RECT 114.270 295.720 117.570 298.365 ;
        RECT 118.410 295.720 121.250 298.365 ;
        RECT 122.090 295.720 125.390 298.365 ;
        RECT 126.230 295.720 129.530 298.365 ;
        RECT 130.370 295.720 133.210 298.365 ;
        RECT 134.050 295.720 137.350 298.365 ;
        RECT 138.190 295.720 141.490 298.365 ;
        RECT 142.330 295.720 145.170 298.365 ;
        RECT 146.010 295.720 149.310 298.365 ;
        RECT 150.150 295.720 153.450 298.365 ;
        RECT 154.290 295.720 157.590 298.365 ;
        RECT 158.430 295.720 161.270 298.365 ;
        RECT 162.110 295.720 165.410 298.365 ;
        RECT 166.250 295.720 169.550 298.365 ;
        RECT 170.390 295.720 173.230 298.365 ;
        RECT 174.070 295.720 177.370 298.365 ;
        RECT 178.210 295.720 181.510 298.365 ;
        RECT 182.350 295.720 185.190 298.365 ;
        RECT 186.030 295.720 189.330 298.365 ;
        RECT 190.170 295.720 193.470 298.365 ;
        RECT 194.310 295.720 197.150 298.365 ;
        RECT 197.990 295.720 201.290 298.365 ;
        RECT 202.130 295.720 205.430 298.365 ;
        RECT 206.270 295.720 209.570 298.365 ;
        RECT 210.410 295.720 213.250 298.365 ;
        RECT 214.090 295.720 217.390 298.365 ;
        RECT 218.230 295.720 221.530 298.365 ;
        RECT 222.370 295.720 225.210 298.365 ;
        RECT 226.050 295.720 229.350 298.365 ;
        RECT 230.190 295.720 233.490 298.365 ;
        RECT 234.330 295.720 237.170 298.365 ;
        RECT 238.010 295.720 241.310 298.365 ;
        RECT 242.150 295.720 245.450 298.365 ;
        RECT 246.290 295.720 249.130 298.365 ;
        RECT 249.970 295.720 253.270 298.365 ;
        RECT 254.110 295.720 257.410 298.365 ;
        RECT 258.250 295.720 261.550 298.365 ;
        RECT 262.390 295.720 265.230 298.365 ;
        RECT 266.070 295.720 269.370 298.365 ;
        RECT 270.210 295.720 273.510 298.365 ;
        RECT 274.350 295.720 277.190 298.365 ;
        RECT 278.030 295.720 281.330 298.365 ;
        RECT 282.170 295.720 285.470 298.365 ;
        RECT 286.310 295.720 289.150 298.365 ;
        RECT 289.990 295.720 293.290 298.365 ;
        RECT 294.130 295.720 297.430 298.365 ;
        RECT 1.940 4.280 297.980 295.720 ;
        RECT 1.940 0.835 2.110 4.280 ;
        RECT 2.950 0.835 6.710 4.280 ;
        RECT 7.550 0.835 11.310 4.280 ;
        RECT 12.150 0.835 15.910 4.280 ;
        RECT 16.750 0.835 20.510 4.280 ;
        RECT 21.350 0.835 25.110 4.280 ;
        RECT 25.950 0.835 30.170 4.280 ;
        RECT 31.010 0.835 34.770 4.280 ;
        RECT 35.610 0.835 39.370 4.280 ;
        RECT 40.210 0.835 43.970 4.280 ;
        RECT 44.810 0.835 48.570 4.280 ;
        RECT 49.410 0.835 53.630 4.280 ;
        RECT 54.470 0.835 58.230 4.280 ;
        RECT 59.070 0.835 62.830 4.280 ;
        RECT 63.670 0.835 67.430 4.280 ;
        RECT 68.270 0.835 72.030 4.280 ;
        RECT 72.870 0.835 77.090 4.280 ;
        RECT 77.930 0.835 81.690 4.280 ;
        RECT 82.530 0.835 86.290 4.280 ;
        RECT 87.130 0.835 90.890 4.280 ;
        RECT 91.730 0.835 95.490 4.280 ;
        RECT 96.330 0.835 100.090 4.280 ;
        RECT 100.930 0.835 105.150 4.280 ;
        RECT 105.990 0.835 109.750 4.280 ;
        RECT 110.590 0.835 114.350 4.280 ;
        RECT 115.190 0.835 118.950 4.280 ;
        RECT 119.790 0.835 123.550 4.280 ;
        RECT 124.390 0.835 128.610 4.280 ;
        RECT 129.450 0.835 133.210 4.280 ;
        RECT 134.050 0.835 137.810 4.280 ;
        RECT 138.650 0.835 142.410 4.280 ;
        RECT 143.250 0.835 147.010 4.280 ;
        RECT 147.850 0.835 152.070 4.280 ;
        RECT 152.910 0.835 156.670 4.280 ;
        RECT 157.510 0.835 161.270 4.280 ;
        RECT 162.110 0.835 165.870 4.280 ;
        RECT 166.710 0.835 170.470 4.280 ;
        RECT 171.310 0.835 175.070 4.280 ;
        RECT 175.910 0.835 180.130 4.280 ;
        RECT 180.970 0.835 184.730 4.280 ;
        RECT 185.570 0.835 189.330 4.280 ;
        RECT 190.170 0.835 193.930 4.280 ;
        RECT 194.770 0.835 198.530 4.280 ;
        RECT 199.370 0.835 203.590 4.280 ;
        RECT 204.430 0.835 208.190 4.280 ;
        RECT 209.030 0.835 212.790 4.280 ;
        RECT 213.630 0.835 217.390 4.280 ;
        RECT 218.230 0.835 221.990 4.280 ;
        RECT 222.830 0.835 227.050 4.280 ;
        RECT 227.890 0.835 231.650 4.280 ;
        RECT 232.490 0.835 236.250 4.280 ;
        RECT 237.090 0.835 240.850 4.280 ;
        RECT 241.690 0.835 245.450 4.280 ;
        RECT 246.290 0.835 250.050 4.280 ;
        RECT 250.890 0.835 255.110 4.280 ;
        RECT 255.950 0.835 259.710 4.280 ;
        RECT 260.550 0.835 264.310 4.280 ;
        RECT 265.150 0.835 268.910 4.280 ;
        RECT 269.750 0.835 273.510 4.280 ;
        RECT 274.350 0.835 278.570 4.280 ;
        RECT 279.410 0.835 283.170 4.280 ;
        RECT 284.010 0.835 287.770 4.280 ;
        RECT 288.610 0.835 292.370 4.280 ;
        RECT 293.210 0.835 296.970 4.280 ;
        RECT 297.810 0.835 297.980 4.280 ;
      LAYER met3 ;
        RECT 4.000 298.200 295.600 298.345 ;
        RECT 4.400 297.480 295.600 298.200 ;
        RECT 4.400 296.800 296.000 297.480 ;
        RECT 4.000 296.160 296.000 296.800 ;
        RECT 4.000 294.760 295.600 296.160 ;
        RECT 4.000 293.440 296.000 294.760 ;
        RECT 4.400 292.040 295.600 293.440 ;
        RECT 4.000 290.720 296.000 292.040 ;
        RECT 4.000 289.320 295.600 290.720 ;
        RECT 4.000 288.680 296.000 289.320 ;
        RECT 4.400 288.000 296.000 288.680 ;
        RECT 4.400 287.280 295.600 288.000 ;
        RECT 4.000 286.600 295.600 287.280 ;
        RECT 4.000 285.280 296.000 286.600 ;
        RECT 4.000 283.920 295.600 285.280 ;
        RECT 4.400 283.880 295.600 283.920 ;
        RECT 4.400 282.560 296.000 283.880 ;
        RECT 4.400 282.520 295.600 282.560 ;
        RECT 4.000 281.160 295.600 282.520 ;
        RECT 4.000 280.520 296.000 281.160 ;
        RECT 4.000 279.160 295.600 280.520 ;
        RECT 4.400 279.120 295.600 279.160 ;
        RECT 4.400 277.800 296.000 279.120 ;
        RECT 4.400 277.760 295.600 277.800 ;
        RECT 4.000 276.400 295.600 277.760 ;
        RECT 4.000 275.080 296.000 276.400 ;
        RECT 4.000 274.400 295.600 275.080 ;
        RECT 4.400 273.680 295.600 274.400 ;
        RECT 4.400 273.000 296.000 273.680 ;
        RECT 4.000 272.360 296.000 273.000 ;
        RECT 4.000 270.960 295.600 272.360 ;
        RECT 4.000 269.640 296.000 270.960 ;
        RECT 4.400 268.240 295.600 269.640 ;
        RECT 4.000 266.920 296.000 268.240 ;
        RECT 4.000 265.520 295.600 266.920 ;
        RECT 4.000 264.880 296.000 265.520 ;
        RECT 4.400 264.200 296.000 264.880 ;
        RECT 4.400 263.480 295.600 264.200 ;
        RECT 4.000 262.800 295.600 263.480 ;
        RECT 4.000 261.480 296.000 262.800 ;
        RECT 4.000 260.120 295.600 261.480 ;
        RECT 4.400 260.080 295.600 260.120 ;
        RECT 4.400 259.440 296.000 260.080 ;
        RECT 4.400 258.720 295.600 259.440 ;
        RECT 4.000 258.040 295.600 258.720 ;
        RECT 4.000 256.720 296.000 258.040 ;
        RECT 4.000 256.040 295.600 256.720 ;
        RECT 4.400 255.320 295.600 256.040 ;
        RECT 4.400 254.640 296.000 255.320 ;
        RECT 4.000 254.000 296.000 254.640 ;
        RECT 4.000 252.600 295.600 254.000 ;
        RECT 4.000 251.280 296.000 252.600 ;
        RECT 4.400 249.880 295.600 251.280 ;
        RECT 4.000 248.560 296.000 249.880 ;
        RECT 4.000 247.160 295.600 248.560 ;
        RECT 4.000 246.520 296.000 247.160 ;
        RECT 4.400 245.840 296.000 246.520 ;
        RECT 4.400 245.120 295.600 245.840 ;
        RECT 4.000 244.440 295.600 245.120 ;
        RECT 4.000 243.120 296.000 244.440 ;
        RECT 4.000 241.760 295.600 243.120 ;
        RECT 4.400 241.720 295.600 241.760 ;
        RECT 4.400 241.080 296.000 241.720 ;
        RECT 4.400 240.360 295.600 241.080 ;
        RECT 4.000 239.680 295.600 240.360 ;
        RECT 4.000 238.360 296.000 239.680 ;
        RECT 4.000 237.000 295.600 238.360 ;
        RECT 4.400 236.960 295.600 237.000 ;
        RECT 4.400 235.640 296.000 236.960 ;
        RECT 4.400 235.600 295.600 235.640 ;
        RECT 4.000 234.240 295.600 235.600 ;
        RECT 4.000 232.920 296.000 234.240 ;
        RECT 4.000 232.240 295.600 232.920 ;
        RECT 4.400 231.520 295.600 232.240 ;
        RECT 4.400 230.840 296.000 231.520 ;
        RECT 4.000 230.200 296.000 230.840 ;
        RECT 4.000 228.800 295.600 230.200 ;
        RECT 4.000 227.480 296.000 228.800 ;
        RECT 4.400 226.080 295.600 227.480 ;
        RECT 4.000 224.760 296.000 226.080 ;
        RECT 4.000 223.360 295.600 224.760 ;
        RECT 4.000 222.720 296.000 223.360 ;
        RECT 4.400 222.040 296.000 222.720 ;
        RECT 4.400 221.320 295.600 222.040 ;
        RECT 4.000 220.640 295.600 221.320 ;
        RECT 4.000 220.000 296.000 220.640 ;
        RECT 4.000 218.600 295.600 220.000 ;
        RECT 4.000 217.960 296.000 218.600 ;
        RECT 4.400 217.280 296.000 217.960 ;
        RECT 4.400 216.560 295.600 217.280 ;
        RECT 4.000 215.880 295.600 216.560 ;
        RECT 4.000 214.560 296.000 215.880 ;
        RECT 4.000 213.880 295.600 214.560 ;
        RECT 4.400 213.160 295.600 213.880 ;
        RECT 4.400 212.480 296.000 213.160 ;
        RECT 4.000 211.840 296.000 212.480 ;
        RECT 4.000 210.440 295.600 211.840 ;
        RECT 4.000 209.120 296.000 210.440 ;
        RECT 4.400 207.720 295.600 209.120 ;
        RECT 4.000 206.400 296.000 207.720 ;
        RECT 4.000 205.000 295.600 206.400 ;
        RECT 4.000 204.360 296.000 205.000 ;
        RECT 4.400 203.680 296.000 204.360 ;
        RECT 4.400 202.960 295.600 203.680 ;
        RECT 4.000 202.280 295.600 202.960 ;
        RECT 4.000 201.640 296.000 202.280 ;
        RECT 4.000 200.240 295.600 201.640 ;
        RECT 4.000 199.600 296.000 200.240 ;
        RECT 4.400 198.920 296.000 199.600 ;
        RECT 4.400 198.200 295.600 198.920 ;
        RECT 4.000 197.520 295.600 198.200 ;
        RECT 4.000 196.200 296.000 197.520 ;
        RECT 4.000 194.840 295.600 196.200 ;
        RECT 4.400 194.800 295.600 194.840 ;
        RECT 4.400 193.480 296.000 194.800 ;
        RECT 4.400 193.440 295.600 193.480 ;
        RECT 4.000 192.080 295.600 193.440 ;
        RECT 4.000 190.760 296.000 192.080 ;
        RECT 4.000 190.080 295.600 190.760 ;
        RECT 4.400 189.360 295.600 190.080 ;
        RECT 4.400 188.680 296.000 189.360 ;
        RECT 4.000 188.040 296.000 188.680 ;
        RECT 4.000 186.640 295.600 188.040 ;
        RECT 4.000 185.320 296.000 186.640 ;
        RECT 4.400 183.920 295.600 185.320 ;
        RECT 4.000 182.600 296.000 183.920 ;
        RECT 4.000 181.200 295.600 182.600 ;
        RECT 4.000 180.560 296.000 181.200 ;
        RECT 4.400 179.160 295.600 180.560 ;
        RECT 4.000 177.840 296.000 179.160 ;
        RECT 4.000 176.440 295.600 177.840 ;
        RECT 4.000 175.800 296.000 176.440 ;
        RECT 4.400 175.120 296.000 175.800 ;
        RECT 4.400 174.400 295.600 175.120 ;
        RECT 4.000 173.720 295.600 174.400 ;
        RECT 4.000 172.400 296.000 173.720 ;
        RECT 4.000 171.720 295.600 172.400 ;
        RECT 4.400 171.000 295.600 171.720 ;
        RECT 4.400 170.320 296.000 171.000 ;
        RECT 4.000 169.680 296.000 170.320 ;
        RECT 4.000 168.280 295.600 169.680 ;
        RECT 4.000 166.960 296.000 168.280 ;
        RECT 4.400 165.560 295.600 166.960 ;
        RECT 4.000 164.240 296.000 165.560 ;
        RECT 4.000 162.840 295.600 164.240 ;
        RECT 4.000 162.200 296.000 162.840 ;
        RECT 4.400 161.520 296.000 162.200 ;
        RECT 4.400 160.800 295.600 161.520 ;
        RECT 4.000 160.120 295.600 160.800 ;
        RECT 4.000 159.480 296.000 160.120 ;
        RECT 4.000 158.080 295.600 159.480 ;
        RECT 4.000 157.440 296.000 158.080 ;
        RECT 4.400 156.760 296.000 157.440 ;
        RECT 4.400 156.040 295.600 156.760 ;
        RECT 4.000 155.360 295.600 156.040 ;
        RECT 4.000 154.040 296.000 155.360 ;
        RECT 4.000 152.680 295.600 154.040 ;
        RECT 4.400 152.640 295.600 152.680 ;
        RECT 4.400 151.320 296.000 152.640 ;
        RECT 4.400 151.280 295.600 151.320 ;
        RECT 4.000 149.920 295.600 151.280 ;
        RECT 4.000 148.600 296.000 149.920 ;
        RECT 4.000 147.920 295.600 148.600 ;
        RECT 4.400 147.200 295.600 147.920 ;
        RECT 4.400 146.520 296.000 147.200 ;
        RECT 4.000 145.880 296.000 146.520 ;
        RECT 4.000 144.480 295.600 145.880 ;
        RECT 4.000 143.160 296.000 144.480 ;
        RECT 4.400 141.760 295.600 143.160 ;
        RECT 4.000 141.120 296.000 141.760 ;
        RECT 4.000 139.720 295.600 141.120 ;
        RECT 4.000 138.400 296.000 139.720 ;
        RECT 4.400 137.000 295.600 138.400 ;
        RECT 4.000 135.680 296.000 137.000 ;
        RECT 4.000 134.280 295.600 135.680 ;
        RECT 4.000 133.640 296.000 134.280 ;
        RECT 4.400 132.960 296.000 133.640 ;
        RECT 4.400 132.240 295.600 132.960 ;
        RECT 4.000 131.560 295.600 132.240 ;
        RECT 4.000 130.240 296.000 131.560 ;
        RECT 4.000 129.560 295.600 130.240 ;
        RECT 4.400 128.840 295.600 129.560 ;
        RECT 4.400 128.160 296.000 128.840 ;
        RECT 4.000 127.520 296.000 128.160 ;
        RECT 4.000 126.120 295.600 127.520 ;
        RECT 4.000 124.800 296.000 126.120 ;
        RECT 4.400 123.400 295.600 124.800 ;
        RECT 4.000 122.080 296.000 123.400 ;
        RECT 4.000 120.680 295.600 122.080 ;
        RECT 4.000 120.040 296.000 120.680 ;
        RECT 4.400 118.640 295.600 120.040 ;
        RECT 4.000 117.320 296.000 118.640 ;
        RECT 4.000 115.920 295.600 117.320 ;
        RECT 4.000 115.280 296.000 115.920 ;
        RECT 4.400 114.600 296.000 115.280 ;
        RECT 4.400 113.880 295.600 114.600 ;
        RECT 4.000 113.200 295.600 113.880 ;
        RECT 4.000 111.880 296.000 113.200 ;
        RECT 4.000 110.520 295.600 111.880 ;
        RECT 4.400 110.480 295.600 110.520 ;
        RECT 4.400 109.160 296.000 110.480 ;
        RECT 4.400 109.120 295.600 109.160 ;
        RECT 4.000 107.760 295.600 109.120 ;
        RECT 4.000 106.440 296.000 107.760 ;
        RECT 4.000 105.760 295.600 106.440 ;
        RECT 4.400 105.040 295.600 105.760 ;
        RECT 4.400 104.360 296.000 105.040 ;
        RECT 4.000 103.720 296.000 104.360 ;
        RECT 4.000 102.320 295.600 103.720 ;
        RECT 4.000 101.680 296.000 102.320 ;
        RECT 4.000 101.000 295.600 101.680 ;
        RECT 4.400 100.280 295.600 101.000 ;
        RECT 4.400 99.600 296.000 100.280 ;
        RECT 4.000 98.960 296.000 99.600 ;
        RECT 4.000 97.560 295.600 98.960 ;
        RECT 4.000 96.240 296.000 97.560 ;
        RECT 4.400 94.840 295.600 96.240 ;
        RECT 4.000 93.520 296.000 94.840 ;
        RECT 4.000 92.120 295.600 93.520 ;
        RECT 4.000 91.480 296.000 92.120 ;
        RECT 4.400 90.800 296.000 91.480 ;
        RECT 4.400 90.080 295.600 90.800 ;
        RECT 4.000 89.400 295.600 90.080 ;
        RECT 4.000 88.080 296.000 89.400 ;
        RECT 4.000 87.400 295.600 88.080 ;
        RECT 4.400 86.680 295.600 87.400 ;
        RECT 4.400 86.000 296.000 86.680 ;
        RECT 4.000 85.360 296.000 86.000 ;
        RECT 4.000 83.960 295.600 85.360 ;
        RECT 4.000 82.640 296.000 83.960 ;
        RECT 4.400 81.240 295.600 82.640 ;
        RECT 4.000 80.600 296.000 81.240 ;
        RECT 4.000 79.200 295.600 80.600 ;
        RECT 4.000 77.880 296.000 79.200 ;
        RECT 4.400 76.480 295.600 77.880 ;
        RECT 4.000 75.160 296.000 76.480 ;
        RECT 4.000 73.760 295.600 75.160 ;
        RECT 4.000 73.120 296.000 73.760 ;
        RECT 4.400 72.440 296.000 73.120 ;
        RECT 4.400 71.720 295.600 72.440 ;
        RECT 4.000 71.040 295.600 71.720 ;
        RECT 4.000 69.720 296.000 71.040 ;
        RECT 4.000 68.360 295.600 69.720 ;
        RECT 4.400 68.320 295.600 68.360 ;
        RECT 4.400 67.000 296.000 68.320 ;
        RECT 4.400 66.960 295.600 67.000 ;
        RECT 4.000 65.600 295.600 66.960 ;
        RECT 4.000 64.280 296.000 65.600 ;
        RECT 4.000 63.600 295.600 64.280 ;
        RECT 4.400 62.880 295.600 63.600 ;
        RECT 4.400 62.200 296.000 62.880 ;
        RECT 4.000 61.560 296.000 62.200 ;
        RECT 4.000 60.160 295.600 61.560 ;
        RECT 4.000 59.520 296.000 60.160 ;
        RECT 4.000 58.840 295.600 59.520 ;
        RECT 4.400 58.120 295.600 58.840 ;
        RECT 4.400 57.440 296.000 58.120 ;
        RECT 4.000 56.800 296.000 57.440 ;
        RECT 4.000 55.400 295.600 56.800 ;
        RECT 4.000 54.080 296.000 55.400 ;
        RECT 4.400 52.680 295.600 54.080 ;
        RECT 4.000 51.360 296.000 52.680 ;
        RECT 4.000 49.960 295.600 51.360 ;
        RECT 4.000 49.320 296.000 49.960 ;
        RECT 4.400 48.640 296.000 49.320 ;
        RECT 4.400 47.920 295.600 48.640 ;
        RECT 4.000 47.240 295.600 47.920 ;
        RECT 4.000 45.920 296.000 47.240 ;
        RECT 4.000 45.240 295.600 45.920 ;
        RECT 4.400 44.520 295.600 45.240 ;
        RECT 4.400 43.840 296.000 44.520 ;
        RECT 4.000 43.200 296.000 43.840 ;
        RECT 4.000 41.800 295.600 43.200 ;
        RECT 4.000 41.160 296.000 41.800 ;
        RECT 4.000 40.480 295.600 41.160 ;
        RECT 4.400 39.760 295.600 40.480 ;
        RECT 4.400 39.080 296.000 39.760 ;
        RECT 4.000 38.440 296.000 39.080 ;
        RECT 4.000 37.040 295.600 38.440 ;
        RECT 4.000 35.720 296.000 37.040 ;
        RECT 4.400 34.320 295.600 35.720 ;
        RECT 4.000 33.000 296.000 34.320 ;
        RECT 4.000 31.600 295.600 33.000 ;
        RECT 4.000 30.960 296.000 31.600 ;
        RECT 4.400 30.280 296.000 30.960 ;
        RECT 4.400 29.560 295.600 30.280 ;
        RECT 4.000 28.880 295.600 29.560 ;
        RECT 4.000 27.560 296.000 28.880 ;
        RECT 4.000 26.200 295.600 27.560 ;
        RECT 4.400 26.160 295.600 26.200 ;
        RECT 4.400 24.840 296.000 26.160 ;
        RECT 4.400 24.800 295.600 24.840 ;
        RECT 4.000 23.440 295.600 24.800 ;
        RECT 4.000 22.120 296.000 23.440 ;
        RECT 4.000 21.440 295.600 22.120 ;
        RECT 4.400 20.720 295.600 21.440 ;
        RECT 4.400 20.080 296.000 20.720 ;
        RECT 4.400 20.040 295.600 20.080 ;
        RECT 4.000 18.680 295.600 20.040 ;
        RECT 4.000 17.360 296.000 18.680 ;
        RECT 4.000 16.680 295.600 17.360 ;
        RECT 4.400 15.960 295.600 16.680 ;
        RECT 4.400 15.280 296.000 15.960 ;
        RECT 4.000 14.640 296.000 15.280 ;
        RECT 4.000 13.240 295.600 14.640 ;
        RECT 4.000 11.920 296.000 13.240 ;
        RECT 4.400 10.520 295.600 11.920 ;
        RECT 4.000 9.200 296.000 10.520 ;
        RECT 4.000 7.800 295.600 9.200 ;
        RECT 4.000 7.160 296.000 7.800 ;
        RECT 4.400 6.480 296.000 7.160 ;
        RECT 4.400 5.760 295.600 6.480 ;
        RECT 4.000 5.080 295.600 5.760 ;
        RECT 4.000 3.760 296.000 5.080 ;
        RECT 4.000 3.080 295.600 3.760 ;
        RECT 4.400 2.360 295.600 3.080 ;
        RECT 4.400 1.720 296.000 2.360 ;
        RECT 4.400 1.680 295.600 1.720 ;
        RECT 4.000 0.855 295.600 1.680 ;
  END
END wrapped_rgb_mixer
END LIBRARY

