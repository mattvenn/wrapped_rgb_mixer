// This is the unpowered netlist.
module wrapped_rgb_mixer (active,
    wb_clk_i,
    io_in,
    io_oeb,
    io_out,
    la1_data_in,
    la1_data_out,
    la1_oenb);
 input active;
 input wb_clk_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [31:0] la1_data_in;
 output [31:0] la1_data_out;
 input [31:0] la1_oenb;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire clknet_0_wb_clk_i;
 wire \rgb_mixer0.debounce0_a.button_hist[0] ;
 wire \rgb_mixer0.debounce0_a.button_hist[1] ;
 wire \rgb_mixer0.debounce0_a.button_hist[2] ;
 wire \rgb_mixer0.debounce0_a.button_hist[3] ;
 wire \rgb_mixer0.debounce0_a.button_hist[4] ;
 wire \rgb_mixer0.debounce0_a.button_hist[5] ;
 wire \rgb_mixer0.debounce0_a.button_hist[6] ;
 wire \rgb_mixer0.debounce0_a.button_hist[7] ;
 wire \rgb_mixer0.debounce0_a.debounced ;
 wire \rgb_mixer0.debounce0_b.button_hist[0] ;
 wire \rgb_mixer0.debounce0_b.button_hist[1] ;
 wire \rgb_mixer0.debounce0_b.button_hist[2] ;
 wire \rgb_mixer0.debounce0_b.button_hist[3] ;
 wire \rgb_mixer0.debounce0_b.button_hist[4] ;
 wire \rgb_mixer0.debounce0_b.button_hist[5] ;
 wire \rgb_mixer0.debounce0_b.button_hist[6] ;
 wire \rgb_mixer0.debounce0_b.button_hist[7] ;
 wire \rgb_mixer0.debounce0_b.debounced ;
 wire \rgb_mixer0.debounce1_a.button_hist[0] ;
 wire \rgb_mixer0.debounce1_a.button_hist[1] ;
 wire \rgb_mixer0.debounce1_a.button_hist[2] ;
 wire \rgb_mixer0.debounce1_a.button_hist[3] ;
 wire \rgb_mixer0.debounce1_a.button_hist[4] ;
 wire \rgb_mixer0.debounce1_a.button_hist[5] ;
 wire \rgb_mixer0.debounce1_a.button_hist[6] ;
 wire \rgb_mixer0.debounce1_a.button_hist[7] ;
 wire \rgb_mixer0.debounce1_a.debounced ;
 wire \rgb_mixer0.debounce1_b.button_hist[0] ;
 wire \rgb_mixer0.debounce1_b.button_hist[1] ;
 wire \rgb_mixer0.debounce1_b.button_hist[2] ;
 wire \rgb_mixer0.debounce1_b.button_hist[3] ;
 wire \rgb_mixer0.debounce1_b.button_hist[4] ;
 wire \rgb_mixer0.debounce1_b.button_hist[5] ;
 wire \rgb_mixer0.debounce1_b.button_hist[6] ;
 wire \rgb_mixer0.debounce1_b.button_hist[7] ;
 wire \rgb_mixer0.debounce1_b.debounced ;
 wire \rgb_mixer0.debounce2_a.button_hist[0] ;
 wire \rgb_mixer0.debounce2_a.button_hist[1] ;
 wire \rgb_mixer0.debounce2_a.button_hist[2] ;
 wire \rgb_mixer0.debounce2_a.button_hist[3] ;
 wire \rgb_mixer0.debounce2_a.button_hist[4] ;
 wire \rgb_mixer0.debounce2_a.button_hist[5] ;
 wire \rgb_mixer0.debounce2_a.button_hist[6] ;
 wire \rgb_mixer0.debounce2_a.button_hist[7] ;
 wire \rgb_mixer0.debounce2_a.debounced ;
 wire \rgb_mixer0.debounce2_b.button_hist[0] ;
 wire \rgb_mixer0.debounce2_b.button_hist[1] ;
 wire \rgb_mixer0.debounce2_b.button_hist[2] ;
 wire \rgb_mixer0.debounce2_b.button_hist[3] ;
 wire \rgb_mixer0.debounce2_b.button_hist[4] ;
 wire \rgb_mixer0.debounce2_b.button_hist[5] ;
 wire \rgb_mixer0.debounce2_b.button_hist[6] ;
 wire \rgb_mixer0.debounce2_b.button_hist[7] ;
 wire \rgb_mixer0.debounce2_b.debounced ;
 wire \rgb_mixer0.enc0[0] ;
 wire \rgb_mixer0.enc0[1] ;
 wire \rgb_mixer0.enc0[2] ;
 wire \rgb_mixer0.enc0[3] ;
 wire \rgb_mixer0.enc0[4] ;
 wire \rgb_mixer0.enc0[5] ;
 wire \rgb_mixer0.enc0[6] ;
 wire \rgb_mixer0.enc0[7] ;
 wire \rgb_mixer0.enc1[0] ;
 wire \rgb_mixer0.enc1[1] ;
 wire \rgb_mixer0.enc1[2] ;
 wire \rgb_mixer0.enc1[3] ;
 wire \rgb_mixer0.enc1[4] ;
 wire \rgb_mixer0.enc1[5] ;
 wire \rgb_mixer0.enc1[6] ;
 wire \rgb_mixer0.enc1[7] ;
 wire \rgb_mixer0.enc2[0] ;
 wire \rgb_mixer0.enc2[1] ;
 wire \rgb_mixer0.enc2[2] ;
 wire \rgb_mixer0.enc2[3] ;
 wire \rgb_mixer0.enc2[4] ;
 wire \rgb_mixer0.enc2[5] ;
 wire \rgb_mixer0.enc2[6] ;
 wire \rgb_mixer0.enc2[7] ;
 wire \rgb_mixer0.encoder0.old_a ;
 wire \rgb_mixer0.encoder0.old_b ;
 wire \rgb_mixer0.encoder1.old_a ;
 wire \rgb_mixer0.encoder1.old_b ;
 wire \rgb_mixer0.encoder2.old_a ;
 wire \rgb_mixer0.encoder2.old_b ;
 wire \rgb_mixer0.pwm0.count[0] ;
 wire \rgb_mixer0.pwm0.count[1] ;
 wire \rgb_mixer0.pwm0.count[2] ;
 wire \rgb_mixer0.pwm0.count[3] ;
 wire \rgb_mixer0.pwm0.count[4] ;
 wire \rgb_mixer0.pwm0.count[5] ;
 wire \rgb_mixer0.pwm0.count[6] ;
 wire \rgb_mixer0.pwm0.count[7] ;
 wire \rgb_mixer0.pwm0.out ;
 wire \rgb_mixer0.pwm1.count[0] ;
 wire \rgb_mixer0.pwm1.count[1] ;
 wire \rgb_mixer0.pwm1.count[2] ;
 wire \rgb_mixer0.pwm1.count[3] ;
 wire \rgb_mixer0.pwm1.count[4] ;
 wire \rgb_mixer0.pwm1.count[5] ;
 wire \rgb_mixer0.pwm1.count[6] ;
 wire \rgb_mixer0.pwm1.count[7] ;
 wire \rgb_mixer0.pwm1.out ;
 wire \rgb_mixer0.pwm2.count[0] ;
 wire \rgb_mixer0.pwm2.count[1] ;
 wire \rgb_mixer0.pwm2.count[2] ;
 wire \rgb_mixer0.pwm2.count[3] ;
 wire \rgb_mixer0.pwm2.count[4] ;
 wire \rgb_mixer0.pwm2.count[5] ;
 wire \rgb_mixer0.pwm2.count[6] ;
 wire \rgb_mixer0.pwm2.count[7] ;
 wire \rgb_mixer0.pwm2.out ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire clknet_3_0__leaf_wb_clk_i;
 wire clknet_3_1__leaf_wb_clk_i;
 wire clknet_3_2__leaf_wb_clk_i;
 wire clknet_3_3__leaf_wb_clk_i;
 wire clknet_3_4__leaf_wb_clk_i;
 wire clknet_3_5__leaf_wb_clk_i;
 wire clknet_3_6__leaf_wb_clk_i;
 wire clknet_3_7__leaf_wb_clk_i;

 sky130_fd_sc_hd__clkbuf_8 _0668_ (.A(net1),
    .X(_0108_));
 sky130_fd_sc_hd__buf_8 _0669_ (.A(_0108_),
    .X(_0109_));
 sky130_fd_sc_hd__buf_8 _0670_ (.A(_0109_),
    .X(_0110_));
 sky130_fd_sc_hd__inv_2 _0671_ (.A(_0110_),
    .Y(_0455_));
 sky130_fd_sc_hd__inv_2 _0672_ (.A(_0110_),
    .Y(_0456_));
 sky130_fd_sc_hd__inv_2 _0673_ (.A(_0110_),
    .Y(_0457_));
 sky130_fd_sc_hd__inv_2 _0674_ (.A(_0110_),
    .Y(_0458_));
 sky130_fd_sc_hd__inv_2 _0675_ (.A(_0110_),
    .Y(_0464_));
 sky130_fd_sc_hd__inv_2 _0676_ (.A(_0110_),
    .Y(_0463_));
 sky130_fd_sc_hd__inv_2 _0677_ (.A(_0110_),
    .Y(_0465_));
 sky130_fd_sc_hd__inv_2 _0678_ (.A(_0110_),
    .Y(_0462_));
 sky130_fd_sc_hd__inv_2 _0679_ (.A(_0110_),
    .Y(_0466_));
 sky130_fd_sc_hd__inv_2 _0680_ (.A(_0110_),
    .Y(_0461_));
 sky130_fd_sc_hd__buf_8 _0681_ (.A(_0109_),
    .X(_0111_));
 sky130_fd_sc_hd__inv_2 _0682_ (.A(_0111_),
    .Y(_0467_));
 sky130_fd_sc_hd__inv_2 _0683_ (.A(_0111_),
    .Y(_0460_));
 sky130_fd_sc_hd__inv_2 _0684_ (.A(_0111_),
    .Y(_0468_));
 sky130_fd_sc_hd__inv_2 _0685_ (.A(_0111_),
    .Y(_0469_));
 sky130_fd_sc_hd__inv_2 _0686_ (.A(_0111_),
    .Y(_0470_));
 sky130_fd_sc_hd__inv_2 _0687_ (.A(_0111_),
    .Y(_0471_));
 sky130_fd_sc_hd__inv_2 _0688_ (.A(_0111_),
    .Y(_0472_));
 sky130_fd_sc_hd__inv_2 _0689_ (.A(_0111_),
    .Y(_0473_));
 sky130_fd_sc_hd__inv_2 _0690_ (.A(_0111_),
    .Y(_0474_));
 sky130_fd_sc_hd__inv_2 _0691_ (.A(_0111_),
    .Y(_0475_));
 sky130_fd_sc_hd__buf_8 _0692_ (.A(_0108_),
    .X(_0112_));
 sky130_fd_sc_hd__inv_2 _0693_ (.A(_0112_),
    .Y(_0481_));
 sky130_fd_sc_hd__inv_2 _0694_ (.A(_0112_),
    .Y(_0480_));
 sky130_fd_sc_hd__inv_2 _0695_ (.A(_0112_),
    .Y(_0482_));
 sky130_fd_sc_hd__inv_2 _0696_ (.A(_0112_),
    .Y(_0479_));
 sky130_fd_sc_hd__inv_2 _0697_ (.A(_0112_),
    .Y(_0483_));
 sky130_fd_sc_hd__inv_2 _0698_ (.A(_0112_),
    .Y(_0478_));
 sky130_fd_sc_hd__inv_2 _0699_ (.A(_0112_),
    .Y(_0484_));
 sky130_fd_sc_hd__inv_2 _0700_ (.A(_0112_),
    .Y(_0477_));
 sky130_fd_sc_hd__inv_2 _0701_ (.A(_0112_),
    .Y(_0485_));
 sky130_fd_sc_hd__inv_2 _0702_ (.A(_0112_),
    .Y(_0486_));
 sky130_fd_sc_hd__buf_8 _0703_ (.A(_0108_),
    .X(_0113_));
 sky130_fd_sc_hd__inv_2 _0704_ (.A(_0113_),
    .Y(_0488_));
 sky130_fd_sc_hd__inv_2 _0705_ (.A(_0113_),
    .Y(_0489_));
 sky130_fd_sc_hd__inv_2 _0706_ (.A(_0113_),
    .Y(_0490_));
 sky130_fd_sc_hd__inv_2 _0707_ (.A(_0113_),
    .Y(_0491_));
 sky130_fd_sc_hd__inv_2 _0708_ (.A(_0113_),
    .Y(_0492_));
 sky130_fd_sc_hd__inv_2 _0709_ (.A(_0113_),
    .Y(_0493_));
 sky130_fd_sc_hd__inv_2 _0710_ (.A(_0113_),
    .Y(_0499_));
 sky130_fd_sc_hd__inv_2 _0711_ (.A(_0113_),
    .Y(_0498_));
 sky130_fd_sc_hd__inv_2 _0712_ (.A(_0113_),
    .Y(_0500_));
 sky130_fd_sc_hd__inv_2 _0713_ (.A(_0113_),
    .Y(_0497_));
 sky130_fd_sc_hd__buf_8 _0714_ (.A(_0108_),
    .X(_0114_));
 sky130_fd_sc_hd__inv_2 _0715_ (.A(_0114_),
    .Y(_0501_));
 sky130_fd_sc_hd__inv_2 _0716_ (.A(_0114_),
    .Y(_0496_));
 sky130_fd_sc_hd__inv_2 _0717_ (.A(_0114_),
    .Y(_0502_));
 sky130_fd_sc_hd__inv_2 _0718_ (.A(_0114_),
    .Y(_0495_));
 sky130_fd_sc_hd__inv_2 _0719_ (.A(_0114_),
    .Y(_0503_));
 sky130_fd_sc_hd__inv_2 _0720_ (.A(_0114_),
    .Y(_0504_));
 sky130_fd_sc_hd__inv_2 _0721_ (.A(_0114_),
    .Y(_0505_));
 sky130_fd_sc_hd__inv_2 _0722_ (.A(_0114_),
    .Y(_0506_));
 sky130_fd_sc_hd__inv_2 _0723_ (.A(_0114_),
    .Y(_0507_));
 sky130_fd_sc_hd__inv_2 _0724_ (.A(_0114_),
    .Y(_0508_));
 sky130_fd_sc_hd__buf_8 _0725_ (.A(_0108_),
    .X(_0115_));
 sky130_fd_sc_hd__inv_2 _0726_ (.A(_0115_),
    .Y(_0509_));
 sky130_fd_sc_hd__inv_2 _0727_ (.A(_0115_),
    .Y(_0510_));
 sky130_fd_sc_hd__inv_2 _0728_ (.A(_0115_),
    .Y(_0516_));
 sky130_fd_sc_hd__inv_2 _0729_ (.A(_0115_),
    .Y(_0515_));
 sky130_fd_sc_hd__inv_2 _0730_ (.A(_0115_),
    .Y(_0517_));
 sky130_fd_sc_hd__inv_2 _0731_ (.A(_0115_),
    .Y(_0514_));
 sky130_fd_sc_hd__inv_2 _0732_ (.A(_0115_),
    .Y(_0518_));
 sky130_fd_sc_hd__inv_2 _0733_ (.A(_0115_),
    .Y(_0513_));
 sky130_fd_sc_hd__inv_2 _0734_ (.A(_0115_),
    .Y(_0519_));
 sky130_fd_sc_hd__inv_2 _0735_ (.A(_0115_),
    .Y(_0512_));
 sky130_fd_sc_hd__buf_8 _0736_ (.A(_0108_),
    .X(_0116_));
 sky130_fd_sc_hd__inv_2 _0737_ (.A(_0116_),
    .Y(_0520_));
 sky130_fd_sc_hd__inv_2 _0738_ (.A(_0116_),
    .Y(_0521_));
 sky130_fd_sc_hd__inv_2 _0739_ (.A(_0116_),
    .Y(_0522_));
 sky130_fd_sc_hd__inv_2 _0740_ (.A(_0116_),
    .Y(_0523_));
 sky130_fd_sc_hd__inv_2 _0741_ (.A(_0116_),
    .Y(_0524_));
 sky130_fd_sc_hd__inv_2 _0742_ (.A(_0116_),
    .Y(_0526_));
 sky130_fd_sc_hd__inv_2 _0743_ (.A(_0116_),
    .Y(_0527_));
 sky130_fd_sc_hd__inv_2 _0744_ (.A(_0116_),
    .Y(_0528_));
 sky130_fd_sc_hd__inv_2 _0745_ (.A(_0116_),
    .Y(_0534_));
 sky130_fd_sc_hd__inv_2 _0746_ (.A(_0116_),
    .Y(_0533_));
 sky130_fd_sc_hd__buf_6 _0747_ (.A(_0108_),
    .X(_0117_));
 sky130_fd_sc_hd__inv_2 _0748_ (.A(_0117_),
    .Y(_0535_));
 sky130_fd_sc_hd__inv_2 _0749_ (.A(_0117_),
    .Y(_0532_));
 sky130_fd_sc_hd__inv_2 _0750_ (.A(_0117_),
    .Y(_0536_));
 sky130_fd_sc_hd__inv_2 _0751_ (.A(_0117_),
    .Y(_0531_));
 sky130_fd_sc_hd__inv_2 _0752_ (.A(_0117_),
    .Y(_0537_));
 sky130_fd_sc_hd__inv_2 _0753_ (.A(_0117_),
    .Y(_0530_));
 sky130_fd_sc_hd__inv_2 _0754_ (.A(_0117_),
    .Y(_0538_));
 sky130_fd_sc_hd__inv_2 _0755_ (.A(_0117_),
    .Y(_0539_));
 sky130_fd_sc_hd__inv_2 _0756_ (.A(_0117_),
    .Y(_0540_));
 sky130_fd_sc_hd__inv_2 _0757_ (.A(_0117_),
    .Y(_0541_));
 sky130_fd_sc_hd__buf_8 _0758_ (.A(_0108_),
    .X(_0118_));
 sky130_fd_sc_hd__inv_2 _0759_ (.A(_0118_),
    .Y(_0542_));
 sky130_fd_sc_hd__inv_2 _0760_ (.A(_0118_),
    .Y(_0543_));
 sky130_fd_sc_hd__inv_2 _0761_ (.A(_0118_),
    .Y(_0544_));
 sky130_fd_sc_hd__inv_2 _0762_ (.A(_0118_),
    .Y(_0545_));
 sky130_fd_sc_hd__inv_2 _0763_ (.A(_0118_),
    .Y(_0546_));
 sky130_fd_sc_hd__inv_2 _0764_ (.A(_0118_),
    .Y(_0547_));
 sky130_fd_sc_hd__inv_2 _0765_ (.A(_0118_),
    .Y(_0548_));
 sky130_fd_sc_hd__inv_2 _0766_ (.A(_0118_),
    .Y(_0549_));
 sky130_fd_sc_hd__inv_2 _0767_ (.A(_0118_),
    .Y(_0550_));
 sky130_fd_sc_hd__inv_2 _0768_ (.A(_0118_),
    .Y(_0459_));
 sky130_fd_sc_hd__buf_8 _0769_ (.A(_0108_),
    .X(_0119_));
 sky130_fd_sc_hd__inv_2 _0770_ (.A(_0119_),
    .Y(_0476_));
 sky130_fd_sc_hd__inv_2 _0771_ (.A(_0119_),
    .Y(_0494_));
 sky130_fd_sc_hd__inv_2 _0772_ (.A(_0119_),
    .Y(_0511_));
 sky130_fd_sc_hd__inv_2 _0773_ (.A(_0119_),
    .Y(_0529_));
 sky130_fd_sc_hd__inv_2 _0774_ (.A(_0119_),
    .Y(_0551_));
 sky130_fd_sc_hd__inv_2 _0775_ (.A(_0119_),
    .Y(_0552_));
 sky130_fd_sc_hd__inv_2 _0776_ (.A(_0119_),
    .Y(_0553_));
 sky130_fd_sc_hd__inv_2 _0777_ (.A(_0119_),
    .Y(_0554_));
 sky130_fd_sc_hd__inv_2 _0778_ (.A(_0119_),
    .Y(_0555_));
 sky130_fd_sc_hd__inv_2 _0779_ (.A(_0119_),
    .Y(_0556_));
 sky130_fd_sc_hd__inv_2 _0780_ (.A(_0109_),
    .Y(_0557_));
 sky130_fd_sc_hd__inv_2 _0781_ (.A(_0109_),
    .Y(_0558_));
 sky130_fd_sc_hd__inv_2 _0782_ (.A(_0109_),
    .Y(_0559_));
 sky130_fd_sc_hd__inv_2 _0783_ (.A(_0109_),
    .Y(_0560_));
 sky130_fd_sc_hd__inv_2 _0784_ (.A(_0109_),
    .Y(_0561_));
 sky130_fd_sc_hd__inv_2 _0785_ (.A(_0109_),
    .Y(_0562_));
 sky130_fd_sc_hd__inv_2 _0786_ (.A(_0109_),
    .Y(_0525_));
 sky130_fd_sc_hd__inv_2 _0787_ (.A(_0109_),
    .Y(_0487_));
 sky130_fd_sc_hd__clkinv_2 _0788_ (.A(net8),
    .Y(_0120_));
 sky130_fd_sc_hd__buf_2 _0789_ (.A(_0120_),
    .X(_0121_));
 sky130_fd_sc_hd__or2b_1 _0790_ (.A(\rgb_mixer0.enc2[7] ),
    .B_N(\rgb_mixer0.pwm2.count[7] ),
    .X(_0122_));
 sky130_fd_sc_hd__inv_2 _0791_ (.A(\rgb_mixer0.pwm2.count[7] ),
    .Y(_0123_));
 sky130_fd_sc_hd__inv_2 _0792_ (.A(\rgb_mixer0.pwm2.count[6] ),
    .Y(_0124_));
 sky130_fd_sc_hd__inv_2 _0793_ (.A(\rgb_mixer0.pwm2.count[5] ),
    .Y(_0125_));
 sky130_fd_sc_hd__inv_2 _0794_ (.A(\rgb_mixer0.pwm2.count[4] ),
    .Y(_0126_));
 sky130_fd_sc_hd__inv_2 _0795_ (.A(\rgb_mixer0.pwm2.count[3] ),
    .Y(_0127_));
 sky130_fd_sc_hd__o22a_1 _0796_ (.A1(\rgb_mixer0.enc2[4] ),
    .A2(_0126_),
    .B1(_0127_),
    .B2(\rgb_mixer0.enc2[3] ),
    .X(_0128_));
 sky130_fd_sc_hd__inv_2 _0797_ (.A(\rgb_mixer0.pwm2.count[2] ),
    .Y(_0129_));
 sky130_fd_sc_hd__inv_2 _0798_ (.A(\rgb_mixer0.pwm2.count[1] ),
    .Y(_0130_));
 sky130_fd_sc_hd__o22a_1 _0799_ (.A1(\rgb_mixer0.enc2[2] ),
    .A2(_0129_),
    .B1(_0130_),
    .B2(\rgb_mixer0.enc2[1] ),
    .X(_0131_));
 sky130_fd_sc_hd__inv_2 _0800_ (.A(\rgb_mixer0.enc2[0] ),
    .Y(_0132_));
 sky130_fd_sc_hd__nand2_1 _0801_ (.A(_0132_),
    .B(\rgb_mixer0.pwm2.count[0] ),
    .Y(_0133_));
 sky130_fd_sc_hd__o21ai_1 _0802_ (.A1(_0132_),
    .A2(\rgb_mixer0.pwm2.count[0] ),
    .B1(_0122_),
    .Y(_0134_));
 sky130_fd_sc_hd__a22o_1 _0803_ (.A1(\rgb_mixer0.enc2[1] ),
    .A2(_0130_),
    .B1(_0133_),
    .B2(_0134_),
    .X(_0135_));
 sky130_fd_sc_hd__a22o_1 _0804_ (.A1(\rgb_mixer0.enc2[3] ),
    .A2(_0127_),
    .B1(_0129_),
    .B2(\rgb_mixer0.enc2[2] ),
    .X(_0136_));
 sky130_fd_sc_hd__a21o_1 _0805_ (.A1(_0131_),
    .A2(_0135_),
    .B1(_0136_),
    .X(_0137_));
 sky130_fd_sc_hd__a22o_1 _0806_ (.A1(\rgb_mixer0.enc2[5] ),
    .A2(_0125_),
    .B1(_0126_),
    .B2(\rgb_mixer0.enc2[4] ),
    .X(_0138_));
 sky130_fd_sc_hd__a21o_1 _0807_ (.A1(_0128_),
    .A2(_0137_),
    .B1(_0138_),
    .X(_0139_));
 sky130_fd_sc_hd__o221a_1 _0808_ (.A1(\rgb_mixer0.enc2[6] ),
    .A2(_0124_),
    .B1(_0125_),
    .B2(\rgb_mixer0.enc2[5] ),
    .C1(_0139_),
    .X(_0140_));
 sky130_fd_sc_hd__a221o_1 _0809_ (.A1(\rgb_mixer0.enc2[7] ),
    .A2(_0123_),
    .B1(_0124_),
    .B2(\rgb_mixer0.enc2[6] ),
    .C1(_0140_),
    .X(_0141_));
 sky130_fd_sc_hd__and3_1 _0810_ (.A(_0121_),
    .B(_0122_),
    .C(_0141_),
    .X(_0142_));
 sky130_fd_sc_hd__clkbuf_1 _0811_ (.A(_0142_),
    .X(\rgb_mixer0.pwm2.out ));
 sky130_fd_sc_hd__or2b_1 _0812_ (.A(\rgb_mixer0.enc1[7] ),
    .B_N(\rgb_mixer0.pwm1.count[7] ),
    .X(_0143_));
 sky130_fd_sc_hd__inv_2 _0813_ (.A(\rgb_mixer0.pwm1.count[7] ),
    .Y(_0144_));
 sky130_fd_sc_hd__inv_2 _0814_ (.A(\rgb_mixer0.pwm1.count[6] ),
    .Y(_0145_));
 sky130_fd_sc_hd__and2b_1 _0815_ (.A_N(\rgb_mixer0.pwm1.count[5] ),
    .B(\rgb_mixer0.enc1[5] ),
    .X(_0146_));
 sky130_fd_sc_hd__inv_2 _0816_ (.A(\rgb_mixer0.pwm1.count[4] ),
    .Y(_0147_));
 sky130_fd_sc_hd__inv_2 _0817_ (.A(\rgb_mixer0.pwm1.count[3] ),
    .Y(_0148_));
 sky130_fd_sc_hd__o22a_1 _0818_ (.A1(\rgb_mixer0.enc1[4] ),
    .A2(_0147_),
    .B1(_0148_),
    .B2(\rgb_mixer0.enc1[3] ),
    .X(_0149_));
 sky130_fd_sc_hd__inv_2 _0819_ (.A(\rgb_mixer0.pwm1.count[2] ),
    .Y(_0150_));
 sky130_fd_sc_hd__inv_2 _0820_ (.A(\rgb_mixer0.pwm1.count[1] ),
    .Y(_0151_));
 sky130_fd_sc_hd__o22a_1 _0821_ (.A1(\rgb_mixer0.enc1[2] ),
    .A2(_0150_),
    .B1(_0151_),
    .B2(\rgb_mixer0.enc1[1] ),
    .X(_0152_));
 sky130_fd_sc_hd__inv_2 _0822_ (.A(\rgb_mixer0.enc1[0] ),
    .Y(_0153_));
 sky130_fd_sc_hd__nand2_1 _0823_ (.A(_0153_),
    .B(\rgb_mixer0.pwm1.count[0] ),
    .Y(_0154_));
 sky130_fd_sc_hd__o21ai_1 _0824_ (.A1(_0153_),
    .A2(\rgb_mixer0.pwm1.count[0] ),
    .B1(_0143_),
    .Y(_0155_));
 sky130_fd_sc_hd__a22o_1 _0825_ (.A1(\rgb_mixer0.enc1[1] ),
    .A2(_0151_),
    .B1(_0154_),
    .B2(_0155_),
    .X(_0156_));
 sky130_fd_sc_hd__a22o_1 _0826_ (.A1(\rgb_mixer0.enc1[3] ),
    .A2(_0148_),
    .B1(_0150_),
    .B2(\rgb_mixer0.enc1[2] ),
    .X(_0157_));
 sky130_fd_sc_hd__a21o_1 _0827_ (.A1(_0152_),
    .A2(_0156_),
    .B1(_0157_),
    .X(_0158_));
 sky130_fd_sc_hd__a22o_1 _0828_ (.A1(\rgb_mixer0.enc1[4] ),
    .A2(_0147_),
    .B1(_0149_),
    .B2(_0158_),
    .X(_0159_));
 sky130_fd_sc_hd__or2b_1 _0829_ (.A(\rgb_mixer0.enc1[5] ),
    .B_N(\rgb_mixer0.pwm1.count[5] ),
    .X(_0160_));
 sky130_fd_sc_hd__o221a_1 _0830_ (.A1(\rgb_mixer0.enc1[6] ),
    .A2(_0145_),
    .B1(_0146_),
    .B2(_0159_),
    .C1(_0160_),
    .X(_0161_));
 sky130_fd_sc_hd__a221o_1 _0831_ (.A1(\rgb_mixer0.enc1[7] ),
    .A2(_0144_),
    .B1(_0145_),
    .B2(\rgb_mixer0.enc1[6] ),
    .C1(_0161_),
    .X(_0162_));
 sky130_fd_sc_hd__and3_1 _0832_ (.A(_0121_),
    .B(_0143_),
    .C(_0162_),
    .X(_0163_));
 sky130_fd_sc_hd__clkbuf_1 _0833_ (.A(_0163_),
    .X(\rgb_mixer0.pwm1.out ));
 sky130_fd_sc_hd__or2b_1 _0834_ (.A(\rgb_mixer0.enc0[7] ),
    .B_N(\rgb_mixer0.pwm0.count[7] ),
    .X(_0164_));
 sky130_fd_sc_hd__inv_2 _0835_ (.A(\rgb_mixer0.pwm0.count[7] ),
    .Y(_0165_));
 sky130_fd_sc_hd__inv_2 _0836_ (.A(\rgb_mixer0.pwm0.count[6] ),
    .Y(_0166_));
 sky130_fd_sc_hd__inv_2 _0837_ (.A(\rgb_mixer0.pwm0.count[5] ),
    .Y(_0167_));
 sky130_fd_sc_hd__inv_2 _0838_ (.A(\rgb_mixer0.pwm0.count[4] ),
    .Y(_0168_));
 sky130_fd_sc_hd__inv_2 _0839_ (.A(\rgb_mixer0.pwm0.count[3] ),
    .Y(_0169_));
 sky130_fd_sc_hd__o22a_1 _0840_ (.A1(\rgb_mixer0.enc0[4] ),
    .A2(_0168_),
    .B1(_0169_),
    .B2(\rgb_mixer0.enc0[3] ),
    .X(_0170_));
 sky130_fd_sc_hd__inv_2 _0841_ (.A(\rgb_mixer0.pwm0.count[2] ),
    .Y(_0171_));
 sky130_fd_sc_hd__inv_2 _0842_ (.A(\rgb_mixer0.pwm0.count[1] ),
    .Y(_0172_));
 sky130_fd_sc_hd__o22a_1 _0843_ (.A1(\rgb_mixer0.enc0[2] ),
    .A2(_0171_),
    .B1(_0172_),
    .B2(\rgb_mixer0.enc0[1] ),
    .X(_0173_));
 sky130_fd_sc_hd__inv_2 _0844_ (.A(\rgb_mixer0.enc0[0] ),
    .Y(_0174_));
 sky130_fd_sc_hd__nand2_1 _0845_ (.A(_0174_),
    .B(\rgb_mixer0.pwm0.count[0] ),
    .Y(_0175_));
 sky130_fd_sc_hd__o21ai_1 _0846_ (.A1(_0174_),
    .A2(\rgb_mixer0.pwm0.count[0] ),
    .B1(_0164_),
    .Y(_0176_));
 sky130_fd_sc_hd__a22o_1 _0847_ (.A1(\rgb_mixer0.enc0[1] ),
    .A2(_0172_),
    .B1(_0175_),
    .B2(_0176_),
    .X(_0177_));
 sky130_fd_sc_hd__a22o_1 _0848_ (.A1(\rgb_mixer0.enc0[3] ),
    .A2(_0169_),
    .B1(_0171_),
    .B2(\rgb_mixer0.enc0[2] ),
    .X(_0178_));
 sky130_fd_sc_hd__a21o_1 _0849_ (.A1(_0173_),
    .A2(_0177_),
    .B1(_0178_),
    .X(_0179_));
 sky130_fd_sc_hd__a22o_1 _0850_ (.A1(\rgb_mixer0.enc0[5] ),
    .A2(_0167_),
    .B1(_0168_),
    .B2(\rgb_mixer0.enc0[4] ),
    .X(_0180_));
 sky130_fd_sc_hd__a21o_1 _0851_ (.A1(_0170_),
    .A2(_0179_),
    .B1(_0180_),
    .X(_0181_));
 sky130_fd_sc_hd__o221a_1 _0852_ (.A1(\rgb_mixer0.enc0[6] ),
    .A2(_0166_),
    .B1(_0167_),
    .B2(\rgb_mixer0.enc0[5] ),
    .C1(_0181_),
    .X(_0182_));
 sky130_fd_sc_hd__a221o_1 _0853_ (.A1(\rgb_mixer0.enc0[7] ),
    .A2(_0165_),
    .B1(_0166_),
    .B2(\rgb_mixer0.enc0[6] ),
    .C1(_0182_),
    .X(_0183_));
 sky130_fd_sc_hd__and3_1 _0854_ (.A(_0121_),
    .B(_0164_),
    .C(_0183_),
    .X(_0184_));
 sky130_fd_sc_hd__clkbuf_1 _0855_ (.A(_0184_),
    .X(\rgb_mixer0.pwm0.out ));
 sky130_fd_sc_hd__clkbuf_4 _0856_ (.A(net8),
    .X(_0185_));
 sky130_fd_sc_hd__nor2_1 _0857_ (.A(_0185_),
    .B(\rgb_mixer0.pwm2.count[0] ),
    .Y(_0000_));
 sky130_fd_sc_hd__clkbuf_4 _0858_ (.A(net8),
    .X(_0186_));
 sky130_fd_sc_hd__a21oi_1 _0859_ (.A1(\rgb_mixer0.pwm2.count[1] ),
    .A2(\rgb_mixer0.pwm2.count[0] ),
    .B1(_0186_),
    .Y(_0187_));
 sky130_fd_sc_hd__o21a_1 _0860_ (.A1(\rgb_mixer0.pwm2.count[1] ),
    .A2(\rgb_mixer0.pwm2.count[0] ),
    .B1(_0187_),
    .X(_0001_));
 sky130_fd_sc_hd__a21oi_1 _0861_ (.A1(\rgb_mixer0.pwm2.count[1] ),
    .A2(\rgb_mixer0.pwm2.count[0] ),
    .B1(\rgb_mixer0.pwm2.count[2] ),
    .Y(_0188_));
 sky130_fd_sc_hd__and3_1 _0862_ (.A(\rgb_mixer0.pwm2.count[2] ),
    .B(\rgb_mixer0.pwm2.count[1] ),
    .C(\rgb_mixer0.pwm2.count[0] ),
    .X(_0189_));
 sky130_fd_sc_hd__nor3_1 _0863_ (.A(_0185_),
    .B(_0188_),
    .C(_0189_),
    .Y(_0002_));
 sky130_fd_sc_hd__and2_1 _0864_ (.A(\rgb_mixer0.pwm2.count[3] ),
    .B(_0189_),
    .X(_0190_));
 sky130_fd_sc_hd__clkbuf_4 _0865_ (.A(_0121_),
    .X(_0191_));
 sky130_fd_sc_hd__o21ai_1 _0866_ (.A1(\rgb_mixer0.pwm2.count[3] ),
    .A2(_0189_),
    .B1(_0191_),
    .Y(_0192_));
 sky130_fd_sc_hd__nor2_1 _0867_ (.A(_0190_),
    .B(_0192_),
    .Y(_0003_));
 sky130_fd_sc_hd__a21oi_1 _0868_ (.A1(\rgb_mixer0.pwm2.count[4] ),
    .A2(_0190_),
    .B1(_0186_),
    .Y(_0193_));
 sky130_fd_sc_hd__o21a_1 _0869_ (.A1(\rgb_mixer0.pwm2.count[4] ),
    .A2(_0190_),
    .B1(_0193_),
    .X(_0004_));
 sky130_fd_sc_hd__a21oi_1 _0870_ (.A1(\rgb_mixer0.pwm2.count[4] ),
    .A2(_0190_),
    .B1(\rgb_mixer0.pwm2.count[5] ),
    .Y(_0194_));
 sky130_fd_sc_hd__and3_1 _0871_ (.A(\rgb_mixer0.pwm2.count[5] ),
    .B(\rgb_mixer0.pwm2.count[4] ),
    .C(_0190_),
    .X(_0195_));
 sky130_fd_sc_hd__nor3_1 _0872_ (.A(_0185_),
    .B(_0194_),
    .C(_0195_),
    .Y(_0005_));
 sky130_fd_sc_hd__and2_1 _0873_ (.A(\rgb_mixer0.pwm2.count[6] ),
    .B(_0195_),
    .X(_0196_));
 sky130_fd_sc_hd__o21ai_1 _0874_ (.A1(\rgb_mixer0.pwm2.count[6] ),
    .A2(_0195_),
    .B1(_0191_),
    .Y(_0197_));
 sky130_fd_sc_hd__nor2_1 _0875_ (.A(_0196_),
    .B(_0197_),
    .Y(_0006_));
 sky130_fd_sc_hd__a21oi_1 _0876_ (.A1(\rgb_mixer0.pwm2.count[7] ),
    .A2(_0196_),
    .B1(_0186_),
    .Y(_0198_));
 sky130_fd_sc_hd__o21a_1 _0877_ (.A1(\rgb_mixer0.pwm2.count[7] ),
    .A2(_0196_),
    .B1(_0198_),
    .X(_0007_));
 sky130_fd_sc_hd__nor2_1 _0878_ (.A(_0185_),
    .B(\rgb_mixer0.pwm1.count[0] ),
    .Y(_0008_));
 sky130_fd_sc_hd__a21oi_1 _0879_ (.A1(\rgb_mixer0.pwm1.count[1] ),
    .A2(\rgb_mixer0.pwm1.count[0] ),
    .B1(_0186_),
    .Y(_0199_));
 sky130_fd_sc_hd__o21a_1 _0880_ (.A1(\rgb_mixer0.pwm1.count[1] ),
    .A2(\rgb_mixer0.pwm1.count[0] ),
    .B1(_0199_),
    .X(_0009_));
 sky130_fd_sc_hd__a21oi_1 _0881_ (.A1(\rgb_mixer0.pwm1.count[1] ),
    .A2(\rgb_mixer0.pwm1.count[0] ),
    .B1(\rgb_mixer0.pwm1.count[2] ),
    .Y(_0200_));
 sky130_fd_sc_hd__and3_1 _0882_ (.A(\rgb_mixer0.pwm1.count[2] ),
    .B(\rgb_mixer0.pwm1.count[1] ),
    .C(\rgb_mixer0.pwm1.count[0] ),
    .X(_0201_));
 sky130_fd_sc_hd__nor3_1 _0883_ (.A(_0185_),
    .B(_0200_),
    .C(_0201_),
    .Y(_0010_));
 sky130_fd_sc_hd__and2_1 _0884_ (.A(\rgb_mixer0.pwm1.count[3] ),
    .B(_0201_),
    .X(_0202_));
 sky130_fd_sc_hd__o21ai_1 _0885_ (.A1(\rgb_mixer0.pwm1.count[3] ),
    .A2(_0201_),
    .B1(_0191_),
    .Y(_0203_));
 sky130_fd_sc_hd__nor2_1 _0886_ (.A(_0202_),
    .B(_0203_),
    .Y(_0011_));
 sky130_fd_sc_hd__and3_1 _0887_ (.A(\rgb_mixer0.pwm1.count[4] ),
    .B(\rgb_mixer0.pwm1.count[3] ),
    .C(_0201_),
    .X(_0204_));
 sky130_fd_sc_hd__o21ai_1 _0888_ (.A1(\rgb_mixer0.pwm1.count[4] ),
    .A2(_0202_),
    .B1(_0191_),
    .Y(_0205_));
 sky130_fd_sc_hd__nor2_1 _0889_ (.A(_0204_),
    .B(_0205_),
    .Y(_0012_));
 sky130_fd_sc_hd__and2_1 _0890_ (.A(\rgb_mixer0.pwm1.count[5] ),
    .B(_0204_),
    .X(_0206_));
 sky130_fd_sc_hd__nor2_1 _0891_ (.A(net8),
    .B(_0206_),
    .Y(_0207_));
 sky130_fd_sc_hd__o21a_1 _0892_ (.A1(\rgb_mixer0.pwm1.count[5] ),
    .A2(_0204_),
    .B1(_0207_),
    .X(_0013_));
 sky130_fd_sc_hd__and3_1 _0893_ (.A(\rgb_mixer0.pwm1.count[6] ),
    .B(\rgb_mixer0.pwm1.count[5] ),
    .C(_0204_),
    .X(_0208_));
 sky130_fd_sc_hd__o21ai_1 _0894_ (.A1(\rgb_mixer0.pwm1.count[6] ),
    .A2(_0206_),
    .B1(_0191_),
    .Y(_0209_));
 sky130_fd_sc_hd__nor2_1 _0895_ (.A(_0208_),
    .B(_0209_),
    .Y(_0014_));
 sky130_fd_sc_hd__a21oi_1 _0896_ (.A1(\rgb_mixer0.pwm1.count[7] ),
    .A2(_0208_),
    .B1(_0186_),
    .Y(_0210_));
 sky130_fd_sc_hd__o21a_1 _0897_ (.A1(\rgb_mixer0.pwm1.count[7] ),
    .A2(_0208_),
    .B1(_0210_),
    .X(_0015_));
 sky130_fd_sc_hd__nor2_1 _0898_ (.A(_0185_),
    .B(\rgb_mixer0.pwm0.count[0] ),
    .Y(_0016_));
 sky130_fd_sc_hd__a21oi_1 _0899_ (.A1(\rgb_mixer0.pwm0.count[1] ),
    .A2(\rgb_mixer0.pwm0.count[0] ),
    .B1(_0186_),
    .Y(_0211_));
 sky130_fd_sc_hd__o21a_1 _0900_ (.A1(\rgb_mixer0.pwm0.count[1] ),
    .A2(\rgb_mixer0.pwm0.count[0] ),
    .B1(_0211_),
    .X(_0017_));
 sky130_fd_sc_hd__a21oi_1 _0901_ (.A1(\rgb_mixer0.pwm0.count[1] ),
    .A2(\rgb_mixer0.pwm0.count[0] ),
    .B1(\rgb_mixer0.pwm0.count[2] ),
    .Y(_0212_));
 sky130_fd_sc_hd__and3_1 _0902_ (.A(\rgb_mixer0.pwm0.count[2] ),
    .B(\rgb_mixer0.pwm0.count[1] ),
    .C(\rgb_mixer0.pwm0.count[0] ),
    .X(_0213_));
 sky130_fd_sc_hd__nor3_1 _0903_ (.A(_0185_),
    .B(_0212_),
    .C(_0213_),
    .Y(_0018_));
 sky130_fd_sc_hd__and2_1 _0904_ (.A(\rgb_mixer0.pwm0.count[3] ),
    .B(_0213_),
    .X(_0214_));
 sky130_fd_sc_hd__o21ai_1 _0905_ (.A1(\rgb_mixer0.pwm0.count[3] ),
    .A2(_0213_),
    .B1(_0191_),
    .Y(_0215_));
 sky130_fd_sc_hd__nor2_1 _0906_ (.A(_0214_),
    .B(_0215_),
    .Y(_0019_));
 sky130_fd_sc_hd__a21oi_1 _0907_ (.A1(\rgb_mixer0.pwm0.count[4] ),
    .A2(_0214_),
    .B1(_0186_),
    .Y(_0216_));
 sky130_fd_sc_hd__o21a_1 _0908_ (.A1(\rgb_mixer0.pwm0.count[4] ),
    .A2(_0214_),
    .B1(_0216_),
    .X(_0020_));
 sky130_fd_sc_hd__a21oi_1 _0909_ (.A1(\rgb_mixer0.pwm0.count[4] ),
    .A2(_0214_),
    .B1(\rgb_mixer0.pwm0.count[5] ),
    .Y(_0217_));
 sky130_fd_sc_hd__and3_1 _0910_ (.A(\rgb_mixer0.pwm0.count[5] ),
    .B(\rgb_mixer0.pwm0.count[4] ),
    .C(_0214_),
    .X(_0218_));
 sky130_fd_sc_hd__nor3_1 _0911_ (.A(_0185_),
    .B(_0217_),
    .C(_0218_),
    .Y(_0021_));
 sky130_fd_sc_hd__and2_1 _0912_ (.A(\rgb_mixer0.pwm0.count[6] ),
    .B(_0218_),
    .X(_0219_));
 sky130_fd_sc_hd__o21ai_1 _0913_ (.A1(\rgb_mixer0.pwm0.count[6] ),
    .A2(_0218_),
    .B1(_0191_),
    .Y(_0220_));
 sky130_fd_sc_hd__nor2_1 _0914_ (.A(_0219_),
    .B(_0220_),
    .Y(_0022_));
 sky130_fd_sc_hd__a21oi_1 _0915_ (.A1(\rgb_mixer0.pwm0.count[7] ),
    .A2(_0219_),
    .B1(_0186_),
    .Y(_0221_));
 sky130_fd_sc_hd__o21a_1 _0916_ (.A1(\rgb_mixer0.pwm0.count[7] ),
    .A2(_0219_),
    .B1(_0221_),
    .X(_0023_));
 sky130_fd_sc_hd__and2_1 _0917_ (.A(\rgb_mixer0.debounce2_b.debounced ),
    .B(_0120_),
    .X(_0222_));
 sky130_fd_sc_hd__clkbuf_1 _0918_ (.A(_0222_),
    .X(_0024_));
 sky130_fd_sc_hd__and2b_1 _0919_ (.A_N(\rgb_mixer0.debounce2_a.debounced ),
    .B(\rgb_mixer0.debounce2_b.debounced ),
    .X(_0223_));
 sky130_fd_sc_hd__and2b_1 _0920_ (.A_N(\rgb_mixer0.debounce2_b.debounced ),
    .B(\rgb_mixer0.debounce2_a.debounced ),
    .X(_0224_));
 sky130_fd_sc_hd__and2_1 _0921_ (.A(\rgb_mixer0.encoder2.old_b ),
    .B(\rgb_mixer0.encoder2.old_a ),
    .X(_0225_));
 sky130_fd_sc_hd__nor2_1 _0922_ (.A(\rgb_mixer0.encoder2.old_b ),
    .B(\rgb_mixer0.encoder2.old_a ),
    .Y(_0226_));
 sky130_fd_sc_hd__o22a_2 _0923_ (.A1(_0223_),
    .A2(_0224_),
    .B1(_0225_),
    .B2(_0226_),
    .X(_0227_));
 sky130_fd_sc_hd__buf_2 _0924_ (.A(_0227_),
    .X(_0228_));
 sky130_fd_sc_hd__a21oi_1 _0925_ (.A1(\rgb_mixer0.enc2[0] ),
    .A2(_0227_),
    .B1(_0186_),
    .Y(_0229_));
 sky130_fd_sc_hd__o21a_1 _0926_ (.A1(\rgb_mixer0.enc2[0] ),
    .A2(_0228_),
    .B1(_0229_),
    .X(_0025_));
 sky130_fd_sc_hd__and4b_1 _0927_ (.A_N(\rgb_mixer0.debounce2_b.debounced ),
    .B(\rgb_mixer0.encoder2.old_b ),
    .C(\rgb_mixer0.encoder2.old_a ),
    .D(\rgb_mixer0.debounce2_a.debounced ),
    .X(_0230_));
 sky130_fd_sc_hd__a21o_1 _0928_ (.A1(_0223_),
    .A2(_0226_),
    .B1(_0230_),
    .X(_0231_));
 sky130_fd_sc_hd__clkbuf_4 _0929_ (.A(_0231_),
    .X(_0232_));
 sky130_fd_sc_hd__nor2_1 _0930_ (.A(\rgb_mixer0.enc2[1] ),
    .B(_0232_),
    .Y(_0233_));
 sky130_fd_sc_hd__o221a_1 _0931_ (.A1(_0223_),
    .A2(_0225_),
    .B1(_0226_),
    .B2(_0224_),
    .C1(\rgb_mixer0.enc2[1] ),
    .X(_0234_));
 sky130_fd_sc_hd__nor2_1 _0932_ (.A(_0233_),
    .B(_0234_),
    .Y(_0235_));
 sky130_fd_sc_hd__xnor2_1 _0933_ (.A(\rgb_mixer0.enc2[0] ),
    .B(_0235_),
    .Y(_0236_));
 sky130_fd_sc_hd__nand2_1 _0934_ (.A(_0228_),
    .B(_0236_),
    .Y(_0237_));
 sky130_fd_sc_hd__clkbuf_4 _0935_ (.A(_0121_),
    .X(_0238_));
 sky130_fd_sc_hd__o211a_1 _0936_ (.A1(\rgb_mixer0.enc2[1] ),
    .A2(_0228_),
    .B1(_0237_),
    .C1(_0238_),
    .X(_0026_));
 sky130_fd_sc_hd__a211o_1 _0937_ (.A1(_0223_),
    .A2(_0226_),
    .B1(_0230_),
    .C1(\rgb_mixer0.enc2[1] ),
    .X(_0239_));
 sky130_fd_sc_hd__a21o_1 _0938_ (.A1(\rgb_mixer0.enc2[0] ),
    .A2(_0239_),
    .B1(_0234_),
    .X(_0240_));
 sky130_fd_sc_hd__xor2_1 _0939_ (.A(\rgb_mixer0.enc2[2] ),
    .B(_0231_),
    .X(_0241_));
 sky130_fd_sc_hd__or2_1 _0940_ (.A(_0240_),
    .B(_0241_),
    .X(_0242_));
 sky130_fd_sc_hd__nand2_1 _0941_ (.A(_0240_),
    .B(_0241_),
    .Y(_0243_));
 sky130_fd_sc_hd__a21bo_1 _0942_ (.A1(_0242_),
    .A2(_0243_),
    .B1_N(_0227_),
    .X(_0244_));
 sky130_fd_sc_hd__o211a_1 _0943_ (.A1(\rgb_mixer0.enc2[2] ),
    .A2(_0228_),
    .B1(_0244_),
    .C1(_0238_),
    .X(_0027_));
 sky130_fd_sc_hd__nand2_1 _0944_ (.A(\rgb_mixer0.enc2[2] ),
    .B(_0232_),
    .Y(_0245_));
 sky130_fd_sc_hd__xor2_1 _0945_ (.A(\rgb_mixer0.enc2[3] ),
    .B(_0231_),
    .X(_0246_));
 sky130_fd_sc_hd__and3_1 _0946_ (.A(_0245_),
    .B(_0243_),
    .C(_0246_),
    .X(_0247_));
 sky130_fd_sc_hd__a21o_1 _0947_ (.A1(_0245_),
    .A2(_0243_),
    .B1(_0246_),
    .X(_0248_));
 sky130_fd_sc_hd__nand2_1 _0948_ (.A(_0227_),
    .B(_0248_),
    .Y(_0249_));
 sky130_fd_sc_hd__clkbuf_4 _0949_ (.A(_0121_),
    .X(_0250_));
 sky130_fd_sc_hd__o221a_1 _0950_ (.A1(\rgb_mixer0.enc2[3] ),
    .A2(_0228_),
    .B1(_0247_),
    .B2(_0249_),
    .C1(_0250_),
    .X(_0028_));
 sky130_fd_sc_hd__o21a_1 _0951_ (.A1(\rgb_mixer0.enc2[3] ),
    .A2(\rgb_mixer0.enc2[2] ),
    .B1(_0232_),
    .X(_0251_));
 sky130_fd_sc_hd__a31o_1 _0952_ (.A1(_0240_),
    .A2(_0241_),
    .A3(_0246_),
    .B1(_0251_),
    .X(_0252_));
 sky130_fd_sc_hd__xor2_1 _0953_ (.A(\rgb_mixer0.enc2[4] ),
    .B(_0232_),
    .X(_0253_));
 sky130_fd_sc_hd__or2_1 _0954_ (.A(_0252_),
    .B(_0253_),
    .X(_0254_));
 sky130_fd_sc_hd__nand2_1 _0955_ (.A(_0252_),
    .B(_0253_),
    .Y(_0255_));
 sky130_fd_sc_hd__a21bo_1 _0956_ (.A1(_0254_),
    .A2(_0255_),
    .B1_N(_0227_),
    .X(_0256_));
 sky130_fd_sc_hd__o211a_1 _0957_ (.A1(\rgb_mixer0.enc2[4] ),
    .A2(_0228_),
    .B1(_0256_),
    .C1(_0238_),
    .X(_0029_));
 sky130_fd_sc_hd__xor2_1 _0958_ (.A(\rgb_mixer0.enc2[5] ),
    .B(_0232_),
    .X(_0257_));
 sky130_fd_sc_hd__a21bo_1 _0959_ (.A1(\rgb_mixer0.enc2[4] ),
    .A2(_0232_),
    .B1_N(_0255_),
    .X(_0258_));
 sky130_fd_sc_hd__xnor2_1 _0960_ (.A(_0257_),
    .B(_0258_),
    .Y(_0259_));
 sky130_fd_sc_hd__o21ai_1 _0961_ (.A1(\rgb_mixer0.enc2[5] ),
    .A2(_0227_),
    .B1(_0191_),
    .Y(_0260_));
 sky130_fd_sc_hd__a21oi_1 _0962_ (.A1(_0228_),
    .A2(_0259_),
    .B1(_0260_),
    .Y(_0030_));
 sky130_fd_sc_hd__nor2_1 _0963_ (.A(\rgb_mixer0.enc2[6] ),
    .B(_0232_),
    .Y(_0261_));
 sky130_fd_sc_hd__and2_1 _0964_ (.A(\rgb_mixer0.enc2[6] ),
    .B(_0232_),
    .X(_0262_));
 sky130_fd_sc_hd__nor2_1 _0965_ (.A(_0261_),
    .B(_0262_),
    .Y(_0263_));
 sky130_fd_sc_hd__o21a_1 _0966_ (.A1(\rgb_mixer0.enc2[5] ),
    .A2(\rgb_mixer0.enc2[4] ),
    .B1(_0232_),
    .X(_0264_));
 sky130_fd_sc_hd__a31o_1 _0967_ (.A1(_0252_),
    .A2(_0253_),
    .A3(_0257_),
    .B1(_0264_),
    .X(_0265_));
 sky130_fd_sc_hd__xnor2_1 _0968_ (.A(_0263_),
    .B(_0265_),
    .Y(_0266_));
 sky130_fd_sc_hd__nand2_1 _0969_ (.A(_0228_),
    .B(_0266_),
    .Y(_0267_));
 sky130_fd_sc_hd__o211a_1 _0970_ (.A1(\rgb_mixer0.enc2[6] ),
    .A2(_0228_),
    .B1(_0267_),
    .C1(_0238_),
    .X(_0031_));
 sky130_fd_sc_hd__a21o_1 _0971_ (.A1(_0263_),
    .A2(_0265_),
    .B1(_0262_),
    .X(_0268_));
 sky130_fd_sc_hd__xor2_1 _0972_ (.A(\rgb_mixer0.enc2[7] ),
    .B(_0232_),
    .X(_0269_));
 sky130_fd_sc_hd__xnor2_1 _0973_ (.A(_0268_),
    .B(_0269_),
    .Y(_0270_));
 sky130_fd_sc_hd__o21ai_1 _0974_ (.A1(\rgb_mixer0.enc2[7] ),
    .A2(_0227_),
    .B1(_0191_),
    .Y(_0271_));
 sky130_fd_sc_hd__a21oi_1 _0975_ (.A1(_0228_),
    .A2(_0270_),
    .B1(_0271_),
    .Y(_0032_));
 sky130_fd_sc_hd__clkbuf_4 _0976_ (.A(_0120_),
    .X(_0272_));
 sky130_fd_sc_hd__and2_1 _0977_ (.A(\rgb_mixer0.debounce1_b.debounced ),
    .B(_0272_),
    .X(_0273_));
 sky130_fd_sc_hd__clkbuf_1 _0978_ (.A(_0273_),
    .X(_0033_));
 sky130_fd_sc_hd__and2_1 _0979_ (.A(\rgb_mixer0.debounce2_a.debounced ),
    .B(_0272_),
    .X(_0274_));
 sky130_fd_sc_hd__clkbuf_1 _0980_ (.A(_0274_),
    .X(_0034_));
 sky130_fd_sc_hd__and2b_1 _0981_ (.A_N(\rgb_mixer0.debounce1_a.debounced ),
    .B(\rgb_mixer0.debounce1_b.debounced ),
    .X(_0275_));
 sky130_fd_sc_hd__and2b_1 _0982_ (.A_N(\rgb_mixer0.debounce1_b.debounced ),
    .B(\rgb_mixer0.debounce1_a.debounced ),
    .X(_0276_));
 sky130_fd_sc_hd__and2_1 _0983_ (.A(\rgb_mixer0.encoder1.old_b ),
    .B(\rgb_mixer0.encoder1.old_a ),
    .X(_0277_));
 sky130_fd_sc_hd__nor2_1 _0984_ (.A(\rgb_mixer0.encoder1.old_b ),
    .B(\rgb_mixer0.encoder1.old_a ),
    .Y(_0278_));
 sky130_fd_sc_hd__o22a_2 _0985_ (.A1(_0275_),
    .A2(_0276_),
    .B1(_0277_),
    .B2(_0278_),
    .X(_0279_));
 sky130_fd_sc_hd__buf_2 _0986_ (.A(_0279_),
    .X(_0280_));
 sky130_fd_sc_hd__a21oi_1 _0987_ (.A1(\rgb_mixer0.enc1[0] ),
    .A2(_0279_),
    .B1(_0186_),
    .Y(_0281_));
 sky130_fd_sc_hd__o21a_1 _0988_ (.A1(\rgb_mixer0.enc1[0] ),
    .A2(_0280_),
    .B1(_0281_),
    .X(_0035_));
 sky130_fd_sc_hd__and4b_1 _0989_ (.A_N(\rgb_mixer0.debounce1_b.debounced ),
    .B(\rgb_mixer0.encoder1.old_b ),
    .C(\rgb_mixer0.encoder1.old_a ),
    .D(\rgb_mixer0.debounce1_a.debounced ),
    .X(_0282_));
 sky130_fd_sc_hd__a21o_1 _0990_ (.A1(_0275_),
    .A2(_0278_),
    .B1(_0282_),
    .X(_0283_));
 sky130_fd_sc_hd__buf_2 _0991_ (.A(_0283_),
    .X(_0284_));
 sky130_fd_sc_hd__nor2_1 _0992_ (.A(\rgb_mixer0.enc1[1] ),
    .B(_0284_),
    .Y(_0285_));
 sky130_fd_sc_hd__o221a_1 _0993_ (.A1(_0275_),
    .A2(_0277_),
    .B1(_0278_),
    .B2(_0276_),
    .C1(\rgb_mixer0.enc1[1] ),
    .X(_0286_));
 sky130_fd_sc_hd__nor2_1 _0994_ (.A(_0285_),
    .B(_0286_),
    .Y(_0287_));
 sky130_fd_sc_hd__xnor2_1 _0995_ (.A(\rgb_mixer0.enc1[0] ),
    .B(_0287_),
    .Y(_0288_));
 sky130_fd_sc_hd__nand2_1 _0996_ (.A(_0280_),
    .B(_0288_),
    .Y(_0289_));
 sky130_fd_sc_hd__o211a_1 _0997_ (.A1(\rgb_mixer0.enc1[1] ),
    .A2(_0280_),
    .B1(_0289_),
    .C1(_0238_),
    .X(_0036_));
 sky130_fd_sc_hd__a211o_1 _0998_ (.A1(_0275_),
    .A2(_0278_),
    .B1(_0282_),
    .C1(\rgb_mixer0.enc1[1] ),
    .X(_0290_));
 sky130_fd_sc_hd__a21o_1 _0999_ (.A1(\rgb_mixer0.enc1[0] ),
    .A2(_0290_),
    .B1(_0286_),
    .X(_0291_));
 sky130_fd_sc_hd__xor2_1 _1000_ (.A(\rgb_mixer0.enc1[2] ),
    .B(_0283_),
    .X(_0292_));
 sky130_fd_sc_hd__or2_1 _1001_ (.A(_0291_),
    .B(_0292_),
    .X(_0293_));
 sky130_fd_sc_hd__nand2_1 _1002_ (.A(_0291_),
    .B(_0292_),
    .Y(_0294_));
 sky130_fd_sc_hd__a21bo_1 _1003_ (.A1(_0293_),
    .A2(_0294_),
    .B1_N(_0279_),
    .X(_0295_));
 sky130_fd_sc_hd__o211a_1 _1004_ (.A1(\rgb_mixer0.enc1[2] ),
    .A2(_0280_),
    .B1(_0295_),
    .C1(_0238_),
    .X(_0037_));
 sky130_fd_sc_hd__nand2_1 _1005_ (.A(\rgb_mixer0.enc1[2] ),
    .B(_0284_),
    .Y(_0296_));
 sky130_fd_sc_hd__xor2_1 _1006_ (.A(\rgb_mixer0.enc1[3] ),
    .B(_0283_),
    .X(_0297_));
 sky130_fd_sc_hd__and3_1 _1007_ (.A(_0296_),
    .B(_0294_),
    .C(_0297_),
    .X(_0298_));
 sky130_fd_sc_hd__a21o_1 _1008_ (.A1(_0296_),
    .A2(_0294_),
    .B1(_0297_),
    .X(_0299_));
 sky130_fd_sc_hd__nand2_1 _1009_ (.A(_0279_),
    .B(_0299_),
    .Y(_0300_));
 sky130_fd_sc_hd__o221a_1 _1010_ (.A1(\rgb_mixer0.enc1[3] ),
    .A2(_0280_),
    .B1(_0298_),
    .B2(_0300_),
    .C1(_0250_),
    .X(_0038_));
 sky130_fd_sc_hd__o21a_1 _1011_ (.A1(\rgb_mixer0.enc1[3] ),
    .A2(\rgb_mixer0.enc1[2] ),
    .B1(_0284_),
    .X(_0301_));
 sky130_fd_sc_hd__a31o_1 _1012_ (.A1(_0291_),
    .A2(_0292_),
    .A3(_0297_),
    .B1(_0301_),
    .X(_0302_));
 sky130_fd_sc_hd__xor2_1 _1013_ (.A(\rgb_mixer0.enc1[4] ),
    .B(_0284_),
    .X(_0303_));
 sky130_fd_sc_hd__or2_1 _1014_ (.A(_0302_),
    .B(_0303_),
    .X(_0304_));
 sky130_fd_sc_hd__nand2_1 _1015_ (.A(_0302_),
    .B(_0303_),
    .Y(_0305_));
 sky130_fd_sc_hd__a21bo_1 _1016_ (.A1(_0304_),
    .A2(_0305_),
    .B1_N(_0279_),
    .X(_0306_));
 sky130_fd_sc_hd__o211a_1 _1017_ (.A1(\rgb_mixer0.enc1[4] ),
    .A2(_0280_),
    .B1(_0306_),
    .C1(_0238_),
    .X(_0039_));
 sky130_fd_sc_hd__xor2_1 _1018_ (.A(\rgb_mixer0.enc1[5] ),
    .B(_0284_),
    .X(_0307_));
 sky130_fd_sc_hd__a21bo_1 _1019_ (.A1(\rgb_mixer0.enc1[4] ),
    .A2(_0284_),
    .B1_N(_0305_),
    .X(_0308_));
 sky130_fd_sc_hd__xnor2_1 _1020_ (.A(_0307_),
    .B(_0308_),
    .Y(_0309_));
 sky130_fd_sc_hd__nor2_1 _1021_ (.A(\rgb_mixer0.enc1[5] ),
    .B(_0279_),
    .Y(_0310_));
 sky130_fd_sc_hd__a211oi_1 _1022_ (.A1(_0280_),
    .A2(_0309_),
    .B1(_0310_),
    .C1(_0185_),
    .Y(_0040_));
 sky130_fd_sc_hd__nor2_1 _1023_ (.A(\rgb_mixer0.enc1[6] ),
    .B(_0284_),
    .Y(_0311_));
 sky130_fd_sc_hd__and2_1 _1024_ (.A(\rgb_mixer0.enc1[6] ),
    .B(_0284_),
    .X(_0312_));
 sky130_fd_sc_hd__nor2_1 _1025_ (.A(_0311_),
    .B(_0312_),
    .Y(_0313_));
 sky130_fd_sc_hd__o21a_1 _1026_ (.A1(\rgb_mixer0.enc1[5] ),
    .A2(\rgb_mixer0.enc1[4] ),
    .B1(_0284_),
    .X(_0314_));
 sky130_fd_sc_hd__a31o_1 _1027_ (.A1(_0302_),
    .A2(_0303_),
    .A3(_0307_),
    .B1(_0314_),
    .X(_0315_));
 sky130_fd_sc_hd__xnor2_1 _1028_ (.A(_0313_),
    .B(_0315_),
    .Y(_0316_));
 sky130_fd_sc_hd__nand2_1 _1029_ (.A(_0280_),
    .B(_0316_),
    .Y(_0317_));
 sky130_fd_sc_hd__o211a_1 _1030_ (.A1(\rgb_mixer0.enc1[6] ),
    .A2(_0280_),
    .B1(_0317_),
    .C1(_0238_),
    .X(_0041_));
 sky130_fd_sc_hd__a21o_1 _1031_ (.A1(_0313_),
    .A2(_0315_),
    .B1(_0312_),
    .X(_0318_));
 sky130_fd_sc_hd__xor2_1 _1032_ (.A(\rgb_mixer0.enc1[7] ),
    .B(_0284_),
    .X(_0319_));
 sky130_fd_sc_hd__xnor2_1 _1033_ (.A(_0318_),
    .B(_0319_),
    .Y(_0320_));
 sky130_fd_sc_hd__nor2_1 _1034_ (.A(\rgb_mixer0.enc1[7] ),
    .B(_0279_),
    .Y(_0321_));
 sky130_fd_sc_hd__a211oi_1 _1035_ (.A1(_0280_),
    .A2(_0320_),
    .B1(_0321_),
    .C1(_0185_),
    .Y(_0042_));
 sky130_fd_sc_hd__clkbuf_2 _1036_ (.A(_0121_),
    .X(_0322_));
 sky130_fd_sc_hd__and2_1 _1037_ (.A(\rgb_mixer0.debounce0_b.debounced ),
    .B(_0322_),
    .X(_0323_));
 sky130_fd_sc_hd__clkbuf_1 _1038_ (.A(_0323_),
    .X(_0043_));
 sky130_fd_sc_hd__and2_1 _1039_ (.A(\rgb_mixer0.debounce1_a.debounced ),
    .B(_0120_),
    .X(_0324_));
 sky130_fd_sc_hd__clkbuf_1 _1040_ (.A(_0324_),
    .X(_0044_));
 sky130_fd_sc_hd__and2b_1 _1041_ (.A_N(\rgb_mixer0.debounce0_a.debounced ),
    .B(\rgb_mixer0.debounce0_b.debounced ),
    .X(_0325_));
 sky130_fd_sc_hd__and2b_1 _1042_ (.A_N(\rgb_mixer0.debounce0_b.debounced ),
    .B(\rgb_mixer0.debounce0_a.debounced ),
    .X(_0326_));
 sky130_fd_sc_hd__and2_1 _1043_ (.A(\rgb_mixer0.encoder0.old_b ),
    .B(\rgb_mixer0.encoder0.old_a ),
    .X(_0327_));
 sky130_fd_sc_hd__nor2_1 _1044_ (.A(\rgb_mixer0.encoder0.old_b ),
    .B(\rgb_mixer0.encoder0.old_a ),
    .Y(_0328_));
 sky130_fd_sc_hd__o22a_1 _1045_ (.A1(_0325_),
    .A2(_0326_),
    .B1(_0327_),
    .B2(_0328_),
    .X(_0329_));
 sky130_fd_sc_hd__clkinv_2 _1046_ (.A(_0329_),
    .Y(_0330_));
 sky130_fd_sc_hd__buf_2 _1047_ (.A(_0329_),
    .X(_0331_));
 sky130_fd_sc_hd__a21o_1 _1048_ (.A1(\rgb_mixer0.enc0[0] ),
    .A2(_0331_),
    .B1(net8),
    .X(_0332_));
 sky130_fd_sc_hd__a21oi_1 _1049_ (.A1(_0174_),
    .A2(_0330_),
    .B1(_0332_),
    .Y(_0045_));
 sky130_fd_sc_hd__and4b_1 _1050_ (.A_N(\rgb_mixer0.debounce0_b.debounced ),
    .B(\rgb_mixer0.encoder0.old_b ),
    .C(\rgb_mixer0.encoder0.old_a ),
    .D(\rgb_mixer0.debounce0_a.debounced ),
    .X(_0333_));
 sky130_fd_sc_hd__a21o_1 _1051_ (.A1(_0325_),
    .A2(_0328_),
    .B1(_0333_),
    .X(_0334_));
 sky130_fd_sc_hd__clkbuf_4 _1052_ (.A(_0334_),
    .X(_0335_));
 sky130_fd_sc_hd__nor2_1 _1053_ (.A(\rgb_mixer0.enc0[1] ),
    .B(_0335_),
    .Y(_0336_));
 sky130_fd_sc_hd__o221a_1 _1054_ (.A1(_0325_),
    .A2(_0327_),
    .B1(_0328_),
    .B2(_0326_),
    .C1(\rgb_mixer0.enc0[1] ),
    .X(_0337_));
 sky130_fd_sc_hd__nor2_1 _1055_ (.A(_0336_),
    .B(_0337_),
    .Y(_0338_));
 sky130_fd_sc_hd__or2_1 _1056_ (.A(\rgb_mixer0.enc0[0] ),
    .B(_0338_),
    .X(_0339_));
 sky130_fd_sc_hd__nand2_1 _1057_ (.A(\rgb_mixer0.enc0[0] ),
    .B(_0338_),
    .Y(_0340_));
 sky130_fd_sc_hd__a21o_1 _1058_ (.A1(_0339_),
    .A2(_0340_),
    .B1(_0330_),
    .X(_0341_));
 sky130_fd_sc_hd__o211a_1 _1059_ (.A1(\rgb_mixer0.enc0[1] ),
    .A2(_0331_),
    .B1(_0341_),
    .C1(_0238_),
    .X(_0046_));
 sky130_fd_sc_hd__a211o_1 _1060_ (.A1(_0325_),
    .A2(_0328_),
    .B1(_0333_),
    .C1(\rgb_mixer0.enc0[1] ),
    .X(_0342_));
 sky130_fd_sc_hd__a21o_1 _1061_ (.A1(\rgb_mixer0.enc0[0] ),
    .A2(_0342_),
    .B1(_0337_),
    .X(_0343_));
 sky130_fd_sc_hd__xor2_1 _1062_ (.A(\rgb_mixer0.enc0[2] ),
    .B(_0334_),
    .X(_0344_));
 sky130_fd_sc_hd__or2_1 _1063_ (.A(_0343_),
    .B(_0344_),
    .X(_0345_));
 sky130_fd_sc_hd__nand2_1 _1064_ (.A(_0343_),
    .B(_0344_),
    .Y(_0346_));
 sky130_fd_sc_hd__a21o_1 _1065_ (.A1(_0345_),
    .A2(_0346_),
    .B1(_0330_),
    .X(_0347_));
 sky130_fd_sc_hd__o211a_1 _1066_ (.A1(\rgb_mixer0.enc0[2] ),
    .A2(_0331_),
    .B1(_0347_),
    .C1(_0238_),
    .X(_0047_));
 sky130_fd_sc_hd__nand2_1 _1067_ (.A(\rgb_mixer0.enc0[2] ),
    .B(_0335_),
    .Y(_0348_));
 sky130_fd_sc_hd__xor2_1 _1068_ (.A(\rgb_mixer0.enc0[3] ),
    .B(_0334_),
    .X(_0349_));
 sky130_fd_sc_hd__a21oi_1 _1069_ (.A1(_0348_),
    .A2(_0346_),
    .B1(_0349_),
    .Y(_0350_));
 sky130_fd_sc_hd__a31o_1 _1070_ (.A1(_0348_),
    .A2(_0346_),
    .A3(_0349_),
    .B1(_0330_),
    .X(_0351_));
 sky130_fd_sc_hd__o221a_1 _1071_ (.A1(\rgb_mixer0.enc0[3] ),
    .A2(_0331_),
    .B1(_0350_),
    .B2(_0351_),
    .C1(_0250_),
    .X(_0048_));
 sky130_fd_sc_hd__o21a_1 _1072_ (.A1(\rgb_mixer0.enc0[3] ),
    .A2(\rgb_mixer0.enc0[2] ),
    .B1(_0335_),
    .X(_0352_));
 sky130_fd_sc_hd__a31o_1 _1073_ (.A1(_0343_),
    .A2(_0344_),
    .A3(_0349_),
    .B1(_0352_),
    .X(_0353_));
 sky130_fd_sc_hd__xor2_1 _1074_ (.A(\rgb_mixer0.enc0[4] ),
    .B(_0335_),
    .X(_0354_));
 sky130_fd_sc_hd__or2_1 _1075_ (.A(_0353_),
    .B(_0354_),
    .X(_0355_));
 sky130_fd_sc_hd__nand2_1 _1076_ (.A(_0353_),
    .B(_0354_),
    .Y(_0356_));
 sky130_fd_sc_hd__a21o_1 _1077_ (.A1(_0355_),
    .A2(_0356_),
    .B1(_0330_),
    .X(_0357_));
 sky130_fd_sc_hd__o211a_1 _1078_ (.A1(\rgb_mixer0.enc0[4] ),
    .A2(_0331_),
    .B1(_0357_),
    .C1(_0250_),
    .X(_0049_));
 sky130_fd_sc_hd__xor2_1 _1079_ (.A(\rgb_mixer0.enc0[5] ),
    .B(_0335_),
    .X(_0358_));
 sky130_fd_sc_hd__a21bo_1 _1080_ (.A1(\rgb_mixer0.enc0[4] ),
    .A2(_0335_),
    .B1_N(_0356_),
    .X(_0359_));
 sky130_fd_sc_hd__xnor2_1 _1081_ (.A(_0358_),
    .B(_0359_),
    .Y(_0360_));
 sky130_fd_sc_hd__o21ai_1 _1082_ (.A1(\rgb_mixer0.enc0[5] ),
    .A2(_0331_),
    .B1(_0272_),
    .Y(_0361_));
 sky130_fd_sc_hd__a21oi_1 _1083_ (.A1(_0331_),
    .A2(_0360_),
    .B1(_0361_),
    .Y(_0050_));
 sky130_fd_sc_hd__nor2_1 _1084_ (.A(\rgb_mixer0.enc0[6] ),
    .B(_0335_),
    .Y(_0362_));
 sky130_fd_sc_hd__and2_1 _1085_ (.A(\rgb_mixer0.enc0[6] ),
    .B(_0335_),
    .X(_0363_));
 sky130_fd_sc_hd__nor2_1 _1086_ (.A(_0362_),
    .B(_0363_),
    .Y(_0364_));
 sky130_fd_sc_hd__o21a_1 _1087_ (.A1(\rgb_mixer0.enc0[5] ),
    .A2(\rgb_mixer0.enc0[4] ),
    .B1(_0335_),
    .X(_0365_));
 sky130_fd_sc_hd__a31o_1 _1088_ (.A1(_0353_),
    .A2(_0354_),
    .A3(_0358_),
    .B1(_0365_),
    .X(_0366_));
 sky130_fd_sc_hd__xor2_1 _1089_ (.A(_0364_),
    .B(_0366_),
    .X(_0367_));
 sky130_fd_sc_hd__or2_1 _1090_ (.A(\rgb_mixer0.enc0[6] ),
    .B(_0331_),
    .X(_0368_));
 sky130_fd_sc_hd__o211a_1 _1091_ (.A1(_0330_),
    .A2(_0367_),
    .B1(_0368_),
    .C1(_0250_),
    .X(_0051_));
 sky130_fd_sc_hd__a21o_1 _1092_ (.A1(_0364_),
    .A2(_0366_),
    .B1(_0363_),
    .X(_0369_));
 sky130_fd_sc_hd__xor2_1 _1093_ (.A(\rgb_mixer0.enc0[7] ),
    .B(_0335_),
    .X(_0370_));
 sky130_fd_sc_hd__xnor2_1 _1094_ (.A(_0369_),
    .B(_0370_),
    .Y(_0371_));
 sky130_fd_sc_hd__o21ai_1 _1095_ (.A1(\rgb_mixer0.enc0[7] ),
    .A2(_0331_),
    .B1(_0272_),
    .Y(_0372_));
 sky130_fd_sc_hd__a21oi_1 _1096_ (.A1(_0331_),
    .A2(_0371_),
    .B1(_0372_),
    .Y(_0052_));
 sky130_fd_sc_hd__and2_1 _1097_ (.A(_0272_),
    .B(net5),
    .X(_0373_));
 sky130_fd_sc_hd__clkbuf_1 _1098_ (.A(_0373_),
    .X(_0053_));
 sky130_fd_sc_hd__and2_1 _1099_ (.A(\rgb_mixer0.debounce2_b.button_hist[0] ),
    .B(_0322_),
    .X(_0374_));
 sky130_fd_sc_hd__clkbuf_1 _1100_ (.A(_0374_),
    .X(_0054_));
 sky130_fd_sc_hd__and2_1 _1101_ (.A(\rgb_mixer0.debounce2_b.button_hist[1] ),
    .B(_0322_),
    .X(_0375_));
 sky130_fd_sc_hd__clkbuf_1 _1102_ (.A(_0375_),
    .X(_0055_));
 sky130_fd_sc_hd__and2_1 _1103_ (.A(\rgb_mixer0.debounce2_b.button_hist[2] ),
    .B(_0322_),
    .X(_0376_));
 sky130_fd_sc_hd__clkbuf_1 _1104_ (.A(_0376_),
    .X(_0056_));
 sky130_fd_sc_hd__and2_1 _1105_ (.A(\rgb_mixer0.debounce2_b.button_hist[3] ),
    .B(_0322_),
    .X(_0377_));
 sky130_fd_sc_hd__clkbuf_1 _1106_ (.A(_0377_),
    .X(_0057_));
 sky130_fd_sc_hd__and2_1 _1107_ (.A(\rgb_mixer0.debounce2_b.button_hist[4] ),
    .B(_0322_),
    .X(_0378_));
 sky130_fd_sc_hd__clkbuf_1 _1108_ (.A(_0378_),
    .X(_0058_));
 sky130_fd_sc_hd__and2_1 _1109_ (.A(\rgb_mixer0.debounce2_b.button_hist[5] ),
    .B(_0322_),
    .X(_0379_));
 sky130_fd_sc_hd__clkbuf_1 _1110_ (.A(_0379_),
    .X(_0059_));
 sky130_fd_sc_hd__and2_1 _1111_ (.A(\rgb_mixer0.debounce2_b.button_hist[6] ),
    .B(_0322_),
    .X(_0380_));
 sky130_fd_sc_hd__clkbuf_1 _1112_ (.A(_0380_),
    .X(_0060_));
 sky130_fd_sc_hd__and2_1 _1113_ (.A(\rgb_mixer0.debounce0_a.debounced ),
    .B(_0120_),
    .X(_0381_));
 sky130_fd_sc_hd__clkbuf_1 _1114_ (.A(_0381_),
    .X(_0061_));
 sky130_fd_sc_hd__and4_1 _1115_ (.A(\rgb_mixer0.debounce2_b.button_hist[4] ),
    .B(\rgb_mixer0.debounce2_b.button_hist[5] ),
    .C(\rgb_mixer0.debounce2_b.button_hist[7] ),
    .D(\rgb_mixer0.debounce2_b.button_hist[6] ),
    .X(_0382_));
 sky130_fd_sc_hd__and4_1 _1116_ (.A(\rgb_mixer0.debounce2_b.button_hist[0] ),
    .B(\rgb_mixer0.debounce2_b.button_hist[1] ),
    .C(\rgb_mixer0.debounce2_b.button_hist[2] ),
    .D(\rgb_mixer0.debounce2_b.button_hist[3] ),
    .X(_0383_));
 sky130_fd_sc_hd__or4_1 _1117_ (.A(\rgb_mixer0.debounce2_b.button_hist[0] ),
    .B(\rgb_mixer0.debounce2_b.button_hist[1] ),
    .C(\rgb_mixer0.debounce2_b.button_hist[2] ),
    .D(\rgb_mixer0.debounce2_b.button_hist[3] ),
    .X(_0384_));
 sky130_fd_sc_hd__or4_1 _1118_ (.A(\rgb_mixer0.debounce2_b.button_hist[4] ),
    .B(\rgb_mixer0.debounce2_b.button_hist[5] ),
    .C(\rgb_mixer0.debounce2_b.button_hist[7] ),
    .D(\rgb_mixer0.debounce2_b.button_hist[6] ),
    .X(_0385_));
 sky130_fd_sc_hd__or2_1 _1119_ (.A(_0384_),
    .B(_0385_),
    .X(_0386_));
 sky130_fd_sc_hd__a32o_1 _1120_ (.A1(_0250_),
    .A2(_0382_),
    .A3(_0383_),
    .B1(_0386_),
    .B2(_0024_),
    .X(_0062_));
 sky130_fd_sc_hd__and2_1 _1121_ (.A(_0272_),
    .B(net4),
    .X(_0387_));
 sky130_fd_sc_hd__clkbuf_1 _1122_ (.A(_0387_),
    .X(_0063_));
 sky130_fd_sc_hd__and2_1 _1123_ (.A(\rgb_mixer0.debounce2_a.button_hist[0] ),
    .B(_0120_),
    .X(_0388_));
 sky130_fd_sc_hd__clkbuf_1 _1124_ (.A(_0388_),
    .X(_0064_));
 sky130_fd_sc_hd__and2_1 _1125_ (.A(\rgb_mixer0.debounce2_a.button_hist[1] ),
    .B(_0322_),
    .X(_0389_));
 sky130_fd_sc_hd__clkbuf_1 _1126_ (.A(_0389_),
    .X(_0065_));
 sky130_fd_sc_hd__and2_1 _1127_ (.A(\rgb_mixer0.debounce2_a.button_hist[2] ),
    .B(_0322_),
    .X(_0390_));
 sky130_fd_sc_hd__clkbuf_1 _1128_ (.A(_0390_),
    .X(_0066_));
 sky130_fd_sc_hd__clkbuf_2 _1129_ (.A(_0121_),
    .X(_0391_));
 sky130_fd_sc_hd__and2_1 _1130_ (.A(\rgb_mixer0.debounce2_a.button_hist[3] ),
    .B(_0391_),
    .X(_0392_));
 sky130_fd_sc_hd__clkbuf_1 _1131_ (.A(_0392_),
    .X(_0067_));
 sky130_fd_sc_hd__and2_1 _1132_ (.A(\rgb_mixer0.debounce2_a.button_hist[4] ),
    .B(_0391_),
    .X(_0393_));
 sky130_fd_sc_hd__clkbuf_1 _1133_ (.A(_0393_),
    .X(_0068_));
 sky130_fd_sc_hd__and2_1 _1134_ (.A(\rgb_mixer0.debounce2_a.button_hist[5] ),
    .B(_0391_),
    .X(_0394_));
 sky130_fd_sc_hd__clkbuf_1 _1135_ (.A(_0394_),
    .X(_0069_));
 sky130_fd_sc_hd__and2_1 _1136_ (.A(\rgb_mixer0.debounce2_a.button_hist[6] ),
    .B(_0391_),
    .X(_0395_));
 sky130_fd_sc_hd__clkbuf_1 _1137_ (.A(_0395_),
    .X(_0070_));
 sky130_fd_sc_hd__and4_1 _1138_ (.A(\rgb_mixer0.debounce2_a.button_hist[5] ),
    .B(\rgb_mixer0.debounce2_a.button_hist[4] ),
    .C(\rgb_mixer0.debounce2_a.button_hist[7] ),
    .D(\rgb_mixer0.debounce2_a.button_hist[6] ),
    .X(_0396_));
 sky130_fd_sc_hd__and3_1 _1139_ (.A(\rgb_mixer0.debounce2_a.button_hist[1] ),
    .B(\rgb_mixer0.debounce2_a.button_hist[2] ),
    .C(_0396_),
    .X(_0397_));
 sky130_fd_sc_hd__or3_1 _1140_ (.A(\rgb_mixer0.debounce2_a.button_hist[1] ),
    .B(\rgb_mixer0.debounce2_a.button_hist[0] ),
    .C(\rgb_mixer0.debounce2_a.button_hist[3] ),
    .X(_0398_));
 sky130_fd_sc_hd__or4_1 _1141_ (.A(\rgb_mixer0.debounce2_a.button_hist[5] ),
    .B(\rgb_mixer0.debounce2_a.button_hist[4] ),
    .C(\rgb_mixer0.debounce2_a.button_hist[7] ),
    .D(\rgb_mixer0.debounce2_a.button_hist[6] ),
    .X(_0399_));
 sky130_fd_sc_hd__o31a_1 _1142_ (.A1(\rgb_mixer0.debounce2_a.button_hist[2] ),
    .A2(_0398_),
    .A3(_0399_),
    .B1(\rgb_mixer0.debounce2_a.debounced ),
    .X(_0400_));
 sky130_fd_sc_hd__a32o_1 _1143_ (.A1(\rgb_mixer0.debounce2_a.button_hist[3] ),
    .A2(_0064_),
    .A3(_0397_),
    .B1(_0400_),
    .B2(_0250_),
    .X(_0071_));
 sky130_fd_sc_hd__and2_1 _1144_ (.A(_0272_),
    .B(net3),
    .X(_0401_));
 sky130_fd_sc_hd__clkbuf_1 _1145_ (.A(_0401_),
    .X(_0072_));
 sky130_fd_sc_hd__and2_1 _1146_ (.A(\rgb_mixer0.debounce1_b.button_hist[0] ),
    .B(_0120_),
    .X(_0402_));
 sky130_fd_sc_hd__clkbuf_1 _1147_ (.A(_0402_),
    .X(_0073_));
 sky130_fd_sc_hd__and2_1 _1148_ (.A(\rgb_mixer0.debounce1_b.button_hist[1] ),
    .B(_0391_),
    .X(_0403_));
 sky130_fd_sc_hd__clkbuf_1 _1149_ (.A(_0403_),
    .X(_0074_));
 sky130_fd_sc_hd__and2_1 _1150_ (.A(\rgb_mixer0.debounce1_b.button_hist[2] ),
    .B(_0391_),
    .X(_0404_));
 sky130_fd_sc_hd__clkbuf_1 _1151_ (.A(_0404_),
    .X(_0075_));
 sky130_fd_sc_hd__and2_1 _1152_ (.A(\rgb_mixer0.debounce1_b.button_hist[3] ),
    .B(_0391_),
    .X(_0405_));
 sky130_fd_sc_hd__clkbuf_1 _1153_ (.A(_0405_),
    .X(_0076_));
 sky130_fd_sc_hd__and2_1 _1154_ (.A(\rgb_mixer0.debounce1_b.button_hist[4] ),
    .B(_0391_),
    .X(_0406_));
 sky130_fd_sc_hd__clkbuf_1 _1155_ (.A(_0406_),
    .X(_0077_));
 sky130_fd_sc_hd__and2_1 _1156_ (.A(\rgb_mixer0.debounce1_b.button_hist[5] ),
    .B(_0391_),
    .X(_0407_));
 sky130_fd_sc_hd__clkbuf_1 _1157_ (.A(_0407_),
    .X(_0078_));
 sky130_fd_sc_hd__and2_1 _1158_ (.A(\rgb_mixer0.debounce1_b.button_hist[6] ),
    .B(_0391_),
    .X(_0408_));
 sky130_fd_sc_hd__clkbuf_1 _1159_ (.A(_0408_),
    .X(_0079_));
 sky130_fd_sc_hd__and4_1 _1160_ (.A(\rgb_mixer0.debounce1_b.button_hist[5] ),
    .B(\rgb_mixer0.debounce1_b.button_hist[4] ),
    .C(\rgb_mixer0.debounce1_b.button_hist[7] ),
    .D(\rgb_mixer0.debounce1_b.button_hist[6] ),
    .X(_0409_));
 sky130_fd_sc_hd__and3_1 _1161_ (.A(\rgb_mixer0.debounce1_b.button_hist[1] ),
    .B(\rgb_mixer0.debounce1_b.button_hist[2] ),
    .C(_0409_),
    .X(_0410_));
 sky130_fd_sc_hd__or3_1 _1162_ (.A(\rgb_mixer0.debounce1_b.button_hist[1] ),
    .B(\rgb_mixer0.debounce1_b.button_hist[0] ),
    .C(\rgb_mixer0.debounce1_b.button_hist[3] ),
    .X(_0411_));
 sky130_fd_sc_hd__or4_1 _1163_ (.A(\rgb_mixer0.debounce1_b.button_hist[5] ),
    .B(\rgb_mixer0.debounce1_b.button_hist[4] ),
    .C(\rgb_mixer0.debounce1_b.button_hist[7] ),
    .D(\rgb_mixer0.debounce1_b.button_hist[6] ),
    .X(_0412_));
 sky130_fd_sc_hd__o31a_1 _1164_ (.A1(\rgb_mixer0.debounce1_b.button_hist[2] ),
    .A2(_0411_),
    .A3(_0412_),
    .B1(\rgb_mixer0.debounce1_b.debounced ),
    .X(_0413_));
 sky130_fd_sc_hd__a32o_1 _1165_ (.A1(\rgb_mixer0.debounce1_b.button_hist[3] ),
    .A2(_0073_),
    .A3(_0410_),
    .B1(_0413_),
    .B2(_0250_),
    .X(_0080_));
 sky130_fd_sc_hd__and2_1 _1166_ (.A(_0272_),
    .B(net2),
    .X(_0414_));
 sky130_fd_sc_hd__clkbuf_1 _1167_ (.A(_0414_),
    .X(_0081_));
 sky130_fd_sc_hd__clkbuf_2 _1168_ (.A(_0121_),
    .X(_0415_));
 sky130_fd_sc_hd__and2_1 _1169_ (.A(\rgb_mixer0.debounce1_a.button_hist[0] ),
    .B(_0415_),
    .X(_0416_));
 sky130_fd_sc_hd__clkbuf_1 _1170_ (.A(_0416_),
    .X(_0082_));
 sky130_fd_sc_hd__and2_1 _1171_ (.A(\rgb_mixer0.debounce1_a.button_hist[1] ),
    .B(_0415_),
    .X(_0417_));
 sky130_fd_sc_hd__clkbuf_1 _1172_ (.A(_0417_),
    .X(_0083_));
 sky130_fd_sc_hd__and2_1 _1173_ (.A(\rgb_mixer0.debounce1_a.button_hist[2] ),
    .B(_0415_),
    .X(_0418_));
 sky130_fd_sc_hd__clkbuf_1 _1174_ (.A(_0418_),
    .X(_0084_));
 sky130_fd_sc_hd__and2_1 _1175_ (.A(\rgb_mixer0.debounce1_a.button_hist[3] ),
    .B(_0415_),
    .X(_0419_));
 sky130_fd_sc_hd__clkbuf_1 _1176_ (.A(_0419_),
    .X(_0085_));
 sky130_fd_sc_hd__and2_1 _1177_ (.A(\rgb_mixer0.debounce1_a.button_hist[4] ),
    .B(_0415_),
    .X(_0420_));
 sky130_fd_sc_hd__clkbuf_1 _1178_ (.A(_0420_),
    .X(_0086_));
 sky130_fd_sc_hd__and2_1 _1179_ (.A(\rgb_mixer0.debounce1_a.button_hist[5] ),
    .B(_0415_),
    .X(_0421_));
 sky130_fd_sc_hd__clkbuf_1 _1180_ (.A(_0421_),
    .X(_0087_));
 sky130_fd_sc_hd__and2_1 _1181_ (.A(\rgb_mixer0.debounce1_a.button_hist[6] ),
    .B(_0415_),
    .X(_0422_));
 sky130_fd_sc_hd__clkbuf_1 _1182_ (.A(_0422_),
    .X(_0088_));
 sky130_fd_sc_hd__and4_1 _1183_ (.A(\rgb_mixer0.debounce1_a.button_hist[5] ),
    .B(\rgb_mixer0.debounce1_a.button_hist[4] ),
    .C(\rgb_mixer0.debounce1_a.button_hist[7] ),
    .D(\rgb_mixer0.debounce1_a.button_hist[6] ),
    .X(_0423_));
 sky130_fd_sc_hd__and4_1 _1184_ (.A(\rgb_mixer0.debounce1_a.button_hist[1] ),
    .B(\rgb_mixer0.debounce1_a.button_hist[0] ),
    .C(\rgb_mixer0.debounce1_a.button_hist[3] ),
    .D(\rgb_mixer0.debounce1_a.button_hist[2] ),
    .X(_0424_));
 sky130_fd_sc_hd__or4_1 _1185_ (.A(\rgb_mixer0.debounce1_a.button_hist[5] ),
    .B(\rgb_mixer0.debounce1_a.button_hist[4] ),
    .C(\rgb_mixer0.debounce1_a.button_hist[7] ),
    .D(\rgb_mixer0.debounce1_a.button_hist[6] ),
    .X(_0425_));
 sky130_fd_sc_hd__or3_1 _1186_ (.A(\rgb_mixer0.debounce1_a.button_hist[3] ),
    .B(\rgb_mixer0.debounce1_a.button_hist[2] ),
    .C(_0425_),
    .X(_0426_));
 sky130_fd_sc_hd__o31a_1 _1187_ (.A1(\rgb_mixer0.debounce1_a.button_hist[1] ),
    .A2(\rgb_mixer0.debounce1_a.button_hist[0] ),
    .A3(_0426_),
    .B1(_0044_),
    .X(_0427_));
 sky130_fd_sc_hd__a31o_1 _1188_ (.A1(_0250_),
    .A2(_0423_),
    .A3(_0424_),
    .B1(_0427_),
    .X(_0089_));
 sky130_fd_sc_hd__and2_1 _1189_ (.A(_0272_),
    .B(net7),
    .X(_0428_));
 sky130_fd_sc_hd__clkbuf_1 _1190_ (.A(_0428_),
    .X(_0090_));
 sky130_fd_sc_hd__and2_1 _1191_ (.A(\rgb_mixer0.debounce0_b.button_hist[0] ),
    .B(_0120_),
    .X(_0429_));
 sky130_fd_sc_hd__clkbuf_1 _1192_ (.A(_0429_),
    .X(_0091_));
 sky130_fd_sc_hd__and2_1 _1193_ (.A(\rgb_mixer0.debounce0_b.button_hist[1] ),
    .B(_0415_),
    .X(_0430_));
 sky130_fd_sc_hd__clkbuf_1 _1194_ (.A(_0430_),
    .X(_0092_));
 sky130_fd_sc_hd__and2_1 _1195_ (.A(\rgb_mixer0.debounce0_b.button_hist[2] ),
    .B(_0415_),
    .X(_0431_));
 sky130_fd_sc_hd__clkbuf_1 _1196_ (.A(_0431_),
    .X(_0093_));
 sky130_fd_sc_hd__and2_1 _1197_ (.A(\rgb_mixer0.debounce0_b.button_hist[3] ),
    .B(_0415_),
    .X(_0432_));
 sky130_fd_sc_hd__clkbuf_1 _1198_ (.A(_0432_),
    .X(_0094_));
 sky130_fd_sc_hd__clkbuf_2 _1199_ (.A(_0121_),
    .X(_0433_));
 sky130_fd_sc_hd__and2_1 _1200_ (.A(\rgb_mixer0.debounce0_b.button_hist[4] ),
    .B(_0433_),
    .X(_0434_));
 sky130_fd_sc_hd__clkbuf_1 _1201_ (.A(_0434_),
    .X(_0095_));
 sky130_fd_sc_hd__and2_1 _1202_ (.A(\rgb_mixer0.debounce0_b.button_hist[5] ),
    .B(_0433_),
    .X(_0435_));
 sky130_fd_sc_hd__clkbuf_1 _1203_ (.A(_0435_),
    .X(_0096_));
 sky130_fd_sc_hd__and2_1 _1204_ (.A(\rgb_mixer0.debounce0_b.button_hist[6] ),
    .B(_0433_),
    .X(_0436_));
 sky130_fd_sc_hd__clkbuf_1 _1205_ (.A(_0436_),
    .X(_0097_));
 sky130_fd_sc_hd__and4_1 _1206_ (.A(\rgb_mixer0.debounce0_b.button_hist[5] ),
    .B(\rgb_mixer0.debounce0_b.button_hist[4] ),
    .C(\rgb_mixer0.debounce0_b.button_hist[7] ),
    .D(\rgb_mixer0.debounce0_b.button_hist[6] ),
    .X(_0437_));
 sky130_fd_sc_hd__and3_1 _1207_ (.A(\rgb_mixer0.debounce0_b.button_hist[1] ),
    .B(\rgb_mixer0.debounce0_b.button_hist[2] ),
    .C(_0437_),
    .X(_0438_));
 sky130_fd_sc_hd__or3_1 _1208_ (.A(\rgb_mixer0.debounce0_b.button_hist[1] ),
    .B(\rgb_mixer0.debounce0_b.button_hist[0] ),
    .C(\rgb_mixer0.debounce0_b.button_hist[3] ),
    .X(_0439_));
 sky130_fd_sc_hd__or4_1 _1209_ (.A(\rgb_mixer0.debounce0_b.button_hist[5] ),
    .B(\rgb_mixer0.debounce0_b.button_hist[4] ),
    .C(\rgb_mixer0.debounce0_b.button_hist[7] ),
    .D(\rgb_mixer0.debounce0_b.button_hist[6] ),
    .X(_0440_));
 sky130_fd_sc_hd__o31a_1 _1210_ (.A1(\rgb_mixer0.debounce0_b.button_hist[2] ),
    .A2(_0439_),
    .A3(_0440_),
    .B1(\rgb_mixer0.debounce0_b.debounced ),
    .X(_0441_));
 sky130_fd_sc_hd__a32o_1 _1211_ (.A1(\rgb_mixer0.debounce0_b.button_hist[3] ),
    .A2(_0091_),
    .A3(_0438_),
    .B1(_0441_),
    .B2(_0250_),
    .X(_0098_));
 sky130_fd_sc_hd__and2_1 _1212_ (.A(_0272_),
    .B(net6),
    .X(_0442_));
 sky130_fd_sc_hd__clkbuf_1 _1213_ (.A(_0442_),
    .X(_0099_));
 sky130_fd_sc_hd__and2_1 _1214_ (.A(\rgb_mixer0.debounce0_a.button_hist[0] ),
    .B(_0433_),
    .X(_0443_));
 sky130_fd_sc_hd__clkbuf_1 _1215_ (.A(_0443_),
    .X(_0100_));
 sky130_fd_sc_hd__and2_1 _1216_ (.A(\rgb_mixer0.debounce0_a.button_hist[1] ),
    .B(_0433_),
    .X(_0444_));
 sky130_fd_sc_hd__clkbuf_1 _1217_ (.A(_0444_),
    .X(_0101_));
 sky130_fd_sc_hd__and2_1 _1218_ (.A(\rgb_mixer0.debounce0_a.button_hist[2] ),
    .B(_0433_),
    .X(_0445_));
 sky130_fd_sc_hd__clkbuf_1 _1219_ (.A(_0445_),
    .X(_0102_));
 sky130_fd_sc_hd__and2_1 _1220_ (.A(\rgb_mixer0.debounce0_a.button_hist[3] ),
    .B(_0433_),
    .X(_0446_));
 sky130_fd_sc_hd__clkbuf_1 _1221_ (.A(_0446_),
    .X(_0103_));
 sky130_fd_sc_hd__and2_1 _1222_ (.A(\rgb_mixer0.debounce0_a.button_hist[4] ),
    .B(_0433_),
    .X(_0447_));
 sky130_fd_sc_hd__clkbuf_1 _1223_ (.A(_0447_),
    .X(_0104_));
 sky130_fd_sc_hd__and2_1 _1224_ (.A(\rgb_mixer0.debounce0_a.button_hist[5] ),
    .B(_0433_),
    .X(_0448_));
 sky130_fd_sc_hd__clkbuf_1 _1225_ (.A(_0448_),
    .X(_0105_));
 sky130_fd_sc_hd__and2_1 _1226_ (.A(\rgb_mixer0.debounce0_a.button_hist[6] ),
    .B(_0433_),
    .X(_0449_));
 sky130_fd_sc_hd__clkbuf_1 _1227_ (.A(_0449_),
    .X(_0106_));
 sky130_fd_sc_hd__and4_1 _1228_ (.A(\rgb_mixer0.debounce0_a.button_hist[5] ),
    .B(\rgb_mixer0.debounce0_a.button_hist[4] ),
    .C(\rgb_mixer0.debounce0_a.button_hist[7] ),
    .D(\rgb_mixer0.debounce0_a.button_hist[6] ),
    .X(_0450_));
 sky130_fd_sc_hd__and4_1 _1229_ (.A(\rgb_mixer0.debounce0_a.button_hist[1] ),
    .B(\rgb_mixer0.debounce0_a.button_hist[0] ),
    .C(\rgb_mixer0.debounce0_a.button_hist[3] ),
    .D(\rgb_mixer0.debounce0_a.button_hist[2] ),
    .X(_0451_));
 sky130_fd_sc_hd__or4_1 _1230_ (.A(\rgb_mixer0.debounce0_a.button_hist[1] ),
    .B(\rgb_mixer0.debounce0_a.button_hist[0] ),
    .C(\rgb_mixer0.debounce0_a.button_hist[3] ),
    .D(\rgb_mixer0.debounce0_a.button_hist[2] ),
    .X(_0452_));
 sky130_fd_sc_hd__or4_1 _1231_ (.A(\rgb_mixer0.debounce0_a.button_hist[5] ),
    .B(\rgb_mixer0.debounce0_a.button_hist[4] ),
    .C(\rgb_mixer0.debounce0_a.button_hist[7] ),
    .D(\rgb_mixer0.debounce0_a.button_hist[6] ),
    .X(_0453_));
 sky130_fd_sc_hd__or2_1 _1232_ (.A(_0452_),
    .B(_0453_),
    .X(_0454_));
 sky130_fd_sc_hd__a32o_1 _1233_ (.A1(_0191_),
    .A2(_0450_),
    .A3(_0451_),
    .B1(_0454_),
    .B2(_0061_),
    .X(_0107_));
 sky130_fd_sc_hd__dfxtp_1 _1234_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0000_),
    .Q(\rgb_mixer0.pwm2.count[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1235_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0001_),
    .Q(\rgb_mixer0.pwm2.count[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1236_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0002_),
    .Q(\rgb_mixer0.pwm2.count[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1237_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0003_),
    .Q(\rgb_mixer0.pwm2.count[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1238_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0004_),
    .Q(\rgb_mixer0.pwm2.count[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1239_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0005_),
    .Q(\rgb_mixer0.pwm2.count[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1240_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0006_),
    .Q(\rgb_mixer0.pwm2.count[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1241_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0007_),
    .Q(\rgb_mixer0.pwm2.count[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1242_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0008_),
    .Q(\rgb_mixer0.pwm1.count[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1243_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0009_),
    .Q(\rgb_mixer0.pwm1.count[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1244_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0010_),
    .Q(\rgb_mixer0.pwm1.count[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1245_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0011_),
    .Q(\rgb_mixer0.pwm1.count[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1246_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0012_),
    .Q(\rgb_mixer0.pwm1.count[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1247_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0013_),
    .Q(\rgb_mixer0.pwm1.count[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1248_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0014_),
    .Q(\rgb_mixer0.pwm1.count[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1249_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0015_),
    .Q(\rgb_mixer0.pwm1.count[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1250_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0016_),
    .Q(\rgb_mixer0.pwm0.count[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1251_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0017_),
    .Q(\rgb_mixer0.pwm0.count[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1252_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0018_),
    .Q(\rgb_mixer0.pwm0.count[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1253_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0019_),
    .Q(\rgb_mixer0.pwm0.count[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1254_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0020_),
    .Q(\rgb_mixer0.pwm0.count[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1255_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0021_),
    .Q(\rgb_mixer0.pwm0.count[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1256_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0022_),
    .Q(\rgb_mixer0.pwm0.count[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1257_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0023_),
    .Q(\rgb_mixer0.pwm0.count[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1258_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0024_),
    .Q(\rgb_mixer0.encoder2.old_b ));
 sky130_fd_sc_hd__dfxtp_1 _1259_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0025_),
    .Q(\rgb_mixer0.enc2[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1260_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0026_),
    .Q(\rgb_mixer0.enc2[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1261_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0027_),
    .Q(\rgb_mixer0.enc2[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1262_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0028_),
    .Q(\rgb_mixer0.enc2[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1263_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0029_),
    .Q(\rgb_mixer0.enc2[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1264_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0030_),
    .Q(\rgb_mixer0.enc2[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1265_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0031_),
    .Q(\rgb_mixer0.enc2[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1266_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0032_),
    .Q(\rgb_mixer0.enc2[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1267_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_0033_),
    .Q(\rgb_mixer0.encoder1.old_b ));
 sky130_fd_sc_hd__dfxtp_1 _1268_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_0034_),
    .Q(\rgb_mixer0.encoder2.old_a ));
 sky130_fd_sc_hd__dfxtp_1 _1269_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0035_),
    .Q(\rgb_mixer0.enc1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1270_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0036_),
    .Q(\rgb_mixer0.enc1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1271_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0037_),
    .Q(\rgb_mixer0.enc1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1272_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0038_),
    .Q(\rgb_mixer0.enc1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1273_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0039_),
    .Q(\rgb_mixer0.enc1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1274_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0040_),
    .Q(\rgb_mixer0.enc1[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1275_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0041_),
    .Q(\rgb_mixer0.enc1[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1276_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0042_),
    .Q(\rgb_mixer0.enc1[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1277_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_0043_),
    .Q(\rgb_mixer0.encoder0.old_b ));
 sky130_fd_sc_hd__dfxtp_1 _1278_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_0044_),
    .Q(\rgb_mixer0.encoder1.old_a ));
 sky130_fd_sc_hd__dfxtp_1 _1279_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0045_),
    .Q(\rgb_mixer0.enc0[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1280_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_0046_),
    .Q(\rgb_mixer0.enc0[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1281_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0047_),
    .Q(\rgb_mixer0.enc0[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1282_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_0048_),
    .Q(\rgb_mixer0.enc0[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1283_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0049_),
    .Q(\rgb_mixer0.enc0[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1284_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_0050_),
    .Q(\rgb_mixer0.enc0[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1285_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_0051_),
    .Q(\rgb_mixer0.enc0[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1286_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_0052_),
    .Q(\rgb_mixer0.enc0[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1287_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_0053_),
    .Q(\rgb_mixer0.debounce2_b.button_hist[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1288_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_0054_),
    .Q(\rgb_mixer0.debounce2_b.button_hist[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1289_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_0055_),
    .Q(\rgb_mixer0.debounce2_b.button_hist[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1290_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_0056_),
    .Q(\rgb_mixer0.debounce2_b.button_hist[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1291_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_0057_),
    .Q(\rgb_mixer0.debounce2_b.button_hist[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1292_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0058_),
    .Q(\rgb_mixer0.debounce2_b.button_hist[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1293_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0059_),
    .Q(\rgb_mixer0.debounce2_b.button_hist[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1294_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0060_),
    .Q(\rgb_mixer0.debounce2_b.button_hist[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1295_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_0061_),
    .Q(\rgb_mixer0.encoder0.old_a ));
 sky130_fd_sc_hd__dfxtp_1 _1296_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_0062_),
    .Q(\rgb_mixer0.debounce2_b.debounced ));
 sky130_fd_sc_hd__dfxtp_1 _1297_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_0063_),
    .Q(\rgb_mixer0.debounce2_a.button_hist[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1298_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0064_),
    .Q(\rgb_mixer0.debounce2_a.button_hist[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1299_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0065_),
    .Q(\rgb_mixer0.debounce2_a.button_hist[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1300_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_0066_),
    .Q(\rgb_mixer0.debounce2_a.button_hist[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1301_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_0067_),
    .Q(\rgb_mixer0.debounce2_a.button_hist[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1302_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_0068_),
    .Q(\rgb_mixer0.debounce2_a.button_hist[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1303_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0069_),
    .Q(\rgb_mixer0.debounce2_a.button_hist[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1304_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0070_),
    .Q(\rgb_mixer0.debounce2_a.button_hist[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1305_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_0071_),
    .Q(\rgb_mixer0.debounce2_a.debounced ));
 sky130_fd_sc_hd__dfxtp_1 _1306_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0072_),
    .Q(\rgb_mixer0.debounce1_b.button_hist[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1307_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0073_),
    .Q(\rgb_mixer0.debounce1_b.button_hist[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1308_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0074_),
    .Q(\rgb_mixer0.debounce1_b.button_hist[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1309_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0075_),
    .Q(\rgb_mixer0.debounce1_b.button_hist[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1310_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_0076_),
    .Q(\rgb_mixer0.debounce1_b.button_hist[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1311_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_0077_),
    .Q(\rgb_mixer0.debounce1_b.button_hist[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1312_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0078_),
    .Q(\rgb_mixer0.debounce1_b.button_hist[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1313_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0079_),
    .Q(\rgb_mixer0.debounce1_b.button_hist[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1314_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_0080_),
    .Q(\rgb_mixer0.debounce1_b.debounced ));
 sky130_fd_sc_hd__dfxtp_1 _1315_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0081_),
    .Q(\rgb_mixer0.debounce1_a.button_hist[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1316_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0082_),
    .Q(\rgb_mixer0.debounce1_a.button_hist[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1317_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0083_),
    .Q(\rgb_mixer0.debounce1_a.button_hist[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1318_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0084_),
    .Q(\rgb_mixer0.debounce1_a.button_hist[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1319_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0085_),
    .Q(\rgb_mixer0.debounce1_a.button_hist[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1320_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0086_),
    .Q(\rgb_mixer0.debounce1_a.button_hist[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1321_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0087_),
    .Q(\rgb_mixer0.debounce1_a.button_hist[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1322_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0088_),
    .Q(\rgb_mixer0.debounce1_a.button_hist[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1323_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0089_),
    .Q(\rgb_mixer0.debounce1_a.debounced ));
 sky130_fd_sc_hd__dfxtp_1 _1324_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0090_),
    .Q(\rgb_mixer0.debounce0_b.button_hist[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1325_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0091_),
    .Q(\rgb_mixer0.debounce0_b.button_hist[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1326_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_0092_),
    .Q(\rgb_mixer0.debounce0_b.button_hist[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1327_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0093_),
    .Q(\rgb_mixer0.debounce0_b.button_hist[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1328_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_0094_),
    .Q(\rgb_mixer0.debounce0_b.button_hist[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1329_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_0095_),
    .Q(\rgb_mixer0.debounce0_b.button_hist[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1330_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_0096_),
    .Q(\rgb_mixer0.debounce0_b.button_hist[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1331_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_0097_),
    .Q(\rgb_mixer0.debounce0_b.button_hist[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1332_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_0098_),
    .Q(\rgb_mixer0.debounce0_b.debounced ));
 sky130_fd_sc_hd__dfxtp_1 _1333_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_0099_),
    .Q(\rgb_mixer0.debounce0_a.button_hist[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1334_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_0100_),
    .Q(\rgb_mixer0.debounce0_a.button_hist[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1335_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_0101_),
    .Q(\rgb_mixer0.debounce0_a.button_hist[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1336_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_0102_),
    .Q(\rgb_mixer0.debounce0_a.button_hist[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1337_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_0103_),
    .Q(\rgb_mixer0.debounce0_a.button_hist[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1338_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_0104_),
    .Q(\rgb_mixer0.debounce0_a.button_hist[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1339_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_0105_),
    .Q(\rgb_mixer0.debounce0_a.button_hist[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1340_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_0106_),
    .Q(\rgb_mixer0.debounce0_a.button_hist[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1341_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_0107_),
    .Q(\rgb_mixer0.debounce0_a.debounced ));
 sky130_fd_sc_hd__conb_1 _1448__10 (.LO(net10));
 sky130_fd_sc_hd__conb_1 _1449__11 (.LO(net11));
 sky130_fd_sc_hd__conb_1 _1450__12 (.LO(net12));
 sky130_fd_sc_hd__conb_1 _1451__13 (.LO(net13));
 sky130_fd_sc_hd__conb_1 _1452__14 (.LO(net14));
 sky130_fd_sc_hd__conb_1 _1453__15 (.LO(net15));
 sky130_fd_sc_hd__conb_1 _1454__16 (.LO(net16));
 sky130_fd_sc_hd__conb_1 _1455__17 (.LO(net17));
 sky130_fd_sc_hd__conb_1 _1456__18 (.LO(net18));
 sky130_fd_sc_hd__conb_1 _1457__19 (.LO(net19));
 sky130_fd_sc_hd__conb_1 _1458__20 (.LO(net20));
 sky130_fd_sc_hd__conb_1 _1459__21 (.LO(net21));
 sky130_fd_sc_hd__conb_1 _1460__22 (.LO(net22));
 sky130_fd_sc_hd__conb_1 _1461__23 (.LO(net23));
 sky130_fd_sc_hd__conb_1 _1462__24 (.LO(net24));
 sky130_fd_sc_hd__conb_1 _1463__25 (.LO(net25));
 sky130_fd_sc_hd__conb_1 _1464__26 (.LO(net26));
 sky130_fd_sc_hd__conb_1 _1465__27 (.LO(net27));
 sky130_fd_sc_hd__conb_1 _1466__28 (.LO(net28));
 sky130_fd_sc_hd__conb_1 _1467__29 (.LO(net29));
 sky130_fd_sc_hd__conb_1 _1468__30 (.LO(net30));
 sky130_fd_sc_hd__conb_1 _1469__31 (.LO(net31));
 sky130_fd_sc_hd__conb_1 _1470__32 (.LO(net32));
 sky130_fd_sc_hd__conb_1 _1471__33 (.LO(net33));
 sky130_fd_sc_hd__conb_1 _1472__34 (.LO(net34));
 sky130_fd_sc_hd__conb_1 _1473__35 (.LO(net35));
 sky130_fd_sc_hd__conb_1 _1474__36 (.LO(net36));
 sky130_fd_sc_hd__conb_1 _1475__37 (.LO(net37));
 sky130_fd_sc_hd__conb_1 _1476__38 (.LO(net38));
 sky130_fd_sc_hd__conb_1 _1477__39 (.LO(net39));
 sky130_fd_sc_hd__conb_1 _1478__40 (.LO(net40));
 sky130_fd_sc_hd__conb_1 _1479__41 (.LO(net41));
 sky130_fd_sc_hd__conb_1 _1480__42 (.LO(net42));
 sky130_fd_sc_hd__conb_1 _1481__43 (.LO(net43));
 sky130_fd_sc_hd__conb_1 _1482__44 (.LO(net44));
 sky130_fd_sc_hd__conb_1 _1483__45 (.LO(net45));
 sky130_fd_sc_hd__conb_1 _1484__46 (.LO(net46));
 sky130_fd_sc_hd__conb_1 _1485__47 (.LO(net47));
 sky130_fd_sc_hd__conb_1 _1486__48 (.LO(net48));
 sky130_fd_sc_hd__conb_1 _1487__49 (.LO(net49));
 sky130_fd_sc_hd__conb_1 _1488__50 (.LO(net50));
 sky130_fd_sc_hd__conb_1 _1489__51 (.LO(net51));
 sky130_fd_sc_hd__conb_1 _1490__52 (.LO(net52));
 sky130_fd_sc_hd__conb_1 _1491__53 (.LO(net53));
 sky130_fd_sc_hd__conb_1 _1492__54 (.LO(net54));
 sky130_fd_sc_hd__conb_1 _1496__55 (.LO(net55));
 sky130_fd_sc_hd__conb_1 _1497__56 (.LO(net56));
 sky130_fd_sc_hd__conb_1 _1498__57 (.LO(net57));
 sky130_fd_sc_hd__conb_1 _1499__58 (.LO(net58));
 sky130_fd_sc_hd__conb_1 _1500__59 (.LO(net59));
 sky130_fd_sc_hd__conb_1 _1501__60 (.LO(net60));
 sky130_fd_sc_hd__conb_1 _1502__61 (.LO(net61));
 sky130_fd_sc_hd__conb_1 _1503__62 (.LO(net62));
 sky130_fd_sc_hd__conb_1 _1504__63 (.LO(net63));
 sky130_fd_sc_hd__conb_1 _1505__64 (.LO(net64));
 sky130_fd_sc_hd__conb_1 _1506__65 (.LO(net65));
 sky130_fd_sc_hd__conb_1 _1507__66 (.LO(net66));
 sky130_fd_sc_hd__conb_1 _1508__67 (.LO(net67));
 sky130_fd_sc_hd__conb_1 _1509__68 (.LO(net68));
 sky130_fd_sc_hd__conb_1 _1510__69 (.LO(net69));
 sky130_fd_sc_hd__conb_1 _1511__70 (.LO(net70));
 sky130_fd_sc_hd__conb_1 _1512__71 (.LO(net71));
 sky130_fd_sc_hd__conb_1 _1513__72 (.LO(net72));
 sky130_fd_sc_hd__conb_1 _1514__73 (.LO(net73));
 sky130_fd_sc_hd__conb_1 _1515__74 (.LO(net74));
 sky130_fd_sc_hd__conb_1 _1516__75 (.LO(net75));
 sky130_fd_sc_hd__conb_1 _1517__76 (.LO(net76));
 sky130_fd_sc_hd__conb_1 _1518__77 (.LO(net77));
 sky130_fd_sc_hd__conb_1 _1519__78 (.LO(net78));
 sky130_fd_sc_hd__conb_1 _1520__79 (.LO(net79));
 sky130_fd_sc_hd__conb_1 _1521__80 (.LO(net80));
 sky130_fd_sc_hd__conb_1 _1522__81 (.LO(net81));
 sky130_fd_sc_hd__conb_1 _1523__82 (.LO(net82));
 sky130_fd_sc_hd__conb_1 _1524__83 (.LO(net83));
 sky130_fd_sc_hd__conb_1 _1525__84 (.LO(net84));
 sky130_fd_sc_hd__conb_1 _1526__85 (.LO(net85));
 sky130_fd_sc_hd__conb_1 _1527__86 (.LO(net86));
 sky130_fd_sc_hd__conb_1 _1528__87 (.LO(net87));
 sky130_fd_sc_hd__conb_1 _1529__88 (.LO(net88));
 sky130_fd_sc_hd__conb_1 _1530__89 (.LO(net89));
 sky130_fd_sc_hd__conb_1 _1531__90 (.LO(net90));
 sky130_fd_sc_hd__conb_1 _1532__91 (.LO(net91));
 sky130_fd_sc_hd__conb_1 _1533__92 (.LO(net92));
 sky130_fd_sc_hd__conb_1 _1534__93 (.LO(net93));
 sky130_fd_sc_hd__conb_1 _1535__94 (.LO(net94));
 sky130_fd_sc_hd__conb_1 _1536__95 (.LO(net95));
 sky130_fd_sc_hd__conb_1 _1537__96 (.LO(net96));
 sky130_fd_sc_hd__conb_1 _1538__97 (.LO(net97));
 sky130_fd_sc_hd__conb_1 _1539__98 (.LO(net98));
 sky130_fd_sc_hd__conb_1 _1540__99 (.LO(net99));
 sky130_fd_sc_hd__conb_1 _1541__100 (.LO(net100));
 sky130_fd_sc_hd__conb_1 _1542__101 (.LO(net101));
 sky130_fd_sc_hd__conb_1 _1543__102 (.LO(net102));
 sky130_fd_sc_hd__conb_1 _1544__103 (.LO(net103));
 sky130_fd_sc_hd__conb_1 _1545__104 (.LO(net104));
 sky130_fd_sc_hd__conb_1 _1546__105 (.LO(net105));
 sky130_fd_sc_hd__conb_1 _1547__106 (.LO(net106));
 sky130_fd_sc_hd__conb_1 _1548__107 (.LO(net107));
 sky130_fd_sc_hd__conb_1 _1549__108 (.LO(net108));
 sky130_fd_sc_hd__conb_1 _1550__109 (.LO(net109));
 sky130_fd_sc_hd__conb_1 _1551__110 (.LO(net110));
 sky130_fd_sc_hd__conb_1 _1552__111 (.LO(net111));
 sky130_fd_sc_hd__conb_1 _1553__112 (.LO(net112));
 sky130_fd_sc_hd__conb_1 _1554__113 (.LO(net113));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__ebufn_8 _1447_ (.A(net9),
    .TE_B(_0455_),
    .Z(la1_data_out[0]));
 sky130_fd_sc_hd__ebufn_8 _1448_ (.A(net10),
    .TE_B(_0456_),
    .Z(la1_data_out[1]));
 sky130_fd_sc_hd__ebufn_8 _1449_ (.A(net11),
    .TE_B(_0457_),
    .Z(la1_data_out[2]));
 sky130_fd_sc_hd__ebufn_8 _1450_ (.A(net12),
    .TE_B(_0458_),
    .Z(la1_data_out[3]));
 sky130_fd_sc_hd__ebufn_8 _1451_ (.A(net13),
    .TE_B(_0459_),
    .Z(la1_data_out[4]));
 sky130_fd_sc_hd__ebufn_8 _1452_ (.A(net14),
    .TE_B(_0460_),
    .Z(la1_data_out[5]));
 sky130_fd_sc_hd__ebufn_8 _1453_ (.A(net15),
    .TE_B(_0461_),
    .Z(la1_data_out[6]));
 sky130_fd_sc_hd__ebufn_8 _1454_ (.A(net16),
    .TE_B(_0462_),
    .Z(la1_data_out[7]));
 sky130_fd_sc_hd__ebufn_8 _1455_ (.A(net17),
    .TE_B(_0463_),
    .Z(la1_data_out[8]));
 sky130_fd_sc_hd__ebufn_8 _1456_ (.A(net18),
    .TE_B(_0464_),
    .Z(la1_data_out[9]));
 sky130_fd_sc_hd__ebufn_8 _1457_ (.A(net19),
    .TE_B(_0465_),
    .Z(la1_data_out[10]));
 sky130_fd_sc_hd__ebufn_8 _1458_ (.A(net20),
    .TE_B(_0466_),
    .Z(la1_data_out[11]));
 sky130_fd_sc_hd__ebufn_8 _1459_ (.A(net21),
    .TE_B(_0467_),
    .Z(la1_data_out[12]));
 sky130_fd_sc_hd__ebufn_8 _1460_ (.A(net22),
    .TE_B(_0468_),
    .Z(la1_data_out[13]));
 sky130_fd_sc_hd__ebufn_8 _1461_ (.A(net23),
    .TE_B(_0469_),
    .Z(la1_data_out[14]));
 sky130_fd_sc_hd__ebufn_8 _1462_ (.A(net24),
    .TE_B(_0470_),
    .Z(la1_data_out[15]));
 sky130_fd_sc_hd__ebufn_8 _1463_ (.A(net25),
    .TE_B(_0471_),
    .Z(la1_data_out[16]));
 sky130_fd_sc_hd__ebufn_8 _1464_ (.A(net26),
    .TE_B(_0472_),
    .Z(la1_data_out[17]));
 sky130_fd_sc_hd__ebufn_8 _1465_ (.A(net27),
    .TE_B(_0473_),
    .Z(la1_data_out[18]));
 sky130_fd_sc_hd__ebufn_8 _1466_ (.A(net28),
    .TE_B(_0474_),
    .Z(la1_data_out[19]));
 sky130_fd_sc_hd__ebufn_8 _1467_ (.A(net29),
    .TE_B(_0475_),
    .Z(la1_data_out[20]));
 sky130_fd_sc_hd__ebufn_8 _1468_ (.A(net30),
    .TE_B(_0476_),
    .Z(la1_data_out[21]));
 sky130_fd_sc_hd__ebufn_8 _1469_ (.A(net31),
    .TE_B(_0477_),
    .Z(la1_data_out[22]));
 sky130_fd_sc_hd__ebufn_8 _1470_ (.A(net32),
    .TE_B(_0478_),
    .Z(la1_data_out[23]));
 sky130_fd_sc_hd__ebufn_8 _1471_ (.A(net33),
    .TE_B(_0479_),
    .Z(la1_data_out[24]));
 sky130_fd_sc_hd__ebufn_8 _1472_ (.A(net34),
    .TE_B(_0480_),
    .Z(la1_data_out[25]));
 sky130_fd_sc_hd__ebufn_8 _1473_ (.A(net35),
    .TE_B(_0481_),
    .Z(la1_data_out[26]));
 sky130_fd_sc_hd__ebufn_8 _1474_ (.A(net36),
    .TE_B(_0482_),
    .Z(la1_data_out[27]));
 sky130_fd_sc_hd__ebufn_8 _1475_ (.A(net37),
    .TE_B(_0483_),
    .Z(la1_data_out[28]));
 sky130_fd_sc_hd__ebufn_8 _1476_ (.A(net38),
    .TE_B(_0484_),
    .Z(la1_data_out[29]));
 sky130_fd_sc_hd__ebufn_8 _1477_ (.A(net39),
    .TE_B(_0485_),
    .Z(la1_data_out[30]));
 sky130_fd_sc_hd__ebufn_8 _1478_ (.A(net40),
    .TE_B(_0486_),
    .Z(la1_data_out[31]));
 sky130_fd_sc_hd__ebufn_8 _1479_ (.A(net41),
    .TE_B(_0487_),
    .Z(io_out[0]));
 sky130_fd_sc_hd__ebufn_8 _1480_ (.A(net42),
    .TE_B(_0488_),
    .Z(io_out[1]));
 sky130_fd_sc_hd__ebufn_8 _1481_ (.A(net43),
    .TE_B(_0489_),
    .Z(io_out[2]));
 sky130_fd_sc_hd__ebufn_8 _1482_ (.A(net44),
    .TE_B(_0490_),
    .Z(io_out[3]));
 sky130_fd_sc_hd__ebufn_8 _1483_ (.A(net45),
    .TE_B(_0491_),
    .Z(io_out[4]));
 sky130_fd_sc_hd__ebufn_8 _1484_ (.A(net46),
    .TE_B(_0492_),
    .Z(io_out[5]));
 sky130_fd_sc_hd__ebufn_8 _1485_ (.A(net47),
    .TE_B(_0493_),
    .Z(io_out[6]));
 sky130_fd_sc_hd__ebufn_8 _1486_ (.A(net48),
    .TE_B(_0494_),
    .Z(io_out[7]));
 sky130_fd_sc_hd__ebufn_8 _1487_ (.A(net49),
    .TE_B(_0495_),
    .Z(io_out[8]));
 sky130_fd_sc_hd__ebufn_8 _1488_ (.A(net50),
    .TE_B(_0496_),
    .Z(io_out[9]));
 sky130_fd_sc_hd__ebufn_8 _1489_ (.A(net51),
    .TE_B(_0497_),
    .Z(io_out[10]));
 sky130_fd_sc_hd__ebufn_8 _1490_ (.A(net52),
    .TE_B(_0498_),
    .Z(io_out[11]));
 sky130_fd_sc_hd__ebufn_8 _1491_ (.A(net53),
    .TE_B(_0499_),
    .Z(io_out[12]));
 sky130_fd_sc_hd__ebufn_8 _1492_ (.A(net54),
    .TE_B(_0500_),
    .Z(io_out[13]));
 sky130_fd_sc_hd__ebufn_8 _1493_ (.A(\rgb_mixer0.pwm0.out ),
    .TE_B(_0501_),
    .Z(io_out[14]));
 sky130_fd_sc_hd__ebufn_8 _1494_ (.A(\rgb_mixer0.pwm1.out ),
    .TE_B(_0502_),
    .Z(io_out[15]));
 sky130_fd_sc_hd__ebufn_8 _1495_ (.A(\rgb_mixer0.pwm2.out ),
    .TE_B(_0503_),
    .Z(io_out[16]));
 sky130_fd_sc_hd__ebufn_8 _1496_ (.A(net55),
    .TE_B(_0504_),
    .Z(io_out[17]));
 sky130_fd_sc_hd__ebufn_8 _1497_ (.A(net56),
    .TE_B(_0505_),
    .Z(io_out[18]));
 sky130_fd_sc_hd__ebufn_8 _1498_ (.A(net57),
    .TE_B(_0506_),
    .Z(io_out[19]));
 sky130_fd_sc_hd__ebufn_8 _1499_ (.A(net58),
    .TE_B(_0507_),
    .Z(io_out[20]));
 sky130_fd_sc_hd__ebufn_8 _1500_ (.A(net59),
    .TE_B(_0508_),
    .Z(io_out[21]));
 sky130_fd_sc_hd__ebufn_8 _1501_ (.A(net60),
    .TE_B(_0509_),
    .Z(io_out[22]));
 sky130_fd_sc_hd__ebufn_8 _1502_ (.A(net61),
    .TE_B(_0510_),
    .Z(io_out[23]));
 sky130_fd_sc_hd__ebufn_8 _1503_ (.A(net62),
    .TE_B(_0511_),
    .Z(io_out[24]));
 sky130_fd_sc_hd__ebufn_8 _1504_ (.A(net63),
    .TE_B(_0512_),
    .Z(io_out[25]));
 sky130_fd_sc_hd__ebufn_8 _1505_ (.A(net64),
    .TE_B(_0513_),
    .Z(io_out[26]));
 sky130_fd_sc_hd__ebufn_8 _1506_ (.A(net65),
    .TE_B(_0514_),
    .Z(io_out[27]));
 sky130_fd_sc_hd__ebufn_8 _1507_ (.A(net66),
    .TE_B(_0515_),
    .Z(io_out[28]));
 sky130_fd_sc_hd__ebufn_8 _1508_ (.A(net67),
    .TE_B(_0516_),
    .Z(io_out[29]));
 sky130_fd_sc_hd__ebufn_8 _1509_ (.A(net68),
    .TE_B(_0517_),
    .Z(io_out[30]));
 sky130_fd_sc_hd__ebufn_8 _1510_ (.A(net69),
    .TE_B(_0518_),
    .Z(io_out[31]));
 sky130_fd_sc_hd__ebufn_8 _1511_ (.A(net70),
    .TE_B(_0519_),
    .Z(io_out[32]));
 sky130_fd_sc_hd__ebufn_8 _1512_ (.A(net71),
    .TE_B(_0520_),
    .Z(io_out[33]));
 sky130_fd_sc_hd__ebufn_8 _1513_ (.A(net72),
    .TE_B(_0521_),
    .Z(io_out[34]));
 sky130_fd_sc_hd__ebufn_8 _1514_ (.A(net73),
    .TE_B(_0522_),
    .Z(io_out[35]));
 sky130_fd_sc_hd__ebufn_8 _1515_ (.A(net74),
    .TE_B(_0523_),
    .Z(io_out[36]));
 sky130_fd_sc_hd__ebufn_8 _1516_ (.A(net75),
    .TE_B(_0524_),
    .Z(io_out[37]));
 sky130_fd_sc_hd__ebufn_8 _1517_ (.A(net76),
    .TE_B(_0525_),
    .Z(io_oeb[0]));
 sky130_fd_sc_hd__ebufn_8 _1518_ (.A(net77),
    .TE_B(_0526_),
    .Z(io_oeb[1]));
 sky130_fd_sc_hd__ebufn_8 _1519_ (.A(net78),
    .TE_B(_0527_),
    .Z(io_oeb[2]));
 sky130_fd_sc_hd__ebufn_8 _1520_ (.A(net79),
    .TE_B(_0528_),
    .Z(io_oeb[3]));
 sky130_fd_sc_hd__ebufn_8 _1521_ (.A(net80),
    .TE_B(_0529_),
    .Z(io_oeb[4]));
 sky130_fd_sc_hd__ebufn_8 _1522_ (.A(net81),
    .TE_B(_0530_),
    .Z(io_oeb[5]));
 sky130_fd_sc_hd__ebufn_8 _1523_ (.A(net82),
    .TE_B(_0531_),
    .Z(io_oeb[6]));
 sky130_fd_sc_hd__ebufn_8 _1524_ (.A(net83),
    .TE_B(_0532_),
    .Z(io_oeb[7]));
 sky130_fd_sc_hd__ebufn_8 _1525_ (.A(net84),
    .TE_B(_0533_),
    .Z(io_oeb[8]));
 sky130_fd_sc_hd__ebufn_8 _1526_ (.A(net85),
    .TE_B(_0534_),
    .Z(io_oeb[9]));
 sky130_fd_sc_hd__ebufn_8 _1527_ (.A(net86),
    .TE_B(_0535_),
    .Z(io_oeb[10]));
 sky130_fd_sc_hd__ebufn_8 _1528_ (.A(net87),
    .TE_B(_0536_),
    .Z(io_oeb[11]));
 sky130_fd_sc_hd__ebufn_8 _1529_ (.A(net88),
    .TE_B(_0537_),
    .Z(io_oeb[12]));
 sky130_fd_sc_hd__ebufn_8 _1530_ (.A(net89),
    .TE_B(_0538_),
    .Z(io_oeb[13]));
 sky130_fd_sc_hd__ebufn_8 _1531_ (.A(net90),
    .TE_B(_0539_),
    .Z(io_oeb[14]));
 sky130_fd_sc_hd__ebufn_8 _1532_ (.A(net91),
    .TE_B(_0540_),
    .Z(io_oeb[15]));
 sky130_fd_sc_hd__ebufn_8 _1533_ (.A(net92),
    .TE_B(_0541_),
    .Z(io_oeb[16]));
 sky130_fd_sc_hd__ebufn_8 _1534_ (.A(net93),
    .TE_B(_0542_),
    .Z(io_oeb[17]));
 sky130_fd_sc_hd__ebufn_8 _1535_ (.A(net94),
    .TE_B(_0543_),
    .Z(io_oeb[18]));
 sky130_fd_sc_hd__ebufn_8 _1536_ (.A(net95),
    .TE_B(_0544_),
    .Z(io_oeb[19]));
 sky130_fd_sc_hd__ebufn_8 _1537_ (.A(net96),
    .TE_B(_0545_),
    .Z(io_oeb[20]));
 sky130_fd_sc_hd__ebufn_8 _1538_ (.A(net97),
    .TE_B(_0546_),
    .Z(io_oeb[21]));
 sky130_fd_sc_hd__ebufn_8 _1539_ (.A(net98),
    .TE_B(_0547_),
    .Z(io_oeb[22]));
 sky130_fd_sc_hd__ebufn_8 _1540_ (.A(net99),
    .TE_B(_0548_),
    .Z(io_oeb[23]));
 sky130_fd_sc_hd__ebufn_8 _1541_ (.A(net100),
    .TE_B(_0549_),
    .Z(io_oeb[24]));
 sky130_fd_sc_hd__ebufn_8 _1542_ (.A(net101),
    .TE_B(_0550_),
    .Z(io_oeb[25]));
 sky130_fd_sc_hd__ebufn_8 _1543_ (.A(net102),
    .TE_B(_0551_),
    .Z(io_oeb[26]));
 sky130_fd_sc_hd__ebufn_8 _1544_ (.A(net103),
    .TE_B(_0552_),
    .Z(io_oeb[27]));
 sky130_fd_sc_hd__ebufn_8 _1545_ (.A(net104),
    .TE_B(_0553_),
    .Z(io_oeb[28]));
 sky130_fd_sc_hd__ebufn_8 _1546_ (.A(net105),
    .TE_B(_0554_),
    .Z(io_oeb[29]));
 sky130_fd_sc_hd__ebufn_8 _1547_ (.A(net106),
    .TE_B(_0555_),
    .Z(io_oeb[30]));
 sky130_fd_sc_hd__ebufn_8 _1548_ (.A(net107),
    .TE_B(_0556_),
    .Z(io_oeb[31]));
 sky130_fd_sc_hd__ebufn_8 _1549_ (.A(net108),
    .TE_B(_0557_),
    .Z(io_oeb[32]));
 sky130_fd_sc_hd__ebufn_8 _1550_ (.A(net109),
    .TE_B(_0558_),
    .Z(io_oeb[33]));
 sky130_fd_sc_hd__ebufn_8 _1551_ (.A(net110),
    .TE_B(_0559_),
    .Z(io_oeb[34]));
 sky130_fd_sc_hd__ebufn_8 _1552_ (.A(net111),
    .TE_B(_0560_),
    .Z(io_oeb[35]));
 sky130_fd_sc_hd__ebufn_8 _1553_ (.A(net112),
    .TE_B(_0561_),
    .Z(io_oeb[36]));
 sky130_fd_sc_hd__ebufn_8 _1554_ (.A(net113),
    .TE_B(_0562_),
    .Z(io_oeb[37]));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(active),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(io_in[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(io_in[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(io_in[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(io_in[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(io_in[8]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(io_in[9]),
    .X(net7));
 sky130_fd_sc_hd__buf_2 input8 (.A(la1_data_in[0]),
    .X(net8));
 sky130_fd_sc_hd__conb_1 _1447__9 (.LO(net9));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_4__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_5__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_6__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_7__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0050_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_0102_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_0361_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_0338_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_0445_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(io_in[12]));
 sky130_fd_sc_hd__fill_2 FILLER_0_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_199 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_303 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_226 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_362 ();
endmodule

