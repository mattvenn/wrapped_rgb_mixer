magic
tech sky130A
magscale 1 2
timestamp 1670925203
<< obsli1 >>
rect 1104 2159 34868 39729
<< obsm1 >>
rect 658 1096 35958 40044
<< metal2 >>
rect -10 41200 102 41800
rect 634 41200 746 41800
rect 1278 41200 1390 41800
rect 1922 41200 2034 41800
rect 2566 41200 2678 41800
rect 3210 41200 3322 41800
rect 4498 41200 4610 41800
rect 5142 41200 5254 41800
rect 5786 41200 5898 41800
rect 6430 41200 6542 41800
rect 7074 41200 7186 41800
rect 7718 41200 7830 41800
rect 8362 41200 8474 41800
rect 9006 41200 9118 41800
rect 9650 41200 9762 41800
rect 10938 41200 11050 41800
rect 11582 41200 11694 41800
rect 12226 41200 12338 41800
rect 12870 41200 12982 41800
rect 13514 41200 13626 41800
rect 14158 41200 14270 41800
rect 14802 41200 14914 41800
rect 15446 41200 15558 41800
rect 16090 41200 16202 41800
rect 17378 41200 17490 41800
rect 18022 41200 18134 41800
rect 18666 41200 18778 41800
rect 19310 41200 19422 41800
rect 19954 41200 20066 41800
rect 20598 41200 20710 41800
rect 21242 41200 21354 41800
rect 21886 41200 21998 41800
rect 22530 41200 22642 41800
rect 23818 41200 23930 41800
rect 24462 41200 24574 41800
rect 25106 41200 25218 41800
rect 25750 41200 25862 41800
rect 26394 41200 26506 41800
rect 27038 41200 27150 41800
rect 27682 41200 27794 41800
rect 28326 41200 28438 41800
rect 28970 41200 29082 41800
rect 30258 41200 30370 41800
rect 30902 41200 31014 41800
rect 31546 41200 31658 41800
rect 32190 41200 32302 41800
rect 32834 41200 32946 41800
rect 33478 41200 33590 41800
rect 34122 41200 34234 41800
rect 34766 41200 34878 41800
rect 35410 41200 35522 41800
rect -10 200 102 800
rect 634 200 746 800
rect 1278 200 1390 800
rect 1922 200 2034 800
rect 2566 200 2678 800
rect 3210 200 3322 800
rect 3854 200 3966 800
rect 4498 200 4610 800
rect 5142 200 5254 800
rect 6430 200 6542 800
rect 7074 200 7186 800
rect 7718 200 7830 800
rect 8362 200 8474 800
rect 9006 200 9118 800
rect 9650 200 9762 800
rect 10294 200 10406 800
rect 10938 200 11050 800
rect 11582 200 11694 800
rect 12870 200 12982 800
rect 13514 200 13626 800
rect 14158 200 14270 800
rect 14802 200 14914 800
rect 15446 200 15558 800
rect 16090 200 16202 800
rect 16734 200 16846 800
rect 17378 200 17490 800
rect 18022 200 18134 800
rect 19310 200 19422 800
rect 19954 200 20066 800
rect 20598 200 20710 800
rect 21242 200 21354 800
rect 21886 200 21998 800
rect 22530 200 22642 800
rect 23174 200 23286 800
rect 23818 200 23930 800
rect 24462 200 24574 800
rect 25750 200 25862 800
rect 26394 200 26506 800
rect 27038 200 27150 800
rect 27682 200 27794 800
rect 28326 200 28438 800
rect 28970 200 29082 800
rect 29614 200 29726 800
rect 30258 200 30370 800
rect 30902 200 31014 800
rect 32190 200 32302 800
rect 32834 200 32946 800
rect 33478 200 33590 800
rect 34122 200 34234 800
rect 34766 200 34878 800
rect 35410 200 35522 800
<< obsm2 >>
rect 802 41144 1222 41585
rect 1446 41144 1866 41585
rect 2090 41144 2510 41585
rect 2734 41144 3154 41585
rect 3378 41144 4442 41585
rect 4666 41144 5086 41585
rect 5310 41144 5730 41585
rect 5954 41144 6374 41585
rect 6598 41144 7018 41585
rect 7242 41144 7662 41585
rect 7886 41144 8306 41585
rect 8530 41144 8950 41585
rect 9174 41144 9594 41585
rect 9818 41144 10882 41585
rect 11106 41144 11526 41585
rect 11750 41144 12170 41585
rect 12394 41144 12814 41585
rect 13038 41144 13458 41585
rect 13682 41144 14102 41585
rect 14326 41144 14746 41585
rect 14970 41144 15390 41585
rect 15614 41144 16034 41585
rect 16258 41144 17322 41585
rect 17546 41144 17966 41585
rect 18190 41144 18610 41585
rect 18834 41144 19254 41585
rect 19478 41144 19898 41585
rect 20122 41144 20542 41585
rect 20766 41144 21186 41585
rect 21410 41144 21830 41585
rect 22054 41144 22474 41585
rect 22698 41144 23762 41585
rect 23986 41144 24406 41585
rect 24630 41144 25050 41585
rect 25274 41144 25694 41585
rect 25918 41144 26338 41585
rect 26562 41144 26982 41585
rect 27206 41144 27626 41585
rect 27850 41144 28270 41585
rect 28494 41144 28914 41585
rect 29138 41144 30202 41585
rect 30426 41144 30846 41585
rect 31070 41144 31490 41585
rect 31714 41144 32134 41585
rect 32358 41144 32778 41585
rect 33002 41144 33422 41585
rect 33646 41144 34066 41585
rect 34290 41144 34710 41585
rect 34934 41144 35354 41585
rect 35578 41144 35954 41585
rect 664 856 35954 41144
rect 802 144 1222 856
rect 1446 144 1866 856
rect 2090 144 2510 856
rect 2734 144 3154 856
rect 3378 144 3798 856
rect 4022 144 4442 856
rect 4666 144 5086 856
rect 5310 144 6374 856
rect 6598 144 7018 856
rect 7242 144 7662 856
rect 7886 144 8306 856
rect 8530 144 8950 856
rect 9174 144 9594 856
rect 9818 144 10238 856
rect 10462 144 10882 856
rect 11106 144 11526 856
rect 11750 144 12814 856
rect 13038 144 13458 856
rect 13682 144 14102 856
rect 14326 144 14746 856
rect 14970 144 15390 856
rect 15614 144 16034 856
rect 16258 144 16678 856
rect 16902 144 17322 856
rect 17546 144 17966 856
rect 18190 144 19254 856
rect 19478 144 19898 856
rect 20122 144 20542 856
rect 20766 144 21186 856
rect 21410 144 21830 856
rect 22054 144 22474 856
rect 22698 144 23118 856
rect 23342 144 23762 856
rect 23986 144 24406 856
rect 24630 144 25694 856
rect 25918 144 26338 856
rect 26562 144 26982 856
rect 27206 144 27626 856
rect 27850 144 28270 856
rect 28494 144 28914 856
rect 29138 144 29558 856
rect 29782 144 30202 856
rect 30426 144 30846 856
rect 31070 144 32134 856
rect 32358 144 32778 856
rect 33002 144 33422 856
rect 33646 144 34066 856
rect 34290 144 34710 856
rect 34934 144 35354 856
rect 35578 144 35954 856
rect 664 31 35954 144
<< metal3 >>
rect 200 41428 800 41668
rect 200 40748 800 40988
rect 35200 40748 35800 40988
rect 35200 40068 35800 40308
rect 200 39388 800 39628
rect 35200 39388 35800 39628
rect 200 38708 800 38948
rect 35200 38708 35800 38948
rect 200 38028 800 38268
rect 35200 38028 35800 38268
rect 200 37348 800 37588
rect 35200 37348 35800 37588
rect 200 36668 800 36908
rect 35200 36668 35800 36908
rect 200 35988 800 36228
rect 35200 35988 35800 36228
rect 200 35308 800 35548
rect 200 34628 800 34868
rect 35200 34628 35800 34868
rect 200 33948 800 34188
rect 35200 33948 35800 34188
rect 35200 33268 35800 33508
rect 200 32588 800 32828
rect 35200 32588 35800 32828
rect 200 31908 800 32148
rect 35200 31908 35800 32148
rect 200 31228 800 31468
rect 35200 31228 35800 31468
rect 200 30548 800 30788
rect 35200 30548 35800 30788
rect 200 29868 800 30108
rect 35200 29868 35800 30108
rect 200 29188 800 29428
rect 35200 29188 35800 29428
rect 200 28508 800 28748
rect 200 27828 800 28068
rect 35200 27828 35800 28068
rect 200 27148 800 27388
rect 35200 27148 35800 27388
rect 35200 26468 35800 26708
rect 200 25788 800 26028
rect 35200 25788 35800 26028
rect 200 25108 800 25348
rect 35200 25108 35800 25348
rect 200 24428 800 24668
rect 35200 24428 35800 24668
rect 200 23748 800 23988
rect 35200 23748 35800 23988
rect 200 23068 800 23308
rect 35200 23068 35800 23308
rect 200 22388 800 22628
rect 35200 22388 35800 22628
rect 200 21708 800 21948
rect 200 21028 800 21268
rect 35200 21028 35800 21268
rect 200 20348 800 20588
rect 35200 20348 35800 20588
rect 35200 19668 35800 19908
rect 200 18988 800 19228
rect 35200 18988 35800 19228
rect 200 18308 800 18548
rect 35200 18308 35800 18548
rect 200 17628 800 17868
rect 35200 17628 35800 17868
rect 200 16948 800 17188
rect 35200 16948 35800 17188
rect 200 16268 800 16508
rect 35200 16268 35800 16508
rect 200 15588 800 15828
rect 35200 15588 35800 15828
rect 200 14908 800 15148
rect 200 14228 800 14468
rect 35200 14228 35800 14468
rect 200 13548 800 13788
rect 35200 13548 35800 13788
rect 35200 12868 35800 13108
rect 200 12188 800 12428
rect 35200 12188 35800 12428
rect 200 11508 800 11748
rect 35200 11508 35800 11748
rect 200 10828 800 11068
rect 35200 10828 35800 11068
rect 200 10148 800 10388
rect 35200 10148 35800 10388
rect 200 9468 800 9708
rect 35200 9468 35800 9708
rect 200 8788 800 9028
rect 35200 8788 35800 9028
rect 200 8108 800 8348
rect 200 7428 800 7668
rect 35200 7428 35800 7668
rect 200 6748 800 6988
rect 35200 6748 35800 6988
rect 35200 6068 35800 6308
rect 200 5388 800 5628
rect 35200 5388 35800 5628
rect 200 4708 800 4948
rect 35200 4708 35800 4948
rect 200 4028 800 4268
rect 35200 4028 35800 4268
rect 200 3348 800 3588
rect 35200 3348 35800 3588
rect 200 2668 800 2908
rect 35200 2668 35800 2908
rect 200 1988 800 2228
rect 35200 1988 35800 2228
rect 200 1308 800 1548
rect 200 628 800 868
rect 35200 628 35800 868
rect 35200 -52 35800 188
<< obsm3 >>
rect 880 41348 35959 41581
rect 800 41068 35959 41348
rect 880 40668 35120 41068
rect 35880 40668 35959 41068
rect 800 40388 35959 40668
rect 800 39988 35120 40388
rect 35880 39988 35959 40388
rect 800 39708 35959 39988
rect 880 39308 35120 39708
rect 35880 39308 35959 39708
rect 800 39028 35959 39308
rect 880 38628 35120 39028
rect 35880 38628 35959 39028
rect 800 38348 35959 38628
rect 880 37948 35120 38348
rect 35880 37948 35959 38348
rect 800 37668 35959 37948
rect 880 37268 35120 37668
rect 35880 37268 35959 37668
rect 800 36988 35959 37268
rect 880 36588 35120 36988
rect 35880 36588 35959 36988
rect 800 36308 35959 36588
rect 880 35908 35120 36308
rect 35880 35908 35959 36308
rect 800 35628 35959 35908
rect 880 35228 35959 35628
rect 800 34948 35959 35228
rect 880 34548 35120 34948
rect 35880 34548 35959 34948
rect 800 34268 35959 34548
rect 880 33868 35120 34268
rect 35880 33868 35959 34268
rect 800 33588 35959 33868
rect 800 33188 35120 33588
rect 35880 33188 35959 33588
rect 800 32908 35959 33188
rect 880 32508 35120 32908
rect 35880 32508 35959 32908
rect 800 32228 35959 32508
rect 880 31828 35120 32228
rect 35880 31828 35959 32228
rect 800 31548 35959 31828
rect 880 31148 35120 31548
rect 35880 31148 35959 31548
rect 800 30868 35959 31148
rect 880 30468 35120 30868
rect 35880 30468 35959 30868
rect 800 30188 35959 30468
rect 880 29788 35120 30188
rect 35880 29788 35959 30188
rect 800 29508 35959 29788
rect 880 29108 35120 29508
rect 35880 29108 35959 29508
rect 800 28828 35959 29108
rect 880 28428 35959 28828
rect 800 28148 35959 28428
rect 880 27748 35120 28148
rect 35880 27748 35959 28148
rect 800 27468 35959 27748
rect 880 27068 35120 27468
rect 35880 27068 35959 27468
rect 800 26788 35959 27068
rect 800 26388 35120 26788
rect 35880 26388 35959 26788
rect 800 26108 35959 26388
rect 880 25708 35120 26108
rect 35880 25708 35959 26108
rect 800 25428 35959 25708
rect 880 25028 35120 25428
rect 35880 25028 35959 25428
rect 800 24748 35959 25028
rect 880 24348 35120 24748
rect 35880 24348 35959 24748
rect 800 24068 35959 24348
rect 880 23668 35120 24068
rect 35880 23668 35959 24068
rect 800 23388 35959 23668
rect 880 22988 35120 23388
rect 35880 22988 35959 23388
rect 800 22708 35959 22988
rect 880 22308 35120 22708
rect 35880 22308 35959 22708
rect 800 22028 35959 22308
rect 880 21628 35959 22028
rect 800 21348 35959 21628
rect 880 20948 35120 21348
rect 35880 20948 35959 21348
rect 800 20668 35959 20948
rect 880 20268 35120 20668
rect 35880 20268 35959 20668
rect 800 19988 35959 20268
rect 800 19588 35120 19988
rect 35880 19588 35959 19988
rect 800 19308 35959 19588
rect 880 18908 35120 19308
rect 35880 18908 35959 19308
rect 800 18628 35959 18908
rect 880 18228 35120 18628
rect 35880 18228 35959 18628
rect 800 17948 35959 18228
rect 880 17548 35120 17948
rect 35880 17548 35959 17948
rect 800 17268 35959 17548
rect 880 16868 35120 17268
rect 35880 16868 35959 17268
rect 800 16588 35959 16868
rect 880 16188 35120 16588
rect 35880 16188 35959 16588
rect 800 15908 35959 16188
rect 880 15508 35120 15908
rect 35880 15508 35959 15908
rect 800 15228 35959 15508
rect 880 14828 35959 15228
rect 800 14548 35959 14828
rect 880 14148 35120 14548
rect 35880 14148 35959 14548
rect 800 13868 35959 14148
rect 880 13468 35120 13868
rect 35880 13468 35959 13868
rect 800 13188 35959 13468
rect 800 12788 35120 13188
rect 35880 12788 35959 13188
rect 800 12508 35959 12788
rect 880 12108 35120 12508
rect 35880 12108 35959 12508
rect 800 11828 35959 12108
rect 880 11428 35120 11828
rect 35880 11428 35959 11828
rect 800 11148 35959 11428
rect 880 10748 35120 11148
rect 35880 10748 35959 11148
rect 800 10468 35959 10748
rect 880 10068 35120 10468
rect 35880 10068 35959 10468
rect 800 9788 35959 10068
rect 880 9388 35120 9788
rect 35880 9388 35959 9788
rect 800 9108 35959 9388
rect 880 8708 35120 9108
rect 35880 8708 35959 9108
rect 800 8428 35959 8708
rect 880 8028 35959 8428
rect 800 7748 35959 8028
rect 880 7348 35120 7748
rect 35880 7348 35959 7748
rect 800 7068 35959 7348
rect 880 6668 35120 7068
rect 35880 6668 35959 7068
rect 800 6388 35959 6668
rect 800 5988 35120 6388
rect 35880 5988 35959 6388
rect 800 5708 35959 5988
rect 880 5308 35120 5708
rect 35880 5308 35959 5708
rect 800 5028 35959 5308
rect 880 4628 35120 5028
rect 35880 4628 35959 5028
rect 800 4348 35959 4628
rect 880 3948 35120 4348
rect 35880 3948 35959 4348
rect 800 3668 35959 3948
rect 880 3268 35120 3668
rect 35880 3268 35959 3668
rect 800 2988 35959 3268
rect 880 2588 35120 2988
rect 35880 2588 35959 2988
rect 800 2308 35959 2588
rect 880 1908 35120 2308
rect 35880 1908 35959 2308
rect 800 1628 35959 1908
rect 880 1228 35959 1628
rect 800 948 35959 1228
rect 880 548 35120 948
rect 35880 548 35959 948
rect 800 268 35959 548
rect 800 35 35120 268
rect 35880 35 35959 268
<< metal4 >>
rect 5164 2128 5484 39760
rect 9384 2128 9704 39760
rect 13605 2128 13925 39760
rect 17825 2128 18145 39760
rect 22046 2128 22366 39760
rect 26266 2128 26586 39760
rect 30487 2128 30807 39760
rect 34707 2128 35027 39760
<< obsm4 >>
rect 23427 11731 26186 39405
rect 26666 11731 30407 39405
rect 30887 11731 34165 39405
<< labels >>
rlabel metal3 s 200 35988 800 36228 6 active
port 1 nsew signal input
rlabel metal2 s 11582 200 11694 800 6 io_in[0]
port 2 nsew signal input
rlabel metal2 s 18666 41200 18778 41800 6 io_in[10]
port 3 nsew signal input
rlabel metal3 s 200 38708 800 38948 6 io_in[11]
port 4 nsew signal input
rlabel metal3 s 35200 35988 35800 36228 6 io_in[12]
port 5 nsew signal input
rlabel metal2 s 18022 200 18134 800 6 io_in[13]
port 6 nsew signal input
rlabel metal2 s 11582 41200 11694 41800 6 io_in[14]
port 7 nsew signal input
rlabel metal3 s 35200 37348 35800 37588 6 io_in[15]
port 8 nsew signal input
rlabel metal3 s 35200 6068 35800 6308 6 io_in[16]
port 9 nsew signal input
rlabel metal2 s 5142 41200 5254 41800 6 io_in[17]
port 10 nsew signal input
rlabel metal2 s 6430 41200 6542 41800 6 io_in[18]
port 11 nsew signal input
rlabel metal2 s 33478 200 33590 800 6 io_in[19]
port 12 nsew signal input
rlabel metal3 s 200 12188 800 12428 6 io_in[1]
port 13 nsew signal input
rlabel metal3 s 200 22388 800 22628 6 io_in[20]
port 14 nsew signal input
rlabel metal3 s 200 14908 800 15148 6 io_in[21]
port 15 nsew signal input
rlabel metal3 s 35200 15588 35800 15828 6 io_in[22]
port 16 nsew signal input
rlabel metal2 s 4498 41200 4610 41800 6 io_in[23]
port 17 nsew signal input
rlabel metal2 s 1922 41200 2034 41800 6 io_in[24]
port 18 nsew signal input
rlabel metal2 s 28970 200 29082 800 6 io_in[25]
port 19 nsew signal input
rlabel metal2 s 28326 200 28438 800 6 io_in[26]
port 20 nsew signal input
rlabel metal3 s 35200 11508 35800 11748 6 io_in[27]
port 21 nsew signal input
rlabel metal2 s 25750 200 25862 800 6 io_in[28]
port 22 nsew signal input
rlabel metal2 s 35410 41200 35522 41800 6 io_in[29]
port 23 nsew signal input
rlabel metal2 s 12870 200 12982 800 6 io_in[2]
port 24 nsew signal input
rlabel metal3 s 35200 18308 35800 18548 6 io_in[30]
port 25 nsew signal input
rlabel metal3 s 200 34628 800 34868 6 io_in[31]
port 26 nsew signal input
rlabel metal2 s 23818 200 23930 800 6 io_in[32]
port 27 nsew signal input
rlabel metal3 s 200 20348 800 20588 6 io_in[33]
port 28 nsew signal input
rlabel metal2 s 26394 41200 26506 41800 6 io_in[34]
port 29 nsew signal input
rlabel metal2 s 30902 41200 31014 41800 6 io_in[35]
port 30 nsew signal input
rlabel metal3 s 35200 27148 35800 27388 6 io_in[36]
port 31 nsew signal input
rlabel metal2 s 31546 41200 31658 41800 6 io_in[37]
port 32 nsew signal input
rlabel metal2 s 19310 41200 19422 41800 6 io_in[3]
port 33 nsew signal input
rlabel metal3 s 35200 26468 35800 26708 6 io_in[4]
port 34 nsew signal input
rlabel metal3 s 35200 40068 35800 40308 6 io_in[5]
port 35 nsew signal input
rlabel metal3 s 200 23748 800 23988 6 io_in[6]
port 36 nsew signal input
rlabel metal3 s 200 16268 800 16508 6 io_in[7]
port 37 nsew signal input
rlabel metal3 s 35200 29188 35800 29428 6 io_in[8]
port 38 nsew signal input
rlabel metal2 s 3210 41200 3322 41800 6 io_in[9]
port 39 nsew signal input
rlabel metal2 s 20598 200 20710 800 6 io_oeb[0]
port 40 nsew signal output
rlabel metal3 s 200 13548 800 13788 6 io_oeb[10]
port 41 nsew signal output
rlabel metal3 s 35200 25108 35800 25348 6 io_oeb[11]
port 42 nsew signal output
rlabel metal3 s 35200 14228 35800 14468 6 io_oeb[12]
port 43 nsew signal output
rlabel metal3 s 35200 13548 35800 13788 6 io_oeb[13]
port 44 nsew signal output
rlabel metal3 s 200 3348 800 3588 6 io_oeb[14]
port 45 nsew signal output
rlabel metal2 s 7718 41200 7830 41800 6 io_oeb[15]
port 46 nsew signal output
rlabel metal3 s 35200 4708 35800 4948 6 io_oeb[16]
port 47 nsew signal output
rlabel metal2 s 10294 200 10406 800 6 io_oeb[17]
port 48 nsew signal output
rlabel metal2 s 25106 41200 25218 41800 6 io_oeb[18]
port 49 nsew signal output
rlabel metal2 s 8362 41200 8474 41800 6 io_oeb[19]
port 50 nsew signal output
rlabel metal2 s 30258 200 30370 800 6 io_oeb[1]
port 51 nsew signal output
rlabel metal3 s 35200 19668 35800 19908 6 io_oeb[20]
port 52 nsew signal output
rlabel metal3 s 200 40748 800 40988 6 io_oeb[21]
port 53 nsew signal output
rlabel metal2 s 3854 200 3966 800 6 io_oeb[22]
port 54 nsew signal output
rlabel metal2 s 16090 41200 16202 41800 6 io_oeb[23]
port 55 nsew signal output
rlabel metal2 s 17378 41200 17490 41800 6 io_oeb[24]
port 56 nsew signal output
rlabel metal3 s 35200 628 35800 868 6 io_oeb[25]
port 57 nsew signal output
rlabel metal3 s 35200 33268 35800 33508 6 io_oeb[26]
port 58 nsew signal output
rlabel metal2 s 19954 41200 20066 41800 6 io_oeb[27]
port 59 nsew signal output
rlabel metal2 s 32834 200 32946 800 6 io_oeb[28]
port 60 nsew signal output
rlabel metal3 s 35200 27828 35800 28068 6 io_oeb[29]
port 61 nsew signal output
rlabel metal2 s 28970 41200 29082 41800 6 io_oeb[2]
port 62 nsew signal output
rlabel metal3 s 200 41428 800 41668 6 io_oeb[30]
port 63 nsew signal output
rlabel metal2 s 32190 200 32302 800 6 io_oeb[31]
port 64 nsew signal output
rlabel metal3 s 200 18988 800 19228 6 io_oeb[32]
port 65 nsew signal output
rlabel metal3 s 35200 1988 35800 2228 6 io_oeb[33]
port 66 nsew signal output
rlabel metal2 s 5786 41200 5898 41800 6 io_oeb[34]
port 67 nsew signal output
rlabel metal3 s 200 16948 800 17188 6 io_oeb[35]
port 68 nsew signal output
rlabel metal3 s 200 8788 800 9028 6 io_oeb[36]
port 69 nsew signal output
rlabel metal3 s 200 14228 800 14468 6 io_oeb[37]
port 70 nsew signal output
rlabel metal2 s 19954 200 20066 800 6 io_oeb[3]
port 71 nsew signal output
rlabel metal3 s 35200 3348 35800 3588 6 io_oeb[4]
port 72 nsew signal output
rlabel metal3 s 200 25108 800 25348 6 io_oeb[5]
port 73 nsew signal output
rlabel metal3 s 35200 16948 35800 17188 6 io_oeb[6]
port 74 nsew signal output
rlabel metal2 s 7074 41200 7186 41800 6 io_oeb[7]
port 75 nsew signal output
rlabel metal2 s 3210 200 3322 800 6 io_oeb[8]
port 76 nsew signal output
rlabel metal2 s 8362 200 8474 800 6 io_oeb[9]
port 77 nsew signal output
rlabel metal3 s 35200 39388 35800 39628 6 io_out[0]
port 78 nsew signal output
rlabel metal3 s 35200 24428 35800 24668 6 io_out[10]
port 79 nsew signal output
rlabel metal3 s 200 1988 800 2228 6 io_out[11]
port 80 nsew signal output
rlabel metal3 s 200 5388 800 5628 6 io_out[12]
port 81 nsew signal output
rlabel metal2 s 30902 200 31014 800 6 io_out[13]
port 82 nsew signal output
rlabel metal3 s 35200 33948 35800 34188 6 io_out[14]
port 83 nsew signal output
rlabel metal3 s 200 31908 800 32148 6 io_out[15]
port 84 nsew signal output
rlabel metal3 s 35200 23748 35800 23988 6 io_out[16]
port 85 nsew signal output
rlabel metal2 s 32834 41200 32946 41800 6 io_out[17]
port 86 nsew signal output
rlabel metal3 s 35200 -52 35800 188 6 io_out[18]
port 87 nsew signal output
rlabel metal3 s 200 18308 800 18548 6 io_out[19]
port 88 nsew signal output
rlabel metal2 s 22530 41200 22642 41800 6 io_out[1]
port 89 nsew signal output
rlabel metal2 s 28326 41200 28438 41800 6 io_out[20]
port 90 nsew signal output
rlabel metal3 s 200 31228 800 31468 6 io_out[21]
port 91 nsew signal output
rlabel metal2 s 24462 200 24574 800 6 io_out[22]
port 92 nsew signal output
rlabel metal3 s 35200 20348 35800 20588 6 io_out[23]
port 93 nsew signal output
rlabel metal2 s 21242 200 21354 800 6 io_out[24]
port 94 nsew signal output
rlabel metal2 s 25750 41200 25862 41800 6 io_out[25]
port 95 nsew signal output
rlabel metal3 s 200 4028 800 4268 6 io_out[26]
port 96 nsew signal output
rlabel metal2 s 27038 41200 27150 41800 6 io_out[27]
port 97 nsew signal output
rlabel metal2 s 13514 200 13626 800 6 io_out[28]
port 98 nsew signal output
rlabel metal3 s 35200 4028 35800 4268 6 io_out[29]
port 99 nsew signal output
rlabel metal2 s 5142 200 5254 800 6 io_out[2]
port 100 nsew signal output
rlabel metal3 s 200 4708 800 4948 6 io_out[30]
port 101 nsew signal output
rlabel metal3 s 200 10828 800 11068 6 io_out[31]
port 102 nsew signal output
rlabel metal3 s 200 36668 800 36908 6 io_out[32]
port 103 nsew signal output
rlabel metal3 s 35200 8788 35800 9028 6 io_out[33]
port 104 nsew signal output
rlabel metal3 s 35200 34628 35800 34868 6 io_out[34]
port 105 nsew signal output
rlabel metal3 s 35200 32588 35800 32828 6 io_out[35]
port 106 nsew signal output
rlabel metal2 s 9006 41200 9118 41800 6 io_out[36]
port 107 nsew signal output
rlabel metal3 s 35200 38028 35800 38268 6 io_out[37]
port 108 nsew signal output
rlabel metal3 s 200 33948 800 34188 6 io_out[3]
port 109 nsew signal output
rlabel metal3 s 35200 25788 35800 26028 6 io_out[4]
port 110 nsew signal output
rlabel metal2 s 14802 41200 14914 41800 6 io_out[5]
port 111 nsew signal output
rlabel metal2 s 34122 41200 34234 41800 6 io_out[6]
port 112 nsew signal output
rlabel metal3 s 200 15588 800 15828 6 io_out[7]
port 113 nsew signal output
rlabel metal2 s 14802 200 14914 800 6 io_out[8]
port 114 nsew signal output
rlabel metal3 s 200 11508 800 11748 6 io_out[9]
port 115 nsew signal output
rlabel metal3 s 35200 9468 35800 9708 6 la1_data_in[0]
port 116 nsew signal input
rlabel metal2 s 16734 200 16846 800 6 la1_data_in[10]
port 117 nsew signal input
rlabel metal3 s 35200 7428 35800 7668 6 la1_data_in[11]
port 118 nsew signal input
rlabel metal3 s 200 29188 800 29428 6 la1_data_in[12]
port 119 nsew signal input
rlabel metal2 s 26394 200 26506 800 6 la1_data_in[13]
port 120 nsew signal input
rlabel metal3 s 200 10148 800 10388 6 la1_data_in[14]
port 121 nsew signal input
rlabel metal2 s 9650 41200 9762 41800 6 la1_data_in[15]
port 122 nsew signal input
rlabel metal2 s 21242 41200 21354 41800 6 la1_data_in[16]
port 123 nsew signal input
rlabel metal2 s 15446 41200 15558 41800 6 la1_data_in[17]
port 124 nsew signal input
rlabel metal2 s 34122 200 34234 800 6 la1_data_in[18]
port 125 nsew signal input
rlabel metal2 s 10938 41200 11050 41800 6 la1_data_in[19]
port 126 nsew signal input
rlabel metal2 s 15446 200 15558 800 6 la1_data_in[1]
port 127 nsew signal input
rlabel metal3 s 200 28508 800 28748 6 la1_data_in[20]
port 128 nsew signal input
rlabel metal2 s 34766 41200 34878 41800 6 la1_data_in[21]
port 129 nsew signal input
rlabel metal3 s 35200 10148 35800 10388 6 la1_data_in[22]
port 130 nsew signal input
rlabel metal3 s 200 628 800 868 6 la1_data_in[23]
port 131 nsew signal input
rlabel metal2 s 10938 200 11050 800 6 la1_data_in[24]
port 132 nsew signal input
rlabel metal3 s 200 29868 800 30108 6 la1_data_in[25]
port 133 nsew signal input
rlabel metal3 s 35200 5388 35800 5628 6 la1_data_in[26]
port 134 nsew signal input
rlabel metal2 s 22530 200 22642 800 6 la1_data_in[27]
port 135 nsew signal input
rlabel metal3 s 200 25788 800 26028 6 la1_data_in[28]
port 136 nsew signal input
rlabel metal3 s 200 39388 800 39628 6 la1_data_in[29]
port 137 nsew signal input
rlabel metal2 s 9006 200 9118 800 6 la1_data_in[2]
port 138 nsew signal input
rlabel metal2 s 1278 200 1390 800 6 la1_data_in[30]
port 139 nsew signal input
rlabel metal2 s 29614 200 29726 800 6 la1_data_in[31]
port 140 nsew signal input
rlabel metal3 s 200 24428 800 24668 6 la1_data_in[3]
port 141 nsew signal input
rlabel metal2 s 30258 41200 30370 41800 6 la1_data_in[4]
port 142 nsew signal input
rlabel metal3 s 35200 22388 35800 22628 6 la1_data_in[5]
port 143 nsew signal input
rlabel metal2 s 12226 41200 12338 41800 6 la1_data_in[6]
port 144 nsew signal input
rlabel metal3 s 200 17628 800 17868 6 la1_data_in[7]
port 145 nsew signal input
rlabel metal2 s 12870 41200 12982 41800 6 la1_data_in[8]
port 146 nsew signal input
rlabel metal3 s 200 27148 800 27388 6 la1_data_in[9]
port 147 nsew signal input
rlabel metal2 s 6430 200 6542 800 6 la1_data_out[0]
port 148 nsew signal output
rlabel metal3 s 35200 12188 35800 12428 6 la1_data_out[10]
port 149 nsew signal output
rlabel metal2 s 17378 200 17490 800 6 la1_data_out[11]
port 150 nsew signal output
rlabel metal3 s 35200 38708 35800 38948 6 la1_data_out[12]
port 151 nsew signal output
rlabel metal2 s 634 41200 746 41800 6 la1_data_out[13]
port 152 nsew signal output
rlabel metal2 s 18022 41200 18134 41800 6 la1_data_out[14]
port 153 nsew signal output
rlabel metal3 s 200 1308 800 1548 6 la1_data_out[15]
port 154 nsew signal output
rlabel metal3 s 35200 16268 35800 16508 6 la1_data_out[16]
port 155 nsew signal output
rlabel metal3 s 35200 31228 35800 31468 6 la1_data_out[17]
port 156 nsew signal output
rlabel metal2 s 1278 41200 1390 41800 6 la1_data_out[18]
port 157 nsew signal output
rlabel metal3 s 35200 23068 35800 23308 6 la1_data_out[19]
port 158 nsew signal output
rlabel metal3 s 200 35308 800 35548 6 la1_data_out[1]
port 159 nsew signal output
rlabel metal3 s 200 8108 800 8348 6 la1_data_out[20]
port 160 nsew signal output
rlabel metal3 s 35200 36668 35800 36908 6 la1_data_out[21]
port 161 nsew signal output
rlabel metal2 s 20598 41200 20710 41800 6 la1_data_out[22]
port 162 nsew signal output
rlabel metal2 s 9650 200 9762 800 6 la1_data_out[23]
port 163 nsew signal output
rlabel metal3 s 35200 17628 35800 17868 6 la1_data_out[24]
port 164 nsew signal output
rlabel metal3 s 200 2668 800 2908 6 la1_data_out[25]
port 165 nsew signal output
rlabel metal3 s 35200 6748 35800 6988 6 la1_data_out[26]
port 166 nsew signal output
rlabel metal3 s 200 37348 800 37588 6 la1_data_out[27]
port 167 nsew signal output
rlabel metal2 s 34766 200 34878 800 6 la1_data_out[28]
port 168 nsew signal output
rlabel metal2 s 4498 200 4610 800 6 la1_data_out[29]
port 169 nsew signal output
rlabel metal2 s 16090 200 16202 800 6 la1_data_out[2]
port 170 nsew signal output
rlabel metal3 s 35200 12868 35800 13108 6 la1_data_out[30]
port 171 nsew signal output
rlabel metal3 s 35200 40748 35800 40988 6 la1_data_out[31]
port 172 nsew signal output
rlabel metal3 s 200 7428 800 7668 6 la1_data_out[3]
port 173 nsew signal output
rlabel metal2 s 35410 200 35522 800 6 la1_data_out[4]
port 174 nsew signal output
rlabel metal2 s 2566 200 2678 800 6 la1_data_out[5]
port 175 nsew signal output
rlabel metal3 s 35200 18988 35800 19228 6 la1_data_out[6]
port 176 nsew signal output
rlabel metal2 s 634 200 746 800 6 la1_data_out[7]
port 177 nsew signal output
rlabel metal3 s 35200 31908 35800 32148 6 la1_data_out[8]
port 178 nsew signal output
rlabel metal2 s 33478 41200 33590 41800 6 la1_data_out[9]
port 179 nsew signal output
rlabel metal3 s 35200 2668 35800 2908 6 la1_oenb[0]
port 180 nsew signal input
rlabel metal2 s 32190 41200 32302 41800 6 la1_oenb[10]
port 181 nsew signal input
rlabel metal3 s 200 21708 800 21948 6 la1_oenb[11]
port 182 nsew signal input
rlabel metal3 s 200 23068 800 23308 6 la1_oenb[12]
port 183 nsew signal input
rlabel metal2 s 23174 200 23286 800 6 la1_oenb[13]
port 184 nsew signal input
rlabel metal2 s -10 200 102 800 6 la1_oenb[14]
port 185 nsew signal input
rlabel metal2 s 27682 200 27794 800 6 la1_oenb[15]
port 186 nsew signal input
rlabel metal3 s 200 27828 800 28068 6 la1_oenb[16]
port 187 nsew signal input
rlabel metal2 s -10 41200 102 41800 6 la1_oenb[17]
port 188 nsew signal input
rlabel metal2 s 14158 41200 14270 41800 6 la1_oenb[18]
port 189 nsew signal input
rlabel metal3 s 200 21028 800 21268 6 la1_oenb[19]
port 190 nsew signal input
rlabel metal2 s 7074 200 7186 800 6 la1_oenb[1]
port 191 nsew signal input
rlabel metal2 s 1922 200 2034 800 6 la1_oenb[20]
port 192 nsew signal input
rlabel metal2 s 21886 41200 21998 41800 6 la1_oenb[21]
port 193 nsew signal input
rlabel metal2 s 13514 41200 13626 41800 6 la1_oenb[22]
port 194 nsew signal input
rlabel metal2 s 19310 200 19422 800 6 la1_oenb[23]
port 195 nsew signal input
rlabel metal2 s 27682 41200 27794 41800 6 la1_oenb[24]
port 196 nsew signal input
rlabel metal3 s 35200 10828 35800 11068 6 la1_oenb[25]
port 197 nsew signal input
rlabel metal3 s 200 30548 800 30788 6 la1_oenb[26]
port 198 nsew signal input
rlabel metal3 s 35200 30548 35800 30788 6 la1_oenb[27]
port 199 nsew signal input
rlabel metal2 s 7718 200 7830 800 6 la1_oenb[28]
port 200 nsew signal input
rlabel metal2 s 14158 200 14270 800 6 la1_oenb[29]
port 201 nsew signal input
rlabel metal3 s 200 6748 800 6988 6 la1_oenb[2]
port 202 nsew signal input
rlabel metal3 s 35200 29868 35800 30108 6 la1_oenb[30]
port 203 nsew signal input
rlabel metal2 s 21886 200 21998 800 6 la1_oenb[31]
port 204 nsew signal input
rlabel metal2 s 24462 41200 24574 41800 6 la1_oenb[3]
port 205 nsew signal input
rlabel metal2 s 23818 41200 23930 41800 6 la1_oenb[4]
port 206 nsew signal input
rlabel metal3 s 200 38028 800 38268 6 la1_oenb[5]
port 207 nsew signal input
rlabel metal2 s 2566 41200 2678 41800 6 la1_oenb[6]
port 208 nsew signal input
rlabel metal2 s 27038 200 27150 800 6 la1_oenb[7]
port 209 nsew signal input
rlabel metal3 s 200 9468 800 9708 6 la1_oenb[8]
port 210 nsew signal input
rlabel metal3 s 200 32588 800 32828 6 la1_oenb[9]
port 211 nsew signal input
rlabel metal4 s 5164 2128 5484 39760 6 vccd1
port 212 nsew power bidirectional
rlabel metal4 s 13605 2128 13925 39760 6 vccd1
port 212 nsew power bidirectional
rlabel metal4 s 22046 2128 22366 39760 6 vccd1
port 212 nsew power bidirectional
rlabel metal4 s 30487 2128 30807 39760 6 vccd1
port 212 nsew power bidirectional
rlabel metal4 s 9384 2128 9704 39760 6 vssd1
port 213 nsew ground bidirectional
rlabel metal4 s 17825 2128 18145 39760 6 vssd1
port 213 nsew ground bidirectional
rlabel metal4 s 26266 2128 26586 39760 6 vssd1
port 213 nsew ground bidirectional
rlabel metal4 s 34707 2128 35027 39760 6 vssd1
port 213 nsew ground bidirectional
rlabel metal3 s 35200 21028 35800 21268 6 wb_clk_i
port 214 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 36000 42000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2814108
string GDS_FILE /openlane/designs/wrapped_rgb_mixer/runs/RUN_2022.12.13_09.51.10/results/signoff/wrapped_rgb_mixer.magic.gds
string GDS_START 293796
<< end >>

