VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_rgb_mixer
  CLASS BLOCK ;
  FOREIGN wrapped_rgb_mixer ;
  ORIGIN 0.000 0.000 ;
  SIZE 130.000 BY 210.000 ;
  PIN active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.920 4.000 181.520 ;
    END
  END active
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 4.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 206.000 68.450 210.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.880 4.000 196.480 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 178.200 130.000 178.800 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 4.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 206.000 42.690 210.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 186.360 130.000 186.960 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 31.320 130.000 31.920 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 206.000 19.690 210.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 206.000 24.290 210.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 4.000 64.560 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 4.000 113.520 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 76.200 130.000 76.800 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.650 206.000 16.930 210.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 206.000 9.570 210.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.970 0.000 105.250 4.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 4.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 57.160 130.000 57.760 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 0.000 92.370 4.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 206.000 129.170 210.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.090 0.000 46.370 4.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 91.160 130.000 91.760 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 4.000 174.720 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.570 0.000 86.850 4.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 206.000 96.050 210.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.410 206.000 111.690 210.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 137.400 130.000 138.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 206.000 114.450 210.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 206.000 70.290 210.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 133.320 130.000 133.920 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 201.320 130.000 201.920 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 4.000 121.680 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 144.200 130.000 144.800 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 206.000 14.170 210.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 0.000 73.970 4.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 125.160 130.000 125.760 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 72.120 130.000 72.720 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 69.400 130.000 70.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 4.000 18.320 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 206.000 29.810 210.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 23.160 130.000 23.760 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 0.000 38.090 4.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 206.000 91.450 210.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 206.000 32.570 210.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 99.320 130.000 99.920 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 0.000 15.090 4.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 206.000 60.170 210.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 206.000 62.930 210.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 4.120 130.000 4.720 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 167.320 130.000 167.920 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 206.000 73.050 210.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 0.000 118.130 4.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 140.120 130.000 140.720 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 206.000 106.170 210.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.120 4.000 208.720 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 0.000 115.370 4.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 4.000 98.560 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 8.200 130.000 8.800 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 206.000 22.450 210.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 4.000 87.680 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 4.000 45.520 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 4.000 71.360 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 16.360 130.000 16.960 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 4.000 128.480 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 84.360 130.000 84.960 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 206.000 27.050 210.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 0.000 12.330 4.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 0.000 30.730 4.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 197.240 130.000 197.840 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 121.080 130.000 121.680 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 4.000 30.560 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 4.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 171.400 130.000 172.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 4.000 162.480 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 118.360 130.000 118.960 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 206.000 119.050 210.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 0.040 130.000 0.640 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 4.000 94.480 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 206.000 83.170 210.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 206.000 104.330 210.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.800 4.000 158.400 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 0.000 89.610 4.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 103.400 130.000 104.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 0.000 76.730 4.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 206.000 94.210 210.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 4.000 22.400 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 206.000 98.810 210.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.930 0.000 48.210 4.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 19.080 130.000 19.680 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.330 0.000 20.610 4.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 4.000 56.400 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.000 4.000 185.600 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 42.200 130.000 42.800 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 174.120 130.000 174.720 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 163.240 130.000 163.840 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 206.000 35.330 210.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 190.440 130.000 191.040 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 129.240 130.000 129.840 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 206.000 55.570 210.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 206.000 124.570 210.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 4.000 79.520 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.450 0.000 53.730 4.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 4.000 60.480 ;
    END
  END io_out[9]
  PIN la1_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 46.280 130.000 46.880 ;
    END
  END la1_data_in[0]
  PIN la1_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 4.000 ;
    END
  END la1_data_in[10]
  PIN la1_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 38.120 130.000 38.720 ;
    END
  END la1_data_in[11]
  PIN la1_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.920 4.000 147.520 ;
    END
  END la1_data_in[12]
  PIN la1_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 0.000 94.210 4.000 ;
    END
  END la1_data_in[13]
  PIN la1_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 4.000 52.320 ;
    END
  END la1_data_in[14]
  PIN la1_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 206.000 37.170 210.000 ;
    END
  END la1_data_in[15]
  PIN la1_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 206.000 78.570 210.000 ;
    END
  END la1_data_in[16]
  PIN la1_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 206.000 58.330 210.000 ;
    END
  END la1_data_in[17]
  PIN la1_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END la1_data_in[18]
  PIN la1_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 206.000 39.930 210.000 ;
    END
  END la1_data_in[19]
  PIN la1_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 0.000 56.490 4.000 ;
    END
  END la1_data_in[1]
  PIN la1_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END la1_data_in[20]
  PIN la1_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.050 206.000 127.330 210.000 ;
    END
  END la1_data_in[21]
  PIN la1_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 50.360 130.000 50.960 ;
    END
  END la1_data_in[22]
  PIN la1_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 4.000 3.360 ;
    END
  END la1_data_in[23]
  PIN la1_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 4.000 ;
    END
  END la1_data_in[24]
  PIN la1_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 4.000 151.600 ;
    END
  END la1_data_in[25]
  PIN la1_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 27.240 130.000 27.840 ;
    END
  END la1_data_in[26]
  PIN la1_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 0.000 82.250 4.000 ;
    END
  END la1_data_in[27]
  PIN la1_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 4.000 132.560 ;
    END
  END la1_data_in[28]
  PIN la1_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.960 4.000 200.560 ;
    END
  END la1_data_in[29]
  PIN la1_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 4.000 ;
    END
  END la1_data_in[2]
  PIN la1_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 4.000 ;
    END
  END la1_data_in[30]
  PIN la1_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 0.000 107.090 4.000 ;
    END
  END la1_data_in[31]
  PIN la1_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.800 4.000 124.400 ;
    END
  END la1_data_in[3]
  PIN la1_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.650 206.000 108.930 210.000 ;
    END
  END la1_data_in[4]
  PIN la1_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 110.200 130.000 110.800 ;
    END
  END la1_data_in[5]
  PIN la1_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 206.000 45.450 210.000 ;
    END
  END la1_data_in[6]
  PIN la1_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 4.000 90.400 ;
    END
  END la1_data_in[7]
  PIN la1_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 206.000 47.290 210.000 ;
    END
  END la1_data_in[8]
  PIN la1_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END la1_data_in[9]
  PIN la1_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 0.000 23.370 4.000 ;
    END
  END la1_data_out[0]
  PIN la1_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 61.240 130.000 61.840 ;
    END
  END la1_data_out[10]
  PIN la1_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.570 0.000 63.850 4.000 ;
    END
  END la1_data_out[11]
  PIN la1_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 193.160 130.000 193.760 ;
    END
  END la1_data_out[12]
  PIN la1_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.770 206.000 4.050 210.000 ;
    END
  END la1_data_out[13]
  PIN la1_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 206.000 65.690 210.000 ;
    END
  END la1_data_out[14]
  PIN la1_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END la1_data_out[15]
  PIN la1_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 80.280 130.000 80.880 ;
    END
  END la1_data_out[16]
  PIN la1_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 156.440 130.000 157.040 ;
    END
  END la1_data_out[17]
  PIN la1_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 206.000 6.810 210.000 ;
    END
  END la1_data_out[18]
  PIN la1_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 114.280 130.000 114.880 ;
    END
  END la1_data_out[19]
  PIN la1_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END la1_data_out[1]
  PIN la1_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END la1_data_out[20]
  PIN la1_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 182.280 130.000 182.880 ;
    END
  END la1_data_out[21]
  PIN la1_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.530 206.000 75.810 210.000 ;
    END
  END la1_data_out[22]
  PIN la1_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 4.000 ;
    END
  END la1_data_out[23]
  PIN la1_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 87.080 130.000 87.680 ;
    END
  END la1_data_out[24]
  PIN la1_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 4.000 15.600 ;
    END
  END la1_data_out[25]
  PIN la1_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 34.040 130.000 34.640 ;
    END
  END la1_data_out[26]
  PIN la1_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.080 4.000 189.680 ;
    END
  END la1_data_out[27]
  PIN la1_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.210 0.000 125.490 4.000 ;
    END
  END la1_data_out[28]
  PIN la1_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 0.000 17.850 4.000 ;
    END
  END la1_data_out[29]
  PIN la1_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 4.000 ;
    END
  END la1_data_out[2]
  PIN la1_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 65.320 130.000 65.920 ;
    END
  END la1_data_out[30]
  PIN la1_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 205.400 130.000 206.000 ;
    END
  END la1_data_out[31]
  PIN la1_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 4.000 37.360 ;
    END
  END la1_data_out[3]
  PIN la1_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.970 0.000 128.250 4.000 ;
    END
  END la1_data_out[4]
  PIN la1_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 0.000 10.490 4.000 ;
    END
  END la1_data_out[5]
  PIN la1_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 95.240 130.000 95.840 ;
    END
  END la1_data_out[6]
  PIN la1_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 0.000 2.210 4.000 ;
    END
  END la1_data_out[7]
  PIN la1_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 159.160 130.000 159.760 ;
    END
  END la1_data_out[8]
  PIN la1_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.530 206.000 121.810 210.000 ;
    END
  END la1_data_out[9]
  PIN la1_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 12.280 130.000 12.880 ;
    END
  END la1_oenb[0]
  PIN la1_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930 206.000 117.210 210.000 ;
    END
  END la1_oenb[10]
  PIN la1_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END la1_oenb[11]
  PIN la1_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 4.000 117.600 ;
    END
  END la1_oenb[12]
  PIN la1_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END la1_oenb[13]
  PIN la1_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END la1_oenb[14]
  PIN la1_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.450 0.000 99.730 4.000 ;
    END
  END la1_oenb[15]
  PIN la1_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 4.000 139.360 ;
    END
  END la1_oenb[16]
  PIN la1_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.010 206.000 1.290 210.000 ;
    END
  END la1_oenb[17]
  PIN la1_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 206.000 52.810 210.000 ;
    END
  END la1_oenb[18]
  PIN la1_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 4.000 105.360 ;
    END
  END la1_oenb[19]
  PIN la1_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 4.000 ;
    END
  END la1_oenb[1]
  PIN la1_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 4.000 ;
    END
  END la1_oenb[20]
  PIN la1_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 206.000 81.330 210.000 ;
    END
  END la1_oenb[21]
  PIN la1_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 206.000 50.050 210.000 ;
    END
  END la1_oenb[22]
  PIN la1_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END la1_oenb[23]
  PIN la1_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 206.000 101.570 210.000 ;
    END
  END la1_oenb[24]
  PIN la1_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 53.080 130.000 53.680 ;
    END
  END la1_oenb[25]
  PIN la1_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.080 4.000 155.680 ;
    END
  END la1_oenb[26]
  PIN la1_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 152.360 130.000 152.960 ;
    END
  END la1_oenb[27]
  PIN la1_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 4.000 ;
    END
  END la1_oenb[28]
  PIN la1_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 0.000 50.970 4.000 ;
    END
  END la1_oenb[29]
  PIN la1_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END la1_oenb[2]
  PIN la1_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 148.280 130.000 148.880 ;
    END
  END la1_oenb[30]
  PIN la1_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 4.000 ;
    END
  END la1_oenb[31]
  PIN la1_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 206.000 88.690 210.000 ;
    END
  END la1_oenb[3]
  PIN la1_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 206.000 85.930 210.000 ;
    END
  END la1_oenb[4]
  PIN la1_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.800 4.000 192.400 ;
    END
  END la1_oenb[5]
  PIN la1_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.130 206.000 11.410 210.000 ;
    END
  END la1_oenb[6]
  PIN la1_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END la1_oenb[7]
  PIN la1_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 4.000 49.600 ;
    END
  END la1_oenb[8]
  PIN la1_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.960 4.000 166.560 ;
    END
  END la1_oenb[9]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 24.545 10.640 26.145 198.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 64.195 10.640 65.795 198.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 103.850 10.640 105.450 198.800 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 44.370 10.640 45.970 198.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 84.025 10.640 85.625 198.800 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126.000 106.120 130.000 106.720 ;
    END
  END wb_clk_i
  OBS
      LAYER li1 ;
        RECT 5.520 0.425 129.575 205.615 ;
      LAYER met1 ;
        RECT 1.910 0.380 129.635 205.660 ;
      LAYER met2 ;
        RECT 1.940 205.720 3.490 208.605 ;
        RECT 4.330 205.720 6.250 208.605 ;
        RECT 7.090 205.720 9.010 208.605 ;
        RECT 9.850 205.720 10.850 208.605 ;
        RECT 11.690 205.720 13.610 208.605 ;
        RECT 14.450 205.720 16.370 208.605 ;
        RECT 17.210 205.720 19.130 208.605 ;
        RECT 19.970 205.720 21.890 208.605 ;
        RECT 22.730 205.720 23.730 208.605 ;
        RECT 24.570 205.720 26.490 208.605 ;
        RECT 27.330 205.720 29.250 208.605 ;
        RECT 30.090 205.720 32.010 208.605 ;
        RECT 32.850 205.720 34.770 208.605 ;
        RECT 35.610 205.720 36.610 208.605 ;
        RECT 37.450 205.720 39.370 208.605 ;
        RECT 40.210 205.720 42.130 208.605 ;
        RECT 42.970 205.720 44.890 208.605 ;
        RECT 45.730 205.720 46.730 208.605 ;
        RECT 47.570 205.720 49.490 208.605 ;
        RECT 50.330 205.720 52.250 208.605 ;
        RECT 53.090 205.720 55.010 208.605 ;
        RECT 55.850 205.720 57.770 208.605 ;
        RECT 58.610 205.720 59.610 208.605 ;
        RECT 60.450 205.720 62.370 208.605 ;
        RECT 63.210 205.720 65.130 208.605 ;
        RECT 65.970 205.720 67.890 208.605 ;
        RECT 68.730 205.720 69.730 208.605 ;
        RECT 70.570 205.720 72.490 208.605 ;
        RECT 73.330 205.720 75.250 208.605 ;
        RECT 76.090 205.720 78.010 208.605 ;
        RECT 78.850 205.720 80.770 208.605 ;
        RECT 81.610 205.720 82.610 208.605 ;
        RECT 83.450 205.720 85.370 208.605 ;
        RECT 86.210 205.720 88.130 208.605 ;
        RECT 88.970 205.720 90.890 208.605 ;
        RECT 91.730 205.720 93.650 208.605 ;
        RECT 94.490 205.720 95.490 208.605 ;
        RECT 96.330 205.720 98.250 208.605 ;
        RECT 99.090 205.720 101.010 208.605 ;
        RECT 101.850 205.720 103.770 208.605 ;
        RECT 104.610 205.720 105.610 208.605 ;
        RECT 106.450 205.720 108.370 208.605 ;
        RECT 109.210 205.720 111.130 208.605 ;
        RECT 111.970 205.720 113.890 208.605 ;
        RECT 114.730 205.720 116.650 208.605 ;
        RECT 117.490 205.720 118.490 208.605 ;
        RECT 119.330 205.720 121.250 208.605 ;
        RECT 122.090 205.720 124.010 208.605 ;
        RECT 124.850 205.720 126.770 208.605 ;
        RECT 127.610 205.720 128.610 208.605 ;
        RECT 1.940 4.280 128.710 205.720 ;
        RECT 2.490 0.155 4.410 4.280 ;
        RECT 5.250 0.155 7.170 4.280 ;
        RECT 8.010 0.155 9.930 4.280 ;
        RECT 10.770 0.155 11.770 4.280 ;
        RECT 12.610 0.155 14.530 4.280 ;
        RECT 15.370 0.155 17.290 4.280 ;
        RECT 18.130 0.155 20.050 4.280 ;
        RECT 20.890 0.155 22.810 4.280 ;
        RECT 23.650 0.155 24.650 4.280 ;
        RECT 25.490 0.155 27.410 4.280 ;
        RECT 28.250 0.155 30.170 4.280 ;
        RECT 31.010 0.155 32.930 4.280 ;
        RECT 33.770 0.155 34.770 4.280 ;
        RECT 35.610 0.155 37.530 4.280 ;
        RECT 38.370 0.155 40.290 4.280 ;
        RECT 41.130 0.155 43.050 4.280 ;
        RECT 43.890 0.155 45.810 4.280 ;
        RECT 46.650 0.155 47.650 4.280 ;
        RECT 48.490 0.155 50.410 4.280 ;
        RECT 51.250 0.155 53.170 4.280 ;
        RECT 54.010 0.155 55.930 4.280 ;
        RECT 56.770 0.155 58.690 4.280 ;
        RECT 59.530 0.155 60.530 4.280 ;
        RECT 61.370 0.155 63.290 4.280 ;
        RECT 64.130 0.155 66.050 4.280 ;
        RECT 66.890 0.155 68.810 4.280 ;
        RECT 69.650 0.155 70.650 4.280 ;
        RECT 71.490 0.155 73.410 4.280 ;
        RECT 74.250 0.155 76.170 4.280 ;
        RECT 77.010 0.155 78.930 4.280 ;
        RECT 79.770 0.155 81.690 4.280 ;
        RECT 82.530 0.155 83.530 4.280 ;
        RECT 84.370 0.155 86.290 4.280 ;
        RECT 87.130 0.155 89.050 4.280 ;
        RECT 89.890 0.155 91.810 4.280 ;
        RECT 92.650 0.155 93.650 4.280 ;
        RECT 94.490 0.155 96.410 4.280 ;
        RECT 97.250 0.155 99.170 4.280 ;
        RECT 100.010 0.155 101.930 4.280 ;
        RECT 102.770 0.155 104.690 4.280 ;
        RECT 105.530 0.155 106.530 4.280 ;
        RECT 107.370 0.155 109.290 4.280 ;
        RECT 110.130 0.155 112.050 4.280 ;
        RECT 112.890 0.155 114.810 4.280 ;
        RECT 115.650 0.155 117.570 4.280 ;
        RECT 118.410 0.155 119.410 4.280 ;
        RECT 120.250 0.155 122.170 4.280 ;
        RECT 123.010 0.155 124.930 4.280 ;
        RECT 125.770 0.155 127.690 4.280 ;
        RECT 128.530 0.155 128.710 4.280 ;
      LAYER met3 ;
        RECT 4.400 207.720 128.735 208.585 ;
        RECT 4.000 206.400 128.735 207.720 ;
        RECT 4.000 205.040 125.600 206.400 ;
        RECT 4.400 205.000 125.600 205.040 ;
        RECT 4.400 203.640 128.735 205.000 ;
        RECT 4.000 202.320 128.735 203.640 ;
        RECT 4.000 200.960 125.600 202.320 ;
        RECT 4.400 200.920 125.600 200.960 ;
        RECT 4.400 199.560 128.735 200.920 ;
        RECT 4.000 198.240 128.735 199.560 ;
        RECT 4.000 196.880 125.600 198.240 ;
        RECT 4.400 196.840 125.600 196.880 ;
        RECT 4.400 195.480 128.735 196.840 ;
        RECT 4.000 194.160 128.735 195.480 ;
        RECT 4.000 192.800 125.600 194.160 ;
        RECT 4.400 192.760 125.600 192.800 ;
        RECT 4.400 191.440 128.735 192.760 ;
        RECT 4.400 191.400 125.600 191.440 ;
        RECT 4.000 190.080 125.600 191.400 ;
        RECT 4.400 190.040 125.600 190.080 ;
        RECT 4.400 188.680 128.735 190.040 ;
        RECT 4.000 187.360 128.735 188.680 ;
        RECT 4.000 186.000 125.600 187.360 ;
        RECT 4.400 185.960 125.600 186.000 ;
        RECT 4.400 184.600 128.735 185.960 ;
        RECT 4.000 183.280 128.735 184.600 ;
        RECT 4.000 181.920 125.600 183.280 ;
        RECT 4.400 181.880 125.600 181.920 ;
        RECT 4.400 180.520 128.735 181.880 ;
        RECT 4.000 179.200 128.735 180.520 ;
        RECT 4.000 177.840 125.600 179.200 ;
        RECT 4.400 177.800 125.600 177.840 ;
        RECT 4.400 176.440 128.735 177.800 ;
        RECT 4.000 175.120 128.735 176.440 ;
        RECT 4.400 173.720 125.600 175.120 ;
        RECT 4.000 172.400 128.735 173.720 ;
        RECT 4.000 171.040 125.600 172.400 ;
        RECT 4.400 171.000 125.600 171.040 ;
        RECT 4.400 169.640 128.735 171.000 ;
        RECT 4.000 168.320 128.735 169.640 ;
        RECT 4.000 166.960 125.600 168.320 ;
        RECT 4.400 166.920 125.600 166.960 ;
        RECT 4.400 165.560 128.735 166.920 ;
        RECT 4.000 164.240 128.735 165.560 ;
        RECT 4.000 162.880 125.600 164.240 ;
        RECT 4.400 162.840 125.600 162.880 ;
        RECT 4.400 161.480 128.735 162.840 ;
        RECT 4.000 160.160 128.735 161.480 ;
        RECT 4.000 158.800 125.600 160.160 ;
        RECT 4.400 158.760 125.600 158.800 ;
        RECT 4.400 157.440 128.735 158.760 ;
        RECT 4.400 157.400 125.600 157.440 ;
        RECT 4.000 156.080 125.600 157.400 ;
        RECT 4.400 156.040 125.600 156.080 ;
        RECT 4.400 154.680 128.735 156.040 ;
        RECT 4.000 153.360 128.735 154.680 ;
        RECT 4.000 152.000 125.600 153.360 ;
        RECT 4.400 151.960 125.600 152.000 ;
        RECT 4.400 150.600 128.735 151.960 ;
        RECT 4.000 149.280 128.735 150.600 ;
        RECT 4.000 147.920 125.600 149.280 ;
        RECT 4.400 147.880 125.600 147.920 ;
        RECT 4.400 146.520 128.735 147.880 ;
        RECT 4.000 145.200 128.735 146.520 ;
        RECT 4.000 143.840 125.600 145.200 ;
        RECT 4.400 143.800 125.600 143.840 ;
        RECT 4.400 142.440 128.735 143.800 ;
        RECT 4.000 141.120 128.735 142.440 ;
        RECT 4.000 139.760 125.600 141.120 ;
        RECT 4.400 139.720 125.600 139.760 ;
        RECT 4.400 138.400 128.735 139.720 ;
        RECT 4.400 138.360 125.600 138.400 ;
        RECT 4.000 137.040 125.600 138.360 ;
        RECT 4.400 137.000 125.600 137.040 ;
        RECT 4.400 135.640 128.735 137.000 ;
        RECT 4.000 134.320 128.735 135.640 ;
        RECT 4.000 132.960 125.600 134.320 ;
        RECT 4.400 132.920 125.600 132.960 ;
        RECT 4.400 131.560 128.735 132.920 ;
        RECT 4.000 130.240 128.735 131.560 ;
        RECT 4.000 128.880 125.600 130.240 ;
        RECT 4.400 128.840 125.600 128.880 ;
        RECT 4.400 127.480 128.735 128.840 ;
        RECT 4.000 126.160 128.735 127.480 ;
        RECT 4.000 124.800 125.600 126.160 ;
        RECT 4.400 124.760 125.600 124.800 ;
        RECT 4.400 123.400 128.735 124.760 ;
        RECT 4.000 122.080 128.735 123.400 ;
        RECT 4.400 120.680 125.600 122.080 ;
        RECT 4.000 119.360 128.735 120.680 ;
        RECT 4.000 118.000 125.600 119.360 ;
        RECT 4.400 117.960 125.600 118.000 ;
        RECT 4.400 116.600 128.735 117.960 ;
        RECT 4.000 115.280 128.735 116.600 ;
        RECT 4.000 113.920 125.600 115.280 ;
        RECT 4.400 113.880 125.600 113.920 ;
        RECT 4.400 112.520 128.735 113.880 ;
        RECT 4.000 111.200 128.735 112.520 ;
        RECT 4.000 109.840 125.600 111.200 ;
        RECT 4.400 109.800 125.600 109.840 ;
        RECT 4.400 108.440 128.735 109.800 ;
        RECT 4.000 107.120 128.735 108.440 ;
        RECT 4.000 105.760 125.600 107.120 ;
        RECT 4.400 105.720 125.600 105.760 ;
        RECT 4.400 104.400 128.735 105.720 ;
        RECT 4.400 104.360 125.600 104.400 ;
        RECT 4.000 103.040 125.600 104.360 ;
        RECT 4.400 103.000 125.600 103.040 ;
        RECT 4.400 101.640 128.735 103.000 ;
        RECT 4.000 100.320 128.735 101.640 ;
        RECT 4.000 98.960 125.600 100.320 ;
        RECT 4.400 98.920 125.600 98.960 ;
        RECT 4.400 97.560 128.735 98.920 ;
        RECT 4.000 96.240 128.735 97.560 ;
        RECT 4.000 94.880 125.600 96.240 ;
        RECT 4.400 94.840 125.600 94.880 ;
        RECT 4.400 93.480 128.735 94.840 ;
        RECT 4.000 92.160 128.735 93.480 ;
        RECT 4.000 90.800 125.600 92.160 ;
        RECT 4.400 90.760 125.600 90.800 ;
        RECT 4.400 89.400 128.735 90.760 ;
        RECT 4.000 88.080 128.735 89.400 ;
        RECT 4.400 86.680 125.600 88.080 ;
        RECT 4.000 85.360 128.735 86.680 ;
        RECT 4.000 84.000 125.600 85.360 ;
        RECT 4.400 83.960 125.600 84.000 ;
        RECT 4.400 82.600 128.735 83.960 ;
        RECT 4.000 81.280 128.735 82.600 ;
        RECT 4.000 79.920 125.600 81.280 ;
        RECT 4.400 79.880 125.600 79.920 ;
        RECT 4.400 78.520 128.735 79.880 ;
        RECT 4.000 77.200 128.735 78.520 ;
        RECT 4.000 75.840 125.600 77.200 ;
        RECT 4.400 75.800 125.600 75.840 ;
        RECT 4.400 74.440 128.735 75.800 ;
        RECT 4.000 73.120 128.735 74.440 ;
        RECT 4.000 71.760 125.600 73.120 ;
        RECT 4.400 71.720 125.600 71.760 ;
        RECT 4.400 70.400 128.735 71.720 ;
        RECT 4.400 70.360 125.600 70.400 ;
        RECT 4.000 69.040 125.600 70.360 ;
        RECT 4.400 69.000 125.600 69.040 ;
        RECT 4.400 67.640 128.735 69.000 ;
        RECT 4.000 66.320 128.735 67.640 ;
        RECT 4.000 64.960 125.600 66.320 ;
        RECT 4.400 64.920 125.600 64.960 ;
        RECT 4.400 63.560 128.735 64.920 ;
        RECT 4.000 62.240 128.735 63.560 ;
        RECT 4.000 60.880 125.600 62.240 ;
        RECT 4.400 60.840 125.600 60.880 ;
        RECT 4.400 59.480 128.735 60.840 ;
        RECT 4.000 58.160 128.735 59.480 ;
        RECT 4.000 56.800 125.600 58.160 ;
        RECT 4.400 56.760 125.600 56.800 ;
        RECT 4.400 55.400 128.735 56.760 ;
        RECT 4.000 54.080 128.735 55.400 ;
        RECT 4.000 52.720 125.600 54.080 ;
        RECT 4.400 52.680 125.600 52.720 ;
        RECT 4.400 51.360 128.735 52.680 ;
        RECT 4.400 51.320 125.600 51.360 ;
        RECT 4.000 50.000 125.600 51.320 ;
        RECT 4.400 49.960 125.600 50.000 ;
        RECT 4.400 48.600 128.735 49.960 ;
        RECT 4.000 47.280 128.735 48.600 ;
        RECT 4.000 45.920 125.600 47.280 ;
        RECT 4.400 45.880 125.600 45.920 ;
        RECT 4.400 44.520 128.735 45.880 ;
        RECT 4.000 43.200 128.735 44.520 ;
        RECT 4.000 41.840 125.600 43.200 ;
        RECT 4.400 41.800 125.600 41.840 ;
        RECT 4.400 40.440 128.735 41.800 ;
        RECT 4.000 39.120 128.735 40.440 ;
        RECT 4.000 37.760 125.600 39.120 ;
        RECT 4.400 37.720 125.600 37.760 ;
        RECT 4.400 36.360 128.735 37.720 ;
        RECT 4.000 35.040 128.735 36.360 ;
        RECT 4.400 33.640 125.600 35.040 ;
        RECT 4.000 32.320 128.735 33.640 ;
        RECT 4.000 30.960 125.600 32.320 ;
        RECT 4.400 30.920 125.600 30.960 ;
        RECT 4.400 29.560 128.735 30.920 ;
        RECT 4.000 28.240 128.735 29.560 ;
        RECT 4.000 26.880 125.600 28.240 ;
        RECT 4.400 26.840 125.600 26.880 ;
        RECT 4.400 25.480 128.735 26.840 ;
        RECT 4.000 24.160 128.735 25.480 ;
        RECT 4.000 22.800 125.600 24.160 ;
        RECT 4.400 22.760 125.600 22.800 ;
        RECT 4.400 21.400 128.735 22.760 ;
        RECT 4.000 20.080 128.735 21.400 ;
        RECT 4.000 18.720 125.600 20.080 ;
        RECT 4.400 18.680 125.600 18.720 ;
        RECT 4.400 17.360 128.735 18.680 ;
        RECT 4.400 17.320 125.600 17.360 ;
        RECT 4.000 16.000 125.600 17.320 ;
        RECT 4.400 15.960 125.600 16.000 ;
        RECT 4.400 14.600 128.735 15.960 ;
        RECT 4.000 13.280 128.735 14.600 ;
        RECT 4.000 11.920 125.600 13.280 ;
        RECT 4.400 11.880 125.600 11.920 ;
        RECT 4.400 10.520 128.735 11.880 ;
        RECT 4.000 9.200 128.735 10.520 ;
        RECT 4.000 7.840 125.600 9.200 ;
        RECT 4.400 7.800 125.600 7.840 ;
        RECT 4.400 6.440 128.735 7.800 ;
        RECT 4.000 5.120 128.735 6.440 ;
        RECT 4.000 3.760 125.600 5.120 ;
        RECT 4.400 3.720 125.600 3.760 ;
        RECT 4.400 2.360 128.735 3.720 ;
        RECT 4.000 1.040 128.735 2.360 ;
        RECT 4.000 0.175 125.600 1.040 ;
      LAYER met4 ;
        RECT 43.535 10.640 43.970 198.800 ;
        RECT 46.370 10.640 63.795 198.800 ;
        RECT 66.195 10.640 83.625 198.800 ;
        RECT 86.025 10.640 103.450 198.800 ;
        RECT 105.850 10.640 115.625 198.800 ;
  END
END wrapped_rgb_mixer
END LIBRARY

