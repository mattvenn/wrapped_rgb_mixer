magic
tech sky130A
magscale 1 2
timestamp 1647002827
<< viali >>
rect 7113 39593 7147 39627
rect 7757 39525 7791 39559
rect 4261 39457 4295 39491
rect 8401 39457 8435 39491
rect 10333 39457 10367 39491
rect 11621 39457 11655 39491
rect 11805 39457 11839 39491
rect 12449 39457 12483 39491
rect 15485 39457 15519 39491
rect 19625 39457 19659 39491
rect 19993 39457 20027 39491
rect 22017 39457 22051 39491
rect 22201 39457 22235 39491
rect 23857 39457 23891 39491
rect 24777 39457 24811 39491
rect 26065 39457 26099 39491
rect 1777 39389 1811 39423
rect 2421 39389 2455 39423
rect 3065 39389 3099 39423
rect 3801 39389 3835 39423
rect 9689 39389 9723 39423
rect 10793 39389 10827 39423
rect 14289 39389 14323 39423
rect 16681 39389 16715 39423
rect 17325 39389 17359 39423
rect 18153 39389 18187 39423
rect 19441 39389 19475 39423
rect 24593 39389 24627 39423
rect 3985 39321 4019 39355
rect 14473 39321 14507 39355
rect 17969 39321 18003 39355
rect 27445 39321 27479 39355
rect 27629 39321 27663 39355
rect 1869 39253 1903 39287
rect 2513 39253 2547 39287
rect 3157 39253 3191 39287
rect 10885 39253 10919 39287
rect 16773 39253 16807 39287
rect 17417 39253 17451 39287
rect 18337 39253 18371 39287
rect 9873 39049 9907 39083
rect 1685 38981 1719 39015
rect 3985 38981 4019 39015
rect 11805 38981 11839 39015
rect 17049 38981 17083 39015
rect 17690 38981 17724 39015
rect 20177 38981 20211 39015
rect 22477 38981 22511 39015
rect 26985 38981 27019 39015
rect 27185 38981 27219 39015
rect 7389 38913 7423 38947
rect 8677 38913 8711 38947
rect 9321 38913 9355 38947
rect 9781 38913 9815 38947
rect 10425 38913 10459 38947
rect 11713 38913 11747 38947
rect 12357 38913 12391 38947
rect 12449 38913 12483 38947
rect 13001 38913 13035 38947
rect 15577 38913 15611 38947
rect 16865 38913 16899 38947
rect 17509 38913 17543 38947
rect 19901 38913 19935 38947
rect 19993 38913 20027 38947
rect 20637 38913 20671 38947
rect 20821 38913 20855 38947
rect 22293 38913 22327 38947
rect 24593 38913 24627 38947
rect 27997 38913 28031 38947
rect 1501 38845 1535 38879
rect 2881 38845 2915 38879
rect 3801 38845 3835 38879
rect 4721 38845 4755 38879
rect 13185 38845 13219 38879
rect 13553 38845 13587 38879
rect 16681 38845 16715 38879
rect 18889 38845 18923 38879
rect 23213 38845 23247 38879
rect 24777 38845 24811 38879
rect 26157 38845 26191 38879
rect 8033 38777 8067 38811
rect 6561 38709 6595 38743
rect 10517 38709 10551 38743
rect 15669 38709 15703 38743
rect 21005 38709 21039 38743
rect 27169 38709 27203 38743
rect 27353 38709 27387 38743
rect 28089 38709 28123 38743
rect 8401 38505 8435 38539
rect 13277 38505 13311 38539
rect 18245 38505 18279 38539
rect 23213 38505 23247 38539
rect 7757 38437 7791 38471
rect 9045 38437 9079 38471
rect 14381 38437 14415 38471
rect 15025 38437 15059 38471
rect 1409 38369 1443 38403
rect 1593 38369 1627 38403
rect 2789 38369 2823 38403
rect 4169 38369 4203 38403
rect 4905 38369 4939 38403
rect 5181 38369 5215 38403
rect 9781 38369 9815 38403
rect 10333 38369 10367 38403
rect 10517 38369 10551 38403
rect 11069 38369 11103 38403
rect 15577 38369 15611 38403
rect 15761 38369 15795 38403
rect 16129 38369 16163 38403
rect 17877 38369 17911 38403
rect 19257 38369 19291 38403
rect 20177 38369 20211 38403
rect 20361 38369 20395 38403
rect 20729 38369 20763 38403
rect 23489 38369 23523 38403
rect 26341 38369 26375 38403
rect 27721 38369 27755 38403
rect 4077 38301 4111 38335
rect 4721 38301 4755 38335
rect 9229 38301 9263 38335
rect 9689 38301 9723 38335
rect 13185 38301 13219 38335
rect 14289 38301 14323 38335
rect 14933 38301 14967 38335
rect 18061 38301 18095 38335
rect 19441 38301 19475 38335
rect 22477 38301 22511 38335
rect 23673 38301 23707 38335
rect 24685 38301 24719 38335
rect 24777 38301 24811 38335
rect 24869 38301 24903 38335
rect 25053 38301 25087 38335
rect 25697 38301 25731 38335
rect 25881 38301 25915 38335
rect 22661 38233 22695 38267
rect 22845 38233 22879 38267
rect 25513 38233 25547 38267
rect 26525 38233 26559 38267
rect 19625 38165 19659 38199
rect 23857 38165 23891 38199
rect 24409 38165 24443 38199
rect 19901 37961 19935 37995
rect 1777 37893 1811 37927
rect 4077 37893 4111 37927
rect 6469 37893 6503 37927
rect 16926 37893 16960 37927
rect 24777 37893 24811 37927
rect 26433 37893 26467 37927
rect 27997 37893 28031 37927
rect 6377 37825 6411 37859
rect 8309 37825 8343 37859
rect 8861 37825 8895 37859
rect 9965 37825 9999 37859
rect 11713 37825 11747 37859
rect 12357 37825 12391 37859
rect 14841 37825 14875 37859
rect 15945 37825 15979 37859
rect 18777 37825 18811 37859
rect 20453 37825 20487 37859
rect 20821 37825 20855 37859
rect 21833 37825 21867 37859
rect 24593 37825 24627 37859
rect 27169 37825 27203 37859
rect 1593 37757 1627 37791
rect 2789 37757 2823 37791
rect 3893 37757 3927 37791
rect 4537 37757 4571 37791
rect 9137 37757 9171 37791
rect 10793 37757 10827 37791
rect 11805 37757 11839 37791
rect 12541 37757 12575 37791
rect 12909 37757 12943 37791
rect 14657 37757 14691 37791
rect 15761 37757 15795 37791
rect 16681 37757 16715 37791
rect 18521 37757 18555 37791
rect 22017 37757 22051 37791
rect 22293 37757 22327 37791
rect 27353 37757 27387 37791
rect 27445 37757 27479 37791
rect 7665 37689 7699 37723
rect 16129 37689 16163 37723
rect 8125 37621 8159 37655
rect 15025 37621 15059 37655
rect 18061 37621 18095 37655
rect 26985 37621 27019 37655
rect 28089 37621 28123 37655
rect 6377 37417 6411 37451
rect 7113 37417 7147 37451
rect 7757 37417 7791 37451
rect 17785 37417 17819 37451
rect 18245 37417 18279 37451
rect 25789 37417 25823 37451
rect 8953 37349 8987 37383
rect 9781 37349 9815 37383
rect 13277 37349 13311 37383
rect 1869 37281 1903 37315
rect 5457 37281 5491 37315
rect 11989 37281 12023 37315
rect 12909 37281 12943 37315
rect 16405 37281 16439 37315
rect 26525 37281 26559 37315
rect 1409 37213 1443 37247
rect 3893 37213 3927 37247
rect 5089 37213 5123 37247
rect 8401 37213 8435 37247
rect 9137 37213 9171 37247
rect 9597 37213 9631 37247
rect 10425 37213 10459 37247
rect 11621 37213 11655 37247
rect 13079 37207 13113 37241
rect 14565 37213 14599 37247
rect 18245 37213 18279 37247
rect 18429 37213 18463 37247
rect 18521 37213 18555 37247
rect 19349 37213 19383 37247
rect 20361 37213 20395 37247
rect 21465 37213 21499 37247
rect 21741 37213 21775 37247
rect 22477 37213 22511 37247
rect 24409 37213 24443 37247
rect 24676 37213 24710 37247
rect 26341 37213 26375 37247
rect 28181 37213 28215 37247
rect 1593 37145 1627 37179
rect 4445 37145 4479 37179
rect 10885 37145 10919 37179
rect 14810 37145 14844 37179
rect 16672 37145 16706 37179
rect 19625 37145 19659 37179
rect 20913 37145 20947 37179
rect 22722 37145 22756 37179
rect 8217 37077 8251 37111
rect 15945 37077 15979 37111
rect 18705 37077 18739 37111
rect 23857 37077 23891 37111
rect 1593 36873 1627 36907
rect 2329 36873 2363 36907
rect 9781 36873 9815 36907
rect 15025 36873 15059 36907
rect 15669 36873 15703 36907
rect 16037 36873 16071 36907
rect 18889 36873 18923 36907
rect 22017 36873 22051 36907
rect 22569 36873 22603 36907
rect 24041 36873 24075 36907
rect 27353 36873 27387 36907
rect 4997 36805 5031 36839
rect 9045 36805 9079 36839
rect 12072 36805 12106 36839
rect 1501 36737 1535 36771
rect 2145 36737 2179 36771
rect 3065 36737 3099 36771
rect 4445 36737 4479 36771
rect 5733 36737 5767 36771
rect 7113 36737 7147 36771
rect 7849 36737 7883 36771
rect 8493 36737 8527 36771
rect 8953 36737 8987 36771
rect 9137 36737 9171 36771
rect 9597 36737 9631 36771
rect 9781 36737 9815 36771
rect 10333 36737 10367 36771
rect 10793 36737 10827 36771
rect 13901 36737 13935 36771
rect 15485 36737 15519 36771
rect 15761 36737 15795 36771
rect 15853 36737 15887 36771
rect 16681 36737 16715 36771
rect 16865 36737 16899 36771
rect 17776 36737 17810 36771
rect 19605 36737 19639 36771
rect 21925 36737 21959 36771
rect 22845 36737 22879 36771
rect 22937 36737 22971 36771
rect 23029 36737 23063 36771
rect 23213 36737 23247 36771
rect 23857 36737 23891 36771
rect 24133 36737 24167 36771
rect 24593 36737 24627 36771
rect 26433 36737 26467 36771
rect 27169 36737 27203 36771
rect 27445 36737 27479 36771
rect 27905 36737 27939 36771
rect 3709 36669 3743 36703
rect 11805 36669 11839 36703
rect 13645 36669 13679 36703
rect 17049 36669 17083 36703
rect 17509 36669 17543 36703
rect 19349 36669 19383 36703
rect 24777 36669 24811 36703
rect 26985 36669 27019 36703
rect 28181 36669 28215 36703
rect 8309 36601 8343 36635
rect 13185 36601 13219 36635
rect 28089 36601 28123 36635
rect 20729 36533 20763 36567
rect 23673 36533 23707 36567
rect 27997 36533 28031 36567
rect 1685 36329 1719 36363
rect 3893 36329 3927 36363
rect 4629 36329 4663 36363
rect 5273 36329 5307 36363
rect 6469 36329 6503 36363
rect 7113 36329 7147 36363
rect 9597 36329 9631 36363
rect 11253 36329 11287 36363
rect 23397 36329 23431 36363
rect 25053 36329 25087 36363
rect 7573 36261 7607 36295
rect 8217 36261 8251 36295
rect 8953 36261 8987 36295
rect 10333 36261 10367 36295
rect 15485 36261 15519 36295
rect 22017 36261 22051 36295
rect 25881 36261 25915 36295
rect 3157 36193 3191 36227
rect 10885 36193 10919 36227
rect 11805 36193 11839 36227
rect 14105 36193 14139 36227
rect 16773 36193 16807 36227
rect 23121 36193 23155 36227
rect 24777 36193 24811 36227
rect 24869 36193 24903 36227
rect 26525 36193 26559 36227
rect 28181 36193 28215 36227
rect 2605 36125 2639 36159
rect 3801 36125 3835 36159
rect 7757 36125 7791 36159
rect 8401 36125 8435 36159
rect 9137 36125 9171 36159
rect 9781 36125 9815 36159
rect 10241 36125 10275 36159
rect 11069 36125 11103 36159
rect 15945 36125 15979 36159
rect 16129 36125 16163 36159
rect 19441 36125 19475 36159
rect 20361 36125 20395 36159
rect 21741 36125 21775 36159
rect 21833 36125 21867 36159
rect 22109 36125 22143 36159
rect 22753 36125 22787 36159
rect 23213 36125 23247 36159
rect 25697 36125 25731 36159
rect 26341 36125 26375 36159
rect 12050 36057 12084 36091
rect 14350 36057 14384 36091
rect 17018 36057 17052 36091
rect 19257 36057 19291 36091
rect 19625 36057 19659 36091
rect 20913 36057 20947 36091
rect 25513 36057 25547 36091
rect 13185 35989 13219 36023
rect 16313 35989 16347 36023
rect 18153 35989 18187 36023
rect 19533 35989 19567 36023
rect 19809 35989 19843 36023
rect 21557 35989 21591 36023
rect 24409 35989 24443 36023
rect 3893 35785 3927 35819
rect 8033 35785 8067 35819
rect 8677 35785 8711 35819
rect 9505 35785 9539 35819
rect 12081 35785 12115 35819
rect 17693 35785 17727 35819
rect 18153 35785 18187 35819
rect 21281 35785 21315 35819
rect 22569 35785 22603 35819
rect 24501 35785 24535 35819
rect 27721 35785 27755 35819
rect 12909 35717 12943 35751
rect 18429 35717 18463 35751
rect 18521 35717 18555 35751
rect 18659 35717 18693 35751
rect 25320 35717 25354 35751
rect 27997 35717 28031 35751
rect 3801 35649 3835 35683
rect 4629 35649 4663 35683
rect 6561 35649 6595 35683
rect 7573 35649 7607 35683
rect 8217 35649 8251 35683
rect 8861 35649 8895 35683
rect 9321 35649 9355 35683
rect 9505 35649 9539 35683
rect 9965 35649 9999 35683
rect 10793 35649 10827 35683
rect 11989 35649 12023 35683
rect 12725 35649 12759 35683
rect 13369 35649 13403 35683
rect 13553 35649 13587 35683
rect 14381 35649 14415 35683
rect 15301 35649 15335 35683
rect 15485 35649 15519 35683
rect 15577 35649 15611 35683
rect 16681 35649 16715 35683
rect 17509 35649 17543 35683
rect 18337 35649 18371 35683
rect 18797 35649 18831 35683
rect 20913 35649 20947 35683
rect 21833 35649 21867 35683
rect 22017 35649 22051 35683
rect 22385 35649 22419 35683
rect 23397 35649 23431 35683
rect 24409 35649 24443 35683
rect 25053 35649 25087 35683
rect 26985 35649 27019 35683
rect 27169 35649 27203 35683
rect 27261 35649 27295 35683
rect 27537 35649 27571 35683
rect 1501 35581 1535 35615
rect 1685 35581 1719 35615
rect 2881 35581 2915 35615
rect 10057 35581 10091 35615
rect 10609 35581 10643 35615
rect 14197 35581 14231 35615
rect 17325 35581 17359 35615
rect 19717 35581 19751 35615
rect 20637 35581 20671 35615
rect 21005 35581 21039 35615
rect 21122 35581 21156 35615
rect 22109 35581 22143 35615
rect 22201 35581 22235 35615
rect 23673 35581 23707 35615
rect 27353 35581 27387 35615
rect 5273 35513 5307 35547
rect 20085 35513 20119 35547
rect 20177 35513 20211 35547
rect 26433 35513 26467 35547
rect 10977 35445 11011 35479
rect 13737 35445 13771 35479
rect 14565 35445 14599 35479
rect 15485 35445 15519 35479
rect 15761 35445 15795 35479
rect 16773 35445 16807 35479
rect 23765 35445 23799 35479
rect 23949 35445 23983 35479
rect 1777 35241 1811 35275
rect 3985 35241 4019 35275
rect 4445 35241 4479 35275
rect 6285 35241 6319 35275
rect 9229 35241 9263 35275
rect 11161 35241 11195 35275
rect 11897 35241 11931 35275
rect 25789 35241 25823 35275
rect 5641 35173 5675 35207
rect 12817 35173 12851 35207
rect 14933 35173 14967 35207
rect 17049 35173 17083 35207
rect 17509 35173 17543 35207
rect 18245 35173 18279 35207
rect 19349 35173 19383 35207
rect 12449 35105 12483 35139
rect 14473 35105 14507 35139
rect 15669 35105 15703 35139
rect 19901 35105 19935 35139
rect 23029 35105 23063 35139
rect 24409 35105 24443 35139
rect 24685 35105 24719 35139
rect 26341 35105 26375 35139
rect 28181 35105 28215 35139
rect 1685 35037 1719 35071
rect 2421 35037 2455 35071
rect 3249 35037 3283 35071
rect 4629 35037 4663 35071
rect 5365 35037 5399 35071
rect 5825 35037 5859 35071
rect 6469 35037 6503 35071
rect 7113 35037 7147 35071
rect 7757 35037 7791 35071
rect 8401 35037 8435 35071
rect 9137 35037 9171 35071
rect 9321 35037 9355 35071
rect 9781 35037 9815 35071
rect 9965 35037 9999 35071
rect 10425 35037 10459 35071
rect 11077 35039 11111 35073
rect 12633 35037 12667 35071
rect 13369 35037 13403 35071
rect 14105 35037 14139 35071
rect 14289 35037 14323 35071
rect 14933 35037 14967 35071
rect 15117 35037 15151 35071
rect 15209 35037 15243 35071
rect 17785 35037 17819 35071
rect 18429 35037 18463 35071
rect 18705 35037 18739 35071
rect 19257 35037 19291 35071
rect 21741 35037 21775 35071
rect 21925 35037 21959 35071
rect 22090 35037 22124 35071
rect 22201 35037 22235 35071
rect 22293 35037 22327 35071
rect 22937 35037 22971 35071
rect 25697 35037 25731 35071
rect 11805 34969 11839 35003
rect 15914 34969 15948 35003
rect 17509 34969 17543 35003
rect 20146 34969 20180 35003
rect 26525 34969 26559 35003
rect 2513 34901 2547 34935
rect 7573 34901 7607 34935
rect 8217 34901 8251 34935
rect 9873 34901 9907 34935
rect 10517 34901 10551 34935
rect 13461 34901 13495 34935
rect 17693 34901 17727 34935
rect 18613 34901 18647 34935
rect 21281 34901 21315 34935
rect 23305 34901 23339 34935
rect 9505 34697 9539 34731
rect 10333 34697 10367 34731
rect 17049 34697 17083 34731
rect 24961 34697 24995 34731
rect 1869 34629 1903 34663
rect 11774 34629 11808 34663
rect 18582 34629 18616 34663
rect 20454 34629 20488 34663
rect 21925 34629 21959 34663
rect 22109 34629 22143 34663
rect 26985 34629 27019 34663
rect 1685 34561 1719 34595
rect 7757 34561 7791 34595
rect 8401 34561 8435 34595
rect 9045 34561 9079 34595
rect 9689 34561 9723 34595
rect 10149 34561 10183 34595
rect 10333 34561 10367 34595
rect 10793 34561 10827 34595
rect 13625 34561 13659 34595
rect 15945 34561 15979 34595
rect 16681 34561 16715 34595
rect 16865 34561 16899 34595
rect 17509 34561 17543 34595
rect 17693 34561 17727 34595
rect 18337 34561 18371 34595
rect 20361 34561 20395 34595
rect 20545 34561 20579 34595
rect 20663 34561 20697 34595
rect 20821 34561 20855 34595
rect 22845 34561 22879 34595
rect 23029 34561 23063 34595
rect 23765 34561 23799 34595
rect 24593 34561 24627 34595
rect 24777 34561 24811 34595
rect 25605 34561 25639 34595
rect 27169 34561 27203 34595
rect 27905 34561 27939 34595
rect 28089 34561 28123 34595
rect 28181 34561 28215 34595
rect 2789 34493 2823 34527
rect 11529 34493 11563 34527
rect 13369 34493 13403 34527
rect 15761 34493 15795 34527
rect 22753 34493 22787 34527
rect 22937 34493 22971 34527
rect 23857 34493 23891 34527
rect 25513 34493 25547 34527
rect 27445 34493 27479 34527
rect 7113 34425 7147 34459
rect 8861 34425 8895 34459
rect 10885 34425 10919 34459
rect 16129 34425 16163 34459
rect 17877 34425 17911 34459
rect 19717 34425 19751 34459
rect 24133 34425 24167 34459
rect 25973 34425 26007 34459
rect 27353 34425 27387 34459
rect 27905 34425 27939 34459
rect 4169 34357 4203 34391
rect 7573 34357 7607 34391
rect 8217 34357 8251 34391
rect 12909 34357 12943 34391
rect 14749 34357 14783 34391
rect 20177 34357 20211 34391
rect 22569 34357 22603 34391
rect 11529 34153 11563 34187
rect 12357 34153 12391 34187
rect 13369 34153 13403 34187
rect 16957 34153 16991 34187
rect 18705 34153 18739 34187
rect 24593 34153 24627 34187
rect 6929 34085 6963 34119
rect 8217 34085 8251 34119
rect 13553 34085 13587 34119
rect 18153 34085 18187 34119
rect 22293 34085 22327 34119
rect 22477 34085 22511 34119
rect 23305 34085 23339 34119
rect 24777 34085 24811 34119
rect 1409 34017 1443 34051
rect 2789 34017 2823 34051
rect 19257 34017 19291 34051
rect 22017 34017 22051 34051
rect 23397 34017 23431 34051
rect 25421 34017 25455 34051
rect 25697 34017 25731 34051
rect 26341 34017 26375 34051
rect 28181 34017 28215 34051
rect 7113 33949 7147 33983
rect 7757 33949 7791 33983
rect 8401 33949 8435 33983
rect 9229 33949 9263 33983
rect 9677 33949 9711 33983
rect 9873 33949 9907 33983
rect 10333 33949 10367 33983
rect 10517 33949 10551 33983
rect 11253 33949 11287 33983
rect 11345 33949 11379 33983
rect 11989 33949 12023 33983
rect 12173 33949 12207 33983
rect 13277 33949 13311 33983
rect 13369 33949 13403 33983
rect 14105 33949 14139 33983
rect 14289 33949 14323 33983
rect 14657 33949 14691 33983
rect 15577 33949 15611 33983
rect 17693 33949 17727 33983
rect 21097 33949 21131 33983
rect 23121 33949 23155 33983
rect 25513 33949 25547 33983
rect 25605 33949 25639 33983
rect 1593 33881 1627 33915
rect 9781 33881 9815 33915
rect 10701 33881 10735 33915
rect 13093 33881 13127 33915
rect 14473 33881 14507 33915
rect 15822 33881 15856 33915
rect 17509 33881 17543 33915
rect 18337 33881 18371 33915
rect 19502 33881 19536 33915
rect 21373 33881 21407 33915
rect 24409 33881 24443 33915
rect 24609 33881 24643 33915
rect 26525 33881 26559 33915
rect 7573 33813 7607 33847
rect 9045 33813 9079 33847
rect 14381 33813 14415 33847
rect 18429 33813 18463 33847
rect 18521 33813 18555 33847
rect 20637 33813 20671 33847
rect 22937 33813 22971 33847
rect 25237 33813 25271 33847
rect 1593 33609 1627 33643
rect 2237 33609 2271 33643
rect 9597 33609 9631 33643
rect 21189 33609 21223 33643
rect 28089 33609 28123 33643
rect 17478 33541 17512 33575
rect 20054 33541 20088 33575
rect 1409 33473 1443 33507
rect 2145 33473 2179 33507
rect 8401 33473 8435 33507
rect 9045 33473 9079 33507
rect 9505 33473 9539 33507
rect 9689 33473 9723 33507
rect 10149 33473 10183 33507
rect 10333 33473 10367 33507
rect 10793 33473 10827 33507
rect 10977 33473 11011 33507
rect 11989 33473 12023 33507
rect 12173 33473 12207 33507
rect 12817 33473 12851 33507
rect 13461 33473 13495 33507
rect 13717 33473 13751 33507
rect 17233 33473 17267 33507
rect 19165 33473 19199 33507
rect 19809 33473 19843 33507
rect 22063 33473 22097 33507
rect 22201 33473 22235 33507
rect 22314 33473 22348 33507
rect 22477 33473 22511 33507
rect 23653 33473 23687 33507
rect 23765 33473 23799 33507
rect 23857 33476 23891 33510
rect 24041 33473 24075 33507
rect 27169 33473 27203 33507
rect 27997 33473 28031 33507
rect 7757 33405 7791 33439
rect 12357 33405 12391 33439
rect 12909 33405 12943 33439
rect 15301 33405 15335 33439
rect 24593 33405 24627 33439
rect 24777 33405 24811 33439
rect 26157 33405 26191 33439
rect 27261 33405 27295 33439
rect 8861 33337 8895 33371
rect 10793 33337 10827 33371
rect 14841 33337 14875 33371
rect 15531 33337 15565 33371
rect 18613 33337 18647 33371
rect 19349 33337 19383 33371
rect 8217 33269 8251 33303
rect 10149 33269 10183 33303
rect 21833 33269 21867 33303
rect 23397 33269 23431 33303
rect 27445 33269 27479 33303
rect 1409 33065 1443 33099
rect 8217 33065 8251 33099
rect 12357 33065 12391 33099
rect 17693 33065 17727 33099
rect 18245 33065 18279 33099
rect 9597 32997 9631 33031
rect 22661 32997 22695 33031
rect 14749 32929 14783 32963
rect 15669 32929 15703 32963
rect 23213 32929 23247 32963
rect 25697 32929 25731 32963
rect 25881 32929 25915 32963
rect 26341 32929 26375 32963
rect 28181 32929 28215 32963
rect 1593 32861 1627 32895
rect 7757 32861 7791 32895
rect 8401 32861 8435 32895
rect 9505 32861 9539 32895
rect 9689 32861 9723 32895
rect 10241 32861 10275 32895
rect 10333 32861 10367 32895
rect 10977 32861 11011 32895
rect 13093 32861 13127 32895
rect 13369 32861 13403 32895
rect 14289 32861 14323 32895
rect 14473 32861 14507 32895
rect 17509 32861 17543 32895
rect 18245 32861 18279 32895
rect 18429 32861 18463 32895
rect 18521 32861 18555 32895
rect 19257 32861 19291 32895
rect 19441 32861 19475 32895
rect 20177 32861 20211 32895
rect 21281 32861 21315 32895
rect 21548 32861 21582 32895
rect 23383 32861 23417 32895
rect 24777 32861 24811 32895
rect 24866 32861 24900 32895
rect 24966 32861 25000 32895
rect 25145 32861 25179 32895
rect 25605 32861 25639 32895
rect 11222 32793 11256 32827
rect 12817 32793 12851 32827
rect 13001 32793 13035 32827
rect 14381 32793 14415 32827
rect 14591 32793 14625 32827
rect 15914 32793 15948 32827
rect 20545 32793 20579 32827
rect 26525 32793 26559 32827
rect 10517 32725 10551 32759
rect 13185 32725 13219 32759
rect 14105 32725 14139 32759
rect 17049 32725 17083 32759
rect 18705 32725 18739 32759
rect 19625 32725 19659 32759
rect 19901 32725 19935 32759
rect 23673 32725 23707 32759
rect 24501 32725 24535 32759
rect 25881 32725 25915 32759
rect 7941 32521 7975 32555
rect 9965 32453 9999 32487
rect 17049 32453 17083 32487
rect 18490 32453 18524 32487
rect 21189 32453 21223 32487
rect 7481 32385 7515 32419
rect 8125 32385 8159 32419
rect 8585 32385 8619 32419
rect 8769 32385 8803 32419
rect 9413 32385 9447 32419
rect 10793 32385 10827 32419
rect 11785 32385 11819 32419
rect 13369 32385 13403 32419
rect 13645 32385 13679 32419
rect 14289 32385 14323 32419
rect 14545 32385 14579 32419
rect 16773 32385 16807 32419
rect 16957 32385 16991 32419
rect 17141 32385 17175 32419
rect 18245 32385 18279 32419
rect 20637 32385 20671 32419
rect 21833 32385 21867 32419
rect 22100 32385 22134 32419
rect 23673 32385 23707 32419
rect 23929 32385 23963 32419
rect 25697 32385 25731 32419
rect 27169 32385 27203 32419
rect 27997 32385 28031 32419
rect 1501 32317 1535 32351
rect 1685 32317 1719 32351
rect 2881 32317 2915 32351
rect 10149 32317 10183 32351
rect 10609 32317 10643 32351
rect 11529 32317 11563 32351
rect 13461 32317 13495 32351
rect 25605 32317 25639 32351
rect 27261 32317 27295 32351
rect 8677 32249 8711 32283
rect 23213 32249 23247 32283
rect 25053 32249 25087 32283
rect 7297 32181 7331 32215
rect 9229 32181 9263 32215
rect 10977 32181 11011 32215
rect 12909 32181 12943 32215
rect 13461 32181 13495 32215
rect 13829 32181 13863 32215
rect 15669 32181 15703 32215
rect 17325 32181 17359 32215
rect 19625 32181 19659 32215
rect 25973 32181 26007 32215
rect 27445 32181 27479 32215
rect 28089 32181 28123 32215
rect 1777 31977 1811 32011
rect 7573 31977 7607 32011
rect 15485 31977 15519 32011
rect 18521 31977 18555 32011
rect 20361 31977 20395 32011
rect 22845 31977 22879 32011
rect 23489 31977 23523 32011
rect 9505 31909 9539 31943
rect 10057 31841 10091 31875
rect 16221 31841 16255 31875
rect 26341 31841 26375 31875
rect 28181 31841 28215 31875
rect 2421 31773 2455 31807
rect 6285 31773 6319 31807
rect 6929 31773 6963 31807
rect 7757 31773 7791 31807
rect 8217 31773 8251 31807
rect 8401 31773 8435 31807
rect 9413 31773 9447 31807
rect 10241 31773 10275 31807
rect 11069 31773 11103 31807
rect 11713 31773 11747 31807
rect 14105 31773 14139 31807
rect 14361 31773 14395 31807
rect 20085 31773 20119 31807
rect 20177 31773 20211 31807
rect 20821 31773 20855 31807
rect 21741 31773 21775 31807
rect 23397 31773 23431 31807
rect 24501 31773 24535 31807
rect 24757 31773 24791 31807
rect 8309 31705 8343 31739
rect 10885 31705 10919 31739
rect 11958 31705 11992 31739
rect 16488 31705 16522 31739
rect 18337 31705 18371 31739
rect 19809 31705 19843 31739
rect 19993 31705 20027 31739
rect 21097 31705 21131 31739
rect 22017 31705 22051 31739
rect 22753 31705 22787 31739
rect 26525 31705 26559 31739
rect 6745 31637 6779 31671
rect 10425 31637 10459 31671
rect 11253 31637 11287 31671
rect 13093 31637 13127 31671
rect 17601 31637 17635 31671
rect 18537 31637 18571 31671
rect 18705 31637 18739 31671
rect 23857 31637 23891 31671
rect 25881 31637 25915 31671
rect 7849 31433 7883 31467
rect 10149 31433 10183 31467
rect 14289 31433 14323 31467
rect 21281 31433 21315 31467
rect 26433 31433 26467 31467
rect 26985 31433 27019 31467
rect 27353 31433 27387 31467
rect 28089 31433 28123 31467
rect 14994 31365 15028 31399
rect 17938 31365 17972 31399
rect 21925 31365 21959 31399
rect 24225 31365 24259 31399
rect 24317 31365 24351 31399
rect 1685 31297 1719 31331
rect 6745 31297 6779 31331
rect 7389 31297 7423 31331
rect 8033 31297 8067 31331
rect 8493 31297 8527 31331
rect 9137 31297 9171 31331
rect 9873 31297 9907 31331
rect 9965 31297 9999 31331
rect 10793 31297 10827 31331
rect 11621 31297 11655 31331
rect 11805 31297 11839 31331
rect 12449 31297 12483 31331
rect 13277 31297 13311 31331
rect 13461 31297 13495 31331
rect 14105 31297 14139 31331
rect 14749 31297 14783 31331
rect 16681 31297 16715 31331
rect 16957 31297 16991 31331
rect 20157 31297 20191 31331
rect 23029 31297 23063 31331
rect 23121 31297 23155 31331
rect 23397 31297 23431 31331
rect 24041 31297 24075 31331
rect 24409 31297 24443 31331
rect 25053 31297 25087 31331
rect 25320 31297 25354 31331
rect 27169 31297 27203 31331
rect 27445 31297 27479 31331
rect 27905 31297 27939 31331
rect 28181 31297 28215 31331
rect 1869 31229 1903 31263
rect 2789 31229 2823 31263
rect 10609 31229 10643 31263
rect 12265 31229 12299 31263
rect 13093 31229 13127 31263
rect 13921 31229 13955 31263
rect 16773 31229 16807 31263
rect 17693 31229 17727 31263
rect 19901 31229 19935 31263
rect 6561 31161 6595 31195
rect 9229 31161 9263 31195
rect 22293 31161 22327 31195
rect 23305 31161 23339 31195
rect 7205 31093 7239 31127
rect 8585 31093 8619 31127
rect 10977 31093 11011 31127
rect 12633 31093 12667 31127
rect 16129 31093 16163 31127
rect 16865 31093 16899 31127
rect 17141 31093 17175 31127
rect 19073 31093 19107 31127
rect 22385 31093 22419 31127
rect 22845 31093 22879 31127
rect 24593 31093 24627 31127
rect 27905 31093 27939 31127
rect 2329 30889 2363 30923
rect 6929 30889 6963 30923
rect 7573 30889 7607 30923
rect 15301 30889 15335 30923
rect 19993 30889 20027 30923
rect 20177 30889 20211 30923
rect 24777 30889 24811 30923
rect 8217 30821 8251 30855
rect 9873 30753 9907 30787
rect 14473 30753 14507 30787
rect 19901 30753 19935 30787
rect 26525 30753 26559 30787
rect 28181 30753 28215 30787
rect 2237 30685 2271 30719
rect 7113 30685 7147 30719
rect 7757 30685 7791 30719
rect 8401 30685 8435 30719
rect 9229 30685 9263 30719
rect 10057 30685 10091 30719
rect 10793 30685 10827 30719
rect 10885 30685 10919 30719
rect 12357 30685 12391 30719
rect 12541 30685 12575 30719
rect 13277 30685 13311 30719
rect 13369 30685 13403 30719
rect 14197 30685 14231 30719
rect 14289 30685 14323 30719
rect 14933 30685 14967 30719
rect 15117 30685 15151 30719
rect 15853 30685 15887 30719
rect 17049 30685 17083 30719
rect 17233 30685 17267 30719
rect 17351 30685 17385 30719
rect 17509 30685 17543 30719
rect 18337 30685 18371 30719
rect 18521 30685 18555 30719
rect 19993 30685 20027 30719
rect 20729 30685 20763 30719
rect 20996 30685 21030 30719
rect 22937 30685 22971 30719
rect 23029 30685 23063 30719
rect 23213 30685 23247 30719
rect 23305 30685 23339 30719
rect 24501 30685 24535 30719
rect 24593 30685 24627 30719
rect 25237 30685 25271 30719
rect 25385 30685 25419 30719
rect 25743 30685 25777 30719
rect 26341 30685 26375 30719
rect 11069 30617 11103 30651
rect 11529 30617 11563 30651
rect 11713 30617 11747 30651
rect 11897 30617 11931 30651
rect 16221 30617 16255 30651
rect 16405 30617 16439 30651
rect 17141 30617 17175 30651
rect 19717 30617 19751 30651
rect 25513 30617 25547 30651
rect 25605 30617 25639 30651
rect 9321 30549 9355 30583
rect 10241 30549 10275 30583
rect 12725 30549 12759 30583
rect 13553 30549 13587 30583
rect 16037 30549 16071 30583
rect 16129 30549 16163 30583
rect 16865 30549 16899 30583
rect 18705 30549 18739 30583
rect 22109 30549 22143 30583
rect 22753 30549 22787 30583
rect 25881 30549 25915 30583
rect 8033 30345 8067 30379
rect 15393 30345 15427 30379
rect 23213 30345 23247 30379
rect 25973 30345 26007 30379
rect 10057 30277 10091 30311
rect 10241 30277 10275 30311
rect 10793 30277 10827 30311
rect 11774 30277 11808 30311
rect 14258 30277 14292 30311
rect 16037 30277 16071 30311
rect 17386 30277 17420 30311
rect 19248 30277 19282 30311
rect 6929 30209 6963 30243
rect 7941 30209 7975 30243
rect 8217 30209 8251 30243
rect 8861 30209 8895 30243
rect 9505 30209 9539 30243
rect 13369 30209 13403 30243
rect 14013 30209 14047 30243
rect 15853 30209 15887 30243
rect 16129 30209 16163 30243
rect 18981 30209 19015 30243
rect 20821 30209 20855 30243
rect 20913 30209 20947 30243
rect 21833 30209 21867 30243
rect 22100 30209 22134 30243
rect 23673 30209 23707 30243
rect 25237 30209 25271 30243
rect 25421 30209 25455 30243
rect 25605 30209 25639 30243
rect 25789 30209 25823 30243
rect 26985 30209 27019 30243
rect 27169 30209 27203 30243
rect 27261 30209 27295 30243
rect 27537 30209 27571 30243
rect 10977 30141 11011 30175
rect 11529 30141 11563 30175
rect 17141 30141 17175 30175
rect 21189 30141 21223 30175
rect 23949 30141 23983 30175
rect 25513 30141 25547 30175
rect 27353 30141 27387 30175
rect 7757 30073 7791 30107
rect 13461 30073 13495 30107
rect 6745 30005 6779 30039
rect 7297 30005 7331 30039
rect 7665 30005 7699 30039
rect 8677 30005 8711 30039
rect 9321 30005 9355 30039
rect 12909 30005 12943 30039
rect 15853 30005 15887 30039
rect 18521 30005 18555 30039
rect 20361 30005 20395 30039
rect 21097 30005 21131 30039
rect 21281 30005 21315 30039
rect 27721 30005 27755 30039
rect 9229 29801 9263 29835
rect 18613 29801 18647 29835
rect 23857 29801 23891 29835
rect 25881 29801 25915 29835
rect 8217 29733 8251 29767
rect 13553 29733 13587 29767
rect 16129 29733 16163 29767
rect 14749 29665 14783 29699
rect 16589 29665 16623 29699
rect 21925 29665 21959 29699
rect 24501 29665 24535 29699
rect 26801 29665 26835 29699
rect 1593 29597 1627 29631
rect 7757 29597 7791 29631
rect 8401 29597 8435 29631
rect 9413 29597 9447 29631
rect 10057 29597 10091 29631
rect 10241 29597 10275 29631
rect 10701 29597 10735 29631
rect 11437 29597 11471 29631
rect 11529 29597 11563 29631
rect 11713 29597 11747 29631
rect 12173 29597 12207 29631
rect 14105 29597 14139 29631
rect 14197 29597 14231 29631
rect 19257 29597 19291 29631
rect 19441 29597 19475 29631
rect 20361 29597 20395 29631
rect 23213 29597 23247 29631
rect 23306 29597 23340 29631
rect 23489 29597 23523 29631
rect 23719 29597 23753 29631
rect 24768 29597 24802 29631
rect 26341 29597 26375 29631
rect 9781 29529 9815 29563
rect 12440 29529 12474 29563
rect 14994 29529 15028 29563
rect 16834 29529 16868 29563
rect 18521 29529 18555 29563
rect 20545 29529 20579 29563
rect 23581 29529 23615 29563
rect 26525 29529 26559 29563
rect 7573 29461 7607 29495
rect 10149 29461 10183 29495
rect 10793 29461 10827 29495
rect 17969 29461 18003 29495
rect 19625 29461 19659 29495
rect 27077 29257 27111 29291
rect 11897 29189 11931 29223
rect 15669 29189 15703 29223
rect 27445 29189 27479 29223
rect 1409 29121 1443 29155
rect 8401 29121 8435 29155
rect 9045 29121 9079 29155
rect 9689 29121 9723 29155
rect 10149 29121 10183 29155
rect 10333 29121 10367 29155
rect 10793 29121 10827 29155
rect 12541 29121 12575 29155
rect 12797 29121 12831 29155
rect 14933 29121 14967 29155
rect 15025 29121 15059 29155
rect 15853 29121 15887 29155
rect 15945 29121 15979 29155
rect 16681 29121 16715 29155
rect 17673 29121 17707 29155
rect 19973 29121 20007 29155
rect 22201 29121 22235 29155
rect 23029 29121 23063 29155
rect 23305 29121 23339 29155
rect 24317 29121 24351 29155
rect 24584 29121 24618 29155
rect 26157 29121 26191 29155
rect 26985 29121 27019 29155
rect 27261 29121 27295 29155
rect 27905 29121 27939 29155
rect 1593 29053 1627 29087
rect 2789 29053 2823 29087
rect 17417 29053 17451 29087
rect 19717 29053 19751 29087
rect 22477 29053 22511 29087
rect 27353 29053 27387 29087
rect 7757 28985 7791 29019
rect 8217 28985 8251 29019
rect 12081 28985 12115 29019
rect 16129 28985 16163 29019
rect 18797 28985 18831 29019
rect 25697 28985 25731 29019
rect 28089 28985 28123 29019
rect 8861 28917 8895 28951
rect 9505 28917 9539 28951
rect 10149 28917 10183 28951
rect 10885 28917 10919 28951
rect 13921 28917 13955 28951
rect 15209 28917 15243 28951
rect 15945 28917 15979 28951
rect 16865 28917 16899 28951
rect 21097 28917 21131 28951
rect 22017 28917 22051 28951
rect 22385 28917 22419 28951
rect 26341 28917 26375 28951
rect 1685 28713 1719 28747
rect 10701 28713 10735 28747
rect 17969 28713 18003 28747
rect 23121 28713 23155 28747
rect 16221 28645 16255 28679
rect 11242 28577 11276 28611
rect 13461 28577 13495 28611
rect 15853 28577 15887 28611
rect 16681 28577 16715 28611
rect 28181 28577 28215 28611
rect 1593 28509 1627 28543
rect 8401 28509 8435 28543
rect 9413 28509 9447 28543
rect 9873 28509 9907 28543
rect 10057 28509 10091 28543
rect 11509 28509 11543 28543
rect 13277 28509 13311 28543
rect 13553 28509 13587 28543
rect 14105 28509 14139 28543
rect 14749 28509 14783 28543
rect 14933 28509 14967 28543
rect 16037 28509 16071 28543
rect 17003 28509 17037 28543
rect 17969 28509 18003 28543
rect 18153 28509 18187 28543
rect 18245 28509 18279 28543
rect 20453 28509 20487 28543
rect 20729 28509 20763 28543
rect 21741 28509 21775 28543
rect 23857 28509 23891 28543
rect 24409 28509 24443 28543
rect 26341 28509 26375 28543
rect 9965 28441 9999 28475
rect 10609 28441 10643 28475
rect 15117 28441 15151 28475
rect 19625 28441 19659 28475
rect 19809 28441 19843 28475
rect 21986 28441 22020 28475
rect 23673 28441 23707 28475
rect 24654 28441 24688 28475
rect 26065 28441 26099 28475
rect 26525 28441 26559 28475
rect 8217 28373 8251 28407
rect 9229 28373 9263 28407
rect 12633 28373 12667 28407
rect 13093 28373 13127 28407
rect 14197 28373 14231 28407
rect 18429 28373 18463 28407
rect 19993 28373 20027 28407
rect 25789 28373 25823 28407
rect 8217 28169 8251 28203
rect 12357 28169 12391 28203
rect 13553 28169 13587 28203
rect 15577 28169 15611 28203
rect 28089 28169 28123 28203
rect 10977 28101 11011 28135
rect 14442 28101 14476 28135
rect 17386 28101 17420 28135
rect 21925 28101 21959 28135
rect 26985 28101 27019 28135
rect 8401 28033 8435 28067
rect 9505 28033 9539 28067
rect 10149 28033 10183 28067
rect 10793 28033 10827 28067
rect 12081 28033 12115 28067
rect 12173 28033 12207 28067
rect 13277 28033 13311 28067
rect 13645 28033 13679 28067
rect 13737 28033 13771 28067
rect 18981 28033 19015 28067
rect 19237 28033 19271 28067
rect 21097 28033 21131 28067
rect 21841 28031 21875 28065
rect 22744 28033 22778 28067
rect 24317 28033 24351 28067
rect 25309 28033 25343 28067
rect 27169 28033 27203 28067
rect 27353 28033 27387 28067
rect 27905 28033 27939 28067
rect 10609 27965 10643 27999
rect 13369 27965 13403 27999
rect 14197 27965 14231 27999
rect 17141 27965 17175 27999
rect 20913 27965 20947 27999
rect 22477 27965 22511 27999
rect 25053 27965 25087 27999
rect 27445 27965 27479 27999
rect 9321 27897 9355 27931
rect 18521 27897 18555 27931
rect 20361 27897 20395 27931
rect 9965 27829 9999 27863
rect 13093 27829 13127 27863
rect 21281 27829 21315 27863
rect 23857 27829 23891 27863
rect 24501 27829 24535 27863
rect 26433 27829 26467 27863
rect 13093 27625 13127 27659
rect 13553 27625 13587 27659
rect 23305 27625 23339 27659
rect 8217 27557 8251 27591
rect 9321 27557 9355 27591
rect 17693 27557 17727 27591
rect 25881 27557 25915 27591
rect 13185 27489 13219 27523
rect 16313 27489 16347 27523
rect 18337 27489 18371 27523
rect 18429 27489 18463 27523
rect 26525 27489 26559 27523
rect 8401 27421 8435 27455
rect 9505 27421 9539 27455
rect 10149 27421 10183 27455
rect 10609 27421 10643 27455
rect 10793 27421 10827 27455
rect 11253 27421 11287 27455
rect 13369 27421 13403 27455
rect 14105 27421 14139 27455
rect 18521 27421 18555 27455
rect 18613 27421 18647 27455
rect 22293 27421 22327 27455
rect 22569 27421 22603 27455
rect 24501 27421 24535 27455
rect 26341 27421 26375 27455
rect 11509 27353 11543 27387
rect 13093 27353 13127 27387
rect 14350 27353 14384 27387
rect 16558 27353 16592 27387
rect 19625 27353 19659 27387
rect 22109 27353 22143 27387
rect 23121 27353 23155 27387
rect 24768 27353 24802 27387
rect 28181 27353 28215 27387
rect 9965 27285 9999 27319
rect 10701 27285 10735 27319
rect 12633 27285 12667 27319
rect 15485 27285 15519 27319
rect 18153 27285 18187 27319
rect 20913 27285 20947 27319
rect 22477 27285 22511 27319
rect 23321 27285 23355 27319
rect 23489 27285 23523 27319
rect 18797 27081 18831 27115
rect 25421 27081 25455 27115
rect 11805 27013 11839 27047
rect 12021 27013 12055 27047
rect 17969 27013 18003 27047
rect 19594 27013 19628 27047
rect 27813 27013 27847 27047
rect 10333 26945 10367 26979
rect 10793 26945 10827 26979
rect 10977 26945 11011 26979
rect 12817 26945 12851 26979
rect 12909 26945 12943 26979
rect 13001 26945 13035 26979
rect 13645 26945 13679 26979
rect 13921 26945 13955 26979
rect 14841 26945 14875 26979
rect 15945 26945 15979 26979
rect 16957 26945 16991 26979
rect 17049 26945 17083 26979
rect 17877 26945 17911 26979
rect 18061 26945 18095 26979
rect 18245 26945 18279 26979
rect 18705 26945 18739 26979
rect 22017 26945 22051 26979
rect 22109 26945 22143 26979
rect 22385 26945 22419 26979
rect 22937 26945 22971 26979
rect 23848 26945 23882 26979
rect 25605 26945 25639 26979
rect 25881 26945 25915 26979
rect 27445 26945 27479 26979
rect 10885 26877 10919 26911
rect 13737 26877 13771 26911
rect 15761 26877 15795 26911
rect 19349 26877 19383 26911
rect 23581 26877 23615 26911
rect 9689 26809 9723 26843
rect 12173 26809 12207 26843
rect 12633 26809 12667 26843
rect 13185 26809 13219 26843
rect 15117 26809 15151 26843
rect 17233 26809 17267 26843
rect 17693 26809 17727 26843
rect 23121 26809 23155 26843
rect 25789 26809 25823 26843
rect 9045 26741 9079 26775
rect 10149 26741 10183 26775
rect 11989 26741 12023 26775
rect 13645 26741 13679 26775
rect 14105 26741 14139 26775
rect 15301 26741 15335 26775
rect 16129 26741 16163 26775
rect 20729 26741 20763 26775
rect 21833 26741 21867 26775
rect 22293 26741 22327 26775
rect 24961 26741 24995 26775
rect 10057 26537 10091 26571
rect 13553 26537 13587 26571
rect 14105 26537 14139 26571
rect 18429 26537 18463 26571
rect 19533 26537 19567 26571
rect 21741 26537 21775 26571
rect 23857 26537 23891 26571
rect 24777 26537 24811 26571
rect 24961 26537 24995 26571
rect 25789 26537 25823 26571
rect 15209 26469 15243 26503
rect 17141 26469 17175 26503
rect 22477 26469 22511 26503
rect 12173 26401 12207 26435
rect 14841 26401 14875 26435
rect 15761 26401 15795 26435
rect 18337 26401 18371 26435
rect 21465 26401 21499 26435
rect 23397 26401 23431 26435
rect 23489 26401 23523 26435
rect 26525 26401 26559 26435
rect 28181 26401 28215 26435
rect 9597 26333 9631 26367
rect 10241 26333 10275 26367
rect 10885 26333 10919 26367
rect 11345 26333 11379 26367
rect 11529 26333 11563 26367
rect 14381 26333 14415 26367
rect 16017 26333 16051 26367
rect 17601 26333 17635 26367
rect 17693 26333 17727 26367
rect 18521 26333 18555 26367
rect 19809 26333 19843 26367
rect 19898 26327 19932 26361
rect 19993 26333 20027 26367
rect 20177 26333 20211 26367
rect 21097 26333 21131 26367
rect 23121 26333 23155 26367
rect 23305 26333 23339 26367
rect 23673 26333 23707 26367
rect 25605 26333 25639 26367
rect 25881 26333 25915 26367
rect 26341 26333 26375 26367
rect 24823 26299 24857 26333
rect 12440 26265 12474 26299
rect 14105 26265 14139 26299
rect 18245 26265 18279 26299
rect 21582 26265 21616 26299
rect 22201 26265 22235 26299
rect 24593 26265 24627 26299
rect 10701 26197 10735 26231
rect 11713 26197 11747 26231
rect 14289 26197 14323 26231
rect 15301 26197 15335 26231
rect 18705 26197 18739 26231
rect 21373 26197 21407 26231
rect 22661 26197 22695 26231
rect 25421 26197 25455 26231
rect 9505 25993 9539 26027
rect 10149 25993 10183 26027
rect 21281 25993 21315 26027
rect 27353 25993 27387 26027
rect 28181 25993 28215 26027
rect 15878 25925 15912 25959
rect 18766 25925 18800 25959
rect 27813 25925 27847 25959
rect 28013 25925 28047 25959
rect 9689 25857 9723 25891
rect 10333 25857 10367 25891
rect 10793 25857 10827 25891
rect 10885 25857 10919 25891
rect 11529 25857 11563 25891
rect 11785 25857 11819 25891
rect 13820 25857 13854 25891
rect 15393 25857 15427 25891
rect 16681 25857 16715 25891
rect 16937 25857 16971 25891
rect 18521 25857 18555 25891
rect 20821 25857 20855 25891
rect 21925 25857 21959 25891
rect 22109 25857 22143 25891
rect 22293 25857 22327 25891
rect 22477 25857 22511 25891
rect 23397 25857 23431 25891
rect 24225 25857 24259 25891
rect 24409 25857 24443 25891
rect 25309 25857 25343 25891
rect 27169 25857 27203 25891
rect 13553 25789 13587 25823
rect 15669 25789 15703 25823
rect 15761 25789 15795 25823
rect 22201 25789 22235 25823
rect 23305 25789 23339 25823
rect 25053 25789 25087 25823
rect 26985 25789 27019 25823
rect 12909 25721 12943 25755
rect 16037 25721 16071 25755
rect 21097 25721 21131 25755
rect 26433 25721 26467 25755
rect 14933 25653 14967 25687
rect 18061 25653 18095 25687
rect 19901 25653 19935 25687
rect 22661 25653 22695 25687
rect 23765 25653 23799 25687
rect 24593 25653 24627 25687
rect 27997 25653 28031 25687
rect 9505 25449 9539 25483
rect 21373 25449 21407 25483
rect 23305 25449 23339 25483
rect 24685 25449 24719 25483
rect 12817 25381 12851 25415
rect 18705 25381 18739 25415
rect 10885 25313 10919 25347
rect 11437 25313 11471 25347
rect 15402 25313 15436 25347
rect 16405 25313 16439 25347
rect 19993 25313 20027 25347
rect 23673 25313 23707 25347
rect 28181 25313 28215 25347
rect 9689 25245 9723 25279
rect 10333 25245 10367 25279
rect 10793 25245 10827 25279
rect 10977 25245 11011 25279
rect 14289 25245 14323 25279
rect 14381 25245 14415 25279
rect 14565 25245 14599 25279
rect 14657 25245 14691 25279
rect 15117 25245 15151 25279
rect 15301 25245 15335 25279
rect 15531 25245 15565 25279
rect 15669 25245 15703 25279
rect 16661 25245 16695 25279
rect 18429 25245 18463 25279
rect 18524 25245 18558 25279
rect 19257 25245 19291 25279
rect 22201 25245 22235 25279
rect 22366 25245 22400 25279
rect 22477 25245 22511 25279
rect 22569 25245 22603 25279
rect 23489 25245 23523 25279
rect 23581 25245 23615 25279
rect 23765 25245 23799 25279
rect 24961 25245 24995 25279
rect 25053 25245 25087 25279
rect 25145 25245 25179 25279
rect 25329 25245 25363 25279
rect 26341 25245 26375 25279
rect 11682 25177 11716 25211
rect 13369 25177 13403 25211
rect 13553 25177 13587 25211
rect 20238 25177 20272 25211
rect 26525 25177 26559 25211
rect 10149 25109 10183 25143
rect 14105 25109 14139 25143
rect 15853 25109 15887 25143
rect 17785 25109 17819 25143
rect 19441 25109 19475 25143
rect 22017 25109 22051 25143
rect 13093 24905 13127 24939
rect 13737 24905 13771 24939
rect 17049 24905 17083 24939
rect 26341 24905 26375 24939
rect 14381 24837 14415 24871
rect 19441 24837 19475 24871
rect 22569 24837 22603 24871
rect 23673 24837 23707 24871
rect 10333 24769 10367 24803
rect 10793 24769 10827 24803
rect 10977 24769 11011 24803
rect 12081 24769 12115 24803
rect 12909 24769 12943 24803
rect 13645 24769 13679 24803
rect 15025 24769 15059 24803
rect 15209 24769 15243 24803
rect 15301 24769 15335 24803
rect 15577 24769 15611 24803
rect 16865 24769 16899 24803
rect 17141 24769 17175 24803
rect 17601 24769 17635 24803
rect 18245 24769 18279 24803
rect 18429 24769 18463 24803
rect 19257 24769 19291 24803
rect 20453 24769 20487 24803
rect 20637 24769 20671 24803
rect 21097 24769 21131 24803
rect 22385 24769 22419 24803
rect 22661 24769 22695 24803
rect 23857 24769 23891 24803
rect 25145 24769 25179 24803
rect 26157 24769 26191 24803
rect 26433 24769 26467 24803
rect 27169 24769 27203 24803
rect 27997 24769 28031 24803
rect 11897 24701 11931 24735
rect 12725 24701 12759 24735
rect 19073 24701 19107 24735
rect 20269 24701 20303 24735
rect 21189 24701 21223 24735
rect 24133 24701 24167 24735
rect 25053 24701 25087 24735
rect 25513 24701 25547 24735
rect 27077 24701 27111 24735
rect 10149 24633 10183 24667
rect 17693 24633 17727 24667
rect 22201 24633 22235 24667
rect 28089 24633 28123 24667
rect 10793 24565 10827 24599
rect 12265 24565 12299 24599
rect 14473 24565 14507 24599
rect 15485 24565 15519 24599
rect 16681 24565 16715 24599
rect 18613 24565 18647 24599
rect 24041 24565 24075 24599
rect 25973 24565 26007 24599
rect 27537 24565 27571 24599
rect 12633 24361 12667 24395
rect 22569 24361 22603 24395
rect 11437 24293 11471 24327
rect 12081 24293 12115 24327
rect 17417 24293 17451 24327
rect 20637 24293 20671 24327
rect 13369 24225 13403 24259
rect 13553 24225 13587 24259
rect 15117 24225 15151 24259
rect 16037 24225 16071 24259
rect 23121 24225 23155 24259
rect 23581 24225 23615 24259
rect 24585 24225 24619 24259
rect 24685 24225 24719 24259
rect 24869 24225 24903 24259
rect 28181 24225 28215 24259
rect 10241 24157 10275 24191
rect 10701 24157 10735 24191
rect 10885 24157 10919 24191
rect 11345 24157 11379 24191
rect 11529 24157 11563 24191
rect 11989 24157 12023 24191
rect 12173 24157 12207 24191
rect 12817 24157 12851 24191
rect 13277 24157 13311 24191
rect 14473 24157 14507 24191
rect 15301 24157 15335 24191
rect 15577 24157 15611 24191
rect 18337 24157 18371 24191
rect 18426 24157 18460 24191
rect 18521 24157 18555 24191
rect 18705 24157 18739 24191
rect 19257 24157 19291 24191
rect 21189 24157 21223 24191
rect 23213 24157 23247 24191
rect 24777 24157 24811 24191
rect 25605 24157 25639 24191
rect 26341 24157 26375 24191
rect 10793 24089 10827 24123
rect 16282 24089 16316 24123
rect 18061 24089 18095 24123
rect 19502 24089 19536 24123
rect 21456 24089 21490 24123
rect 25421 24089 25455 24123
rect 26525 24089 26559 24123
rect 13553 24021 13587 24055
rect 14565 24021 14599 24055
rect 15485 24021 15519 24055
rect 24409 24021 24443 24055
rect 25789 24021 25823 24055
rect 9689 23817 9723 23851
rect 13835 23817 13869 23851
rect 15761 23817 15795 23851
rect 18521 23817 18555 23851
rect 21833 23817 21867 23851
rect 24501 23817 24535 23851
rect 26433 23817 26467 23851
rect 28089 23817 28123 23851
rect 13185 23749 13219 23783
rect 18981 23749 19015 23783
rect 20913 23749 20947 23783
rect 23581 23749 23615 23783
rect 9505 23681 9539 23715
rect 9689 23681 9723 23715
rect 10149 23681 10183 23715
rect 10333 23681 10367 23715
rect 10793 23681 10827 23715
rect 10977 23681 11011 23715
rect 11805 23681 11839 23715
rect 11989 23681 12023 23715
rect 12449 23681 12483 23715
rect 12633 23681 12667 23715
rect 13093 23681 13127 23715
rect 13277 23681 13311 23715
rect 13737 23681 13771 23715
rect 13921 23681 13955 23715
rect 14013 23681 14047 23715
rect 14565 23681 14599 23715
rect 14749 23681 14783 23715
rect 15393 23681 15427 23715
rect 18153 23681 18187 23715
rect 19165 23681 19199 23715
rect 20269 23681 20303 23715
rect 20453 23681 20487 23715
rect 21097 23681 21131 23715
rect 22109 23681 22143 23715
rect 22201 23681 22235 23715
rect 22293 23681 22327 23715
rect 22477 23681 22511 23715
rect 23397 23681 23431 23715
rect 23673 23681 23707 23715
rect 24317 23681 24351 23715
rect 24593 23681 24627 23715
rect 25053 23681 25087 23715
rect 25320 23681 25354 23715
rect 27169 23681 27203 23715
rect 27997 23681 28031 23715
rect 12541 23613 12575 23647
rect 15301 23613 15335 23647
rect 16681 23613 16715 23647
rect 16957 23613 16991 23647
rect 18061 23613 18095 23647
rect 19349 23613 19383 23647
rect 20085 23613 20119 23647
rect 27261 23613 27295 23647
rect 10793 23545 10827 23579
rect 19257 23545 19291 23579
rect 19441 23545 19475 23579
rect 1961 23477 1995 23511
rect 10241 23477 10275 23511
rect 11805 23477 11839 23511
rect 21281 23477 21315 23511
rect 23213 23477 23247 23511
rect 24133 23477 24167 23511
rect 27445 23477 27479 23511
rect 11345 23273 11379 23307
rect 13461 23273 13495 23307
rect 18245 23273 18279 23307
rect 15485 23205 15519 23239
rect 16129 23205 16163 23239
rect 17785 23205 17819 23239
rect 21925 23205 21959 23239
rect 1409 23137 1443 23171
rect 2789 23137 2823 23171
rect 14105 23137 14139 23171
rect 17325 23137 17359 23171
rect 19993 23137 20027 23171
rect 23673 23137 23707 23171
rect 25605 23137 25639 23171
rect 26341 23137 26375 23171
rect 28181 23137 28215 23171
rect 10701 23069 10735 23103
rect 10885 23069 10919 23103
rect 11345 23069 11379 23103
rect 11529 23069 11563 23103
rect 11989 23069 12023 23103
rect 12173 23069 12207 23103
rect 12633 23069 12667 23103
rect 13369 23069 13403 23103
rect 16405 23069 16439 23103
rect 16497 23069 16531 23103
rect 16589 23069 16623 23103
rect 16785 23069 16819 23103
rect 17417 23069 17451 23103
rect 18429 23069 18463 23103
rect 18705 23069 18739 23103
rect 19533 23069 19567 23103
rect 22109 23069 22143 23103
rect 22293 23069 22327 23103
rect 22385 23069 22419 23103
rect 23489 23069 23523 23103
rect 23581 23069 23615 23103
rect 23765 23069 23799 23103
rect 24409 23069 24443 23103
rect 24501 23069 24535 23103
rect 25513 23069 25547 23103
rect 1593 23001 1627 23035
rect 12081 23001 12115 23035
rect 14372 23001 14406 23035
rect 19257 23001 19291 23035
rect 20260 23001 20294 23035
rect 24685 23001 24719 23035
rect 26525 23001 26559 23035
rect 10793 22933 10827 22967
rect 12725 22933 12759 22967
rect 18613 22933 18647 22967
rect 19355 22933 19389 22967
rect 19441 22933 19475 22967
rect 21373 22933 21407 22967
rect 23305 22933 23339 22967
rect 24409 22933 24443 22967
rect 25145 22933 25179 22967
rect 25789 22933 25823 22967
rect 2513 22729 2547 22763
rect 13461 22729 13495 22763
rect 16129 22729 16163 22763
rect 17877 22729 17911 22763
rect 21833 22729 21867 22763
rect 10885 22661 10919 22695
rect 2421 22593 2455 22627
rect 10793 22593 10827 22627
rect 10977 22593 11011 22627
rect 11989 22593 12023 22627
rect 12633 22593 12667 22627
rect 13277 22593 13311 22627
rect 13553 22593 13587 22627
rect 14105 22593 14139 22627
rect 14933 22593 14967 22627
rect 15209 22593 15243 22627
rect 15761 22593 15795 22627
rect 15945 22593 15979 22627
rect 16681 22593 16715 22627
rect 17509 22593 17543 22627
rect 18613 22593 18647 22627
rect 18880 22593 18914 22627
rect 20637 22593 20671 22627
rect 20729 22593 20763 22627
rect 21005 22593 21039 22627
rect 22017 22593 22051 22627
rect 23213 22593 23247 22627
rect 23305 22593 23339 22627
rect 23397 22593 23431 22627
rect 23581 22593 23615 22627
rect 24225 22593 24259 22627
rect 25309 22593 25343 22627
rect 27169 22593 27203 22627
rect 27997 22593 28031 22627
rect 14289 22525 14323 22559
rect 14749 22525 14783 22559
rect 17601 22525 17635 22559
rect 20913 22525 20947 22559
rect 22293 22525 22327 22559
rect 24133 22525 24167 22559
rect 25053 22525 25087 22559
rect 27077 22525 27111 22559
rect 13277 22457 13311 22491
rect 24593 22457 24627 22491
rect 12081 22389 12115 22423
rect 12725 22389 12759 22423
rect 15117 22389 15151 22423
rect 16773 22389 16807 22423
rect 19993 22389 20027 22423
rect 20453 22389 20487 22423
rect 22201 22389 22235 22423
rect 22937 22389 22971 22423
rect 26433 22389 26467 22423
rect 27445 22389 27479 22423
rect 28089 22389 28123 22423
rect 15393 22185 15427 22219
rect 25697 22185 25731 22219
rect 18061 22117 18095 22151
rect 11989 22049 12023 22083
rect 14545 22049 14579 22083
rect 16109 22049 16143 22083
rect 19257 22049 19291 22083
rect 19625 22049 19659 22083
rect 20085 22049 20119 22083
rect 20453 22049 20487 22083
rect 23857 22049 23891 22083
rect 26525 22049 26559 22083
rect 28181 22049 28215 22083
rect 11253 21981 11287 22015
rect 11621 21981 11655 22015
rect 11897 21981 11931 22015
rect 12081 21981 12115 22015
rect 12633 21981 12667 22015
rect 13369 21981 13403 22015
rect 14657 21981 14691 22015
rect 14749 21959 14783 21993
rect 16313 21981 16347 22015
rect 17693 21981 17727 22015
rect 17877 21981 17911 22015
rect 18153 21981 18187 22015
rect 19441 21981 19475 22015
rect 20545 21981 20579 22015
rect 20913 21981 20947 22015
rect 21005 21981 21039 22015
rect 21741 21981 21775 22015
rect 23673 21981 23707 22015
rect 24685 21981 24719 22015
rect 24777 21981 24811 22015
rect 24869 21981 24903 22015
rect 25053 21981 25087 22015
rect 26341 21981 26375 22015
rect 12817 21913 12851 21947
rect 13553 21913 13587 21947
rect 14473 21913 14507 21947
rect 15209 21913 15243 21947
rect 16037 21913 16071 21947
rect 16773 21913 16807 21947
rect 16957 21913 16991 21947
rect 17141 21913 17175 21947
rect 20269 21913 20303 21947
rect 21986 21913 22020 21947
rect 25513 21913 25547 21947
rect 25729 21913 25763 21947
rect 15409 21845 15443 21879
rect 15577 21845 15611 21879
rect 16221 21845 16255 21879
rect 23121 21845 23155 21879
rect 24409 21845 24443 21879
rect 25881 21845 25915 21879
rect 16957 21641 16991 21675
rect 18521 21641 18555 21675
rect 19073 21641 19107 21675
rect 26985 21641 27019 21675
rect 13369 21573 13403 21607
rect 14105 21573 14139 21607
rect 15669 21573 15703 21607
rect 15853 21573 15887 21607
rect 18981 21573 19015 21607
rect 20361 21573 20395 21607
rect 20561 21573 20595 21607
rect 28089 21573 28123 21607
rect 11805 21505 11839 21539
rect 11989 21505 12023 21539
rect 12449 21505 12483 21539
rect 12633 21505 12667 21539
rect 13185 21505 13219 21539
rect 13921 21505 13955 21539
rect 14841 21505 14875 21539
rect 14933 21505 14967 21539
rect 15025 21505 15059 21539
rect 15209 21505 15243 21539
rect 17133 21505 17167 21539
rect 17417 21505 17451 21539
rect 18153 21505 18187 21539
rect 21833 21505 21867 21539
rect 22017 21505 22051 21539
rect 22201 21505 22235 21539
rect 22293 21505 22327 21539
rect 22753 21505 22787 21539
rect 23020 21505 23054 21539
rect 27169 21505 27203 21539
rect 27905 21505 27939 21539
rect 28181 21505 28215 21539
rect 11897 21437 11931 21471
rect 17233 21437 17267 21471
rect 17325 21437 17359 21471
rect 18061 21437 18095 21471
rect 19349 21437 19383 21471
rect 24593 21437 24627 21471
rect 24777 21437 24811 21471
rect 26157 21437 26191 21471
rect 27445 21437 27479 21471
rect 12541 21369 12575 21403
rect 14565 21301 14599 21335
rect 16037 21301 16071 21335
rect 19257 21301 19291 21335
rect 19349 21301 19383 21335
rect 20545 21301 20579 21335
rect 20729 21301 20763 21335
rect 24133 21301 24167 21335
rect 27353 21301 27387 21335
rect 27905 21301 27939 21335
rect 13369 21097 13403 21131
rect 15485 21097 15519 21131
rect 20177 21097 20211 21131
rect 25513 21097 25547 21131
rect 12081 21029 12115 21063
rect 14105 21029 14139 21063
rect 14841 20961 14875 20995
rect 15209 20961 15243 20995
rect 15301 20961 15335 20995
rect 17785 20961 17819 20995
rect 22753 20931 22787 20965
rect 25237 20961 25271 20995
rect 26525 20961 26559 20995
rect 28181 20961 28215 20995
rect 12081 20893 12115 20927
rect 12265 20893 12299 20927
rect 12725 20893 12759 20927
rect 12909 20893 12943 20927
rect 13369 20893 13403 20927
rect 13547 20893 13581 20927
rect 14381 20893 14415 20927
rect 16497 20893 16531 20927
rect 16589 20893 16623 20927
rect 16681 20893 16715 20927
rect 16865 20893 16899 20927
rect 17693 20893 17727 20927
rect 17969 20893 18003 20927
rect 18521 20893 18555 20927
rect 19533 20893 19567 20927
rect 19626 20893 19660 20927
rect 19901 20893 19935 20927
rect 20039 20893 20073 20927
rect 20637 20893 20671 20927
rect 22477 20893 22511 20927
rect 22569 20893 22603 20927
rect 23397 20893 23431 20927
rect 23581 20893 23615 20927
rect 23670 20903 23704 20937
rect 25145 20893 25179 20927
rect 26341 20893 26375 20927
rect 12817 20825 12851 20859
rect 14105 20825 14139 20859
rect 14289 20825 14323 20859
rect 19809 20825 19843 20859
rect 20904 20825 20938 20859
rect 23213 20825 23247 20859
rect 16221 20757 16255 20791
rect 17325 20757 17359 20791
rect 18613 20757 18647 20791
rect 22017 20757 22051 20791
rect 22753 20757 22787 20791
rect 17325 20553 17359 20587
rect 19717 20553 19751 20587
rect 21189 20553 21223 20587
rect 23305 20553 23339 20587
rect 27629 20553 27663 20587
rect 23029 20485 23063 20519
rect 27353 20485 27387 20519
rect 13369 20417 13403 20451
rect 13636 20417 13670 20451
rect 15485 20417 15519 20451
rect 15577 20417 15611 20451
rect 15669 20417 15703 20451
rect 15853 20417 15887 20451
rect 18337 20417 18371 20451
rect 18604 20417 18638 20451
rect 20361 20417 20395 20451
rect 21097 20417 21131 20451
rect 22017 20417 22051 20451
rect 22753 20417 22787 20451
rect 22937 20417 22971 20451
rect 23121 20417 23155 20451
rect 24501 20417 24535 20451
rect 24593 20417 24627 20451
rect 24869 20417 24903 20451
rect 25329 20417 25363 20451
rect 25513 20417 25547 20451
rect 25605 20417 25639 20451
rect 25881 20417 25915 20451
rect 26065 20417 26099 20451
rect 26985 20417 27019 20451
rect 27078 20417 27112 20451
rect 27261 20417 27295 20451
rect 27450 20417 27484 20451
rect 16681 20349 16715 20383
rect 17049 20349 17083 20383
rect 17141 20349 17175 20383
rect 20637 20349 20671 20383
rect 21833 20349 21867 20383
rect 25697 20349 25731 20383
rect 14749 20281 14783 20315
rect 22201 20281 22235 20315
rect 15209 20213 15243 20247
rect 20177 20213 20211 20247
rect 20545 20213 20579 20247
rect 24317 20213 24351 20247
rect 24777 20213 24811 20247
rect 14565 20009 14599 20043
rect 15485 20009 15519 20043
rect 15669 20009 15703 20043
rect 17693 20009 17727 20043
rect 18613 20009 18647 20043
rect 23121 20009 23155 20043
rect 13461 19941 13495 19975
rect 16313 19873 16347 19907
rect 18429 19873 18463 19907
rect 19441 19873 19475 19907
rect 21281 19873 21315 19907
rect 23581 19873 23615 19907
rect 26525 19873 26559 19907
rect 13369 19805 13403 19839
rect 13553 19805 13587 19839
rect 14381 19805 14415 19839
rect 14657 19805 14691 19839
rect 15117 19805 15151 19839
rect 15485 19805 15519 19839
rect 16569 19805 16603 19839
rect 18337 19805 18371 19839
rect 19708 19805 19742 19839
rect 23305 19805 23339 19839
rect 23397 19805 23431 19839
rect 23673 19805 23707 19839
rect 24409 19805 24443 19839
rect 24676 19805 24710 19839
rect 26341 19805 26375 19839
rect 28181 19805 28215 19839
rect 21548 19737 21582 19771
rect 14197 19669 14231 19703
rect 20821 19669 20855 19703
rect 22661 19669 22695 19703
rect 25789 19669 25823 19703
rect 17785 19465 17819 19499
rect 18889 19465 18923 19499
rect 21097 19465 21131 19499
rect 24133 19465 24167 19499
rect 27445 19465 27479 19499
rect 18521 19397 18555 19431
rect 23857 19397 23891 19431
rect 27997 19397 28031 19431
rect 14473 19329 14507 19363
rect 15393 19329 15427 19363
rect 15485 19329 15519 19363
rect 16865 19329 16899 19363
rect 17693 19329 17727 19363
rect 18337 19329 18371 19363
rect 18613 19329 18647 19363
rect 18705 19329 18739 19363
rect 19349 19329 19383 19363
rect 19533 19329 19567 19363
rect 19717 19329 19751 19363
rect 19901 19329 19935 19363
rect 20821 19329 20855 19363
rect 22569 19329 22603 19363
rect 23581 19329 23615 19363
rect 23765 19329 23799 19363
rect 23949 19329 23983 19363
rect 25053 19329 25087 19363
rect 25320 19329 25354 19363
rect 26985 19329 27019 19363
rect 15117 19261 15151 19295
rect 15301 19261 15335 19295
rect 15577 19261 15611 19295
rect 16957 19261 16991 19295
rect 19625 19261 19659 19295
rect 20085 19261 20119 19295
rect 20913 19261 20947 19295
rect 21097 19261 21131 19295
rect 22293 19261 22327 19295
rect 14565 19125 14599 19159
rect 17141 19125 17175 19159
rect 26433 19125 26467 19159
rect 27077 19125 27111 19159
rect 28089 19125 28123 19159
rect 16405 18921 16439 18955
rect 19625 18921 19659 18955
rect 20269 18921 20303 18955
rect 23765 18921 23799 18955
rect 15577 18853 15611 18887
rect 17969 18853 18003 18887
rect 15117 18785 15151 18819
rect 21189 18785 21223 18819
rect 22569 18785 22603 18819
rect 28181 18785 28215 18819
rect 14381 18717 14415 18751
rect 14473 18717 14507 18751
rect 15209 18717 15243 18751
rect 17141 18717 17175 18751
rect 17233 18717 17267 18751
rect 17417 18717 17451 18751
rect 17509 18717 17543 18751
rect 18245 18717 18279 18751
rect 19441 18717 19475 18751
rect 20913 18717 20947 18751
rect 21005 18717 21039 18751
rect 21741 18717 21775 18751
rect 21925 18717 21959 18751
rect 22017 18717 22051 18751
rect 22477 18717 22511 18751
rect 23673 18717 23707 18751
rect 24869 18717 24903 18751
rect 25237 18717 25271 18751
rect 26341 18717 26375 18751
rect 16313 18649 16347 18683
rect 17969 18649 18003 18683
rect 19257 18649 19291 18683
rect 20085 18649 20119 18683
rect 21189 18649 21223 18683
rect 22753 18649 22787 18683
rect 25053 18649 25087 18683
rect 25145 18649 25179 18683
rect 26525 18649 26559 18683
rect 16957 18581 16991 18615
rect 18153 18581 18187 18615
rect 20285 18581 20319 18615
rect 20453 18581 20487 18615
rect 21839 18581 21873 18615
rect 22477 18581 22511 18615
rect 25421 18581 25455 18615
rect 13737 18377 13771 18411
rect 19165 18377 19199 18411
rect 21189 18377 21223 18411
rect 23121 18377 23155 18411
rect 24501 18377 24535 18411
rect 26985 18377 27019 18411
rect 16773 18309 16807 18343
rect 18797 18309 18831 18343
rect 22753 18309 22787 18343
rect 22953 18309 22987 18343
rect 24133 18309 24167 18343
rect 2329 18241 2363 18275
rect 13645 18241 13679 18275
rect 14289 18241 14323 18275
rect 14556 18241 14590 18275
rect 16681 18241 16715 18275
rect 17325 18241 17359 18275
rect 17509 18241 17543 18275
rect 17693 18241 17727 18275
rect 17877 18241 17911 18275
rect 18061 18241 18095 18275
rect 18521 18241 18555 18275
rect 18614 18241 18648 18275
rect 18889 18241 18923 18275
rect 19027 18241 19061 18275
rect 19809 18241 19843 18275
rect 20076 18241 20110 18275
rect 22017 18241 22051 18275
rect 24317 18241 24351 18275
rect 24593 18241 24627 18275
rect 25053 18241 25087 18275
rect 25320 18241 25354 18275
rect 27169 18241 27203 18275
rect 27905 18241 27939 18275
rect 17601 18173 17635 18207
rect 22293 18173 22327 18207
rect 27445 18173 27479 18207
rect 28181 18173 28215 18207
rect 15669 18105 15703 18139
rect 28089 18105 28123 18139
rect 1869 18037 1903 18071
rect 2421 18037 2455 18071
rect 21833 18037 21867 18071
rect 22201 18037 22235 18071
rect 22937 18037 22971 18071
rect 26433 18037 26467 18071
rect 27353 18037 27387 18071
rect 27997 18037 28031 18071
rect 17233 17833 17267 17867
rect 19441 17833 19475 17867
rect 20453 17833 20487 17867
rect 15393 17765 15427 17799
rect 19625 17765 19659 17799
rect 25789 17765 25823 17799
rect 1409 17697 1443 17731
rect 2789 17697 2823 17731
rect 14933 17697 14967 17731
rect 15853 17697 15887 17731
rect 17693 17697 17727 17731
rect 24409 17697 24443 17731
rect 28181 17697 28215 17731
rect 15025 17629 15059 17663
rect 17969 17629 18003 17663
rect 20085 17629 20119 17663
rect 20255 17629 20289 17663
rect 21005 17629 21039 17663
rect 21272 17629 21306 17663
rect 23581 17629 23615 17663
rect 23765 17629 23799 17663
rect 23857 17629 23891 17663
rect 26341 17629 26375 17663
rect 1593 17561 1627 17595
rect 16098 17561 16132 17595
rect 19257 17561 19291 17595
rect 23397 17561 23431 17595
rect 24654 17561 24688 17595
rect 26525 17561 26559 17595
rect 19457 17493 19491 17527
rect 22385 17493 22419 17527
rect 15669 17289 15703 17323
rect 19349 17289 19383 17323
rect 21189 17289 21223 17323
rect 23213 17289 23247 17323
rect 25513 17221 25547 17255
rect 25713 17221 25747 17255
rect 28089 17221 28123 17255
rect 15853 17153 15887 17187
rect 17969 17153 18003 17187
rect 18236 17153 18270 17187
rect 19809 17153 19843 17187
rect 20076 17153 20110 17187
rect 21833 17153 21867 17187
rect 22100 17153 22134 17187
rect 23673 17153 23707 17187
rect 23929 17153 23963 17187
rect 27169 17153 27203 17187
rect 27813 17153 27847 17187
rect 1409 17085 1443 17119
rect 1593 17085 1627 17119
rect 1869 17085 1903 17119
rect 16129 17085 16163 17119
rect 16681 17085 16715 17119
rect 16957 17085 16991 17119
rect 26985 17085 27019 17119
rect 27905 17085 27939 17119
rect 27813 17017 27847 17051
rect 16037 16949 16071 16983
rect 25053 16949 25087 16983
rect 25697 16949 25731 16983
rect 25881 16949 25915 16983
rect 27353 16949 27387 16983
rect 1777 16745 1811 16779
rect 2513 16745 2547 16779
rect 20453 16745 20487 16779
rect 21465 16745 21499 16779
rect 22109 16745 22143 16779
rect 16681 16609 16715 16643
rect 19809 16609 19843 16643
rect 19993 16609 20027 16643
rect 24501 16609 24535 16643
rect 1685 16551 1719 16585
rect 16037 16541 16071 16575
rect 16129 16541 16163 16575
rect 18521 16541 18555 16575
rect 19717 16541 19751 16575
rect 20453 16541 20487 16575
rect 20637 16541 20671 16575
rect 21465 16541 21499 16575
rect 21649 16541 21683 16575
rect 22385 16541 22419 16575
rect 23397 16541 23431 16575
rect 23581 16541 23615 16575
rect 24768 16541 24802 16575
rect 26341 16541 26375 16575
rect 16948 16473 16982 16507
rect 18613 16473 18647 16507
rect 19993 16473 20027 16507
rect 22109 16473 22143 16507
rect 23765 16473 23799 16507
rect 26525 16473 26559 16507
rect 28181 16473 28215 16507
rect 18061 16405 18095 16439
rect 22293 16405 22327 16439
rect 25881 16405 25915 16439
rect 17049 16201 17083 16235
rect 18153 16201 18187 16235
rect 20177 16201 20211 16235
rect 20913 16201 20947 16235
rect 22201 16201 22235 16235
rect 27537 16201 27571 16235
rect 16865 16133 16899 16167
rect 18429 16133 18463 16167
rect 24777 16133 24811 16167
rect 17141 16065 17175 16099
rect 18153 16065 18187 16099
rect 20085 16065 20119 16099
rect 20269 16065 20303 16099
rect 20821 16065 20855 16099
rect 21005 16065 21039 16099
rect 22017 16065 22051 16099
rect 22201 16065 22235 16099
rect 22661 16065 22695 16099
rect 23305 16065 23339 16099
rect 27445 16065 27479 16099
rect 18245 15997 18279 16031
rect 23581 15997 23615 16031
rect 24593 15997 24627 16031
rect 26157 15997 26191 16031
rect 16865 15929 16899 15963
rect 22753 15929 22787 15963
rect 23397 15929 23431 15963
rect 1593 15861 1627 15895
rect 23489 15861 23523 15895
rect 17141 15657 17175 15691
rect 22937 15657 22971 15691
rect 25145 15657 25179 15691
rect 22477 15589 22511 15623
rect 23857 15589 23891 15623
rect 1409 15521 1443 15555
rect 2789 15521 2823 15555
rect 17141 15453 17175 15487
rect 17325 15453 17359 15487
rect 22937 15453 22971 15487
rect 23121 15453 23155 15487
rect 24685 15453 24719 15487
rect 25421 15453 25455 15487
rect 26341 15453 26375 15487
rect 1593 15385 1627 15419
rect 23673 15385 23707 15419
rect 24409 15385 24443 15419
rect 25145 15385 25179 15419
rect 25329 15385 25363 15419
rect 26525 15385 26559 15419
rect 28181 15385 28215 15419
rect 24507 15317 24541 15351
rect 24593 15317 24627 15351
rect 1685 15113 1719 15147
rect 23765 15113 23799 15147
rect 25053 15113 25087 15147
rect 25697 15113 25731 15147
rect 26341 15113 26375 15147
rect 27169 15113 27203 15147
rect 1593 14977 1627 15011
rect 23673 14977 23707 15011
rect 24501 14977 24535 15011
rect 24961 14977 24995 15011
rect 25605 14977 25639 15011
rect 26249 14977 26283 15011
rect 27077 14977 27111 15011
rect 27721 14977 27755 15011
rect 27997 14909 28031 14943
rect 27905 14841 27939 14875
rect 2421 14773 2455 14807
rect 27813 14773 27847 14807
rect 24961 14569 24995 14603
rect 25697 14569 25731 14603
rect 23857 14501 23891 14535
rect 1409 14433 1443 14467
rect 1869 14433 1903 14467
rect 26341 14433 26375 14467
rect 24869 14365 24903 14399
rect 25605 14365 25639 14399
rect 1593 14297 1627 14331
rect 26525 14297 26559 14331
rect 28181 14297 28215 14331
rect 1869 14025 1903 14059
rect 25789 14025 25823 14059
rect 27169 14025 27203 14059
rect 27813 14025 27847 14059
rect 1777 13889 1811 13923
rect 25237 13889 25271 13923
rect 25697 13889 25731 13923
rect 27077 13889 27111 13923
rect 27721 13889 27755 13923
rect 25605 13481 25639 13515
rect 26065 13481 26099 13515
rect 27169 13481 27203 13515
rect 27905 13481 27939 13515
rect 1593 13277 1627 13311
rect 2421 13277 2455 13311
rect 3065 13277 3099 13311
rect 26065 13277 26099 13311
rect 26249 13277 26283 13311
rect 27353 13277 27387 13311
rect 27813 13277 27847 13311
rect 1685 13141 1719 13175
rect 1593 12869 1627 12903
rect 1409 12801 1443 12835
rect 26433 12801 26467 12835
rect 27445 12801 27479 12835
rect 2789 12733 2823 12767
rect 28089 12733 28123 12767
rect 28089 12393 28123 12427
rect 1409 12257 1443 12291
rect 2789 12257 2823 12291
rect 27445 12189 27479 12223
rect 1593 12121 1627 12155
rect 2513 11849 2547 11883
rect 1777 11713 1811 11747
rect 2421 11713 2455 11747
rect 27261 11713 27295 11747
rect 27997 11713 28031 11747
rect 28181 11577 28215 11611
rect 1869 11509 1903 11543
rect 3249 11509 3283 11543
rect 27353 11509 27387 11543
rect 1409 11169 1443 11203
rect 1593 11169 1627 11203
rect 1869 11169 1903 11203
rect 26341 11169 26375 11203
rect 26525 11169 26559 11203
rect 3985 11101 4019 11135
rect 28181 11033 28215 11067
rect 1501 10625 1535 10659
rect 27813 10625 27847 10659
rect 1685 10557 1719 10591
rect 2881 10557 2915 10591
rect 27353 10421 27387 10455
rect 27905 10421 27939 10455
rect 1961 10217 1995 10251
rect 26525 10081 26559 10115
rect 1869 10013 1903 10047
rect 26341 10013 26375 10047
rect 28181 9945 28215 9979
rect 1593 9537 1627 9571
rect 27261 9537 27295 9571
rect 27721 9537 27755 9571
rect 1685 9333 1719 9367
rect 2421 9333 2455 9367
rect 27813 9333 27847 9367
rect 1409 8993 1443 9027
rect 1593 8993 1627 9027
rect 2789 8993 2823 9027
rect 26341 8993 26375 9027
rect 26525 8993 26559 9027
rect 28181 8993 28215 9027
rect 1869 8449 1903 8483
rect 2513 8449 2547 8483
rect 27905 8313 27939 8347
rect 1961 8245 1995 8279
rect 2605 8245 2639 8279
rect 3341 8245 3375 8279
rect 27261 8245 27295 8279
rect 1409 7905 1443 7939
rect 1593 7905 1627 7939
rect 2789 7905 2823 7939
rect 26341 7905 26375 7939
rect 3985 7837 4019 7871
rect 26525 7769 26559 7803
rect 28181 7769 28215 7803
rect 27813 7497 27847 7531
rect 2145 7429 2179 7463
rect 1961 7361 1995 7395
rect 27721 7361 27755 7395
rect 2973 7293 3007 7327
rect 4445 7157 4479 7191
rect 27261 7157 27295 7191
rect 1409 6817 1443 6851
rect 2881 6817 2915 6851
rect 26341 6817 26375 6851
rect 28181 6817 28215 6851
rect 3801 6749 3835 6783
rect 4629 6749 4663 6783
rect 1593 6681 1627 6715
rect 26525 6681 26559 6715
rect 3893 6613 3927 6647
rect 1961 6409 1995 6443
rect 2605 6409 2639 6443
rect 27905 6409 27939 6443
rect 3617 6341 3651 6375
rect 1961 6273 1995 6307
rect 2513 6273 2547 6307
rect 27169 6273 27203 6307
rect 27813 6273 27847 6307
rect 3433 6205 3467 6239
rect 4537 6205 4571 6239
rect 24593 6205 24627 6239
rect 24777 6205 24811 6239
rect 26065 6205 26099 6239
rect 27261 6069 27295 6103
rect 25237 5865 25271 5899
rect 5917 5797 5951 5831
rect 1409 5729 1443 5763
rect 1869 5729 1903 5763
rect 7205 5729 7239 5763
rect 26341 5729 26375 5763
rect 26525 5729 26559 5763
rect 28181 5729 28215 5763
rect 3801 5661 3835 5695
rect 4629 5661 4663 5695
rect 5273 5661 5307 5695
rect 6561 5661 6595 5695
rect 25881 5661 25915 5695
rect 1593 5593 1627 5627
rect 3893 5525 3927 5559
rect 1501 5321 1535 5355
rect 27905 5321 27939 5355
rect 2237 5253 2271 5287
rect 24777 5253 24811 5287
rect 27261 5253 27295 5287
rect 1409 5185 1443 5219
rect 2053 5185 2087 5219
rect 27169 5185 27203 5219
rect 27813 5185 27847 5219
rect 2789 5117 2823 5151
rect 24593 5117 24627 5151
rect 26157 5117 26191 5151
rect 6561 5049 6595 5083
rect 4537 4981 4571 5015
rect 5181 4981 5215 5015
rect 5825 4981 5859 5015
rect 7205 4981 7239 5015
rect 3801 4641 3835 4675
rect 1777 4573 1811 4607
rect 2421 4573 2455 4607
rect 3065 4573 3099 4607
rect 6285 4573 6319 4607
rect 7297 4573 7331 4607
rect 8125 4573 8159 4607
rect 9229 4573 9263 4607
rect 23857 4573 23891 4607
rect 25881 4573 25915 4607
rect 26341 4573 26375 4607
rect 3157 4505 3191 4539
rect 3985 4505 4019 4539
rect 5641 4505 5675 4539
rect 24869 4505 24903 4539
rect 26525 4505 26559 4539
rect 28181 4505 28215 4539
rect 1869 4437 1903 4471
rect 2513 4437 2547 4471
rect 7389 4437 7423 4471
rect 24961 4437 24995 4471
rect 1593 4165 1627 4199
rect 7389 4165 7423 4199
rect 1409 4097 1443 4131
rect 3709 4097 3743 4131
rect 9505 4097 9539 4131
rect 27169 4097 27203 4131
rect 27537 4097 27571 4131
rect 1869 4029 1903 4063
rect 3893 4029 3927 4063
rect 4169 4029 4203 4063
rect 7205 4029 7239 4063
rect 8217 4029 8251 4063
rect 13001 4029 13035 4063
rect 13185 4029 13219 4063
rect 13553 4029 13587 4063
rect 17509 4029 17543 4063
rect 17693 4029 17727 4063
rect 18061 4029 18095 4063
rect 23489 4029 23523 4063
rect 23673 4029 23707 4063
rect 25329 4029 25363 4063
rect 6745 3893 6779 3927
rect 9597 3893 9631 3927
rect 10333 3893 10367 3927
rect 15853 3893 15887 3927
rect 23029 3893 23063 3927
rect 25973 3893 26007 3927
rect 12541 3689 12575 3723
rect 13093 3689 13127 3723
rect 19257 3689 19291 3723
rect 23121 3689 23155 3723
rect 23857 3689 23891 3723
rect 1409 3553 1443 3587
rect 1593 3553 1627 3587
rect 3893 3553 3927 3587
rect 5365 3553 5399 3587
rect 5917 3553 5951 3587
rect 9137 3553 9171 3587
rect 9321 3553 9355 3587
rect 9689 3553 9723 3587
rect 15669 3553 15703 3587
rect 16129 3553 16163 3587
rect 25145 3553 25179 3587
rect 26157 3553 26191 3587
rect 3801 3485 3835 3519
rect 4721 3485 4755 3519
rect 7665 3485 7699 3519
rect 11897 3485 11931 3519
rect 13001 3485 13035 3519
rect 14473 3485 14507 3519
rect 18705 3485 18739 3519
rect 19441 3485 19475 3519
rect 19993 3485 20027 3519
rect 20821 3485 20855 3519
rect 21649 3485 21683 3519
rect 22109 3485 22143 3519
rect 23029 3485 23063 3519
rect 24501 3485 24535 3519
rect 27813 3485 27847 3519
rect 3249 3417 3283 3451
rect 5549 3417 5583 3451
rect 15853 3417 15887 3451
rect 24593 3417 24627 3451
rect 25329 3417 25363 3451
rect 4813 3349 4847 3383
rect 7757 3349 7791 3383
rect 20085 3349 20119 3383
rect 22201 3349 22235 3383
rect 27905 3349 27939 3383
rect 5457 3145 5491 3179
rect 27721 3145 27755 3179
rect 2513 3077 2547 3111
rect 7113 3077 7147 3111
rect 17693 3077 17727 3111
rect 22109 3077 22143 3111
rect 24777 3077 24811 3111
rect 1685 3009 1719 3043
rect 2329 3009 2363 3043
rect 4629 3009 4663 3043
rect 5365 3009 5399 3043
rect 6929 3009 6963 3043
rect 9689 3009 9723 3043
rect 11713 3009 11747 3043
rect 14197 3009 14231 3043
rect 17601 3009 17635 3043
rect 18245 3009 18279 3043
rect 18889 3009 18923 3043
rect 21925 3009 21959 3043
rect 26433 3009 26467 3043
rect 26985 3009 27019 3043
rect 27629 3009 27663 3043
rect 2789 2941 2823 2975
rect 7389 2941 7423 2975
rect 11897 2941 11931 2975
rect 12265 2941 12299 2975
rect 14381 2941 14415 2975
rect 14749 2941 14783 2975
rect 18337 2941 18371 2975
rect 19073 2941 19107 2975
rect 19349 2941 19383 2975
rect 22569 2941 22603 2975
rect 24593 2941 24627 2975
rect 27077 2941 27111 2975
rect 1777 2805 1811 2839
rect 4721 2805 4755 2839
rect 9781 2805 9815 2839
rect 11989 2601 12023 2635
rect 14473 2601 14507 2635
rect 15853 2601 15887 2635
rect 17233 2601 17267 2635
rect 17969 2601 18003 2635
rect 27169 2601 27203 2635
rect 1409 2465 1443 2499
rect 1593 2465 1627 2499
rect 2789 2465 2823 2499
rect 3985 2465 4019 2499
rect 4169 2465 4203 2499
rect 4537 2465 4571 2499
rect 6377 2465 6411 2499
rect 6561 2465 6595 2499
rect 6837 2465 6871 2499
rect 9045 2465 9079 2499
rect 9229 2465 9263 2499
rect 9873 2465 9907 2499
rect 19441 2465 19475 2499
rect 20177 2465 20211 2499
rect 22017 2465 22051 2499
rect 24593 2465 24627 2499
rect 24777 2465 24811 2499
rect 27905 2465 27939 2499
rect 11897 2397 11931 2431
rect 14381 2397 14415 2431
rect 15761 2397 15795 2431
rect 19257 2397 19291 2431
rect 27813 2397 27847 2431
rect 17141 2329 17175 2363
rect 22201 2329 22235 2363
rect 23857 2329 23891 2363
rect 26433 2329 26467 2363
<< metal1 >>
rect 9030 40808 9036 40860
rect 9088 40848 9094 40860
rect 23566 40848 23572 40860
rect 9088 40820 23572 40848
rect 9088 40808 9094 40820
rect 23566 40808 23572 40820
rect 23624 40808 23630 40860
rect 8846 40740 8852 40792
rect 8904 40780 8910 40792
rect 15930 40780 15936 40792
rect 8904 40752 15936 40780
rect 8904 40740 8910 40752
rect 15930 40740 15936 40752
rect 15988 40740 15994 40792
rect 7558 40672 7564 40724
rect 7616 40712 7622 40724
rect 13906 40712 13912 40724
rect 7616 40684 13912 40712
rect 7616 40672 7622 40684
rect 13906 40672 13912 40684
rect 13964 40672 13970 40724
rect 7650 40604 7656 40656
rect 7708 40644 7714 40656
rect 20346 40644 20352 40656
rect 7708 40616 20352 40644
rect 7708 40604 7714 40616
rect 20346 40604 20352 40616
rect 20404 40604 20410 40656
rect 7466 40536 7472 40588
rect 7524 40576 7530 40588
rect 23934 40576 23940 40588
rect 7524 40548 23940 40576
rect 7524 40536 7530 40548
rect 23934 40536 23940 40548
rect 23992 40536 23998 40588
rect 8938 40468 8944 40520
rect 8996 40508 9002 40520
rect 26878 40508 26884 40520
rect 8996 40480 26884 40508
rect 8996 40468 9002 40480
rect 26878 40468 26884 40480
rect 26936 40468 26942 40520
rect 7374 40400 7380 40452
rect 7432 40440 7438 40452
rect 22278 40440 22284 40452
rect 7432 40412 22284 40440
rect 7432 40400 7438 40412
rect 22278 40400 22284 40412
rect 22336 40400 22342 40452
rect 7190 40332 7196 40384
rect 7248 40372 7254 40384
rect 22002 40372 22008 40384
rect 7248 40344 22008 40372
rect 7248 40332 7254 40344
rect 22002 40332 22008 40344
rect 22060 40332 22066 40384
rect 9306 40264 9312 40316
rect 9364 40304 9370 40316
rect 23658 40304 23664 40316
rect 9364 40276 23664 40304
rect 9364 40264 9370 40276
rect 23658 40264 23664 40276
rect 23716 40264 23722 40316
rect 10318 40196 10324 40248
rect 10376 40236 10382 40248
rect 26326 40236 26332 40248
rect 10376 40208 26332 40236
rect 10376 40196 10382 40208
rect 26326 40196 26332 40208
rect 26384 40196 26390 40248
rect 9858 40128 9864 40180
rect 9916 40168 9922 40180
rect 9916 40140 12575 40168
rect 9916 40128 9922 40140
rect 8386 40060 8392 40112
rect 8444 40100 8450 40112
rect 11054 40100 11060 40112
rect 8444 40072 11060 40100
rect 8444 40060 8450 40072
rect 11054 40060 11060 40072
rect 11112 40060 11118 40112
rect 12547 40100 12575 40140
rect 12618 40128 12624 40180
rect 12676 40168 12682 40180
rect 24762 40168 24768 40180
rect 12676 40140 24768 40168
rect 12676 40128 12682 40140
rect 24762 40128 24768 40140
rect 24820 40128 24826 40180
rect 13078 40100 13084 40112
rect 12547 40072 13084 40100
rect 13078 40060 13084 40072
rect 13136 40060 13142 40112
rect 16574 40060 16580 40112
rect 16632 40100 16638 40112
rect 16632 40072 17080 40100
rect 16632 40060 16638 40072
rect 7926 39992 7932 40044
rect 7984 40032 7990 40044
rect 16942 40032 16948 40044
rect 7984 40004 16948 40032
rect 7984 39992 7990 40004
rect 16942 39992 16948 40004
rect 17000 39992 17006 40044
rect 17052 40032 17080 40072
rect 18046 40060 18052 40112
rect 18104 40100 18110 40112
rect 18874 40100 18880 40112
rect 18104 40072 18880 40100
rect 18104 40060 18110 40072
rect 18874 40060 18880 40072
rect 18932 40060 18938 40112
rect 21266 40032 21272 40044
rect 17052 40004 21272 40032
rect 21266 39992 21272 40004
rect 21324 39992 21330 40044
rect 9674 39924 9680 39976
rect 9732 39964 9738 39976
rect 9732 39936 12664 39964
rect 9732 39924 9738 39936
rect 8478 39856 8484 39908
rect 8536 39896 8542 39908
rect 11882 39896 11888 39908
rect 8536 39868 11888 39896
rect 8536 39856 8542 39868
rect 11882 39856 11888 39868
rect 11940 39896 11946 39908
rect 12434 39896 12440 39908
rect 11940 39868 12440 39896
rect 11940 39856 11946 39868
rect 12434 39856 12440 39868
rect 12492 39856 12498 39908
rect 12636 39896 12664 39936
rect 12710 39924 12716 39976
rect 12768 39964 12774 39976
rect 22186 39964 22192 39976
rect 12768 39936 22192 39964
rect 12768 39924 12774 39936
rect 22186 39924 22192 39936
rect 22244 39924 22250 39976
rect 12986 39896 12992 39908
rect 12636 39868 12992 39896
rect 12986 39856 12992 39868
rect 13044 39856 13050 39908
rect 13998 39856 14004 39908
rect 14056 39896 14062 39908
rect 16574 39896 16580 39908
rect 14056 39868 16580 39896
rect 14056 39856 14062 39868
rect 16574 39856 16580 39868
rect 16632 39856 16638 39908
rect 16666 39856 16672 39908
rect 16724 39896 16730 39908
rect 20806 39896 20812 39908
rect 16724 39868 20812 39896
rect 16724 39856 16730 39868
rect 20806 39856 20812 39868
rect 20864 39856 20870 39908
rect 6638 39788 6644 39840
rect 6696 39828 6702 39840
rect 14274 39828 14280 39840
rect 6696 39800 14280 39828
rect 6696 39788 6702 39800
rect 14274 39788 14280 39800
rect 14332 39788 14338 39840
rect 15562 39788 15568 39840
rect 15620 39828 15626 39840
rect 23474 39828 23480 39840
rect 15620 39800 23480 39828
rect 15620 39788 15626 39800
rect 23474 39788 23480 39800
rect 23532 39788 23538 39840
rect 1104 39738 28888 39760
rect 1104 39686 5582 39738
rect 5634 39686 5646 39738
rect 5698 39686 5710 39738
rect 5762 39686 5774 39738
rect 5826 39686 5838 39738
rect 5890 39686 14846 39738
rect 14898 39686 14910 39738
rect 14962 39686 14974 39738
rect 15026 39686 15038 39738
rect 15090 39686 15102 39738
rect 15154 39686 24110 39738
rect 24162 39686 24174 39738
rect 24226 39686 24238 39738
rect 24290 39686 24302 39738
rect 24354 39686 24366 39738
rect 24418 39686 28888 39738
rect 1104 39664 28888 39686
rect 7098 39624 7104 39636
rect 7059 39596 7104 39624
rect 7098 39584 7104 39596
rect 7156 39584 7162 39636
rect 10870 39624 10876 39636
rect 7208 39596 10876 39624
rect 5442 39556 5448 39568
rect 3712 39528 5448 39556
rect 1762 39420 1768 39432
rect 1723 39392 1768 39420
rect 1762 39380 1768 39392
rect 1820 39380 1826 39432
rect 2406 39420 2412 39432
rect 2367 39392 2412 39420
rect 2406 39380 2412 39392
rect 2464 39380 2470 39432
rect 3053 39423 3111 39429
rect 3053 39389 3065 39423
rect 3099 39420 3111 39423
rect 3712 39420 3740 39528
rect 5442 39516 5448 39528
rect 5500 39516 5506 39568
rect 7006 39516 7012 39568
rect 7064 39556 7070 39568
rect 7208 39556 7236 39596
rect 10870 39584 10876 39596
rect 10928 39584 10934 39636
rect 11054 39584 11060 39636
rect 11112 39624 11118 39636
rect 17494 39624 17500 39636
rect 11112 39596 17500 39624
rect 11112 39584 11118 39596
rect 17494 39584 17500 39596
rect 17552 39584 17558 39636
rect 7064 39528 7236 39556
rect 7745 39559 7803 39565
rect 7064 39516 7070 39528
rect 7745 39525 7757 39559
rect 7791 39556 7803 39559
rect 20162 39556 20168 39568
rect 7791 39528 20168 39556
rect 7791 39525 7803 39528
rect 7745 39519 7803 39525
rect 20162 39516 20168 39528
rect 20220 39516 20226 39568
rect 4154 39448 4160 39500
rect 4212 39488 4218 39500
rect 4249 39491 4307 39497
rect 4249 39488 4261 39491
rect 4212 39460 4261 39488
rect 4212 39448 4218 39460
rect 4249 39457 4261 39460
rect 4295 39457 4307 39491
rect 4249 39451 4307 39457
rect 8389 39491 8447 39497
rect 8389 39457 8401 39491
rect 8435 39488 8447 39491
rect 10134 39488 10140 39500
rect 8435 39460 10140 39488
rect 8435 39457 8447 39460
rect 8389 39451 8447 39457
rect 10134 39448 10140 39460
rect 10192 39448 10198 39500
rect 10318 39488 10324 39500
rect 10279 39460 10324 39488
rect 10318 39448 10324 39460
rect 10376 39448 10382 39500
rect 10686 39448 10692 39500
rect 10744 39488 10750 39500
rect 11609 39491 11667 39497
rect 11609 39488 11621 39491
rect 10744 39460 11621 39488
rect 10744 39448 10750 39460
rect 11609 39457 11621 39460
rect 11655 39457 11667 39491
rect 11790 39488 11796 39500
rect 11751 39460 11796 39488
rect 11609 39451 11667 39457
rect 11790 39448 11796 39460
rect 11848 39448 11854 39500
rect 12250 39448 12256 39500
rect 12308 39488 12314 39500
rect 12437 39491 12495 39497
rect 12437 39488 12449 39491
rect 12308 39460 12449 39488
rect 12308 39448 12314 39460
rect 12437 39457 12449 39460
rect 12483 39457 12495 39491
rect 12437 39451 12495 39457
rect 12526 39448 12532 39500
rect 12584 39488 12590 39500
rect 14090 39488 14096 39500
rect 12584 39460 14096 39488
rect 12584 39448 12590 39460
rect 14090 39448 14096 39460
rect 14148 39448 14154 39500
rect 15470 39488 15476 39500
rect 15431 39460 15476 39488
rect 15470 39448 15476 39460
rect 15528 39448 15534 39500
rect 15654 39448 15660 39500
rect 15712 39488 15718 39500
rect 19613 39491 19671 39497
rect 19613 39488 19625 39491
rect 15712 39460 19625 39488
rect 15712 39448 15718 39460
rect 19613 39457 19625 39460
rect 19659 39457 19671 39491
rect 19978 39488 19984 39500
rect 19939 39460 19984 39488
rect 19613 39451 19671 39457
rect 19978 39448 19984 39460
rect 20036 39448 20042 39500
rect 22002 39488 22008 39500
rect 21963 39460 22008 39488
rect 22002 39448 22008 39460
rect 22060 39448 22066 39500
rect 22186 39488 22192 39500
rect 22147 39460 22192 39488
rect 22186 39448 22192 39460
rect 22244 39448 22250 39500
rect 23842 39488 23848 39500
rect 23803 39460 23848 39488
rect 23842 39448 23848 39460
rect 23900 39448 23906 39500
rect 24762 39488 24768 39500
rect 24723 39460 24768 39488
rect 24762 39448 24768 39460
rect 24820 39448 24826 39500
rect 26050 39488 26056 39500
rect 26011 39460 26056 39488
rect 26050 39448 26056 39460
rect 26108 39448 26114 39500
rect 3099 39392 3740 39420
rect 3789 39423 3847 39429
rect 3099 39389 3111 39392
rect 3053 39383 3111 39389
rect 3789 39389 3801 39423
rect 3835 39389 3847 39423
rect 3789 39383 3847 39389
rect 1670 39244 1676 39296
rect 1728 39284 1734 39296
rect 1857 39287 1915 39293
rect 1857 39284 1869 39287
rect 1728 39256 1869 39284
rect 1728 39244 1734 39256
rect 1857 39253 1869 39256
rect 1903 39253 1915 39287
rect 2498 39284 2504 39296
rect 2459 39256 2504 39284
rect 1857 39247 1915 39253
rect 2498 39244 2504 39256
rect 2556 39244 2562 39296
rect 3142 39284 3148 39296
rect 3103 39256 3148 39284
rect 3142 39244 3148 39256
rect 3200 39244 3206 39296
rect 3804 39284 3832 39383
rect 9674 39380 9680 39432
rect 9732 39420 9738 39432
rect 9732 39392 9777 39420
rect 9732 39380 9738 39392
rect 10042 39380 10048 39432
rect 10100 39420 10106 39432
rect 10778 39420 10784 39432
rect 10100 39392 10784 39420
rect 10100 39380 10106 39392
rect 10778 39380 10784 39392
rect 10836 39380 10842 39432
rect 10870 39380 10876 39432
rect 10928 39420 10934 39432
rect 14274 39420 14280 39432
rect 10928 39392 11652 39420
rect 14235 39392 14280 39420
rect 10928 39380 10934 39392
rect 3970 39352 3976 39364
rect 3931 39324 3976 39352
rect 3970 39312 3976 39324
rect 4028 39312 4034 39364
rect 9766 39312 9772 39364
rect 9824 39352 9830 39364
rect 11514 39352 11520 39364
rect 9824 39324 11520 39352
rect 9824 39312 9830 39324
rect 11514 39312 11520 39324
rect 11572 39312 11578 39364
rect 11624 39352 11652 39392
rect 14274 39380 14280 39392
rect 14332 39380 14338 39432
rect 16666 39420 16672 39432
rect 16491 39392 16672 39420
rect 13998 39352 14004 39364
rect 11624 39324 14004 39352
rect 13998 39312 14004 39324
rect 14056 39312 14062 39364
rect 14458 39352 14464 39364
rect 14419 39324 14464 39352
rect 14458 39312 14464 39324
rect 14516 39312 14522 39364
rect 14550 39312 14556 39364
rect 14608 39352 14614 39364
rect 16491 39352 16519 39392
rect 16666 39380 16672 39392
rect 16724 39380 16730 39432
rect 17313 39423 17371 39429
rect 17313 39389 17325 39423
rect 17359 39389 17371 39423
rect 17313 39383 17371 39389
rect 17328 39352 17356 39383
rect 17586 39380 17592 39432
rect 17644 39420 17650 39432
rect 18141 39423 18199 39429
rect 18141 39420 18153 39423
rect 17644 39392 18153 39420
rect 17644 39380 17650 39392
rect 18141 39389 18153 39392
rect 18187 39389 18199 39423
rect 18141 39383 18199 39389
rect 19334 39380 19340 39432
rect 19392 39420 19398 39432
rect 19429 39423 19487 39429
rect 19429 39420 19441 39423
rect 19392 39392 19441 39420
rect 19392 39380 19398 39392
rect 19429 39389 19441 39392
rect 19475 39389 19487 39423
rect 24578 39420 24584 39432
rect 24539 39392 24584 39420
rect 19429 39383 19487 39389
rect 24578 39380 24584 39392
rect 24636 39380 24642 39432
rect 14608 39324 16519 39352
rect 16592 39324 17816 39352
rect 14608 39312 14614 39324
rect 5258 39284 5264 39296
rect 3804 39256 5264 39284
rect 5258 39244 5264 39256
rect 5316 39244 5322 39296
rect 7098 39244 7104 39296
rect 7156 39284 7162 39296
rect 10686 39284 10692 39296
rect 7156 39256 10692 39284
rect 7156 39244 7162 39256
rect 10686 39244 10692 39256
rect 10744 39244 10750 39296
rect 10873 39287 10931 39293
rect 10873 39253 10885 39287
rect 10919 39284 10931 39287
rect 12342 39284 12348 39296
rect 10919 39256 12348 39284
rect 10919 39253 10931 39256
rect 10873 39247 10931 39253
rect 12342 39244 12348 39256
rect 12400 39244 12406 39296
rect 12802 39244 12808 39296
rect 12860 39284 12866 39296
rect 16592 39284 16620 39324
rect 12860 39256 16620 39284
rect 16761 39287 16819 39293
rect 12860 39244 12866 39256
rect 16761 39253 16773 39287
rect 16807 39284 16819 39287
rect 17310 39284 17316 39296
rect 16807 39256 17316 39284
rect 16807 39253 16819 39256
rect 16761 39247 16819 39253
rect 17310 39244 17316 39256
rect 17368 39244 17374 39296
rect 17405 39287 17463 39293
rect 17405 39253 17417 39287
rect 17451 39284 17463 39287
rect 17678 39284 17684 39296
rect 17451 39256 17684 39284
rect 17451 39253 17463 39256
rect 17405 39247 17463 39253
rect 17678 39244 17684 39256
rect 17736 39244 17742 39296
rect 17788 39284 17816 39324
rect 17862 39312 17868 39364
rect 17920 39352 17926 39364
rect 17957 39355 18015 39361
rect 17957 39352 17969 39355
rect 17920 39324 17969 39352
rect 17920 39312 17926 39324
rect 17957 39321 17969 39324
rect 18003 39321 18015 39355
rect 18966 39352 18972 39364
rect 17957 39315 18015 39321
rect 18064 39324 18972 39352
rect 18064 39284 18092 39324
rect 18966 39312 18972 39324
rect 19024 39312 19030 39364
rect 26786 39312 26792 39364
rect 26844 39352 26850 39364
rect 27433 39355 27491 39361
rect 27433 39352 27445 39355
rect 26844 39324 27445 39352
rect 26844 39312 26850 39324
rect 27433 39321 27445 39324
rect 27479 39321 27491 39355
rect 27614 39352 27620 39364
rect 27575 39324 27620 39352
rect 27433 39315 27491 39321
rect 27614 39312 27620 39324
rect 27672 39312 27678 39364
rect 17788 39256 18092 39284
rect 18325 39287 18383 39293
rect 18325 39253 18337 39287
rect 18371 39284 18383 39287
rect 18598 39284 18604 39296
rect 18371 39256 18604 39284
rect 18371 39253 18383 39256
rect 18325 39247 18383 39253
rect 18598 39244 18604 39256
rect 18656 39244 18662 39296
rect 19886 39244 19892 39296
rect 19944 39284 19950 39296
rect 20990 39284 20996 39296
rect 19944 39256 20996 39284
rect 19944 39244 19950 39256
rect 20990 39244 20996 39256
rect 21048 39244 21054 39296
rect 1104 39194 28888 39216
rect 1104 39142 10214 39194
rect 10266 39142 10278 39194
rect 10330 39142 10342 39194
rect 10394 39142 10406 39194
rect 10458 39142 10470 39194
rect 10522 39142 19478 39194
rect 19530 39142 19542 39194
rect 19594 39142 19606 39194
rect 19658 39142 19670 39194
rect 19722 39142 19734 39194
rect 19786 39142 28888 39194
rect 1104 39120 28888 39142
rect 9861 39083 9919 39089
rect 9861 39049 9873 39083
rect 9907 39080 9919 39083
rect 14458 39080 14464 39092
rect 9907 39052 14464 39080
rect 9907 39049 9919 39052
rect 9861 39043 9919 39049
rect 14458 39040 14464 39052
rect 14516 39040 14522 39092
rect 14550 39040 14556 39092
rect 14608 39080 14614 39092
rect 15286 39080 15292 39092
rect 14608 39052 15292 39080
rect 14608 39040 14614 39052
rect 15286 39040 15292 39052
rect 15344 39040 15350 39092
rect 15470 39040 15476 39092
rect 15528 39080 15534 39092
rect 15528 39052 17908 39080
rect 15528 39040 15534 39052
rect 1670 39012 1676 39024
rect 1631 38984 1676 39012
rect 1670 38972 1676 38984
rect 1728 38972 1734 39024
rect 3142 38972 3148 39024
rect 3200 39012 3206 39024
rect 3973 39015 4031 39021
rect 3973 39012 3985 39015
rect 3200 38984 3985 39012
rect 3200 38972 3206 38984
rect 3973 38981 3985 38984
rect 4019 38981 4031 39015
rect 10870 39012 10876 39024
rect 3973 38975 4031 38981
rect 9968 38984 10876 39012
rect 7374 38944 7380 38956
rect 7335 38916 7380 38944
rect 7374 38904 7380 38916
rect 7432 38904 7438 38956
rect 8662 38944 8668 38956
rect 8623 38916 8668 38944
rect 8662 38904 8668 38916
rect 8720 38904 8726 38956
rect 9306 38944 9312 38956
rect 9267 38916 9312 38944
rect 9306 38904 9312 38916
rect 9364 38904 9370 38956
rect 9769 38947 9827 38953
rect 9769 38913 9781 38947
rect 9815 38944 9827 38947
rect 9968 38944 9996 38984
rect 10870 38972 10876 38984
rect 10928 38972 10934 39024
rect 11793 39015 11851 39021
rect 11793 38981 11805 39015
rect 11839 39012 11851 39015
rect 15654 39012 15660 39024
rect 11839 38984 15660 39012
rect 11839 38981 11851 38984
rect 11793 38975 11851 38981
rect 15654 38972 15660 38984
rect 15712 38972 15718 39024
rect 16758 39012 16764 39024
rect 16132 38984 16764 39012
rect 9815 38916 9996 38944
rect 9815 38913 9827 38916
rect 9769 38907 9827 38913
rect 10226 38904 10232 38956
rect 10284 38944 10290 38956
rect 10413 38947 10471 38953
rect 10413 38944 10425 38947
rect 10284 38916 10425 38944
rect 10284 38904 10290 38916
rect 10413 38913 10425 38916
rect 10459 38913 10471 38947
rect 10413 38907 10471 38913
rect 11701 38947 11759 38953
rect 11701 38913 11713 38947
rect 11747 38944 11759 38947
rect 11882 38944 11888 38956
rect 11747 38916 11888 38944
rect 11747 38913 11759 38916
rect 11701 38907 11759 38913
rect 11882 38904 11888 38916
rect 11940 38904 11946 38956
rect 12345 38947 12403 38953
rect 12345 38913 12357 38947
rect 12391 38913 12403 38947
rect 12345 38907 12403 38913
rect 12437 38947 12495 38953
rect 12437 38913 12449 38947
rect 12483 38944 12495 38947
rect 12710 38944 12716 38956
rect 12483 38916 12716 38944
rect 12483 38913 12495 38916
rect 12437 38907 12495 38913
rect 1486 38876 1492 38888
rect 1447 38848 1492 38876
rect 1486 38836 1492 38848
rect 1544 38836 1550 38888
rect 2866 38876 2872 38888
rect 2827 38848 2872 38876
rect 2866 38836 2872 38848
rect 2924 38836 2930 38888
rect 3789 38879 3847 38885
rect 3789 38845 3801 38879
rect 3835 38876 3847 38879
rect 4614 38876 4620 38888
rect 3835 38848 4620 38876
rect 3835 38845 3847 38848
rect 3789 38839 3847 38845
rect 4614 38836 4620 38848
rect 4672 38836 4678 38888
rect 4706 38836 4712 38888
rect 4764 38876 4770 38888
rect 4764 38848 4809 38876
rect 4764 38836 4770 38848
rect 8570 38836 8576 38888
rect 8628 38876 8634 38888
rect 9214 38876 9220 38888
rect 8628 38848 9220 38876
rect 8628 38836 8634 38848
rect 9214 38836 9220 38848
rect 9272 38836 9278 38888
rect 10318 38836 10324 38888
rect 10376 38876 10382 38888
rect 12360 38876 12388 38907
rect 12710 38904 12716 38916
rect 12768 38904 12774 38956
rect 12986 38944 12992 38956
rect 12947 38916 12992 38944
rect 12986 38904 12992 38916
rect 13044 38904 13050 38956
rect 14642 38904 14648 38956
rect 14700 38944 14706 38956
rect 15562 38944 15568 38956
rect 14700 38916 15568 38944
rect 14700 38904 14706 38916
rect 15562 38904 15568 38916
rect 15620 38904 15626 38956
rect 13170 38876 13176 38888
rect 10376 38848 12388 38876
rect 13131 38848 13176 38876
rect 10376 38836 10382 38848
rect 13170 38836 13176 38848
rect 13228 38836 13234 38888
rect 13538 38876 13544 38888
rect 13499 38848 13544 38876
rect 13538 38836 13544 38848
rect 13596 38836 13602 38888
rect 14090 38836 14096 38888
rect 14148 38876 14154 38888
rect 16132 38876 16160 38984
rect 16758 38972 16764 38984
rect 16816 38972 16822 39024
rect 16942 38972 16948 39024
rect 17000 39012 17006 39024
rect 17037 39015 17095 39021
rect 17037 39012 17049 39015
rect 17000 38984 17049 39012
rect 17000 38972 17006 38984
rect 17037 38981 17049 38984
rect 17083 38981 17095 39015
rect 17037 38975 17095 38981
rect 17678 38972 17684 39024
rect 17736 39012 17742 39024
rect 17880 39012 17908 39052
rect 18414 39040 18420 39092
rect 18472 39080 18478 39092
rect 18472 39052 22094 39080
rect 18472 39040 18478 39052
rect 18322 39012 18328 39024
rect 17736 38984 17778 39012
rect 17880 38984 18328 39012
rect 17736 38972 17742 38984
rect 18322 38972 18328 38984
rect 18380 38972 18386 39024
rect 18874 38972 18880 39024
rect 18932 38972 18938 39024
rect 20070 39012 20076 39024
rect 19904 38984 20076 39012
rect 16482 38904 16488 38956
rect 16540 38944 16546 38956
rect 16853 38947 16911 38953
rect 16853 38944 16865 38947
rect 16540 38916 16865 38944
rect 16540 38904 16546 38916
rect 16853 38913 16865 38916
rect 16899 38913 16911 38947
rect 17494 38944 17500 38956
rect 17455 38916 17500 38944
rect 16853 38907 16911 38913
rect 17494 38904 17500 38916
rect 17552 38904 17558 38956
rect 18892 38885 18920 38972
rect 19904 38953 19932 38984
rect 20070 38972 20076 38984
rect 20128 38972 20134 39024
rect 20165 39015 20223 39021
rect 20165 38981 20177 39015
rect 20211 39012 20223 39015
rect 20346 39012 20352 39024
rect 20211 38984 20352 39012
rect 20211 38981 20223 38984
rect 20165 38975 20223 38981
rect 20346 38972 20352 38984
rect 20404 38972 20410 39024
rect 22066 39012 22094 39052
rect 22465 39015 22523 39021
rect 22465 39012 22477 39015
rect 22066 38984 22477 39012
rect 22465 38981 22477 38984
rect 22511 38981 22523 39015
rect 26970 39012 26976 39024
rect 26931 38984 26976 39012
rect 22465 38975 22523 38981
rect 26970 38972 26976 38984
rect 27028 38972 27034 39024
rect 27154 38972 27160 39024
rect 27212 39021 27218 39024
rect 27212 39015 27231 39021
rect 27219 38981 27231 39015
rect 27212 38975 27231 38981
rect 27212 38972 27218 38975
rect 19889 38947 19947 38953
rect 19889 38913 19901 38947
rect 19935 38913 19947 38947
rect 19889 38907 19947 38913
rect 19981 38947 20039 38953
rect 19981 38913 19993 38947
rect 20027 38944 20039 38947
rect 20027 38916 20116 38944
rect 20027 38913 20039 38916
rect 19981 38907 20039 38913
rect 14148 38848 16160 38876
rect 16669 38879 16727 38885
rect 14148 38836 14154 38848
rect 16669 38845 16681 38879
rect 16715 38845 16727 38879
rect 16669 38839 16727 38845
rect 18877 38879 18935 38885
rect 18877 38845 18889 38879
rect 18923 38845 18935 38879
rect 18877 38839 18935 38845
rect 1670 38768 1676 38820
rect 1728 38808 1734 38820
rect 2406 38808 2412 38820
rect 1728 38780 2412 38808
rect 1728 38768 1734 38780
rect 2406 38768 2412 38780
rect 2464 38808 2470 38820
rect 8018 38808 8024 38820
rect 2464 38780 7880 38808
rect 7979 38780 8024 38808
rect 2464 38768 2470 38780
rect 6546 38740 6552 38752
rect 6507 38712 6552 38740
rect 6546 38700 6552 38712
rect 6604 38700 6610 38752
rect 7852 38740 7880 38780
rect 8018 38768 8024 38780
rect 8076 38768 8082 38820
rect 11330 38768 11336 38820
rect 11388 38808 11394 38820
rect 13262 38808 13268 38820
rect 11388 38780 13268 38808
rect 11388 38768 11394 38780
rect 13262 38768 13268 38780
rect 13320 38768 13326 38820
rect 13354 38768 13360 38820
rect 13412 38808 13418 38820
rect 16206 38808 16212 38820
rect 13412 38780 16212 38808
rect 13412 38768 13418 38780
rect 16206 38768 16212 38780
rect 16264 38768 16270 38820
rect 16684 38808 16712 38839
rect 19058 38836 19064 38888
rect 19116 38876 19122 38888
rect 19794 38876 19800 38888
rect 19116 38848 19800 38876
rect 19116 38836 19122 38848
rect 19794 38836 19800 38848
rect 19852 38836 19858 38888
rect 16684 38780 17724 38808
rect 9122 38740 9128 38752
rect 7852 38712 9128 38740
rect 9122 38700 9128 38712
rect 9180 38700 9186 38752
rect 9214 38700 9220 38752
rect 9272 38740 9278 38752
rect 10318 38740 10324 38752
rect 9272 38712 10324 38740
rect 9272 38700 9278 38712
rect 10318 38700 10324 38712
rect 10376 38700 10382 38752
rect 10502 38700 10508 38752
rect 10560 38740 10566 38752
rect 10560 38712 10605 38740
rect 10560 38700 10566 38712
rect 11238 38700 11244 38752
rect 11296 38740 11302 38752
rect 12526 38740 12532 38752
rect 11296 38712 12532 38740
rect 11296 38700 11302 38712
rect 12526 38700 12532 38712
rect 12584 38700 12590 38752
rect 13078 38700 13084 38752
rect 13136 38740 13142 38752
rect 15470 38740 15476 38752
rect 13136 38712 15476 38740
rect 13136 38700 13142 38712
rect 15470 38700 15476 38712
rect 15528 38700 15534 38752
rect 15657 38743 15715 38749
rect 15657 38709 15669 38743
rect 15703 38740 15715 38743
rect 15746 38740 15752 38752
rect 15703 38712 15752 38740
rect 15703 38709 15715 38712
rect 15657 38703 15715 38709
rect 15746 38700 15752 38712
rect 15804 38700 15810 38752
rect 16298 38700 16304 38752
rect 16356 38740 16362 38752
rect 17586 38740 17592 38752
rect 16356 38712 17592 38740
rect 16356 38700 16362 38712
rect 17586 38700 17592 38712
rect 17644 38700 17650 38752
rect 17696 38740 17724 38780
rect 18322 38768 18328 38820
rect 18380 38808 18386 38820
rect 20088 38808 20116 38916
rect 20254 38904 20260 38956
rect 20312 38944 20318 38956
rect 20625 38947 20683 38953
rect 20625 38944 20637 38947
rect 20312 38916 20637 38944
rect 20312 38904 20318 38916
rect 20625 38913 20637 38916
rect 20671 38913 20683 38947
rect 20625 38907 20683 38913
rect 20714 38904 20720 38956
rect 20772 38944 20778 38956
rect 20809 38947 20867 38953
rect 20809 38944 20821 38947
rect 20772 38916 20821 38944
rect 20772 38904 20778 38916
rect 20809 38913 20821 38916
rect 20855 38913 20867 38947
rect 22278 38944 22284 38956
rect 22239 38916 22284 38944
rect 20809 38907 20867 38913
rect 22278 38904 22284 38916
rect 22336 38904 22342 38956
rect 23658 38904 23664 38956
rect 23716 38944 23722 38956
rect 24581 38947 24639 38953
rect 24581 38944 24593 38947
rect 23716 38916 24593 38944
rect 23716 38904 23722 38916
rect 24581 38913 24593 38916
rect 24627 38913 24639 38947
rect 27982 38944 27988 38956
rect 27943 38916 27988 38944
rect 24581 38907 24639 38913
rect 27982 38904 27988 38916
rect 28040 38904 28046 38956
rect 23198 38876 23204 38888
rect 23159 38848 23204 38876
rect 23198 38836 23204 38848
rect 23256 38836 23262 38888
rect 24765 38879 24823 38885
rect 24765 38845 24777 38879
rect 24811 38876 24823 38879
rect 25958 38876 25964 38888
rect 24811 38848 25964 38876
rect 24811 38845 24823 38848
rect 24765 38839 24823 38845
rect 25958 38836 25964 38848
rect 26016 38836 26022 38888
rect 26142 38876 26148 38888
rect 26103 38848 26148 38876
rect 26142 38836 26148 38848
rect 26200 38836 26206 38888
rect 27430 38808 27436 38820
rect 18380 38780 20116 38808
rect 27172 38780 27436 38808
rect 18380 38768 18386 38780
rect 18414 38740 18420 38752
rect 17696 38712 18420 38740
rect 18414 38700 18420 38712
rect 18472 38740 18478 38752
rect 19886 38740 19892 38752
rect 18472 38712 19892 38740
rect 18472 38700 18478 38712
rect 19886 38700 19892 38712
rect 19944 38700 19950 38752
rect 20622 38700 20628 38752
rect 20680 38740 20686 38752
rect 27172 38749 27200 38780
rect 27430 38768 27436 38780
rect 27488 38768 27494 38820
rect 20993 38743 21051 38749
rect 20993 38740 21005 38743
rect 20680 38712 21005 38740
rect 20680 38700 20686 38712
rect 20993 38709 21005 38712
rect 21039 38709 21051 38743
rect 20993 38703 21051 38709
rect 27157 38743 27215 38749
rect 27157 38709 27169 38743
rect 27203 38709 27215 38743
rect 27338 38740 27344 38752
rect 27299 38712 27344 38740
rect 27157 38703 27215 38709
rect 27338 38700 27344 38712
rect 27396 38700 27402 38752
rect 27522 38700 27528 38752
rect 27580 38740 27586 38752
rect 28077 38743 28135 38749
rect 28077 38740 28089 38743
rect 27580 38712 28089 38740
rect 27580 38700 27586 38712
rect 28077 38709 28089 38712
rect 28123 38709 28135 38743
rect 28077 38703 28135 38709
rect 1104 38650 28888 38672
rect 1104 38598 5582 38650
rect 5634 38598 5646 38650
rect 5698 38598 5710 38650
rect 5762 38598 5774 38650
rect 5826 38598 5838 38650
rect 5890 38598 14846 38650
rect 14898 38598 14910 38650
rect 14962 38598 14974 38650
rect 15026 38598 15038 38650
rect 15090 38598 15102 38650
rect 15154 38598 24110 38650
rect 24162 38598 24174 38650
rect 24226 38598 24238 38650
rect 24290 38598 24302 38650
rect 24354 38598 24366 38650
rect 24418 38598 28888 38650
rect 1104 38576 28888 38598
rect 14 38496 20 38548
rect 72 38536 78 38548
rect 1394 38536 1400 38548
rect 72 38508 1400 38536
rect 72 38496 78 38508
rect 1394 38496 1400 38508
rect 1452 38496 1458 38548
rect 3234 38496 3240 38548
rect 3292 38536 3298 38548
rect 4706 38536 4712 38548
rect 3292 38508 4712 38536
rect 3292 38496 3298 38508
rect 4706 38496 4712 38508
rect 4764 38496 4770 38548
rect 8386 38536 8392 38548
rect 8347 38508 8392 38536
rect 8386 38496 8392 38508
rect 8444 38496 8450 38548
rect 9398 38496 9404 38548
rect 9456 38536 9462 38548
rect 9456 38508 12112 38536
rect 9456 38496 9462 38508
rect 6546 38468 6552 38480
rect 1412 38440 6552 38468
rect 1412 38409 1440 38440
rect 6546 38428 6552 38440
rect 6604 38428 6610 38480
rect 7742 38468 7748 38480
rect 7703 38440 7748 38468
rect 7742 38428 7748 38440
rect 7800 38428 7806 38480
rect 9033 38471 9091 38477
rect 9033 38437 9045 38471
rect 9079 38468 9091 38471
rect 12084 38468 12112 38508
rect 12158 38496 12164 38548
rect 12216 38536 12222 38548
rect 12986 38536 12992 38548
rect 12216 38508 12992 38536
rect 12216 38496 12222 38508
rect 12986 38496 12992 38508
rect 13044 38496 13050 38548
rect 13170 38496 13176 38548
rect 13228 38536 13234 38548
rect 13265 38539 13323 38545
rect 13265 38536 13277 38539
rect 13228 38508 13277 38536
rect 13228 38496 13234 38508
rect 13265 38505 13277 38508
rect 13311 38505 13323 38539
rect 18233 38539 18291 38545
rect 18233 38536 18245 38539
rect 13265 38499 13323 38505
rect 13924 38508 18245 38536
rect 13924 38468 13952 38508
rect 18233 38505 18245 38508
rect 18279 38505 18291 38539
rect 18233 38499 18291 38505
rect 18414 38496 18420 38548
rect 18472 38536 18478 38548
rect 23201 38539 23259 38545
rect 18472 38508 23152 38536
rect 18472 38496 18478 38508
rect 9079 38440 12020 38468
rect 12084 38440 13952 38468
rect 14369 38471 14427 38477
rect 9079 38437 9091 38440
rect 9033 38431 9091 38437
rect 1397 38403 1455 38409
rect 1397 38369 1409 38403
rect 1443 38369 1455 38403
rect 1397 38363 1455 38369
rect 1581 38403 1639 38409
rect 1581 38369 1593 38403
rect 1627 38400 1639 38403
rect 2498 38400 2504 38412
rect 1627 38372 2504 38400
rect 1627 38369 1639 38372
rect 1581 38363 1639 38369
rect 2498 38360 2504 38372
rect 2556 38360 2562 38412
rect 2774 38360 2780 38412
rect 2832 38400 2838 38412
rect 4157 38403 4215 38409
rect 2832 38372 2877 38400
rect 2832 38360 2838 38372
rect 4157 38369 4169 38403
rect 4203 38400 4215 38403
rect 4893 38403 4951 38409
rect 4893 38400 4905 38403
rect 4203 38372 4905 38400
rect 4203 38369 4215 38372
rect 4157 38363 4215 38369
rect 4893 38369 4905 38372
rect 4939 38369 4951 38403
rect 5166 38400 5172 38412
rect 5127 38372 5172 38400
rect 4893 38363 4951 38369
rect 5166 38360 5172 38372
rect 5224 38360 5230 38412
rect 5350 38360 5356 38412
rect 5408 38400 5414 38412
rect 8570 38400 8576 38412
rect 5408 38372 8576 38400
rect 5408 38360 5414 38372
rect 8570 38360 8576 38372
rect 8628 38360 8634 38412
rect 9398 38400 9404 38412
rect 9324 38372 9404 38400
rect 4065 38335 4123 38341
rect 4065 38301 4077 38335
rect 4111 38332 4123 38335
rect 4246 38332 4252 38344
rect 4111 38304 4252 38332
rect 4111 38301 4123 38304
rect 4065 38295 4123 38301
rect 4246 38292 4252 38304
rect 4304 38292 4310 38344
rect 4709 38335 4767 38341
rect 4709 38301 4721 38335
rect 4755 38301 4767 38335
rect 4709 38295 4767 38301
rect 9217 38335 9275 38341
rect 9217 38301 9229 38335
rect 9263 38332 9275 38335
rect 9324 38332 9352 38372
rect 9398 38360 9404 38372
rect 9456 38360 9462 38412
rect 9766 38400 9772 38412
rect 9727 38372 9772 38400
rect 9766 38360 9772 38372
rect 9824 38360 9830 38412
rect 10134 38360 10140 38412
rect 10192 38400 10198 38412
rect 10321 38403 10379 38409
rect 10321 38400 10333 38403
rect 10192 38372 10333 38400
rect 10192 38360 10198 38372
rect 10321 38369 10333 38372
rect 10367 38369 10379 38403
rect 10502 38400 10508 38412
rect 10463 38372 10508 38400
rect 10321 38363 10379 38369
rect 10502 38360 10508 38372
rect 10560 38360 10566 38412
rect 10962 38360 10968 38412
rect 11020 38400 11026 38412
rect 11057 38403 11115 38409
rect 11057 38400 11069 38403
rect 11020 38372 11069 38400
rect 11020 38360 11026 38372
rect 11057 38369 11069 38372
rect 11103 38369 11115 38403
rect 11992 38400 12020 38440
rect 14369 38437 14381 38471
rect 14415 38468 14427 38471
rect 14734 38468 14740 38480
rect 14415 38440 14740 38468
rect 14415 38437 14427 38440
rect 14369 38431 14427 38437
rect 14734 38428 14740 38440
rect 14792 38428 14798 38480
rect 15013 38471 15071 38477
rect 15013 38437 15025 38471
rect 15059 38468 15071 38471
rect 23124 38468 23152 38508
rect 23201 38505 23213 38539
rect 23247 38536 23259 38539
rect 23658 38536 23664 38548
rect 23247 38508 23664 38536
rect 23247 38505 23259 38508
rect 23201 38499 23259 38505
rect 23658 38496 23664 38508
rect 23716 38536 23722 38548
rect 26970 38536 26976 38548
rect 23716 38508 26976 38536
rect 23716 38496 23722 38508
rect 26970 38496 26976 38508
rect 27028 38496 27034 38548
rect 15059 38440 20392 38468
rect 23124 38440 25728 38468
rect 15059 38437 15071 38440
rect 15013 38431 15071 38437
rect 11992 38372 12572 38400
rect 11057 38363 11115 38369
rect 9263 38304 9352 38332
rect 9263 38301 9275 38304
rect 9217 38295 9275 38301
rect 1946 38224 1952 38276
rect 2004 38264 2010 38276
rect 2866 38264 2872 38276
rect 2004 38236 2872 38264
rect 2004 38224 2010 38236
rect 2866 38224 2872 38236
rect 2924 38224 2930 38276
rect 4724 38264 4752 38295
rect 9490 38292 9496 38344
rect 9548 38332 9554 38344
rect 9677 38335 9735 38341
rect 9677 38332 9689 38335
rect 9548 38304 9689 38332
rect 9548 38292 9554 38304
rect 9677 38301 9689 38304
rect 9723 38332 9735 38335
rect 10042 38332 10048 38344
rect 9723 38304 10048 38332
rect 9723 38301 9735 38304
rect 9677 38295 9735 38301
rect 10042 38292 10048 38304
rect 10100 38292 10106 38344
rect 11790 38292 11796 38344
rect 11848 38332 11854 38344
rect 12158 38332 12164 38344
rect 11848 38304 12164 38332
rect 11848 38292 11854 38304
rect 12158 38292 12164 38304
rect 12216 38292 12222 38344
rect 12544 38332 12572 38372
rect 12618 38360 12624 38412
rect 12676 38400 12682 38412
rect 15378 38400 15384 38412
rect 12676 38372 15384 38400
rect 12676 38360 12682 38372
rect 15378 38360 15384 38372
rect 15436 38360 15442 38412
rect 15562 38400 15568 38412
rect 15523 38372 15568 38400
rect 15562 38360 15568 38372
rect 15620 38360 15626 38412
rect 15746 38400 15752 38412
rect 15707 38372 15752 38400
rect 15746 38360 15752 38372
rect 15804 38360 15810 38412
rect 16114 38400 16120 38412
rect 16075 38372 16120 38400
rect 16114 38360 16120 38372
rect 16172 38360 16178 38412
rect 16482 38360 16488 38412
rect 16540 38400 16546 38412
rect 17862 38400 17868 38412
rect 16540 38372 17356 38400
rect 17823 38372 17868 38400
rect 16540 38360 16546 38372
rect 12802 38332 12808 38344
rect 12544 38304 12808 38332
rect 12802 38292 12808 38304
rect 12860 38292 12866 38344
rect 13170 38332 13176 38344
rect 13131 38304 13176 38332
rect 13170 38292 13176 38304
rect 13228 38292 13234 38344
rect 13262 38292 13268 38344
rect 13320 38332 13326 38344
rect 14277 38335 14335 38341
rect 14277 38332 14289 38335
rect 13320 38304 14289 38332
rect 13320 38292 13326 38304
rect 14277 38301 14289 38304
rect 14323 38332 14335 38335
rect 14826 38332 14832 38344
rect 14323 38304 14832 38332
rect 14323 38301 14335 38304
rect 14277 38295 14335 38301
rect 14826 38292 14832 38304
rect 14884 38292 14890 38344
rect 14921 38335 14979 38341
rect 14921 38301 14933 38335
rect 14967 38332 14979 38335
rect 15470 38332 15476 38344
rect 14967 38304 15476 38332
rect 14967 38301 14979 38304
rect 14921 38295 14979 38301
rect 15470 38292 15476 38304
rect 15528 38292 15534 38344
rect 17328 38332 17356 38372
rect 17862 38360 17868 38372
rect 17920 38360 17926 38412
rect 18690 38360 18696 38412
rect 18748 38400 18754 38412
rect 19245 38403 19303 38409
rect 19245 38400 19257 38403
rect 18748 38372 19257 38400
rect 18748 38360 18754 38372
rect 19245 38369 19257 38372
rect 19291 38369 19303 38403
rect 20162 38400 20168 38412
rect 20123 38372 20168 38400
rect 19245 38363 19303 38369
rect 20162 38360 20168 38372
rect 20220 38360 20226 38412
rect 20364 38409 20392 38440
rect 20349 38403 20407 38409
rect 20349 38369 20361 38403
rect 20395 38369 20407 38403
rect 20349 38363 20407 38369
rect 20530 38360 20536 38412
rect 20588 38400 20594 38412
rect 20717 38403 20775 38409
rect 20717 38400 20729 38403
rect 20588 38372 20729 38400
rect 20588 38360 20594 38372
rect 20717 38369 20729 38372
rect 20763 38369 20775 38403
rect 22922 38400 22928 38412
rect 20717 38363 20775 38369
rect 22480 38372 22928 38400
rect 18049 38335 18107 38341
rect 18049 38332 18061 38335
rect 17328 38304 18061 38332
rect 18049 38301 18061 38304
rect 18095 38332 18107 38335
rect 19429 38335 19487 38341
rect 19429 38332 19441 38335
rect 18095 38304 19441 38332
rect 18095 38301 18107 38304
rect 18049 38295 18107 38301
rect 19429 38301 19441 38304
rect 19475 38301 19487 38335
rect 19429 38295 19487 38301
rect 21542 38292 21548 38344
rect 21600 38332 21606 38344
rect 22480 38341 22508 38372
rect 22922 38360 22928 38372
rect 22980 38360 22986 38412
rect 23477 38403 23535 38409
rect 23477 38369 23489 38403
rect 23523 38400 23535 38403
rect 23842 38400 23848 38412
rect 23523 38372 23848 38400
rect 23523 38369 23535 38372
rect 23477 38363 23535 38369
rect 23842 38360 23848 38372
rect 23900 38360 23906 38412
rect 22465 38335 22523 38341
rect 22465 38332 22477 38335
rect 21600 38304 22477 38332
rect 21600 38292 21606 38304
rect 22465 38301 22477 38304
rect 22511 38301 22523 38335
rect 23658 38332 23664 38344
rect 22465 38295 22523 38301
rect 22756 38304 23664 38332
rect 5166 38264 5172 38276
rect 4724 38236 5172 38264
rect 5166 38224 5172 38236
rect 5224 38224 5230 38276
rect 6362 38224 6368 38276
rect 6420 38264 6426 38276
rect 8478 38264 8484 38276
rect 6420 38236 8484 38264
rect 6420 38224 6426 38236
rect 8478 38224 8484 38236
rect 8536 38224 8542 38276
rect 9122 38224 9128 38276
rect 9180 38264 9186 38276
rect 9180 38236 14504 38264
rect 9180 38224 9186 38236
rect 10042 38156 10048 38208
rect 10100 38196 10106 38208
rect 11790 38196 11796 38208
rect 10100 38168 11796 38196
rect 10100 38156 10106 38168
rect 11790 38156 11796 38168
rect 11848 38156 11854 38208
rect 11974 38156 11980 38208
rect 12032 38196 12038 38208
rect 13170 38196 13176 38208
rect 12032 38168 13176 38196
rect 12032 38156 12038 38168
rect 13170 38156 13176 38168
rect 13228 38156 13234 38208
rect 14476 38196 14504 38236
rect 14734 38224 14740 38276
rect 14792 38264 14798 38276
rect 22002 38264 22008 38276
rect 14792 38236 22008 38264
rect 14792 38224 14798 38236
rect 22002 38224 22008 38236
rect 22060 38224 22066 38276
rect 22278 38224 22284 38276
rect 22336 38264 22342 38276
rect 22649 38267 22707 38273
rect 22649 38264 22661 38267
rect 22336 38236 22661 38264
rect 22336 38224 22342 38236
rect 22649 38233 22661 38236
rect 22695 38233 22707 38267
rect 22649 38227 22707 38233
rect 18230 38196 18236 38208
rect 14476 38168 18236 38196
rect 18230 38156 18236 38168
rect 18288 38156 18294 38208
rect 18322 38156 18328 38208
rect 18380 38196 18386 38208
rect 19613 38199 19671 38205
rect 19613 38196 19625 38199
rect 18380 38168 19625 38196
rect 18380 38156 18386 38168
rect 19613 38165 19625 38168
rect 19659 38165 19671 38199
rect 19613 38159 19671 38165
rect 20898 38156 20904 38208
rect 20956 38196 20962 38208
rect 22756 38196 22784 38304
rect 23658 38292 23664 38304
rect 23716 38292 23722 38344
rect 24587 38332 24615 38440
rect 24673 38335 24731 38341
rect 24673 38332 24685 38335
rect 24587 38304 24685 38332
rect 24673 38301 24685 38304
rect 24719 38301 24731 38335
rect 24673 38295 24731 38301
rect 24765 38335 24823 38341
rect 24765 38301 24777 38335
rect 24811 38301 24823 38335
rect 24765 38295 24823 38301
rect 22833 38267 22891 38273
rect 22833 38233 22845 38267
rect 22879 38264 22891 38267
rect 23750 38264 23756 38276
rect 22879 38236 23756 38264
rect 22879 38233 22891 38236
rect 22833 38227 22891 38233
rect 23750 38224 23756 38236
rect 23808 38224 23814 38276
rect 24780 38264 24808 38295
rect 24854 38292 24860 38344
rect 24912 38332 24918 38344
rect 25038 38332 25044 38344
rect 24912 38304 24957 38332
rect 24999 38304 25044 38332
rect 24912 38292 24918 38304
rect 25038 38292 25044 38304
rect 25096 38292 25102 38344
rect 25590 38292 25596 38344
rect 25648 38332 25654 38344
rect 25700 38341 25728 38440
rect 26326 38400 26332 38412
rect 26287 38372 26332 38400
rect 26326 38360 26332 38372
rect 26384 38360 26390 38412
rect 27706 38400 27712 38412
rect 27667 38372 27712 38400
rect 27706 38360 27712 38372
rect 27764 38360 27770 38412
rect 25685 38335 25743 38341
rect 25685 38332 25697 38335
rect 25648 38304 25697 38332
rect 25648 38292 25654 38304
rect 25685 38301 25697 38304
rect 25731 38301 25743 38335
rect 25866 38332 25872 38344
rect 25827 38304 25872 38332
rect 25685 38295 25743 38301
rect 25866 38292 25872 38304
rect 25924 38292 25930 38344
rect 24946 38264 24952 38276
rect 24780 38236 24952 38264
rect 24946 38224 24952 38236
rect 25004 38224 25010 38276
rect 25501 38267 25559 38273
rect 25501 38233 25513 38267
rect 25547 38233 25559 38267
rect 25501 38227 25559 38233
rect 20956 38168 22784 38196
rect 20956 38156 20962 38168
rect 22922 38156 22928 38208
rect 22980 38196 22986 38208
rect 23842 38196 23848 38208
rect 22980 38168 23848 38196
rect 22980 38156 22986 38168
rect 23842 38156 23848 38168
rect 23900 38156 23906 38208
rect 24397 38199 24455 38205
rect 24397 38165 24409 38199
rect 24443 38196 24455 38199
rect 24670 38196 24676 38208
rect 24443 38168 24676 38196
rect 24443 38165 24455 38168
rect 24397 38159 24455 38165
rect 24670 38156 24676 38168
rect 24728 38156 24734 38208
rect 24762 38156 24768 38208
rect 24820 38196 24826 38208
rect 25516 38196 25544 38227
rect 25774 38224 25780 38276
rect 25832 38264 25838 38276
rect 26513 38267 26571 38273
rect 26513 38264 26525 38267
rect 25832 38236 26525 38264
rect 25832 38224 25838 38236
rect 26513 38233 26525 38236
rect 26559 38233 26571 38267
rect 26513 38227 26571 38233
rect 24820 38168 25544 38196
rect 24820 38156 24826 38168
rect 1104 38106 28888 38128
rect 1104 38054 10214 38106
rect 10266 38054 10278 38106
rect 10330 38054 10342 38106
rect 10394 38054 10406 38106
rect 10458 38054 10470 38106
rect 10522 38054 19478 38106
rect 19530 38054 19542 38106
rect 19594 38054 19606 38106
rect 19658 38054 19670 38106
rect 19722 38054 19734 38106
rect 19786 38054 28888 38106
rect 1104 38032 28888 38054
rect 18322 37992 18328 38004
rect 8312 37964 18328 37992
rect 1765 37927 1823 37933
rect 1765 37893 1777 37927
rect 1811 37924 1823 37927
rect 3786 37924 3792 37936
rect 1811 37896 3792 37924
rect 1811 37893 1823 37896
rect 1765 37887 1823 37893
rect 3786 37884 3792 37896
rect 3844 37884 3850 37936
rect 4065 37927 4123 37933
rect 4065 37893 4077 37927
rect 4111 37924 4123 37927
rect 6457 37927 6515 37933
rect 6457 37924 6469 37927
rect 4111 37896 6469 37924
rect 4111 37893 4123 37896
rect 4065 37887 4123 37893
rect 6457 37893 6469 37896
rect 6503 37893 6515 37927
rect 6457 37887 6515 37893
rect 6362 37856 6368 37868
rect 6323 37828 6368 37856
rect 6362 37816 6368 37828
rect 6420 37816 6426 37868
rect 8312 37865 8340 37964
rect 18322 37952 18328 37964
rect 18380 37952 18386 38004
rect 19886 37992 19892 38004
rect 19847 37964 19892 37992
rect 19886 37952 19892 37964
rect 19944 37952 19950 38004
rect 23382 37952 23388 38004
rect 23440 37992 23446 38004
rect 25038 37992 25044 38004
rect 23440 37964 25044 37992
rect 23440 37952 23446 37964
rect 25038 37952 25044 37964
rect 25096 37952 25102 38004
rect 25130 37952 25136 38004
rect 25188 37992 25194 38004
rect 25188 37964 28028 37992
rect 25188 37952 25194 37964
rect 28000 37936 28028 37964
rect 8404 37896 11836 37924
rect 8297 37859 8355 37865
rect 8297 37825 8309 37859
rect 8343 37825 8355 37859
rect 8297 37819 8355 37825
rect 1581 37791 1639 37797
rect 1581 37757 1593 37791
rect 1627 37757 1639 37791
rect 1581 37751 1639 37757
rect 1596 37720 1624 37751
rect 2774 37748 2780 37800
rect 2832 37788 2838 37800
rect 3878 37788 3884 37800
rect 2832 37760 2877 37788
rect 3839 37760 3884 37788
rect 2832 37748 2838 37760
rect 3878 37748 3884 37760
rect 3936 37748 3942 37800
rect 4522 37788 4528 37800
rect 4483 37760 4528 37788
rect 4522 37748 4528 37760
rect 4580 37748 4586 37800
rect 6914 37748 6920 37800
rect 6972 37788 6978 37800
rect 8404 37788 8432 37896
rect 8849 37859 8907 37865
rect 8849 37825 8861 37859
rect 8895 37856 8907 37859
rect 9766 37856 9772 37868
rect 8895 37828 9772 37856
rect 8895 37825 8907 37828
rect 8849 37819 8907 37825
rect 9766 37816 9772 37828
rect 9824 37856 9830 37868
rect 9953 37859 10011 37865
rect 9953 37856 9965 37859
rect 9824 37828 9965 37856
rect 9824 37816 9830 37828
rect 9953 37825 9965 37828
rect 9999 37856 10011 37859
rect 10410 37856 10416 37868
rect 9999 37828 10416 37856
rect 9999 37825 10011 37828
rect 9953 37819 10011 37825
rect 10410 37816 10416 37828
rect 10468 37816 10474 37868
rect 10502 37816 10508 37868
rect 10560 37856 10566 37868
rect 11054 37856 11060 37868
rect 10560 37828 11060 37856
rect 10560 37816 10566 37828
rect 11054 37816 11060 37828
rect 11112 37816 11118 37868
rect 11238 37816 11244 37868
rect 11296 37856 11302 37868
rect 11422 37856 11428 37868
rect 11296 37828 11428 37856
rect 11296 37816 11302 37828
rect 11422 37816 11428 37828
rect 11480 37816 11486 37868
rect 11514 37816 11520 37868
rect 11572 37856 11578 37868
rect 11701 37859 11759 37865
rect 11701 37856 11713 37859
rect 11572 37828 11713 37856
rect 11572 37816 11578 37828
rect 11701 37825 11713 37828
rect 11747 37825 11759 37859
rect 11808 37856 11836 37896
rect 11882 37884 11888 37936
rect 11940 37924 11946 37936
rect 12618 37924 12624 37936
rect 11940 37896 12624 37924
rect 11940 37884 11946 37896
rect 12618 37884 12624 37896
rect 12676 37884 12682 37936
rect 12802 37884 12808 37936
rect 12860 37924 12866 37936
rect 16914 37927 16972 37933
rect 16914 37924 16926 37927
rect 12860 37896 16926 37924
rect 12860 37884 12866 37896
rect 16914 37893 16926 37896
rect 16960 37893 16972 37927
rect 24765 37927 24823 37933
rect 24765 37924 24777 37927
rect 16914 37887 16972 37893
rect 17021 37896 24777 37924
rect 12345 37859 12403 37865
rect 12345 37856 12357 37859
rect 11808 37828 12357 37856
rect 11701 37819 11759 37825
rect 12345 37825 12357 37828
rect 12391 37825 12403 37859
rect 12345 37819 12403 37825
rect 14366 37816 14372 37868
rect 14424 37856 14430 37868
rect 14829 37859 14887 37865
rect 14829 37856 14841 37859
rect 14424 37828 14841 37856
rect 14424 37816 14430 37828
rect 14829 37825 14841 37828
rect 14875 37825 14887 37859
rect 14829 37819 14887 37825
rect 15933 37859 15991 37865
rect 15933 37825 15945 37859
rect 15979 37856 15991 37859
rect 15979 37828 16160 37856
rect 15979 37825 15991 37828
rect 15933 37819 15991 37825
rect 9122 37788 9128 37800
rect 6972 37760 8432 37788
rect 9083 37760 9128 37788
rect 6972 37748 6978 37760
rect 9122 37748 9128 37760
rect 9180 37748 9186 37800
rect 9306 37748 9312 37800
rect 9364 37788 9370 37800
rect 10042 37788 10048 37800
rect 9364 37760 10048 37788
rect 9364 37748 9370 37760
rect 10042 37748 10048 37760
rect 10100 37748 10106 37800
rect 10134 37748 10140 37800
rect 10192 37788 10198 37800
rect 10781 37791 10839 37797
rect 10781 37788 10793 37791
rect 10192 37760 10793 37788
rect 10192 37748 10198 37760
rect 10781 37757 10793 37760
rect 10827 37788 10839 37791
rect 11606 37788 11612 37800
rect 10827 37760 11612 37788
rect 10827 37757 10839 37760
rect 10781 37751 10839 37757
rect 11606 37748 11612 37760
rect 11664 37748 11670 37800
rect 11793 37791 11851 37797
rect 11793 37757 11805 37791
rect 11839 37788 11851 37791
rect 11974 37788 11980 37800
rect 11839 37760 11980 37788
rect 11839 37757 11851 37760
rect 11793 37751 11851 37757
rect 11974 37748 11980 37760
rect 12032 37748 12038 37800
rect 12158 37748 12164 37800
rect 12216 37788 12222 37800
rect 12529 37791 12587 37797
rect 12529 37788 12541 37791
rect 12216 37760 12541 37788
rect 12216 37748 12222 37760
rect 12529 37757 12541 37760
rect 12575 37757 12587 37791
rect 12894 37788 12900 37800
rect 12855 37760 12900 37788
rect 12529 37751 12587 37757
rect 12894 37748 12900 37760
rect 12952 37748 12958 37800
rect 12986 37748 12992 37800
rect 13044 37788 13050 37800
rect 13446 37788 13452 37800
rect 13044 37760 13452 37788
rect 13044 37748 13050 37760
rect 13446 37748 13452 37760
rect 13504 37748 13510 37800
rect 14642 37788 14648 37800
rect 14603 37760 14648 37788
rect 14642 37748 14648 37760
rect 14700 37748 14706 37800
rect 15746 37788 15752 37800
rect 15707 37760 15752 37788
rect 15746 37748 15752 37760
rect 15804 37748 15810 37800
rect 16132 37788 16160 37828
rect 16206 37816 16212 37868
rect 16264 37856 16270 37868
rect 17021 37856 17049 37896
rect 24765 37893 24777 37896
rect 24811 37893 24823 37927
rect 24765 37887 24823 37893
rect 26421 37927 26479 37933
rect 26421 37893 26433 37927
rect 26467 37924 26479 37927
rect 27062 37924 27068 37936
rect 26467 37896 27068 37924
rect 26467 37893 26479 37896
rect 26421 37887 26479 37893
rect 27062 37884 27068 37896
rect 27120 37884 27126 37936
rect 27982 37924 27988 37936
rect 27943 37896 27988 37924
rect 27982 37884 27988 37896
rect 28040 37884 28046 37936
rect 16264 37828 17049 37856
rect 16264 37816 16270 37828
rect 17310 37816 17316 37868
rect 17368 37856 17374 37868
rect 18765 37859 18823 37865
rect 18765 37856 18777 37859
rect 17368 37828 18777 37856
rect 17368 37816 17374 37828
rect 18765 37825 18777 37828
rect 18811 37825 18823 37859
rect 18765 37819 18823 37825
rect 19058 37816 19064 37868
rect 19116 37856 19122 37868
rect 19116 37828 19564 37856
rect 19116 37816 19122 37828
rect 16482 37788 16488 37800
rect 16132 37760 16488 37788
rect 16482 37748 16488 37760
rect 16540 37748 16546 37800
rect 16669 37791 16727 37797
rect 16669 37757 16681 37791
rect 16715 37757 16727 37791
rect 16669 37751 16727 37757
rect 18509 37791 18567 37797
rect 18509 37757 18521 37791
rect 18555 37757 18567 37791
rect 18509 37751 18567 37757
rect 4430 37720 4436 37732
rect 1596 37692 4436 37720
rect 4430 37680 4436 37692
rect 4488 37680 4494 37732
rect 7653 37723 7711 37729
rect 7653 37689 7665 37723
rect 7699 37720 7711 37723
rect 8294 37720 8300 37732
rect 7699 37692 8300 37720
rect 7699 37689 7711 37692
rect 7653 37683 7711 37689
rect 8294 37680 8300 37692
rect 8352 37680 8358 37732
rect 8478 37680 8484 37732
rect 8536 37720 8542 37732
rect 16117 37723 16175 37729
rect 16117 37720 16129 37723
rect 8536 37692 16129 37720
rect 8536 37680 8542 37692
rect 16117 37689 16129 37692
rect 16163 37689 16175 37723
rect 16117 37683 16175 37689
rect 16390 37680 16396 37732
rect 16448 37720 16454 37732
rect 16684 37720 16712 37751
rect 18414 37720 18420 37732
rect 16448 37692 16712 37720
rect 17604 37692 18420 37720
rect 16448 37680 16454 37692
rect 8110 37652 8116 37664
rect 8071 37624 8116 37652
rect 8110 37612 8116 37624
rect 8168 37612 8174 37664
rect 8386 37612 8392 37664
rect 8444 37652 8450 37664
rect 15013 37655 15071 37661
rect 15013 37652 15025 37655
rect 8444 37624 15025 37652
rect 8444 37612 8450 37624
rect 15013 37621 15025 37624
rect 15059 37621 15071 37655
rect 15013 37615 15071 37621
rect 15194 37612 15200 37664
rect 15252 37652 15258 37664
rect 17604 37652 17632 37692
rect 18414 37680 18420 37692
rect 18472 37680 18478 37732
rect 18046 37652 18052 37664
rect 15252 37624 17632 37652
rect 18007 37624 18052 37652
rect 15252 37612 15258 37624
rect 18046 37612 18052 37624
rect 18104 37612 18110 37664
rect 18524 37652 18552 37751
rect 19150 37652 19156 37664
rect 18524 37624 19156 37652
rect 19150 37612 19156 37624
rect 19208 37612 19214 37664
rect 19536 37652 19564 37828
rect 20346 37816 20352 37868
rect 20404 37856 20410 37868
rect 20441 37859 20499 37865
rect 20441 37856 20453 37859
rect 20404 37828 20453 37856
rect 20404 37816 20410 37828
rect 20441 37825 20453 37828
rect 20487 37825 20499 37859
rect 20806 37856 20812 37868
rect 20767 37828 20812 37856
rect 20441 37819 20499 37825
rect 20806 37816 20812 37828
rect 20864 37816 20870 37868
rect 21818 37856 21824 37868
rect 21779 37828 21824 37856
rect 21818 37816 21824 37828
rect 21876 37816 21882 37868
rect 24578 37856 24584 37868
rect 24539 37828 24584 37856
rect 24578 37816 24584 37828
rect 24636 37816 24642 37868
rect 26786 37816 26792 37868
rect 26844 37856 26850 37868
rect 27157 37859 27215 37865
rect 27157 37856 27169 37859
rect 26844 37828 27169 37856
rect 26844 37816 26850 37828
rect 27157 37825 27169 37828
rect 27203 37825 27215 37859
rect 27157 37819 27215 37825
rect 19978 37748 19984 37800
rect 20036 37788 20042 37800
rect 21634 37788 21640 37800
rect 20036 37760 21640 37788
rect 20036 37748 20042 37760
rect 21634 37748 21640 37760
rect 21692 37748 21698 37800
rect 22002 37788 22008 37800
rect 21963 37760 22008 37788
rect 22002 37748 22008 37760
rect 22060 37748 22066 37800
rect 22281 37791 22339 37797
rect 22281 37757 22293 37791
rect 22327 37757 22339 37791
rect 22281 37751 22339 37757
rect 19610 37680 19616 37732
rect 19668 37720 19674 37732
rect 21726 37720 21732 37732
rect 19668 37692 21732 37720
rect 19668 37680 19674 37692
rect 21726 37680 21732 37692
rect 21784 37680 21790 37732
rect 21910 37680 21916 37732
rect 21968 37720 21974 37732
rect 22296 37720 22324 37751
rect 23842 37748 23848 37800
rect 23900 37788 23906 37800
rect 25038 37788 25044 37800
rect 23900 37760 25044 37788
rect 23900 37748 23906 37760
rect 25038 37748 25044 37760
rect 25096 37748 25102 37800
rect 25590 37748 25596 37800
rect 25648 37788 25654 37800
rect 27341 37791 27399 37797
rect 27341 37788 27353 37791
rect 25648 37760 27353 37788
rect 25648 37748 25654 37760
rect 27341 37757 27353 37760
rect 27387 37757 27399 37791
rect 27341 37751 27399 37757
rect 27433 37791 27491 37797
rect 27433 37757 27445 37791
rect 27479 37757 27491 37791
rect 27433 37751 27491 37757
rect 21968 37692 22324 37720
rect 21968 37680 21974 37692
rect 26418 37680 26424 37732
rect 26476 37720 26482 37732
rect 27448 37720 27476 37751
rect 26476 37692 27476 37720
rect 26476 37680 26482 37692
rect 20438 37652 20444 37664
rect 19536 37624 20444 37652
rect 20438 37612 20444 37624
rect 20496 37612 20502 37664
rect 20806 37612 20812 37664
rect 20864 37652 20870 37664
rect 22922 37652 22928 37664
rect 20864 37624 22928 37652
rect 20864 37612 20870 37624
rect 22922 37612 22928 37624
rect 22980 37612 22986 37664
rect 25682 37612 25688 37664
rect 25740 37652 25746 37664
rect 26973 37655 27031 37661
rect 26973 37652 26985 37655
rect 25740 37624 26985 37652
rect 25740 37612 25746 37624
rect 26973 37621 26985 37624
rect 27019 37621 27031 37655
rect 28074 37652 28080 37664
rect 28035 37624 28080 37652
rect 26973 37615 27031 37621
rect 28074 37612 28080 37624
rect 28132 37612 28138 37664
rect 1104 37562 28888 37584
rect 1104 37510 5582 37562
rect 5634 37510 5646 37562
rect 5698 37510 5710 37562
rect 5762 37510 5774 37562
rect 5826 37510 5838 37562
rect 5890 37510 14846 37562
rect 14898 37510 14910 37562
rect 14962 37510 14974 37562
rect 15026 37510 15038 37562
rect 15090 37510 15102 37562
rect 15154 37510 24110 37562
rect 24162 37510 24174 37562
rect 24226 37510 24238 37562
rect 24290 37510 24302 37562
rect 24354 37510 24366 37562
rect 24418 37510 28888 37562
rect 1104 37488 28888 37510
rect 3878 37408 3884 37460
rect 3936 37448 3942 37460
rect 6365 37451 6423 37457
rect 6365 37448 6377 37451
rect 3936 37420 6377 37448
rect 3936 37408 3942 37420
rect 6365 37417 6377 37420
rect 6411 37417 6423 37451
rect 6365 37411 6423 37417
rect 7101 37451 7159 37457
rect 7101 37417 7113 37451
rect 7147 37448 7159 37451
rect 7190 37448 7196 37460
rect 7147 37420 7196 37448
rect 7147 37417 7159 37420
rect 7101 37411 7159 37417
rect 7190 37408 7196 37420
rect 7248 37408 7254 37460
rect 7745 37451 7803 37457
rect 7745 37417 7757 37451
rect 7791 37448 7803 37451
rect 7834 37448 7840 37460
rect 7791 37420 7840 37448
rect 7791 37417 7803 37420
rect 7745 37411 7803 37417
rect 7834 37408 7840 37420
rect 7892 37408 7898 37460
rect 8110 37408 8116 37460
rect 8168 37448 8174 37460
rect 17310 37448 17316 37460
rect 8168 37420 17316 37448
rect 8168 37408 8174 37420
rect 17310 37408 17316 37420
rect 17368 37408 17374 37460
rect 17773 37451 17831 37457
rect 17773 37417 17785 37451
rect 17819 37448 17831 37451
rect 17862 37448 17868 37460
rect 17819 37420 17868 37448
rect 17819 37417 17831 37420
rect 17773 37411 17831 37417
rect 17862 37408 17868 37420
rect 17920 37448 17926 37460
rect 18233 37451 18291 37457
rect 18233 37448 18245 37451
rect 17920 37420 18245 37448
rect 17920 37408 17926 37420
rect 18233 37417 18245 37420
rect 18279 37417 18291 37451
rect 18233 37411 18291 37417
rect 18322 37408 18328 37460
rect 18380 37448 18386 37460
rect 25406 37448 25412 37460
rect 18380 37420 25412 37448
rect 18380 37408 18386 37420
rect 25406 37408 25412 37420
rect 25464 37408 25470 37460
rect 25590 37408 25596 37460
rect 25648 37448 25654 37460
rect 25777 37451 25835 37457
rect 25777 37448 25789 37451
rect 25648 37420 25789 37448
rect 25648 37408 25654 37420
rect 25777 37417 25789 37420
rect 25823 37417 25835 37451
rect 25777 37411 25835 37417
rect 8941 37383 8999 37389
rect 8941 37349 8953 37383
rect 8987 37349 8999 37383
rect 8941 37343 8999 37349
rect 1854 37312 1860 37324
rect 1815 37284 1860 37312
rect 1854 37272 1860 37284
rect 1912 37272 1918 37324
rect 5442 37312 5448 37324
rect 5403 37284 5448 37312
rect 5442 37272 5448 37284
rect 5500 37272 5506 37324
rect 8956 37312 8984 37343
rect 9582 37340 9588 37392
rect 9640 37380 9646 37392
rect 9766 37380 9772 37392
rect 9640 37352 9772 37380
rect 9640 37340 9646 37352
rect 9766 37340 9772 37352
rect 9824 37340 9830 37392
rect 11422 37380 11428 37392
rect 10152 37352 11428 37380
rect 10152 37312 10180 37352
rect 11422 37340 11428 37352
rect 11480 37340 11486 37392
rect 11514 37340 11520 37392
rect 11572 37380 11578 37392
rect 12710 37380 12716 37392
rect 11572 37352 12716 37380
rect 11572 37340 11578 37352
rect 12710 37340 12716 37352
rect 12768 37340 12774 37392
rect 13265 37383 13323 37389
rect 13265 37380 13277 37383
rect 12820 37352 13277 37380
rect 11974 37312 11980 37324
rect 8956 37284 10180 37312
rect 10244 37284 11861 37312
rect 11935 37284 11980 37312
rect 1397 37247 1455 37253
rect 1397 37213 1409 37247
rect 1443 37213 1455 37247
rect 1397 37207 1455 37213
rect 3881 37247 3939 37253
rect 3881 37213 3893 37247
rect 3927 37244 3939 37247
rect 4338 37244 4344 37256
rect 3927 37216 4344 37244
rect 3927 37213 3939 37216
rect 3881 37207 3939 37213
rect 1412 37108 1440 37207
rect 4338 37204 4344 37216
rect 4396 37244 4402 37256
rect 5077 37247 5135 37253
rect 5077 37244 5089 37247
rect 4396 37216 5089 37244
rect 4396 37204 4402 37216
rect 5077 37213 5089 37216
rect 5123 37213 5135 37247
rect 5077 37207 5135 37213
rect 8110 37204 8116 37256
rect 8168 37244 8174 37256
rect 8389 37247 8447 37253
rect 8389 37244 8401 37247
rect 8168 37216 8401 37244
rect 8168 37204 8174 37216
rect 8389 37213 8401 37216
rect 8435 37213 8447 37247
rect 9122 37244 9128 37256
rect 9083 37216 9128 37244
rect 8389 37207 8447 37213
rect 9122 37204 9128 37216
rect 9180 37204 9186 37256
rect 9585 37247 9643 37253
rect 9585 37213 9597 37247
rect 9631 37244 9643 37247
rect 9674 37244 9680 37256
rect 9631 37216 9680 37244
rect 9631 37213 9643 37216
rect 9585 37207 9643 37213
rect 9674 37204 9680 37216
rect 9732 37204 9738 37256
rect 9766 37204 9772 37256
rect 9824 37244 9830 37256
rect 10244 37244 10272 37284
rect 10410 37244 10416 37256
rect 9824 37216 10272 37244
rect 10371 37216 10416 37244
rect 9824 37204 9830 37216
rect 10410 37204 10416 37216
rect 10468 37244 10474 37256
rect 11609 37247 11667 37253
rect 11609 37244 11621 37247
rect 10468 37216 11621 37244
rect 10468 37204 10474 37216
rect 11609 37213 11621 37216
rect 11655 37213 11667 37247
rect 11833 37244 11861 37284
rect 11974 37272 11980 37284
rect 12032 37272 12038 37324
rect 12526 37312 12532 37324
rect 12084 37284 12532 37312
rect 12084 37244 12112 37284
rect 12526 37272 12532 37284
rect 12584 37272 12590 37324
rect 12820 37312 12848 37352
rect 13265 37349 13277 37352
rect 13311 37349 13323 37383
rect 21358 37380 21364 37392
rect 13265 37343 13323 37349
rect 17420 37352 21364 37380
rect 12636 37284 12848 37312
rect 12897 37315 12955 37321
rect 12636 37244 12664 37284
rect 12897 37281 12909 37315
rect 12943 37312 12955 37315
rect 12986 37312 12992 37324
rect 12943 37284 12992 37312
rect 12943 37281 12955 37284
rect 12897 37275 12955 37281
rect 12986 37272 12992 37284
rect 13044 37312 13050 37324
rect 14182 37312 14188 37324
rect 13044 37284 14188 37312
rect 13044 37272 13050 37284
rect 14182 37272 14188 37284
rect 14240 37272 14246 37324
rect 16390 37312 16396 37324
rect 16351 37284 16396 37312
rect 16390 37272 16396 37284
rect 16448 37272 16454 37324
rect 13067 37244 13125 37247
rect 11833 37216 12112 37244
rect 12176 37216 12664 37244
rect 12912 37241 13125 37244
rect 12912 37216 13079 37241
rect 11609 37207 11667 37213
rect 1578 37176 1584 37188
rect 1539 37148 1584 37176
rect 1578 37136 1584 37148
rect 1636 37136 1642 37188
rect 4246 37136 4252 37188
rect 4304 37176 4310 37188
rect 4433 37179 4491 37185
rect 4433 37176 4445 37179
rect 4304 37148 4445 37176
rect 4304 37136 4310 37148
rect 4433 37145 4445 37148
rect 4479 37176 4491 37179
rect 4706 37176 4712 37188
rect 4479 37148 4712 37176
rect 4479 37145 4491 37148
rect 4433 37139 4491 37145
rect 4706 37136 4712 37148
rect 4764 37176 4770 37188
rect 10686 37176 10692 37188
rect 4764 37148 10692 37176
rect 4764 37136 4770 37148
rect 10686 37136 10692 37148
rect 10744 37136 10750 37188
rect 10870 37176 10876 37188
rect 10831 37148 10876 37176
rect 10870 37136 10876 37148
rect 10928 37136 10934 37188
rect 11054 37136 11060 37188
rect 11112 37176 11118 37188
rect 12176 37176 12204 37216
rect 11112 37148 12204 37176
rect 11112 37136 11118 37148
rect 12250 37136 12256 37188
rect 12308 37176 12314 37188
rect 12912 37176 12940 37216
rect 13067 37207 13079 37216
rect 13113 37207 13125 37241
rect 13067 37201 13125 37207
rect 13630 37204 13636 37256
rect 13688 37244 13694 37256
rect 14090 37244 14096 37256
rect 13688 37216 14096 37244
rect 13688 37204 13694 37216
rect 14090 37204 14096 37216
rect 14148 37244 14154 37256
rect 14553 37247 14611 37253
rect 14553 37244 14565 37247
rect 14148 37216 14565 37244
rect 14148 37204 14154 37216
rect 14553 37213 14565 37216
rect 14599 37244 14611 37247
rect 16408 37244 16436 37272
rect 14599 37216 16436 37244
rect 16546 37216 16804 37244
rect 14599 37213 14611 37216
rect 14553 37207 14611 37213
rect 12308 37148 12940 37176
rect 12308 37136 12314 37148
rect 13722 37136 13728 37188
rect 13780 37176 13786 37188
rect 14798 37179 14856 37185
rect 14798 37176 14810 37179
rect 13780 37148 14810 37176
rect 13780 37136 13786 37148
rect 14798 37145 14810 37148
rect 14844 37145 14856 37179
rect 16546 37176 16574 37216
rect 14798 37139 14856 37145
rect 15672 37148 16574 37176
rect 16660 37179 16718 37185
rect 3878 37108 3884 37120
rect 1412 37080 3884 37108
rect 3878 37068 3884 37080
rect 3936 37068 3942 37120
rect 8205 37111 8263 37117
rect 8205 37077 8217 37111
rect 8251 37108 8263 37111
rect 13078 37108 13084 37120
rect 8251 37080 13084 37108
rect 8251 37077 8263 37080
rect 8205 37071 8263 37077
rect 13078 37068 13084 37080
rect 13136 37068 13142 37120
rect 13262 37068 13268 37120
rect 13320 37108 13326 37120
rect 15672 37108 15700 37148
rect 16660 37145 16672 37179
rect 16706 37145 16718 37179
rect 16776 37176 16804 37216
rect 16942 37204 16948 37256
rect 17000 37244 17006 37256
rect 17420 37244 17448 37352
rect 21358 37340 21364 37352
rect 21416 37380 21422 37392
rect 21416 37352 21588 37380
rect 21416 37340 21422 37352
rect 18046 37272 18052 37324
rect 18104 37312 18110 37324
rect 18104 37284 18552 37312
rect 18104 37272 18110 37284
rect 17000 37216 17448 37244
rect 17000 37204 17006 37216
rect 18138 37204 18144 37256
rect 18196 37244 18202 37256
rect 18233 37247 18291 37253
rect 18233 37244 18245 37247
rect 18196 37216 18245 37244
rect 18196 37204 18202 37216
rect 18233 37213 18245 37216
rect 18279 37213 18291 37247
rect 18233 37207 18291 37213
rect 18322 37204 18328 37256
rect 18380 37244 18386 37256
rect 18524 37253 18552 37284
rect 19352 37284 21128 37312
rect 18417 37247 18475 37253
rect 18417 37244 18429 37247
rect 18380 37216 18429 37244
rect 18380 37204 18386 37216
rect 18417 37213 18429 37216
rect 18463 37213 18475 37247
rect 18417 37207 18475 37213
rect 18509 37247 18567 37253
rect 18509 37213 18521 37247
rect 18555 37244 18567 37247
rect 18690 37244 18696 37256
rect 18555 37216 18696 37244
rect 18555 37213 18567 37216
rect 18509 37207 18567 37213
rect 18690 37204 18696 37216
rect 18748 37204 18754 37256
rect 19352 37253 19380 37284
rect 20364 37256 20392 37284
rect 19337 37247 19395 37253
rect 19337 37213 19349 37247
rect 19383 37213 19395 37247
rect 20346 37244 20352 37256
rect 19337 37207 19395 37213
rect 19444 37216 19748 37244
rect 20259 37216 20352 37244
rect 19444 37176 19472 37216
rect 19610 37176 19616 37188
rect 16776 37148 19472 37176
rect 19571 37148 19616 37176
rect 16660 37139 16718 37145
rect 13320 37080 15700 37108
rect 13320 37068 13326 37080
rect 15746 37068 15752 37120
rect 15804 37108 15810 37120
rect 15933 37111 15991 37117
rect 15933 37108 15945 37111
rect 15804 37080 15945 37108
rect 15804 37068 15810 37080
rect 15933 37077 15945 37080
rect 15979 37077 15991 37111
rect 15933 37071 15991 37077
rect 16022 37068 16028 37120
rect 16080 37108 16086 37120
rect 16675 37108 16703 37139
rect 19610 37136 19616 37148
rect 19668 37136 19674 37188
rect 19720 37176 19748 37216
rect 20346 37204 20352 37216
rect 20404 37204 20410 37256
rect 21100 37244 21128 37284
rect 21450 37244 21456 37256
rect 20456 37216 21036 37244
rect 21100 37216 21456 37244
rect 20456 37176 20484 37216
rect 20898 37176 20904 37188
rect 19720 37148 20484 37176
rect 20859 37148 20904 37176
rect 20898 37136 20904 37148
rect 20956 37136 20962 37188
rect 21008 37176 21036 37216
rect 21450 37204 21456 37216
rect 21508 37204 21514 37256
rect 21560 37244 21588 37352
rect 23474 37272 23480 37324
rect 23532 37312 23538 37324
rect 23842 37312 23848 37324
rect 23532 37284 23848 37312
rect 23532 37272 23538 37284
rect 23842 37272 23848 37284
rect 23900 37272 23906 37324
rect 26510 37312 26516 37324
rect 26471 37284 26516 37312
rect 26510 37272 26516 37284
rect 26568 37272 26574 37324
rect 21729 37247 21787 37253
rect 21729 37244 21741 37247
rect 21560 37216 21741 37244
rect 21729 37213 21741 37216
rect 21775 37213 21787 37247
rect 21729 37207 21787 37213
rect 22465 37247 22523 37253
rect 22465 37213 22477 37247
rect 22511 37244 22523 37247
rect 24397 37247 24455 37253
rect 24397 37244 24409 37247
rect 22511 37216 24409 37244
rect 22511 37213 22523 37216
rect 22465 37207 22523 37213
rect 24397 37213 24409 37216
rect 24443 37244 24455 37247
rect 24486 37244 24492 37256
rect 24443 37216 24492 37244
rect 24443 37213 24455 37216
rect 24397 37207 24455 37213
rect 22002 37176 22008 37188
rect 21008 37148 22008 37176
rect 22002 37136 22008 37148
rect 22060 37136 22066 37188
rect 16080 37080 16703 37108
rect 16080 37068 16086 37080
rect 17954 37068 17960 37120
rect 18012 37108 18018 37120
rect 18693 37111 18751 37117
rect 18693 37108 18705 37111
rect 18012 37080 18705 37108
rect 18012 37068 18018 37080
rect 18693 37077 18705 37080
rect 18739 37077 18751 37111
rect 18693 37071 18751 37077
rect 19150 37068 19156 37120
rect 19208 37108 19214 37120
rect 22480 37108 22508 37207
rect 24486 37204 24492 37216
rect 24544 37204 24550 37256
rect 24670 37253 24676 37256
rect 24664 37244 24676 37253
rect 24631 37216 24676 37244
rect 24664 37207 24676 37216
rect 24670 37204 24676 37207
rect 24728 37204 24734 37256
rect 26234 37204 26240 37256
rect 26292 37244 26298 37256
rect 26329 37247 26387 37253
rect 26329 37244 26341 37247
rect 26292 37216 26341 37244
rect 26292 37204 26298 37216
rect 26329 37213 26341 37216
rect 26375 37213 26387 37247
rect 28166 37244 28172 37256
rect 28127 37216 28172 37244
rect 26329 37207 26387 37213
rect 28166 37204 28172 37216
rect 28224 37204 28230 37256
rect 22554 37136 22560 37188
rect 22612 37176 22618 37188
rect 22710 37179 22768 37185
rect 22710 37176 22722 37179
rect 22612 37148 22722 37176
rect 22612 37136 22618 37148
rect 22710 37145 22722 37148
rect 22756 37145 22768 37179
rect 22710 37139 22768 37145
rect 22830 37136 22836 37188
rect 22888 37176 22894 37188
rect 22888 37148 23980 37176
rect 22888 37136 22894 37148
rect 19208 37080 22508 37108
rect 19208 37068 19214 37080
rect 23106 37068 23112 37120
rect 23164 37108 23170 37120
rect 23658 37108 23664 37120
rect 23164 37080 23664 37108
rect 23164 37068 23170 37080
rect 23658 37068 23664 37080
rect 23716 37108 23722 37120
rect 23845 37111 23903 37117
rect 23845 37108 23857 37111
rect 23716 37080 23857 37108
rect 23716 37068 23722 37080
rect 23845 37077 23857 37080
rect 23891 37077 23903 37111
rect 23952 37108 23980 37148
rect 28074 37108 28080 37120
rect 23952 37080 28080 37108
rect 23845 37071 23903 37077
rect 28074 37068 28080 37080
rect 28132 37068 28138 37120
rect 1104 37018 28888 37040
rect 1104 36966 10214 37018
rect 10266 36966 10278 37018
rect 10330 36966 10342 37018
rect 10394 36966 10406 37018
rect 10458 36966 10470 37018
rect 10522 36966 19478 37018
rect 19530 36966 19542 37018
rect 19594 36966 19606 37018
rect 19658 36966 19670 37018
rect 19722 36966 19734 37018
rect 19786 36966 28888 37018
rect 1104 36944 28888 36966
rect 1578 36904 1584 36916
rect 1539 36876 1584 36904
rect 1578 36864 1584 36876
rect 1636 36864 1642 36916
rect 2317 36907 2375 36913
rect 2317 36873 2329 36907
rect 2363 36904 2375 36907
rect 2590 36904 2596 36916
rect 2363 36876 2596 36904
rect 2363 36873 2375 36876
rect 2317 36867 2375 36873
rect 2590 36864 2596 36876
rect 2648 36904 2654 36916
rect 9674 36904 9680 36916
rect 2648 36876 2774 36904
rect 2648 36864 2654 36876
rect 1489 36771 1547 36777
rect 1489 36737 1501 36771
rect 1535 36768 1547 36771
rect 1578 36768 1584 36780
rect 1535 36740 1584 36768
rect 1535 36737 1547 36740
rect 1489 36731 1547 36737
rect 1578 36728 1584 36740
rect 1636 36728 1642 36780
rect 2133 36771 2191 36777
rect 2133 36737 2145 36771
rect 2179 36737 2191 36771
rect 2746 36768 2774 36876
rect 7760 36876 9680 36904
rect 4982 36836 4988 36848
rect 4895 36808 4988 36836
rect 4982 36796 4988 36808
rect 5040 36836 5046 36848
rect 5350 36836 5356 36848
rect 5040 36808 5356 36836
rect 5040 36796 5046 36808
rect 5350 36796 5356 36808
rect 5408 36796 5414 36848
rect 3053 36771 3111 36777
rect 3053 36768 3065 36771
rect 2746 36740 3065 36768
rect 2133 36731 2191 36737
rect 3053 36737 3065 36740
rect 3099 36768 3111 36771
rect 4338 36768 4344 36780
rect 3099 36740 4344 36768
rect 3099 36737 3111 36740
rect 3053 36731 3111 36737
rect 2038 36592 2044 36644
rect 2096 36632 2102 36644
rect 2148 36632 2176 36731
rect 4338 36728 4344 36740
rect 4396 36768 4402 36780
rect 4433 36771 4491 36777
rect 4433 36768 4445 36771
rect 4396 36740 4445 36768
rect 4396 36728 4402 36740
rect 4433 36737 4445 36740
rect 4479 36737 4491 36771
rect 4433 36731 4491 36737
rect 5166 36728 5172 36780
rect 5224 36768 5230 36780
rect 5721 36771 5779 36777
rect 5721 36768 5733 36771
rect 5224 36740 5733 36768
rect 5224 36728 5230 36740
rect 5721 36737 5733 36740
rect 5767 36737 5779 36771
rect 5721 36731 5779 36737
rect 7101 36771 7159 36777
rect 7101 36737 7113 36771
rect 7147 36768 7159 36771
rect 7282 36768 7288 36780
rect 7147 36740 7288 36768
rect 7147 36737 7159 36740
rect 7101 36731 7159 36737
rect 7282 36728 7288 36740
rect 7340 36728 7346 36780
rect 3694 36700 3700 36712
rect 3655 36672 3700 36700
rect 3694 36660 3700 36672
rect 3752 36660 3758 36712
rect 7760 36632 7788 36876
rect 9674 36864 9680 36876
rect 9732 36864 9738 36916
rect 9769 36907 9827 36913
rect 9769 36873 9781 36907
rect 9815 36904 9827 36907
rect 12434 36904 12440 36916
rect 9815 36876 12440 36904
rect 9815 36873 9827 36876
rect 9769 36867 9827 36873
rect 12434 36864 12440 36876
rect 12492 36864 12498 36916
rect 12526 36864 12532 36916
rect 12584 36904 12590 36916
rect 12584 36876 14136 36904
rect 12584 36864 12590 36876
rect 8846 36796 8852 36848
rect 8904 36836 8910 36848
rect 9033 36839 9091 36845
rect 9033 36836 9045 36839
rect 8904 36808 9045 36836
rect 8904 36796 8910 36808
rect 9033 36805 9045 36808
rect 9079 36805 9091 36839
rect 11054 36836 11060 36848
rect 9033 36799 9091 36805
rect 9600 36808 11060 36836
rect 7837 36771 7895 36777
rect 7837 36737 7849 36771
rect 7883 36768 7895 36771
rect 8202 36768 8208 36780
rect 7883 36740 8208 36768
rect 7883 36737 7895 36740
rect 7837 36731 7895 36737
rect 8202 36728 8208 36740
rect 8260 36728 8266 36780
rect 8478 36768 8484 36780
rect 8439 36740 8484 36768
rect 8478 36728 8484 36740
rect 8536 36728 8542 36780
rect 8938 36768 8944 36780
rect 8899 36740 8944 36768
rect 8938 36728 8944 36740
rect 8996 36728 9002 36780
rect 9125 36771 9183 36777
rect 9125 36737 9137 36771
rect 9171 36768 9183 36771
rect 9214 36768 9220 36780
rect 9171 36740 9220 36768
rect 9171 36737 9183 36740
rect 9125 36731 9183 36737
rect 7926 36660 7932 36712
rect 7984 36700 7990 36712
rect 9140 36700 9168 36731
rect 9214 36728 9220 36740
rect 9272 36728 9278 36780
rect 9600 36777 9628 36808
rect 11054 36796 11060 36808
rect 11112 36796 11118 36848
rect 12060 36839 12118 36845
rect 12060 36805 12072 36839
rect 12106 36836 12118 36839
rect 12158 36836 12164 36848
rect 12106 36808 12164 36836
rect 12106 36805 12118 36808
rect 12060 36799 12118 36805
rect 12158 36796 12164 36808
rect 12216 36796 12222 36848
rect 12618 36796 12624 36848
rect 12676 36836 12682 36848
rect 13262 36836 13268 36848
rect 12676 36808 13268 36836
rect 12676 36796 12682 36808
rect 13262 36796 13268 36808
rect 13320 36796 13326 36848
rect 14108 36836 14136 36876
rect 14642 36864 14648 36916
rect 14700 36904 14706 36916
rect 15010 36904 15016 36916
rect 14700 36876 15016 36904
rect 14700 36864 14706 36876
rect 15010 36864 15016 36876
rect 15068 36864 15074 36916
rect 15470 36864 15476 36916
rect 15528 36904 15534 36916
rect 15657 36907 15715 36913
rect 15657 36904 15669 36907
rect 15528 36876 15669 36904
rect 15528 36864 15534 36876
rect 15657 36873 15669 36876
rect 15703 36873 15715 36907
rect 15657 36867 15715 36873
rect 16025 36907 16083 36913
rect 16025 36873 16037 36907
rect 16071 36904 16083 36907
rect 18138 36904 18144 36916
rect 16071 36876 18144 36904
rect 16071 36873 16083 36876
rect 16025 36867 16083 36873
rect 18138 36864 18144 36876
rect 18196 36864 18202 36916
rect 18877 36907 18935 36913
rect 18877 36873 18889 36907
rect 18923 36904 18935 36907
rect 20162 36904 20168 36916
rect 18923 36876 20168 36904
rect 18923 36873 18935 36876
rect 18877 36867 18935 36873
rect 20162 36864 20168 36876
rect 20220 36864 20226 36916
rect 21450 36864 21456 36916
rect 21508 36904 21514 36916
rect 22005 36907 22063 36913
rect 22005 36904 22017 36907
rect 21508 36876 22017 36904
rect 21508 36864 21514 36876
rect 22005 36873 22017 36876
rect 22051 36873 22063 36907
rect 22370 36904 22376 36916
rect 22005 36867 22063 36873
rect 22112 36876 22376 36904
rect 22112 36836 22140 36876
rect 22370 36864 22376 36876
rect 22428 36864 22434 36916
rect 22554 36904 22560 36916
rect 22515 36876 22560 36904
rect 22554 36864 22560 36876
rect 22612 36864 22618 36916
rect 22646 36864 22652 36916
rect 22704 36904 22710 36916
rect 24029 36907 24087 36913
rect 24029 36904 24041 36907
rect 22704 36876 24041 36904
rect 22704 36864 22710 36876
rect 24029 36873 24041 36876
rect 24075 36873 24087 36907
rect 24029 36867 24087 36873
rect 24118 36864 24124 36916
rect 24176 36904 24182 36916
rect 26418 36904 26424 36916
rect 24176 36876 26424 36904
rect 24176 36864 24182 36876
rect 26418 36864 26424 36876
rect 26476 36864 26482 36916
rect 26970 36864 26976 36916
rect 27028 36904 27034 36916
rect 27341 36907 27399 36913
rect 27341 36904 27353 36907
rect 27028 36876 27353 36904
rect 27028 36864 27034 36876
rect 27341 36873 27353 36876
rect 27387 36873 27399 36907
rect 27341 36867 27399 36873
rect 23290 36836 23296 36848
rect 13464 36808 14044 36836
rect 14108 36808 22140 36836
rect 22940 36808 23296 36836
rect 9585 36771 9643 36777
rect 9585 36737 9597 36771
rect 9631 36737 9643 36771
rect 9766 36768 9772 36780
rect 9727 36740 9772 36768
rect 9585 36731 9643 36737
rect 9766 36728 9772 36740
rect 9824 36728 9830 36780
rect 10042 36728 10048 36780
rect 10100 36768 10106 36780
rect 10321 36771 10379 36777
rect 10321 36768 10333 36771
rect 10100 36740 10333 36768
rect 10100 36728 10106 36740
rect 10321 36737 10333 36740
rect 10367 36737 10379 36771
rect 10321 36731 10379 36737
rect 10410 36728 10416 36780
rect 10468 36768 10474 36780
rect 10778 36768 10784 36780
rect 10468 36740 10640 36768
rect 10739 36740 10784 36768
rect 10468 36728 10474 36740
rect 7984 36672 9168 36700
rect 7984 36660 7990 36672
rect 9398 36660 9404 36712
rect 9456 36700 9462 36712
rect 10612 36700 10640 36740
rect 10778 36728 10784 36740
rect 10836 36728 10842 36780
rect 10962 36728 10968 36780
rect 11020 36768 11026 36780
rect 11422 36768 11428 36780
rect 11020 36740 11428 36768
rect 11020 36728 11026 36740
rect 11422 36728 11428 36740
rect 11480 36728 11486 36780
rect 13464 36768 13492 36808
rect 11716 36740 13492 36768
rect 11514 36700 11520 36712
rect 9456 36672 10548 36700
rect 10612 36672 11520 36700
rect 9456 36660 9462 36672
rect 2096 36604 7788 36632
rect 8297 36635 8355 36641
rect 2096 36592 2102 36604
rect 8297 36601 8309 36635
rect 8343 36632 8355 36635
rect 10520 36632 10548 36672
rect 11514 36660 11520 36672
rect 11572 36660 11578 36712
rect 11606 36632 11612 36644
rect 8343 36604 10464 36632
rect 10520 36604 11612 36632
rect 8343 36601 8355 36604
rect 8297 36595 8355 36601
rect 8110 36524 8116 36576
rect 8168 36564 8174 36576
rect 10318 36564 10324 36576
rect 8168 36536 10324 36564
rect 8168 36524 8174 36536
rect 10318 36524 10324 36536
rect 10376 36524 10382 36576
rect 10436 36564 10464 36604
rect 11606 36592 11612 36604
rect 11664 36592 11670 36644
rect 11716 36564 11744 36740
rect 13538 36728 13544 36780
rect 13596 36768 13602 36780
rect 13889 36771 13947 36777
rect 13889 36768 13901 36771
rect 13596 36740 13901 36768
rect 13596 36728 13602 36740
rect 13889 36737 13901 36740
rect 13935 36737 13947 36771
rect 14016 36768 14044 36808
rect 14016 36740 14688 36768
rect 13889 36731 13947 36737
rect 11793 36703 11851 36709
rect 11793 36669 11805 36703
rect 11839 36669 11851 36703
rect 13630 36700 13636 36712
rect 11793 36663 11851 36669
rect 12800 36672 13636 36700
rect 11815 36576 11843 36663
rect 10436 36536 11744 36564
rect 11790 36524 11796 36576
rect 11848 36564 11854 36576
rect 12800 36564 12828 36672
rect 13630 36660 13636 36672
rect 13688 36660 13694 36712
rect 14660 36700 14688 36740
rect 15010 36728 15016 36780
rect 15068 36768 15074 36780
rect 15473 36771 15531 36777
rect 15473 36768 15485 36771
rect 15068 36740 15485 36768
rect 15068 36728 15074 36740
rect 15473 36737 15485 36740
rect 15519 36768 15531 36771
rect 15562 36768 15568 36780
rect 15519 36740 15568 36768
rect 15519 36737 15531 36740
rect 15473 36731 15531 36737
rect 15562 36728 15568 36740
rect 15620 36728 15626 36780
rect 15746 36768 15752 36780
rect 15707 36740 15752 36768
rect 15746 36728 15752 36740
rect 15804 36728 15810 36780
rect 15838 36728 15844 36780
rect 15896 36768 15902 36780
rect 16669 36771 16727 36777
rect 16669 36768 16681 36771
rect 15896 36740 16681 36768
rect 15896 36728 15902 36740
rect 16669 36737 16681 36740
rect 16715 36737 16727 36771
rect 16669 36731 16727 36737
rect 16853 36771 16911 36777
rect 16853 36737 16865 36771
rect 16899 36737 16911 36771
rect 16853 36731 16911 36737
rect 17764 36771 17822 36777
rect 17764 36737 17776 36771
rect 17810 36768 17822 36771
rect 18046 36768 18052 36780
rect 17810 36740 18052 36768
rect 17810 36737 17822 36740
rect 17764 36731 17822 36737
rect 16022 36700 16028 36712
rect 14660 36672 16028 36700
rect 16022 36660 16028 36672
rect 16080 36660 16086 36712
rect 16206 36660 16212 36712
rect 16264 36700 16270 36712
rect 16868 36700 16896 36731
rect 18046 36728 18052 36740
rect 18104 36728 18110 36780
rect 19058 36728 19064 36780
rect 19116 36768 19122 36780
rect 19593 36771 19651 36777
rect 19593 36768 19605 36771
rect 19116 36740 19605 36768
rect 19116 36728 19122 36740
rect 19593 36737 19605 36740
rect 19639 36737 19651 36771
rect 19593 36731 19651 36737
rect 20898 36728 20904 36780
rect 20956 36768 20962 36780
rect 21450 36768 21456 36780
rect 20956 36740 21456 36768
rect 20956 36728 20962 36740
rect 21450 36728 21456 36740
rect 21508 36728 21514 36780
rect 21910 36768 21916 36780
rect 21871 36740 21916 36768
rect 21910 36728 21916 36740
rect 21968 36728 21974 36780
rect 22940 36777 22968 36808
rect 23290 36796 23296 36808
rect 23348 36836 23354 36848
rect 24946 36836 24952 36848
rect 23348 36808 24952 36836
rect 23348 36796 23354 36808
rect 24946 36796 24952 36808
rect 25004 36796 25010 36848
rect 28350 36836 28356 36848
rect 27080 36808 28356 36836
rect 22833 36771 22891 36777
rect 22833 36737 22845 36771
rect 22879 36737 22891 36771
rect 22833 36731 22891 36737
rect 22925 36771 22983 36777
rect 22925 36737 22937 36771
rect 22971 36737 22983 36771
rect 22925 36731 22983 36737
rect 17034 36700 17040 36712
rect 16264 36672 16896 36700
rect 16995 36672 17040 36700
rect 16264 36660 16270 36672
rect 17034 36660 17040 36672
rect 17092 36660 17098 36712
rect 17497 36703 17555 36709
rect 17497 36669 17509 36703
rect 17543 36669 17555 36703
rect 17497 36663 17555 36669
rect 13078 36592 13084 36644
rect 13136 36632 13142 36644
rect 13173 36635 13231 36641
rect 13173 36632 13185 36635
rect 13136 36604 13185 36632
rect 13136 36592 13142 36604
rect 13173 36601 13185 36604
rect 13219 36601 13231 36635
rect 13173 36595 13231 36601
rect 16390 36592 16396 36644
rect 16448 36632 16454 36644
rect 17512 36632 17540 36663
rect 19150 36660 19156 36712
rect 19208 36700 19214 36712
rect 19337 36703 19395 36709
rect 19337 36700 19349 36703
rect 19208 36672 19349 36700
rect 19208 36660 19214 36672
rect 19337 36669 19349 36672
rect 19383 36669 19395 36703
rect 19337 36663 19395 36669
rect 20806 36660 20812 36712
rect 20864 36700 20870 36712
rect 22848 36700 22876 36731
rect 23014 36728 23020 36780
rect 23072 36768 23078 36780
rect 23201 36771 23259 36777
rect 23072 36740 23117 36768
rect 23072 36728 23078 36740
rect 23201 36737 23213 36771
rect 23247 36737 23259 36771
rect 23201 36731 23259 36737
rect 23106 36700 23112 36712
rect 20864 36672 23112 36700
rect 20864 36660 20870 36672
rect 23106 36660 23112 36672
rect 23164 36660 23170 36712
rect 23216 36700 23244 36731
rect 23474 36728 23480 36780
rect 23532 36768 23538 36780
rect 23845 36771 23903 36777
rect 23845 36768 23857 36771
rect 23532 36740 23857 36768
rect 23532 36728 23538 36740
rect 23845 36737 23857 36740
rect 23891 36737 23903 36771
rect 24118 36768 24124 36780
rect 24079 36740 24124 36768
rect 23845 36731 23903 36737
rect 24118 36728 24124 36740
rect 24176 36728 24182 36780
rect 24578 36768 24584 36780
rect 24539 36740 24584 36768
rect 24578 36728 24584 36740
rect 24636 36728 24642 36780
rect 26421 36771 26479 36777
rect 26421 36737 26433 36771
rect 26467 36768 26479 36771
rect 27080 36768 27108 36808
rect 28350 36796 28356 36808
rect 28408 36796 28414 36848
rect 26467 36740 27108 36768
rect 26467 36737 26479 36740
rect 26421 36731 26479 36737
rect 27154 36728 27160 36780
rect 27212 36768 27218 36780
rect 27430 36768 27436 36780
rect 27212 36740 27257 36768
rect 27391 36740 27436 36768
rect 27212 36728 27218 36740
rect 27430 36728 27436 36740
rect 27488 36728 27494 36780
rect 27893 36771 27951 36777
rect 27893 36737 27905 36771
rect 27939 36737 27951 36771
rect 27893 36731 27951 36737
rect 23382 36700 23388 36712
rect 23216 36672 23388 36700
rect 23382 36660 23388 36672
rect 23440 36700 23446 36712
rect 23658 36700 23664 36712
rect 23440 36672 23664 36700
rect 23440 36660 23446 36672
rect 23658 36660 23664 36672
rect 23716 36660 23722 36712
rect 24765 36703 24823 36709
rect 24765 36669 24777 36703
rect 24811 36669 24823 36703
rect 24765 36663 24823 36669
rect 16448 36604 17540 36632
rect 16448 36592 16454 36604
rect 18506 36592 18512 36644
rect 18564 36632 18570 36644
rect 19242 36632 19248 36644
rect 18564 36604 19248 36632
rect 18564 36592 18570 36604
rect 19242 36592 19248 36604
rect 19300 36592 19306 36644
rect 21542 36632 21548 36644
rect 20640 36604 21548 36632
rect 11848 36536 12828 36564
rect 11848 36524 11854 36536
rect 13446 36524 13452 36576
rect 13504 36564 13510 36576
rect 20640 36564 20668 36604
rect 21542 36592 21548 36604
rect 21600 36592 21606 36644
rect 21818 36592 21824 36644
rect 21876 36632 21882 36644
rect 24780 36632 24808 36663
rect 26878 36660 26884 36712
rect 26936 36700 26942 36712
rect 26973 36703 27031 36709
rect 26973 36700 26985 36703
rect 26936 36672 26985 36700
rect 26936 36660 26942 36672
rect 26973 36669 26985 36672
rect 27019 36669 27031 36703
rect 26973 36663 27031 36669
rect 27062 36660 27068 36712
rect 27120 36700 27126 36712
rect 27908 36700 27936 36731
rect 27120 36672 27936 36700
rect 28169 36703 28227 36709
rect 27120 36660 27126 36672
rect 28169 36669 28181 36703
rect 28215 36700 28227 36703
rect 28350 36700 28356 36712
rect 28215 36672 28356 36700
rect 28215 36669 28227 36672
rect 28169 36663 28227 36669
rect 28350 36660 28356 36672
rect 28408 36660 28414 36712
rect 21876 36604 24808 36632
rect 21876 36592 21882 36604
rect 27614 36592 27620 36644
rect 27672 36632 27678 36644
rect 28077 36635 28135 36641
rect 28077 36632 28089 36635
rect 27672 36604 28089 36632
rect 27672 36592 27678 36604
rect 28077 36601 28089 36604
rect 28123 36601 28135 36635
rect 28077 36595 28135 36601
rect 13504 36536 20668 36564
rect 20717 36567 20775 36573
rect 13504 36524 13510 36536
rect 20717 36533 20729 36567
rect 20763 36564 20775 36567
rect 20806 36564 20812 36576
rect 20763 36536 20812 36564
rect 20763 36533 20775 36536
rect 20717 36527 20775 36533
rect 20806 36524 20812 36536
rect 20864 36524 20870 36576
rect 23661 36567 23719 36573
rect 23661 36533 23673 36567
rect 23707 36564 23719 36567
rect 24762 36564 24768 36576
rect 23707 36536 24768 36564
rect 23707 36533 23719 36536
rect 23661 36527 23719 36533
rect 24762 36524 24768 36536
rect 24820 36524 24826 36576
rect 27890 36524 27896 36576
rect 27948 36564 27954 36576
rect 27985 36567 28043 36573
rect 27985 36564 27997 36567
rect 27948 36536 27997 36564
rect 27948 36524 27954 36536
rect 27985 36533 27997 36536
rect 28031 36533 28043 36567
rect 27985 36527 28043 36533
rect 1104 36474 28888 36496
rect 1104 36422 5582 36474
rect 5634 36422 5646 36474
rect 5698 36422 5710 36474
rect 5762 36422 5774 36474
rect 5826 36422 5838 36474
rect 5890 36422 14846 36474
rect 14898 36422 14910 36474
rect 14962 36422 14974 36474
rect 15026 36422 15038 36474
rect 15090 36422 15102 36474
rect 15154 36422 24110 36474
rect 24162 36422 24174 36474
rect 24226 36422 24238 36474
rect 24290 36422 24302 36474
rect 24354 36422 24366 36474
rect 24418 36422 28888 36474
rect 1104 36400 28888 36422
rect 1486 36320 1492 36372
rect 1544 36360 1550 36372
rect 1673 36363 1731 36369
rect 1673 36360 1685 36363
rect 1544 36332 1685 36360
rect 1544 36320 1550 36332
rect 1673 36329 1685 36332
rect 1719 36329 1731 36363
rect 1673 36323 1731 36329
rect 3881 36363 3939 36369
rect 3881 36329 3893 36363
rect 3927 36360 3939 36363
rect 3970 36360 3976 36372
rect 3927 36332 3976 36360
rect 3927 36329 3939 36332
rect 3881 36323 3939 36329
rect 3970 36320 3976 36332
rect 4028 36320 4034 36372
rect 4614 36360 4620 36372
rect 4575 36332 4620 36360
rect 4614 36320 4620 36332
rect 4672 36320 4678 36372
rect 5258 36360 5264 36372
rect 5219 36332 5264 36360
rect 5258 36320 5264 36332
rect 5316 36320 5322 36372
rect 6457 36363 6515 36369
rect 6457 36329 6469 36363
rect 6503 36360 6515 36363
rect 6914 36360 6920 36372
rect 6503 36332 6920 36360
rect 6503 36329 6515 36332
rect 6457 36323 6515 36329
rect 6914 36320 6920 36332
rect 6972 36320 6978 36372
rect 7098 36360 7104 36372
rect 7059 36332 7104 36360
rect 7098 36320 7104 36332
rect 7156 36320 7162 36372
rect 9306 36360 9312 36372
rect 7484 36332 9312 36360
rect 6730 36252 6736 36304
rect 6788 36292 6794 36304
rect 7484 36292 7512 36332
rect 9306 36320 9312 36332
rect 9364 36320 9370 36372
rect 9582 36360 9588 36372
rect 9543 36332 9588 36360
rect 9582 36320 9588 36332
rect 9640 36320 9646 36372
rect 11241 36363 11299 36369
rect 11241 36360 11253 36363
rect 10152 36332 11253 36360
rect 6788 36264 7512 36292
rect 6788 36252 6794 36264
rect 7558 36252 7564 36304
rect 7616 36292 7622 36304
rect 8205 36295 8263 36301
rect 7616 36264 7661 36292
rect 7616 36252 7622 36264
rect 8205 36261 8217 36295
rect 8251 36261 8263 36295
rect 8938 36292 8944 36304
rect 8899 36264 8944 36292
rect 8205 36255 8263 36261
rect 1578 36184 1584 36236
rect 1636 36224 1642 36236
rect 3145 36227 3203 36233
rect 3145 36224 3157 36227
rect 1636 36196 3157 36224
rect 1636 36184 1642 36196
rect 3145 36193 3157 36196
rect 3191 36224 3203 36227
rect 6362 36224 6368 36236
rect 3191 36196 6368 36224
rect 3191 36193 3203 36196
rect 3145 36187 3203 36193
rect 6362 36184 6368 36196
rect 6420 36184 6426 36236
rect 8220 36224 8248 36255
rect 8938 36252 8944 36264
rect 8996 36252 9002 36304
rect 9122 36252 9128 36304
rect 9180 36292 9186 36304
rect 10152 36292 10180 36332
rect 11241 36329 11253 36332
rect 11287 36329 11299 36363
rect 13630 36360 13636 36372
rect 11241 36323 11299 36329
rect 11833 36332 13636 36360
rect 9180 36264 10180 36292
rect 10321 36295 10379 36301
rect 9180 36252 9186 36264
rect 10321 36261 10333 36295
rect 10367 36292 10379 36295
rect 10594 36292 10600 36304
rect 10367 36264 10600 36292
rect 10367 36261 10379 36264
rect 10321 36255 10379 36261
rect 10594 36252 10600 36264
rect 10652 36252 10658 36304
rect 11833 36292 11861 36332
rect 13630 36320 13636 36332
rect 13688 36320 13694 36372
rect 13722 36320 13728 36372
rect 13780 36360 13786 36372
rect 14366 36360 14372 36372
rect 13780 36332 14372 36360
rect 13780 36320 13786 36332
rect 14366 36320 14372 36332
rect 14424 36320 14430 36372
rect 14458 36320 14464 36372
rect 14516 36360 14522 36372
rect 15378 36360 15384 36372
rect 14516 36332 15384 36360
rect 14516 36320 14522 36332
rect 15378 36320 15384 36332
rect 15436 36320 15442 36372
rect 15930 36320 15936 36372
rect 15988 36360 15994 36372
rect 15988 36332 17721 36360
rect 15988 36320 15994 36332
rect 10704 36264 11861 36292
rect 10704 36224 10732 36264
rect 12986 36252 12992 36304
rect 13044 36292 13050 36304
rect 13998 36292 14004 36304
rect 13044 36264 14004 36292
rect 13044 36252 13050 36264
rect 13998 36252 14004 36264
rect 14056 36252 14062 36304
rect 15286 36252 15292 36304
rect 15344 36292 15350 36304
rect 15473 36295 15531 36301
rect 15473 36292 15485 36295
rect 15344 36264 15485 36292
rect 15344 36252 15350 36264
rect 15473 36261 15485 36264
rect 15519 36292 15531 36295
rect 15838 36292 15844 36304
rect 15519 36264 15844 36292
rect 15519 36261 15531 36264
rect 15473 36255 15531 36261
rect 15838 36252 15844 36264
rect 15896 36252 15902 36304
rect 17693 36292 17721 36332
rect 17862 36320 17868 36372
rect 17920 36360 17926 36372
rect 17920 36332 19104 36360
rect 17920 36320 17926 36332
rect 18874 36292 18880 36304
rect 17693 36264 18880 36292
rect 18874 36252 18880 36264
rect 18932 36252 18938 36304
rect 19076 36292 19104 36332
rect 19518 36320 19524 36372
rect 19576 36360 19582 36372
rect 19576 36332 22968 36360
rect 19576 36320 19582 36332
rect 21818 36292 21824 36304
rect 19076 36264 21824 36292
rect 21818 36252 21824 36264
rect 21876 36252 21882 36304
rect 22002 36292 22008 36304
rect 21963 36264 22008 36292
rect 22002 36252 22008 36264
rect 22060 36252 22066 36304
rect 22940 36292 22968 36332
rect 23014 36320 23020 36372
rect 23072 36360 23078 36372
rect 23385 36363 23443 36369
rect 23385 36360 23397 36363
rect 23072 36332 23397 36360
rect 23072 36320 23078 36332
rect 23385 36329 23397 36332
rect 23431 36329 23443 36363
rect 23385 36323 23443 36329
rect 23566 36320 23572 36372
rect 23624 36360 23630 36372
rect 24670 36360 24676 36372
rect 23624 36332 24676 36360
rect 23624 36320 23630 36332
rect 24670 36320 24676 36332
rect 24728 36320 24734 36372
rect 24854 36320 24860 36372
rect 24912 36360 24918 36372
rect 25041 36363 25099 36369
rect 25041 36360 25053 36363
rect 24912 36332 25053 36360
rect 24912 36320 24918 36332
rect 25041 36329 25053 36332
rect 25087 36329 25099 36363
rect 27430 36360 27436 36372
rect 25041 36323 25099 36329
rect 25746 36332 27436 36360
rect 25746 36292 25774 36332
rect 27430 36320 27436 36332
rect 27488 36320 27494 36372
rect 25866 36292 25872 36304
rect 22940 36264 25774 36292
rect 25827 36264 25872 36292
rect 8220 36196 10732 36224
rect 10778 36184 10784 36236
rect 10836 36224 10842 36236
rect 10873 36227 10931 36233
rect 10873 36224 10885 36227
rect 10836 36196 10885 36224
rect 10836 36184 10842 36196
rect 10873 36193 10885 36196
rect 10919 36193 10931 36227
rect 11790 36224 11796 36236
rect 11751 36196 11796 36224
rect 10873 36187 10931 36193
rect 11790 36184 11796 36196
rect 11848 36184 11854 36236
rect 14090 36224 14096 36236
rect 14051 36196 14096 36224
rect 14090 36184 14096 36196
rect 14148 36184 14154 36236
rect 15654 36184 15660 36236
rect 15712 36224 15718 36236
rect 16390 36224 16396 36236
rect 15712 36196 16396 36224
rect 15712 36184 15718 36196
rect 16390 36184 16396 36196
rect 16448 36224 16454 36236
rect 16761 36227 16819 36233
rect 16761 36224 16773 36227
rect 16448 36196 16773 36224
rect 16448 36184 16454 36196
rect 16761 36193 16773 36196
rect 16807 36193 16819 36227
rect 18506 36224 18512 36236
rect 16761 36187 16819 36193
rect 17779 36196 18512 36224
rect 2590 36156 2596 36168
rect 2551 36128 2596 36156
rect 2590 36116 2596 36128
rect 2648 36116 2654 36168
rect 3694 36116 3700 36168
rect 3752 36156 3758 36168
rect 3789 36159 3847 36165
rect 3789 36156 3801 36159
rect 3752 36128 3801 36156
rect 3752 36116 3758 36128
rect 3789 36125 3801 36128
rect 3835 36125 3847 36159
rect 3789 36119 3847 36125
rect 7745 36159 7803 36165
rect 7745 36125 7757 36159
rect 7791 36156 7803 36159
rect 7834 36156 7840 36168
rect 7791 36128 7840 36156
rect 7791 36125 7803 36128
rect 7745 36119 7803 36125
rect 7834 36116 7840 36128
rect 7892 36116 7898 36168
rect 8386 36156 8392 36168
rect 8347 36128 8392 36156
rect 8386 36116 8392 36128
rect 8444 36116 8450 36168
rect 9125 36159 9183 36165
rect 9125 36125 9137 36159
rect 9171 36125 9183 36159
rect 9766 36156 9772 36168
rect 9727 36128 9772 36156
rect 9125 36119 9183 36125
rect 9140 36020 9168 36119
rect 9766 36116 9772 36128
rect 9824 36116 9830 36168
rect 10229 36159 10287 36165
rect 10229 36125 10241 36159
rect 10275 36156 10287 36159
rect 10962 36156 10968 36168
rect 10275 36128 10968 36156
rect 10275 36125 10287 36128
rect 10229 36119 10287 36125
rect 10962 36116 10968 36128
rect 11020 36116 11026 36168
rect 11054 36116 11060 36168
rect 11112 36156 11118 36168
rect 11112 36128 11157 36156
rect 11539 36128 12434 36156
rect 11112 36116 11118 36128
rect 9214 36048 9220 36100
rect 9272 36088 9278 36100
rect 11539 36088 11567 36128
rect 9272 36060 11567 36088
rect 9272 36048 9278 36060
rect 11606 36048 11612 36100
rect 11664 36088 11670 36100
rect 12038 36091 12096 36097
rect 12038 36088 12050 36091
rect 11664 36060 12050 36088
rect 11664 36048 11670 36060
rect 12038 36057 12050 36060
rect 12084 36057 12096 36091
rect 12406 36088 12434 36128
rect 12986 36116 12992 36168
rect 13044 36156 13050 36168
rect 14108 36156 14136 36184
rect 13044 36128 14136 36156
rect 13044 36116 13050 36128
rect 14182 36116 14188 36168
rect 14240 36156 14246 36168
rect 15933 36159 15991 36165
rect 15933 36156 15945 36159
rect 14240 36128 15945 36156
rect 14240 36116 14246 36128
rect 15933 36125 15945 36128
rect 15979 36125 15991 36159
rect 16114 36156 16120 36168
rect 16075 36128 16120 36156
rect 15933 36119 15991 36125
rect 16114 36116 16120 36128
rect 16172 36116 16178 36168
rect 16206 36116 16212 36168
rect 16264 36156 16270 36168
rect 17779 36156 17807 36196
rect 18506 36184 18512 36196
rect 18564 36184 18570 36236
rect 19518 36224 19524 36236
rect 18892 36196 19196 36224
rect 18892 36190 18920 36196
rect 18800 36162 18920 36190
rect 18800 36156 18828 36162
rect 16264 36128 17807 36156
rect 17926 36128 18828 36156
rect 19168 36156 19196 36196
rect 19352 36196 19524 36224
rect 19352 36158 19380 36196
rect 19518 36184 19524 36196
rect 19576 36184 19582 36236
rect 19610 36184 19616 36236
rect 19668 36224 19674 36236
rect 23109 36227 23167 36233
rect 19668 36196 23060 36224
rect 19668 36184 19674 36196
rect 19260 36156 19380 36158
rect 19168 36130 19380 36156
rect 19429 36159 19487 36165
rect 19168 36128 19288 36130
rect 16264 36116 16270 36128
rect 12406 36060 13584 36088
rect 12038 36051 12096 36057
rect 9950 36020 9956 36032
rect 9140 35992 9956 36020
rect 9950 35980 9956 35992
rect 10008 35980 10014 36032
rect 10042 35980 10048 36032
rect 10100 36020 10106 36032
rect 10870 36020 10876 36032
rect 10100 35992 10876 36020
rect 10100 35980 10106 35992
rect 10870 35980 10876 35992
rect 10928 35980 10934 36032
rect 10962 35980 10968 36032
rect 11020 36020 11026 36032
rect 12158 36020 12164 36032
rect 11020 35992 12164 36020
rect 11020 35980 11026 35992
rect 12158 35980 12164 35992
rect 12216 35980 12222 36032
rect 12434 35980 12440 36032
rect 12492 36020 12498 36032
rect 13173 36023 13231 36029
rect 13173 36020 13185 36023
rect 12492 35992 13185 36020
rect 12492 35980 12498 35992
rect 13173 35989 13185 35992
rect 13219 35989 13231 36023
rect 13556 36020 13584 36060
rect 13630 36048 13636 36100
rect 13688 36088 13694 36100
rect 14338 36091 14396 36097
rect 14338 36088 14350 36091
rect 13688 36060 14350 36088
rect 13688 36048 13694 36060
rect 14338 36057 14350 36060
rect 14384 36057 14396 36091
rect 17006 36091 17064 36097
rect 17006 36088 17018 36091
rect 14338 36051 14396 36057
rect 14445 36060 17018 36088
rect 13814 36020 13820 36032
rect 13556 35992 13820 36020
rect 13173 35983 13231 35989
rect 13814 35980 13820 35992
rect 13872 35980 13878 36032
rect 13906 35980 13912 36032
rect 13964 36020 13970 36032
rect 14445 36020 14473 36060
rect 17006 36057 17018 36060
rect 17052 36057 17064 36091
rect 17006 36051 17064 36057
rect 17218 36048 17224 36100
rect 17276 36088 17282 36100
rect 17926 36088 17954 36128
rect 19429 36125 19441 36159
rect 19475 36125 19487 36159
rect 20346 36156 20352 36168
rect 20307 36128 20352 36156
rect 19429 36119 19487 36125
rect 17276 36060 17954 36088
rect 17276 36048 17282 36060
rect 18690 36048 18696 36100
rect 18748 36088 18754 36100
rect 19245 36091 19303 36097
rect 19245 36088 19257 36091
rect 18748 36060 19257 36088
rect 18748 36048 18754 36060
rect 19245 36057 19257 36060
rect 19291 36057 19303 36091
rect 19245 36051 19303 36057
rect 19334 36048 19340 36100
rect 19392 36088 19398 36100
rect 19444 36088 19472 36119
rect 20346 36116 20352 36128
rect 20404 36116 20410 36168
rect 21542 36156 21548 36168
rect 20456 36128 21548 36156
rect 19392 36060 19472 36088
rect 19613 36091 19671 36097
rect 19392 36048 19398 36060
rect 19613 36057 19625 36091
rect 19659 36088 19671 36091
rect 19886 36088 19892 36100
rect 19659 36060 19892 36088
rect 19659 36057 19671 36060
rect 19613 36051 19671 36057
rect 19886 36048 19892 36060
rect 19944 36048 19950 36100
rect 19978 36048 19984 36100
rect 20036 36088 20042 36100
rect 20456 36088 20484 36128
rect 21542 36116 21548 36128
rect 21600 36116 21606 36168
rect 21729 36159 21787 36165
rect 21729 36125 21741 36159
rect 21775 36125 21787 36159
rect 21729 36119 21787 36125
rect 21821 36159 21879 36165
rect 21821 36125 21833 36159
rect 21867 36156 21879 36159
rect 21910 36156 21916 36168
rect 21867 36128 21916 36156
rect 21867 36125 21879 36128
rect 21821 36119 21879 36125
rect 20036 36060 20484 36088
rect 20901 36091 20959 36097
rect 20036 36048 20042 36060
rect 20901 36057 20913 36091
rect 20947 36088 20959 36091
rect 21174 36088 21180 36100
rect 20947 36060 21180 36088
rect 20947 36057 20959 36060
rect 20901 36051 20959 36057
rect 21174 36048 21180 36060
rect 21232 36048 21238 36100
rect 21744 36088 21772 36119
rect 21910 36116 21916 36128
rect 21968 36116 21974 36168
rect 22097 36159 22155 36165
rect 22097 36125 22109 36159
rect 22143 36156 22155 36159
rect 22278 36156 22284 36168
rect 22143 36128 22284 36156
rect 22143 36125 22155 36128
rect 22097 36119 22155 36125
rect 22278 36116 22284 36128
rect 22336 36156 22342 36168
rect 22646 36156 22652 36168
rect 22336 36128 22652 36156
rect 22336 36116 22342 36128
rect 22646 36116 22652 36128
rect 22704 36116 22710 36168
rect 22741 36159 22799 36165
rect 22741 36125 22753 36159
rect 22787 36156 22799 36159
rect 22830 36156 22836 36168
rect 22787 36128 22836 36156
rect 22787 36125 22799 36128
rect 22741 36119 22799 36125
rect 22830 36116 22836 36128
rect 22888 36116 22894 36168
rect 22554 36088 22560 36100
rect 21744 36060 22560 36088
rect 22554 36048 22560 36060
rect 22612 36048 22618 36100
rect 23032 36088 23060 36196
rect 23109 36193 23121 36227
rect 23155 36224 23167 36227
rect 23382 36224 23388 36236
rect 23155 36196 23388 36224
rect 23155 36193 23167 36196
rect 23109 36187 23167 36193
rect 23382 36184 23388 36196
rect 23440 36184 23446 36236
rect 23750 36184 23756 36236
rect 23808 36224 23814 36236
rect 24872 36233 24900 36264
rect 25866 36252 25872 36264
rect 25924 36252 25930 36304
rect 24765 36227 24823 36233
rect 24765 36224 24777 36227
rect 23808 36196 24777 36224
rect 23808 36184 23814 36196
rect 24765 36193 24777 36196
rect 24811 36193 24823 36227
rect 24765 36187 24823 36193
rect 24857 36227 24915 36233
rect 24857 36193 24869 36227
rect 24903 36193 24915 36227
rect 24857 36187 24915 36193
rect 25222 36184 25228 36236
rect 25280 36224 25286 36236
rect 26513 36227 26571 36233
rect 26513 36224 26525 36227
rect 25280 36196 26525 36224
rect 25280 36184 25286 36196
rect 26513 36193 26525 36196
rect 26559 36193 26571 36227
rect 28166 36224 28172 36236
rect 28127 36196 28172 36224
rect 26513 36187 26571 36193
rect 28166 36184 28172 36196
rect 28224 36184 28230 36236
rect 23198 36156 23204 36168
rect 23159 36128 23204 36156
rect 23198 36116 23204 36128
rect 23256 36116 23262 36168
rect 25590 36116 25596 36168
rect 25648 36156 25654 36168
rect 25685 36159 25743 36165
rect 25685 36156 25697 36159
rect 25648 36128 25697 36156
rect 25648 36116 25654 36128
rect 25685 36125 25697 36128
rect 25731 36125 25743 36159
rect 26326 36156 26332 36168
rect 26287 36128 26332 36156
rect 25685 36119 25743 36125
rect 26326 36116 26332 36128
rect 26384 36116 26390 36168
rect 23032 36060 25452 36088
rect 13964 35992 14473 36020
rect 13964 35980 13970 35992
rect 14550 35980 14556 36032
rect 14608 36020 14614 36032
rect 16301 36023 16359 36029
rect 16301 36020 16313 36023
rect 14608 35992 16313 36020
rect 14608 35980 14614 35992
rect 16301 35989 16313 35992
rect 16347 35989 16359 36023
rect 16301 35983 16359 35989
rect 16666 35980 16672 36032
rect 16724 36020 16730 36032
rect 17770 36020 17776 36032
rect 16724 35992 17776 36020
rect 16724 35980 16730 35992
rect 17770 35980 17776 35992
rect 17828 35980 17834 36032
rect 18141 36023 18199 36029
rect 18141 35989 18153 36023
rect 18187 36020 18199 36023
rect 18322 36020 18328 36032
rect 18187 35992 18328 36020
rect 18187 35989 18199 35992
rect 18141 35983 18199 35989
rect 18322 35980 18328 35992
rect 18380 36020 18386 36032
rect 19521 36023 19579 36029
rect 19521 36020 19533 36023
rect 18380 35992 19533 36020
rect 18380 35980 18386 35992
rect 19521 35989 19533 35992
rect 19567 35989 19579 36023
rect 19521 35983 19579 35989
rect 19797 36023 19855 36029
rect 19797 35989 19809 36023
rect 19843 36020 19855 36023
rect 20806 36020 20812 36032
rect 19843 35992 20812 36020
rect 19843 35989 19855 35992
rect 19797 35983 19855 35989
rect 20806 35980 20812 35992
rect 20864 35980 20870 36032
rect 21545 36023 21603 36029
rect 21545 35989 21557 36023
rect 21591 36020 21603 36023
rect 22738 36020 22744 36032
rect 21591 35992 22744 36020
rect 21591 35989 21603 35992
rect 21545 35983 21603 35989
rect 22738 35980 22744 35992
rect 22796 35980 22802 36032
rect 23750 35980 23756 36032
rect 23808 36020 23814 36032
rect 24397 36023 24455 36029
rect 24397 36020 24409 36023
rect 23808 35992 24409 36020
rect 23808 35980 23814 35992
rect 24397 35989 24409 35992
rect 24443 36020 24455 36023
rect 25130 36020 25136 36032
rect 24443 35992 25136 36020
rect 24443 35989 24455 35992
rect 24397 35983 24455 35989
rect 25130 35980 25136 35992
rect 25188 35980 25194 36032
rect 25424 36020 25452 36060
rect 25498 36048 25504 36100
rect 25556 36088 25562 36100
rect 25556 36060 25601 36088
rect 25556 36048 25562 36060
rect 27246 36020 27252 36032
rect 25424 35992 27252 36020
rect 27246 35980 27252 35992
rect 27304 35980 27310 36032
rect 1104 35930 28888 35952
rect 1104 35878 10214 35930
rect 10266 35878 10278 35930
rect 10330 35878 10342 35930
rect 10394 35878 10406 35930
rect 10458 35878 10470 35930
rect 10522 35878 19478 35930
rect 19530 35878 19542 35930
rect 19594 35878 19606 35930
rect 19658 35878 19670 35930
rect 19722 35878 19734 35930
rect 19786 35878 28888 35930
rect 1104 35856 28888 35878
rect 3786 35776 3792 35828
rect 3844 35816 3850 35828
rect 3881 35819 3939 35825
rect 3881 35816 3893 35819
rect 3844 35788 3893 35816
rect 3844 35776 3850 35788
rect 3881 35785 3893 35788
rect 3927 35785 3939 35819
rect 8018 35816 8024 35828
rect 7979 35788 8024 35816
rect 3881 35779 3939 35785
rect 8018 35776 8024 35788
rect 8076 35776 8082 35828
rect 8665 35819 8723 35825
rect 8665 35785 8677 35819
rect 8711 35816 8723 35819
rect 9214 35816 9220 35828
rect 8711 35788 9220 35816
rect 8711 35785 8723 35788
rect 8665 35779 8723 35785
rect 9214 35776 9220 35788
rect 9272 35776 9278 35828
rect 9493 35819 9551 35825
rect 9493 35785 9505 35819
rect 9539 35816 9551 35819
rect 11974 35816 11980 35828
rect 9539 35788 11980 35816
rect 9539 35785 9551 35788
rect 9493 35779 9551 35785
rect 11974 35776 11980 35788
rect 12032 35776 12038 35828
rect 12069 35819 12127 35825
rect 12069 35785 12081 35819
rect 12115 35816 12127 35819
rect 12342 35816 12348 35828
rect 12115 35788 12348 35816
rect 12115 35785 12127 35788
rect 12069 35779 12127 35785
rect 12342 35776 12348 35788
rect 12400 35776 12406 35828
rect 12443 35788 13768 35816
rect 7374 35748 7380 35760
rect 3804 35720 7380 35748
rect 3804 35689 3832 35720
rect 7374 35708 7380 35720
rect 7432 35708 7438 35760
rect 7668 35720 10180 35748
rect 3789 35683 3847 35689
rect 3789 35649 3801 35683
rect 3835 35649 3847 35683
rect 3789 35643 3847 35649
rect 4430 35640 4436 35692
rect 4488 35680 4494 35692
rect 4617 35683 4675 35689
rect 4617 35680 4629 35683
rect 4488 35652 4629 35680
rect 4488 35640 4494 35652
rect 4617 35649 4629 35652
rect 4663 35649 4675 35683
rect 4617 35643 4675 35649
rect 6549 35683 6607 35689
rect 6549 35649 6561 35683
rect 6595 35680 6607 35683
rect 6638 35680 6644 35692
rect 6595 35652 6644 35680
rect 6595 35649 6607 35652
rect 6549 35643 6607 35649
rect 6638 35640 6644 35652
rect 6696 35640 6702 35692
rect 7558 35680 7564 35692
rect 7519 35652 7564 35680
rect 7558 35640 7564 35652
rect 7616 35640 7622 35692
rect 1489 35615 1547 35621
rect 1489 35581 1501 35615
rect 1535 35581 1547 35615
rect 1489 35575 1547 35581
rect 1673 35615 1731 35621
rect 1673 35581 1685 35615
rect 1719 35612 1731 35615
rect 1762 35612 1768 35624
rect 1719 35584 1768 35612
rect 1719 35581 1731 35584
rect 1673 35575 1731 35581
rect 1504 35544 1532 35575
rect 1762 35572 1768 35584
rect 1820 35572 1826 35624
rect 2866 35612 2872 35624
rect 2827 35584 2872 35612
rect 2866 35572 2872 35584
rect 2924 35572 2930 35624
rect 4522 35572 4528 35624
rect 4580 35612 4586 35624
rect 7668 35612 7696 35720
rect 8202 35680 8208 35692
rect 8163 35652 8208 35680
rect 8202 35640 8208 35652
rect 8260 35640 8266 35692
rect 8849 35683 8907 35689
rect 8849 35649 8861 35683
rect 8895 35649 8907 35683
rect 9306 35680 9312 35692
rect 9267 35652 9312 35680
rect 8849 35643 8907 35649
rect 4580 35584 7696 35612
rect 4580 35572 4586 35584
rect 5261 35547 5319 35553
rect 5261 35544 5273 35547
rect 1504 35516 5273 35544
rect 5261 35513 5273 35516
rect 5307 35513 5319 35547
rect 5261 35507 5319 35513
rect 5902 35504 5908 35556
rect 5960 35544 5966 35556
rect 8754 35544 8760 35556
rect 5960 35516 8760 35544
rect 5960 35504 5966 35516
rect 8754 35504 8760 35516
rect 8812 35504 8818 35556
rect 8864 35544 8892 35643
rect 9306 35640 9312 35652
rect 9364 35640 9370 35692
rect 9490 35680 9496 35692
rect 9451 35652 9496 35680
rect 9490 35640 9496 35652
rect 9548 35640 9554 35692
rect 9950 35682 9956 35692
rect 9692 35680 9956 35682
rect 9600 35654 9956 35680
rect 9600 35652 9720 35654
rect 9030 35572 9036 35624
rect 9088 35612 9094 35624
rect 9600 35612 9628 35652
rect 9950 35640 9956 35654
rect 10008 35680 10014 35692
rect 10008 35652 10101 35680
rect 10008 35640 10014 35652
rect 9088 35584 9628 35612
rect 9088 35572 9094 35584
rect 9858 35572 9864 35624
rect 9916 35612 9922 35624
rect 10045 35615 10103 35621
rect 10045 35612 10057 35615
rect 9916 35584 10057 35612
rect 9916 35572 9922 35584
rect 10045 35581 10057 35584
rect 10091 35581 10103 35615
rect 10152 35612 10180 35720
rect 10226 35708 10232 35760
rect 10284 35748 10290 35760
rect 10284 35720 10916 35748
rect 10284 35708 10290 35720
rect 10781 35683 10839 35689
rect 10781 35680 10793 35683
rect 10428 35652 10793 35680
rect 10428 35612 10456 35652
rect 10781 35649 10793 35652
rect 10827 35649 10839 35683
rect 10888 35680 10916 35720
rect 11054 35708 11060 35760
rect 11112 35748 11118 35760
rect 12443 35748 12471 35788
rect 11112 35720 12471 35748
rect 11112 35708 11118 35720
rect 12618 35708 12624 35760
rect 12676 35748 12682 35760
rect 12802 35748 12808 35760
rect 12676 35720 12808 35748
rect 12676 35708 12682 35720
rect 12802 35708 12808 35720
rect 12860 35708 12866 35760
rect 12897 35751 12955 35757
rect 12897 35717 12909 35751
rect 12943 35748 12955 35751
rect 12986 35748 12992 35760
rect 12943 35720 12992 35748
rect 12943 35717 12955 35720
rect 12897 35711 12955 35717
rect 12986 35708 12992 35720
rect 13044 35748 13050 35760
rect 13262 35748 13268 35760
rect 13044 35720 13268 35748
rect 13044 35708 13050 35720
rect 13262 35708 13268 35720
rect 13320 35708 13326 35760
rect 13630 35748 13636 35760
rect 13556 35720 13636 35748
rect 11422 35680 11428 35692
rect 10888 35678 11120 35680
rect 11164 35678 11428 35680
rect 10888 35652 11428 35678
rect 11092 35650 11192 35652
rect 10781 35643 10839 35649
rect 11422 35640 11428 35652
rect 11480 35640 11486 35692
rect 11977 35683 12035 35689
rect 11977 35649 11989 35683
rect 12023 35682 12035 35683
rect 12250 35682 12256 35692
rect 12023 35654 12256 35682
rect 12023 35649 12035 35654
rect 11977 35643 12035 35649
rect 12250 35640 12256 35654
rect 12308 35640 12314 35692
rect 12342 35640 12348 35692
rect 12400 35680 12406 35692
rect 12713 35683 12771 35689
rect 12713 35680 12725 35683
rect 12400 35652 12725 35680
rect 12400 35640 12406 35652
rect 12713 35649 12725 35652
rect 12759 35649 12771 35683
rect 12713 35643 12771 35649
rect 13078 35640 13084 35692
rect 13136 35680 13142 35692
rect 13357 35683 13415 35689
rect 13357 35680 13369 35683
rect 13136 35652 13369 35680
rect 13136 35640 13142 35652
rect 13357 35649 13369 35652
rect 13403 35678 13415 35683
rect 13446 35678 13452 35692
rect 13403 35650 13452 35678
rect 13403 35649 13415 35650
rect 13357 35643 13415 35649
rect 13446 35640 13452 35650
rect 13504 35640 13510 35692
rect 13556 35689 13584 35720
rect 13630 35708 13636 35720
rect 13688 35708 13694 35760
rect 13740 35748 13768 35788
rect 13906 35776 13912 35828
rect 13964 35816 13970 35828
rect 15194 35816 15200 35828
rect 13964 35788 15200 35816
rect 13964 35776 13970 35788
rect 15194 35776 15200 35788
rect 15252 35776 15258 35828
rect 16206 35816 16212 35828
rect 15304 35788 16212 35816
rect 15304 35748 15332 35788
rect 16206 35776 16212 35788
rect 16264 35776 16270 35828
rect 16758 35776 16764 35828
rect 16816 35816 16822 35828
rect 17681 35819 17739 35825
rect 17681 35816 17693 35819
rect 16816 35788 17693 35816
rect 16816 35776 16822 35788
rect 17681 35785 17693 35788
rect 17727 35785 17739 35819
rect 17681 35779 17739 35785
rect 18046 35776 18052 35828
rect 18104 35816 18110 35828
rect 18141 35819 18199 35825
rect 18141 35816 18153 35819
rect 18104 35788 18153 35816
rect 18104 35776 18110 35788
rect 18141 35785 18153 35788
rect 18187 35785 18199 35819
rect 18141 35779 18199 35785
rect 18322 35776 18328 35828
rect 18380 35816 18386 35828
rect 18380 35788 18552 35816
rect 18380 35776 18386 35788
rect 15746 35748 15752 35760
rect 13740 35720 15332 35748
rect 15488 35720 15752 35748
rect 13541 35683 13599 35689
rect 13541 35649 13553 35683
rect 13587 35649 13599 35683
rect 13541 35643 13599 35649
rect 13786 35652 14320 35680
rect 10152 35584 10456 35612
rect 10597 35615 10655 35621
rect 10045 35575 10103 35581
rect 10597 35581 10609 35615
rect 10643 35612 10655 35615
rect 10870 35612 10876 35624
rect 10643 35584 10876 35612
rect 10643 35581 10655 35584
rect 10597 35575 10655 35581
rect 10870 35572 10876 35584
rect 10928 35612 10934 35624
rect 11790 35612 11796 35624
rect 10928 35584 11796 35612
rect 10928 35572 10934 35584
rect 11790 35572 11796 35584
rect 11848 35612 11854 35624
rect 12066 35612 12072 35624
rect 11848 35584 12072 35612
rect 11848 35572 11854 35584
rect 12066 35572 12072 35584
rect 12124 35572 12130 35624
rect 12158 35572 12164 35624
rect 12216 35612 12222 35624
rect 13786 35612 13814 35652
rect 14182 35612 14188 35624
rect 12216 35584 13492 35612
rect 12216 35572 12222 35584
rect 13464 35556 13492 35584
rect 13542 35584 13814 35612
rect 14143 35584 14188 35612
rect 13262 35544 13268 35556
rect 8864 35516 13268 35544
rect 13262 35504 13268 35516
rect 13320 35504 13326 35556
rect 13446 35504 13452 35556
rect 13504 35504 13510 35556
rect 3418 35436 3424 35488
rect 3476 35476 3482 35488
rect 10226 35476 10232 35488
rect 3476 35448 10232 35476
rect 3476 35436 3482 35448
rect 10226 35436 10232 35448
rect 10284 35436 10290 35488
rect 10318 35436 10324 35488
rect 10376 35476 10382 35488
rect 10965 35479 11023 35485
rect 10965 35476 10977 35479
rect 10376 35448 10977 35476
rect 10376 35436 10382 35448
rect 10965 35445 10977 35448
rect 11011 35445 11023 35479
rect 10965 35439 11023 35445
rect 11514 35436 11520 35488
rect 11572 35476 11578 35488
rect 12710 35476 12716 35488
rect 11572 35448 12716 35476
rect 11572 35436 11578 35448
rect 12710 35436 12716 35448
rect 12768 35436 12774 35488
rect 12802 35436 12808 35488
rect 12860 35476 12866 35488
rect 13542 35476 13570 35584
rect 14182 35572 14188 35584
rect 14240 35572 14246 35624
rect 14292 35612 14320 35652
rect 14366 35640 14372 35692
rect 14424 35680 14430 35692
rect 15286 35680 15292 35692
rect 14424 35652 14469 35680
rect 15247 35652 15292 35680
rect 14424 35640 14430 35652
rect 15286 35640 15292 35652
rect 15344 35640 15350 35692
rect 15488 35689 15516 35720
rect 15746 35708 15752 35720
rect 15804 35708 15810 35760
rect 15930 35708 15936 35760
rect 15988 35748 15994 35760
rect 17218 35748 17224 35760
rect 15988 35720 17224 35748
rect 15988 35708 15994 35720
rect 17218 35708 17224 35720
rect 17276 35708 17282 35760
rect 18414 35748 18420 35760
rect 18375 35720 18420 35748
rect 18414 35708 18420 35720
rect 18472 35708 18478 35760
rect 18524 35757 18552 35788
rect 18874 35776 18880 35828
rect 18932 35776 18938 35828
rect 20806 35816 20812 35828
rect 19444 35788 20812 35816
rect 18690 35757 18696 35760
rect 18509 35751 18567 35757
rect 18509 35717 18521 35751
rect 18555 35717 18567 35751
rect 18509 35711 18567 35717
rect 18647 35751 18696 35757
rect 18647 35717 18659 35751
rect 18693 35717 18696 35751
rect 18647 35711 18696 35717
rect 18690 35708 18696 35711
rect 18748 35708 18754 35760
rect 15473 35683 15531 35689
rect 15473 35649 15485 35683
rect 15519 35649 15531 35683
rect 15473 35643 15531 35649
rect 15562 35640 15568 35692
rect 15620 35680 15626 35692
rect 16666 35680 16672 35692
rect 15620 35652 15665 35680
rect 16627 35652 16672 35680
rect 15620 35640 15626 35652
rect 16666 35640 16672 35652
rect 16724 35640 16730 35692
rect 17497 35683 17555 35689
rect 17236 35652 17448 35680
rect 17236 35612 17264 35652
rect 14292 35584 17264 35612
rect 17313 35615 17371 35621
rect 17313 35581 17325 35615
rect 17359 35612 17371 35615
rect 17420 35612 17448 35652
rect 17497 35649 17509 35683
rect 17543 35680 17555 35683
rect 17678 35680 17684 35692
rect 17543 35652 17684 35680
rect 17543 35649 17555 35652
rect 17497 35643 17555 35649
rect 17678 35640 17684 35652
rect 17736 35640 17742 35692
rect 18138 35640 18144 35692
rect 18196 35680 18202 35692
rect 18325 35683 18383 35689
rect 18325 35680 18337 35683
rect 18196 35652 18337 35680
rect 18196 35640 18202 35652
rect 18325 35649 18337 35652
rect 18371 35649 18383 35683
rect 18325 35643 18383 35649
rect 18785 35683 18843 35689
rect 18785 35649 18797 35683
rect 18831 35678 18843 35683
rect 18892 35678 18920 35776
rect 19444 35760 19472 35788
rect 20806 35776 20812 35788
rect 20864 35776 20870 35828
rect 21269 35819 21327 35825
rect 21269 35785 21281 35819
rect 21315 35785 21327 35819
rect 21269 35779 21327 35785
rect 19058 35708 19064 35760
rect 19116 35748 19122 35760
rect 19242 35748 19248 35760
rect 19116 35720 19248 35748
rect 19116 35708 19122 35720
rect 19242 35708 19248 35720
rect 19300 35708 19306 35760
rect 19426 35708 19432 35760
rect 19484 35708 19490 35760
rect 19610 35748 19616 35760
rect 19597 35708 19616 35748
rect 19668 35708 19674 35760
rect 19794 35708 19800 35760
rect 19852 35748 19858 35760
rect 20530 35748 20536 35760
rect 19852 35720 20536 35748
rect 19852 35708 19858 35720
rect 20530 35708 20536 35720
rect 20588 35708 20594 35760
rect 21284 35748 21312 35779
rect 22094 35776 22100 35828
rect 22152 35816 22158 35828
rect 22557 35819 22615 35825
rect 22557 35816 22569 35819
rect 22152 35788 22569 35816
rect 22152 35776 22158 35788
rect 22557 35785 22569 35788
rect 22603 35785 22615 35819
rect 22557 35779 22615 35785
rect 23842 35776 23848 35828
rect 23900 35816 23906 35828
rect 24489 35819 24547 35825
rect 23900 35788 24440 35816
rect 23900 35776 23906 35788
rect 21542 35748 21548 35760
rect 21284 35720 21548 35748
rect 21542 35708 21548 35720
rect 21600 35708 21606 35760
rect 24412 35748 24440 35788
rect 24489 35785 24501 35819
rect 24535 35816 24547 35819
rect 25222 35816 25228 35828
rect 24535 35788 25228 35816
rect 24535 35785 24547 35788
rect 24489 35779 24547 35785
rect 25222 35776 25228 35788
rect 25280 35776 25286 35828
rect 27709 35819 27767 35825
rect 27709 35816 27721 35819
rect 25323 35788 27721 35816
rect 24578 35748 24584 35760
rect 24412 35720 24584 35748
rect 19597 35702 19625 35708
rect 18831 35650 18920 35678
rect 18831 35649 18843 35650
rect 18785 35643 18843 35649
rect 19334 35640 19340 35692
rect 19392 35680 19398 35692
rect 19536 35682 19625 35702
rect 19505 35680 19625 35682
rect 20898 35680 20904 35692
rect 19392 35674 19625 35680
rect 19392 35654 19564 35674
rect 19392 35652 19533 35654
rect 20859 35652 20904 35680
rect 19392 35640 19398 35652
rect 20898 35640 20904 35652
rect 20956 35640 20962 35692
rect 21821 35683 21879 35689
rect 21821 35649 21833 35683
rect 21867 35649 21879 35683
rect 21821 35643 21879 35649
rect 17359 35581 17382 35612
rect 17420 35584 18276 35612
rect 17313 35575 17382 35581
rect 13630 35504 13636 35556
rect 13688 35544 13694 35556
rect 13688 35516 15516 35544
rect 13688 35504 13694 35516
rect 15488 35488 15516 35516
rect 15562 35504 15568 35556
rect 15620 35544 15626 35556
rect 17218 35544 17224 35556
rect 15620 35516 17224 35544
rect 15620 35504 15626 35516
rect 17218 35504 17224 35516
rect 17276 35504 17282 35556
rect 17354 35544 17382 35575
rect 18248 35544 18276 35584
rect 18800 35584 19268 35612
rect 18800 35544 18828 35584
rect 17354 35516 18000 35544
rect 18248 35516 18828 35544
rect 19240 35544 19268 35584
rect 19518 35572 19524 35624
rect 19576 35612 19582 35624
rect 19705 35615 19763 35621
rect 19705 35612 19717 35615
rect 19576 35584 19717 35612
rect 19576 35572 19582 35584
rect 19705 35581 19717 35584
rect 19751 35581 19763 35615
rect 20346 35612 20352 35624
rect 19705 35575 19763 35581
rect 20160 35584 20352 35612
rect 19978 35544 19984 35556
rect 19240 35516 19984 35544
rect 13722 35476 13728 35488
rect 12860 35448 13570 35476
rect 13683 35448 13728 35476
rect 12860 35436 12866 35448
rect 13722 35436 13728 35448
rect 13780 35436 13786 35488
rect 13998 35436 14004 35488
rect 14056 35476 14062 35488
rect 14553 35479 14611 35485
rect 14553 35476 14565 35479
rect 14056 35448 14565 35476
rect 14056 35436 14062 35448
rect 14553 35445 14565 35448
rect 14599 35445 14611 35479
rect 14553 35439 14611 35445
rect 14642 35436 14648 35488
rect 14700 35476 14706 35488
rect 15286 35476 15292 35488
rect 14700 35448 15292 35476
rect 14700 35436 14706 35448
rect 15286 35436 15292 35448
rect 15344 35436 15350 35488
rect 15470 35476 15476 35488
rect 15431 35448 15476 35476
rect 15470 35436 15476 35448
rect 15528 35436 15534 35488
rect 15749 35479 15807 35485
rect 15749 35445 15761 35479
rect 15795 35476 15807 35479
rect 16298 35476 16304 35488
rect 15795 35448 16304 35476
rect 15795 35445 15807 35448
rect 15749 35439 15807 35445
rect 16298 35436 16304 35448
rect 16356 35436 16362 35488
rect 16761 35479 16819 35485
rect 16761 35445 16773 35479
rect 16807 35476 16819 35479
rect 17862 35476 17868 35488
rect 16807 35448 17868 35476
rect 16807 35445 16819 35448
rect 16761 35439 16819 35445
rect 17862 35436 17868 35448
rect 17920 35436 17926 35488
rect 17972 35476 18000 35516
rect 19978 35504 19984 35516
rect 20036 35504 20042 35556
rect 20160 35553 20188 35584
rect 20346 35572 20352 35584
rect 20404 35572 20410 35624
rect 20625 35615 20683 35621
rect 20625 35581 20637 35615
rect 20671 35581 20683 35615
rect 20625 35575 20683 35581
rect 20073 35547 20131 35553
rect 20073 35513 20085 35547
rect 20119 35513 20131 35547
rect 20160 35547 20223 35553
rect 20160 35516 20177 35547
rect 20073 35507 20131 35513
rect 20165 35513 20177 35516
rect 20211 35513 20223 35547
rect 20165 35507 20223 35513
rect 19886 35476 19892 35488
rect 17972 35448 19892 35476
rect 19886 35436 19892 35448
rect 19944 35476 19950 35488
rect 20088 35476 20116 35507
rect 20640 35476 20668 35575
rect 20806 35572 20812 35624
rect 20864 35612 20870 35624
rect 20993 35615 21051 35621
rect 20993 35612 21005 35615
rect 20864 35584 21005 35612
rect 20864 35572 20870 35584
rect 20993 35581 21005 35584
rect 21039 35581 21051 35615
rect 20993 35575 21051 35581
rect 21008 35544 21036 35575
rect 21082 35572 21088 35624
rect 21140 35621 21146 35624
rect 21140 35615 21168 35621
rect 21156 35581 21168 35615
rect 21140 35575 21168 35581
rect 21140 35572 21146 35575
rect 21266 35544 21272 35556
rect 21008 35516 21272 35544
rect 21266 35504 21272 35516
rect 21324 35504 21330 35556
rect 21542 35476 21548 35488
rect 19944 35448 21548 35476
rect 19944 35436 19950 35448
rect 21542 35436 21548 35448
rect 21600 35436 21606 35488
rect 21836 35476 21864 35643
rect 21910 35640 21916 35692
rect 21968 35680 21974 35692
rect 22005 35683 22063 35689
rect 22005 35680 22017 35683
rect 21968 35652 22017 35680
rect 21968 35640 21974 35652
rect 22005 35649 22017 35652
rect 22051 35649 22063 35683
rect 22005 35643 22063 35649
rect 22278 35640 22284 35692
rect 22336 35680 22342 35692
rect 22373 35683 22431 35689
rect 22373 35680 22385 35683
rect 22336 35652 22385 35680
rect 22336 35640 22342 35652
rect 22373 35649 22385 35652
rect 22419 35649 22431 35683
rect 22373 35643 22431 35649
rect 22738 35640 22744 35692
rect 22796 35680 22802 35692
rect 23385 35683 23443 35689
rect 23385 35680 23397 35683
rect 22796 35652 23397 35680
rect 22796 35640 22802 35652
rect 23385 35649 23397 35652
rect 23431 35680 23443 35683
rect 23750 35680 23756 35692
rect 23431 35652 23756 35680
rect 23431 35649 23443 35652
rect 23385 35643 23443 35649
rect 23750 35640 23756 35652
rect 23808 35640 23814 35692
rect 24412 35689 24440 35720
rect 24578 35708 24584 35720
rect 24636 35708 24642 35760
rect 25323 35757 25351 35788
rect 27709 35785 27721 35788
rect 27755 35785 27767 35819
rect 27709 35779 27767 35785
rect 25308 35751 25366 35757
rect 25308 35717 25320 35751
rect 25354 35717 25366 35751
rect 27338 35748 27344 35760
rect 25308 35711 25366 35717
rect 27172 35720 27344 35748
rect 24397 35683 24455 35689
rect 24397 35649 24409 35683
rect 24443 35649 24455 35683
rect 24397 35643 24455 35649
rect 24486 35640 24492 35692
rect 24544 35680 24550 35692
rect 25041 35683 25099 35689
rect 25041 35680 25053 35683
rect 24544 35652 25053 35680
rect 24544 35640 24550 35652
rect 25041 35649 25053 35652
rect 25087 35649 25099 35683
rect 26970 35680 26976 35692
rect 26931 35652 26976 35680
rect 25041 35643 25099 35649
rect 26970 35640 26976 35652
rect 27028 35640 27034 35692
rect 27172 35689 27200 35720
rect 27338 35708 27344 35720
rect 27396 35708 27402 35760
rect 27985 35751 28043 35757
rect 27985 35748 27997 35751
rect 27448 35720 27997 35748
rect 27157 35683 27215 35689
rect 27157 35649 27169 35683
rect 27203 35649 27215 35683
rect 27157 35643 27215 35649
rect 27246 35640 27252 35692
rect 27304 35680 27310 35692
rect 27448 35680 27476 35720
rect 27985 35717 27997 35720
rect 28031 35717 28043 35751
rect 27985 35711 28043 35717
rect 27304 35652 27476 35680
rect 27525 35683 27583 35689
rect 27304 35640 27310 35652
rect 27525 35649 27537 35683
rect 27571 35649 27583 35683
rect 27525 35643 27583 35649
rect 22097 35615 22155 35621
rect 22097 35581 22109 35615
rect 22143 35581 22155 35615
rect 22097 35575 22155 35581
rect 22189 35615 22247 35621
rect 22189 35581 22201 35615
rect 22235 35612 22247 35615
rect 22554 35612 22560 35624
rect 22235 35584 22560 35612
rect 22235 35581 22247 35584
rect 22189 35575 22247 35581
rect 22002 35504 22008 35556
rect 22060 35544 22066 35556
rect 22112 35544 22140 35575
rect 22554 35572 22560 35584
rect 22612 35572 22618 35624
rect 23566 35572 23572 35624
rect 23624 35612 23630 35624
rect 23661 35615 23719 35621
rect 23661 35612 23673 35615
rect 23624 35584 23673 35612
rect 23624 35572 23630 35584
rect 23661 35581 23673 35584
rect 23707 35581 23719 35615
rect 23661 35575 23719 35581
rect 27341 35615 27399 35621
rect 27341 35581 27353 35615
rect 27387 35612 27399 35615
rect 27430 35612 27436 35624
rect 27387 35584 27436 35612
rect 27387 35581 27399 35584
rect 27341 35575 27399 35581
rect 27430 35572 27436 35584
rect 27488 35572 27494 35624
rect 22462 35544 22468 35556
rect 22060 35516 22468 35544
rect 22060 35504 22066 35516
rect 22462 35504 22468 35516
rect 22520 35504 22526 35556
rect 22572 35544 22600 35572
rect 23382 35544 23388 35556
rect 22572 35516 23388 35544
rect 23382 35504 23388 35516
rect 23440 35504 23446 35556
rect 24486 35504 24492 35556
rect 24544 35544 24550 35556
rect 24762 35544 24768 35556
rect 24544 35516 24768 35544
rect 24544 35504 24550 35516
rect 24762 35504 24768 35516
rect 24820 35504 24826 35556
rect 26418 35544 26424 35556
rect 26379 35516 26424 35544
rect 26418 35504 26424 35516
rect 26476 35544 26482 35556
rect 27540 35544 27568 35643
rect 26476 35516 27568 35544
rect 26476 35504 26482 35516
rect 22646 35476 22652 35488
rect 21836 35448 22652 35476
rect 22646 35436 22652 35448
rect 22704 35436 22710 35488
rect 22738 35436 22744 35488
rect 22796 35476 22802 35488
rect 23474 35476 23480 35488
rect 22796 35448 23480 35476
rect 22796 35436 22802 35448
rect 23474 35436 23480 35448
rect 23532 35436 23538 35488
rect 23750 35476 23756 35488
rect 23711 35448 23756 35476
rect 23750 35436 23756 35448
rect 23808 35436 23814 35488
rect 23842 35436 23848 35488
rect 23900 35476 23906 35488
rect 23937 35479 23995 35485
rect 23937 35476 23949 35479
rect 23900 35448 23949 35476
rect 23900 35436 23906 35448
rect 23937 35445 23949 35448
rect 23983 35445 23995 35479
rect 23937 35439 23995 35445
rect 25314 35436 25320 35488
rect 25372 35476 25378 35488
rect 27338 35476 27344 35488
rect 25372 35448 27344 35476
rect 25372 35436 25378 35448
rect 27338 35436 27344 35448
rect 27396 35436 27402 35488
rect 1104 35386 28888 35408
rect 1104 35334 5582 35386
rect 5634 35334 5646 35386
rect 5698 35334 5710 35386
rect 5762 35334 5774 35386
rect 5826 35334 5838 35386
rect 5890 35334 14846 35386
rect 14898 35334 14910 35386
rect 14962 35334 14974 35386
rect 15026 35334 15038 35386
rect 15090 35334 15102 35386
rect 15154 35334 24110 35386
rect 24162 35334 24174 35386
rect 24226 35334 24238 35386
rect 24290 35334 24302 35386
rect 24354 35334 24366 35386
rect 24418 35334 28888 35386
rect 1104 35312 28888 35334
rect 1762 35272 1768 35284
rect 1723 35244 1768 35272
rect 1762 35232 1768 35244
rect 1820 35232 1826 35284
rect 3878 35232 3884 35284
rect 3936 35272 3942 35284
rect 3973 35275 4031 35281
rect 3973 35272 3985 35275
rect 3936 35244 3985 35272
rect 3936 35232 3942 35244
rect 3973 35241 3985 35244
rect 4019 35241 4031 35275
rect 3973 35235 4031 35241
rect 4433 35275 4491 35281
rect 4433 35241 4445 35275
rect 4479 35272 4491 35275
rect 4522 35272 4528 35284
rect 4479 35244 4528 35272
rect 4479 35241 4491 35244
rect 4433 35235 4491 35241
rect 4522 35232 4528 35244
rect 4580 35232 4586 35284
rect 6270 35272 6276 35284
rect 6231 35244 6276 35272
rect 6270 35232 6276 35244
rect 6328 35232 6334 35284
rect 9214 35272 9220 35284
rect 9175 35244 9220 35272
rect 9214 35232 9220 35244
rect 9272 35232 9278 35284
rect 9582 35232 9588 35284
rect 9640 35272 9646 35284
rect 10962 35272 10968 35284
rect 9640 35244 10968 35272
rect 9640 35232 9646 35244
rect 10962 35232 10968 35244
rect 11020 35232 11026 35284
rect 11149 35275 11207 35281
rect 11149 35241 11161 35275
rect 11195 35272 11207 35275
rect 11606 35272 11612 35284
rect 11195 35244 11612 35272
rect 11195 35241 11207 35244
rect 11149 35235 11207 35241
rect 11606 35232 11612 35244
rect 11664 35232 11670 35284
rect 11885 35275 11943 35281
rect 11885 35241 11897 35275
rect 11931 35272 11943 35275
rect 11931 35244 18368 35272
rect 11931 35241 11943 35244
rect 11885 35235 11943 35241
rect 5629 35207 5687 35213
rect 5629 35173 5641 35207
rect 5675 35204 5687 35207
rect 5902 35204 5908 35216
rect 5675 35176 5908 35204
rect 5675 35173 5687 35176
rect 5629 35167 5687 35173
rect 5902 35164 5908 35176
rect 5960 35164 5966 35216
rect 8018 35164 8024 35216
rect 8076 35204 8082 35216
rect 10134 35204 10140 35216
rect 8076 35176 10140 35204
rect 8076 35164 8082 35176
rect 10134 35164 10140 35176
rect 10192 35164 10198 35216
rect 10410 35164 10416 35216
rect 10468 35204 10474 35216
rect 11238 35204 11244 35216
rect 10468 35176 11244 35204
rect 10468 35164 10474 35176
rect 11238 35164 11244 35176
rect 11296 35164 11302 35216
rect 11422 35164 11428 35216
rect 11480 35204 11486 35216
rect 12805 35207 12863 35213
rect 12805 35204 12817 35207
rect 11480 35176 12817 35204
rect 11480 35164 11486 35176
rect 12805 35173 12817 35176
rect 12851 35173 12863 35207
rect 12805 35167 12863 35173
rect 13446 35164 13452 35216
rect 13504 35204 13510 35216
rect 14921 35207 14979 35213
rect 13504 35176 14596 35204
rect 13504 35164 13510 35176
rect 7282 35136 7288 35148
rect 2424 35108 7288 35136
rect 2424 35080 2452 35108
rect 7282 35096 7288 35108
rect 7340 35096 7346 35148
rect 8938 35136 8944 35148
rect 7760 35108 8944 35136
rect 1673 35071 1731 35077
rect 1673 35037 1685 35071
rect 1719 35037 1731 35071
rect 2406 35068 2412 35080
rect 2367 35040 2412 35068
rect 1673 35031 1731 35037
rect 1688 35000 1716 35031
rect 2406 35028 2412 35040
rect 2464 35028 2470 35080
rect 3234 35068 3240 35080
rect 3195 35040 3240 35068
rect 3234 35028 3240 35040
rect 3292 35028 3298 35080
rect 4154 35028 4160 35080
rect 4212 35068 4218 35080
rect 4617 35071 4675 35077
rect 4617 35068 4629 35071
rect 4212 35040 4629 35068
rect 4212 35028 4218 35040
rect 4617 35037 4629 35040
rect 4663 35037 4675 35071
rect 4617 35031 4675 35037
rect 5353 35071 5411 35077
rect 5353 35037 5365 35071
rect 5399 35068 5411 35071
rect 5813 35071 5871 35077
rect 5813 35068 5825 35071
rect 5399 35040 5825 35068
rect 5399 35037 5411 35040
rect 5353 35031 5411 35037
rect 5813 35037 5825 35040
rect 5859 35068 5871 35071
rect 5994 35068 6000 35080
rect 5859 35040 6000 35068
rect 5859 35037 5871 35040
rect 5813 35031 5871 35037
rect 5994 35028 6000 35040
rect 6052 35028 6058 35080
rect 6457 35071 6515 35077
rect 6457 35037 6469 35071
rect 6503 35068 6515 35071
rect 6730 35068 6736 35080
rect 6503 35040 6736 35068
rect 6503 35037 6515 35040
rect 6457 35031 6515 35037
rect 6730 35028 6736 35040
rect 6788 35028 6794 35080
rect 7098 35068 7104 35080
rect 7059 35040 7104 35068
rect 7098 35028 7104 35040
rect 7156 35028 7162 35080
rect 7760 35077 7788 35108
rect 8938 35096 8944 35108
rect 8996 35096 9002 35148
rect 12158 35136 12164 35148
rect 9784 35108 12164 35136
rect 7745 35071 7803 35077
rect 7745 35037 7757 35071
rect 7791 35037 7803 35071
rect 8386 35068 8392 35080
rect 8347 35040 8392 35068
rect 7745 35031 7803 35037
rect 8386 35028 8392 35040
rect 8444 35028 8450 35080
rect 9122 35068 9128 35080
rect 9083 35040 9128 35068
rect 9122 35028 9128 35040
rect 9180 35028 9186 35080
rect 9214 35028 9220 35080
rect 9272 35068 9278 35080
rect 9309 35071 9367 35077
rect 9309 35068 9321 35071
rect 9272 35040 9321 35068
rect 9272 35028 9278 35040
rect 9309 35037 9321 35040
rect 9355 35068 9367 35071
rect 9398 35068 9404 35080
rect 9355 35040 9404 35068
rect 9355 35037 9367 35040
rect 9309 35031 9367 35037
rect 9398 35028 9404 35040
rect 9456 35028 9462 35080
rect 9784 35077 9812 35108
rect 12158 35096 12164 35108
rect 12216 35096 12222 35148
rect 12437 35139 12495 35145
rect 12437 35105 12449 35139
rect 12483 35136 12495 35139
rect 12483 35108 12940 35136
rect 12483 35105 12495 35108
rect 12437 35099 12495 35105
rect 12912 35080 12940 35108
rect 12986 35096 12992 35148
rect 13044 35136 13050 35148
rect 14461 35139 14519 35145
rect 14461 35136 14473 35139
rect 13044 35108 14473 35136
rect 13044 35096 13050 35108
rect 14461 35105 14473 35108
rect 14507 35105 14519 35139
rect 14568 35136 14596 35176
rect 14921 35173 14933 35207
rect 14967 35204 14979 35207
rect 15562 35204 15568 35216
rect 14967 35176 15568 35204
rect 14967 35173 14979 35176
rect 14921 35167 14979 35173
rect 15562 35164 15568 35176
rect 15620 35164 15626 35216
rect 16666 35164 16672 35216
rect 16724 35204 16730 35216
rect 17034 35204 17040 35216
rect 16724 35176 17040 35204
rect 16724 35164 16730 35176
rect 17034 35164 17040 35176
rect 17092 35164 17098 35216
rect 17497 35207 17555 35213
rect 17497 35173 17509 35207
rect 17543 35204 17555 35207
rect 17954 35204 17960 35216
rect 17543 35176 17960 35204
rect 17543 35173 17555 35176
rect 17497 35167 17555 35173
rect 17954 35164 17960 35176
rect 18012 35164 18018 35216
rect 18230 35204 18236 35216
rect 18191 35176 18236 35204
rect 18230 35164 18236 35176
rect 18288 35164 18294 35216
rect 18340 35148 18368 35244
rect 18414 35232 18420 35284
rect 18472 35272 18478 35284
rect 18472 35244 22048 35272
rect 18472 35232 18478 35244
rect 18598 35164 18604 35216
rect 18656 35204 18662 35216
rect 19150 35204 19156 35216
rect 18656 35176 19156 35204
rect 18656 35164 18662 35176
rect 19150 35164 19156 35176
rect 19208 35164 19214 35216
rect 19242 35164 19248 35216
rect 19300 35164 19306 35216
rect 19337 35207 19395 35213
rect 19337 35173 19349 35207
rect 19383 35204 19395 35207
rect 19794 35204 19800 35216
rect 19383 35176 19800 35204
rect 19383 35173 19395 35176
rect 19337 35167 19395 35173
rect 19794 35164 19800 35176
rect 19852 35164 19858 35216
rect 15654 35136 15660 35148
rect 14568 35108 15424 35136
rect 15615 35108 15660 35136
rect 14461 35099 14519 35105
rect 9769 35071 9827 35077
rect 9769 35037 9781 35071
rect 9815 35037 9827 35071
rect 9769 35031 9827 35037
rect 9953 35071 10011 35077
rect 9953 35037 9965 35071
rect 9999 35068 10011 35071
rect 10318 35068 10324 35080
rect 9999 35040 10324 35068
rect 9999 35037 10011 35040
rect 9953 35031 10011 35037
rect 10318 35028 10324 35040
rect 10376 35028 10382 35080
rect 10413 35071 10471 35077
rect 10413 35037 10425 35071
rect 10459 35068 10471 35071
rect 11065 35073 11123 35079
rect 10612 35068 10824 35070
rect 10459 35042 11008 35068
rect 10459 35040 10640 35042
rect 10796 35040 11008 35042
rect 10459 35037 10471 35040
rect 10413 35031 10471 35037
rect 2130 35000 2136 35012
rect 1688 34972 2136 35000
rect 2130 34960 2136 34972
rect 2188 35000 2194 35012
rect 3786 35000 3792 35012
rect 2188 34972 3792 35000
rect 2188 34960 2194 34972
rect 3786 34960 3792 34972
rect 3844 34960 3850 35012
rect 7834 34960 7840 35012
rect 7892 35000 7898 35012
rect 10226 35000 10232 35012
rect 7892 34972 10232 35000
rect 7892 34960 7898 34972
rect 10226 34960 10232 34972
rect 10284 34960 10290 35012
rect 10980 35000 11008 35040
rect 11065 35039 11077 35073
rect 11111 35068 11123 35073
rect 11238 35068 11244 35080
rect 11111 35040 11244 35068
rect 11111 35039 11123 35040
rect 11065 35033 11123 35039
rect 11238 35028 11244 35040
rect 11296 35028 11302 35080
rect 11330 35028 11336 35080
rect 11388 35068 11394 35080
rect 12250 35068 12256 35080
rect 11388 35040 12256 35068
rect 11388 35028 11394 35040
rect 12250 35028 12256 35040
rect 12308 35028 12314 35080
rect 12526 35028 12532 35080
rect 12584 35068 12590 35080
rect 12621 35071 12679 35077
rect 12621 35068 12633 35071
rect 12584 35040 12633 35068
rect 12584 35028 12590 35040
rect 12621 35037 12633 35040
rect 12667 35037 12679 35071
rect 12621 35031 12679 35037
rect 12894 35028 12900 35080
rect 12952 35028 12958 35080
rect 13357 35071 13415 35077
rect 13357 35037 13369 35071
rect 13403 35068 13415 35071
rect 13906 35068 13912 35080
rect 13403 35040 13912 35068
rect 13403 35037 13415 35040
rect 13357 35031 13415 35037
rect 13906 35028 13912 35040
rect 13964 35028 13970 35080
rect 14090 35068 14096 35080
rect 14051 35040 14096 35068
rect 14090 35028 14096 35040
rect 14148 35028 14154 35080
rect 14277 35071 14335 35077
rect 14277 35037 14289 35071
rect 14323 35068 14335 35071
rect 14366 35068 14372 35080
rect 14323 35040 14372 35068
rect 14323 35037 14335 35040
rect 14277 35031 14335 35037
rect 14366 35028 14372 35040
rect 14424 35028 14430 35080
rect 14918 35068 14924 35080
rect 14879 35040 14924 35068
rect 14918 35028 14924 35040
rect 14976 35028 14982 35080
rect 15102 35068 15108 35080
rect 15063 35040 15108 35068
rect 15102 35028 15108 35040
rect 15160 35028 15166 35080
rect 15194 35028 15200 35080
rect 15252 35068 15258 35080
rect 15396 35068 15424 35108
rect 15654 35096 15660 35108
rect 15712 35096 15718 35148
rect 17126 35096 17132 35148
rect 17184 35136 17190 35148
rect 17184 35108 17816 35136
rect 17184 35096 17190 35108
rect 17310 35068 17316 35080
rect 15252 35040 15297 35068
rect 15396 35040 17316 35068
rect 15252 35028 15258 35040
rect 17310 35028 17316 35040
rect 17368 35028 17374 35080
rect 17788 35077 17816 35108
rect 18322 35096 18328 35148
rect 18380 35136 18386 35148
rect 19260 35136 19288 35164
rect 22020 35152 22048 35244
rect 22370 35232 22376 35284
rect 22428 35272 22434 35284
rect 22554 35272 22560 35284
rect 22428 35244 22560 35272
rect 22428 35232 22434 35244
rect 22554 35232 22560 35244
rect 22612 35232 22618 35284
rect 22830 35232 22836 35284
rect 22888 35272 22894 35284
rect 25498 35272 25504 35284
rect 22888 35244 25504 35272
rect 22888 35232 22894 35244
rect 25498 35232 25504 35244
rect 25556 35232 25562 35284
rect 25774 35272 25780 35284
rect 25735 35244 25780 35272
rect 25774 35232 25780 35244
rect 25832 35232 25838 35284
rect 26970 35232 26976 35284
rect 27028 35272 27034 35284
rect 27798 35272 27804 35284
rect 27028 35244 27804 35272
rect 27028 35232 27034 35244
rect 27798 35232 27804 35244
rect 27856 35232 27862 35284
rect 27982 35204 27988 35216
rect 22103 35176 24716 35204
rect 22103 35152 22131 35176
rect 19889 35139 19947 35145
rect 19889 35136 19901 35139
rect 18380 35108 19901 35136
rect 18380 35096 18386 35108
rect 19889 35105 19901 35108
rect 19935 35105 19947 35139
rect 22020 35124 22131 35152
rect 22738 35136 22744 35148
rect 19889 35099 19947 35105
rect 22204 35108 22744 35136
rect 17773 35071 17831 35077
rect 17773 35037 17785 35071
rect 17819 35037 17831 35071
rect 17773 35031 17831 35037
rect 18138 35028 18144 35080
rect 18196 35068 18202 35080
rect 18417 35071 18475 35077
rect 18417 35068 18429 35071
rect 18196 35040 18429 35068
rect 18196 35028 18202 35040
rect 18417 35037 18429 35040
rect 18463 35037 18475 35071
rect 18417 35031 18475 35037
rect 18693 35071 18751 35077
rect 18693 35037 18705 35071
rect 18739 35068 18751 35071
rect 18739 35040 18920 35068
rect 18739 35037 18751 35040
rect 18693 35031 18751 35037
rect 11146 35000 11152 35012
rect 10980 34972 11152 35000
rect 11146 34960 11152 34972
rect 11204 34960 11210 35012
rect 11606 34960 11612 35012
rect 11664 35000 11670 35012
rect 11793 35003 11851 35009
rect 11793 35000 11805 35003
rect 11664 34972 11805 35000
rect 11664 34960 11670 34972
rect 11793 34969 11805 34972
rect 11839 34969 11851 35003
rect 11793 34963 11851 34969
rect 11974 34960 11980 35012
rect 12032 35000 12038 35012
rect 14734 35000 14740 35012
rect 12032 34972 14740 35000
rect 12032 34960 12038 34972
rect 14734 34960 14740 34972
rect 14792 34960 14798 35012
rect 15902 35003 15960 35009
rect 15902 35000 15914 35003
rect 14844 34972 15914 35000
rect 1854 34892 1860 34944
rect 1912 34932 1918 34944
rect 2501 34935 2559 34941
rect 2501 34932 2513 34935
rect 1912 34904 2513 34932
rect 1912 34892 1918 34904
rect 2501 34901 2513 34904
rect 2547 34901 2559 34935
rect 7558 34932 7564 34944
rect 7519 34904 7564 34932
rect 2501 34895 2559 34901
rect 7558 34892 7564 34904
rect 7616 34892 7622 34944
rect 8205 34935 8263 34941
rect 8205 34901 8217 34935
rect 8251 34932 8263 34935
rect 8478 34932 8484 34944
rect 8251 34904 8484 34932
rect 8251 34901 8263 34904
rect 8205 34895 8263 34901
rect 8478 34892 8484 34904
rect 8536 34892 8542 34944
rect 9858 34932 9864 34944
rect 9819 34904 9864 34932
rect 9858 34892 9864 34904
rect 9916 34892 9922 34944
rect 10134 34892 10140 34944
rect 10192 34932 10198 34944
rect 10505 34935 10563 34941
rect 10505 34932 10517 34935
rect 10192 34904 10517 34932
rect 10192 34892 10198 34904
rect 10505 34901 10517 34904
rect 10551 34901 10563 34935
rect 10505 34895 10563 34901
rect 10962 34892 10968 34944
rect 11020 34932 11026 34944
rect 12986 34932 12992 34944
rect 11020 34904 12992 34932
rect 11020 34892 11026 34904
rect 12986 34892 12992 34904
rect 13044 34892 13050 34944
rect 13078 34892 13084 34944
rect 13136 34932 13142 34944
rect 13449 34935 13507 34941
rect 13449 34932 13461 34935
rect 13136 34904 13461 34932
rect 13136 34892 13142 34904
rect 13449 34901 13461 34904
rect 13495 34932 13507 34935
rect 13722 34932 13728 34944
rect 13495 34904 13728 34932
rect 13495 34901 13507 34904
rect 13449 34895 13507 34901
rect 13722 34892 13728 34904
rect 13780 34892 13786 34944
rect 13814 34892 13820 34944
rect 13872 34932 13878 34944
rect 14844 34932 14872 34972
rect 15902 34969 15914 34972
rect 15948 34969 15960 35003
rect 15902 34963 15960 34969
rect 16390 34960 16396 35012
rect 16448 35000 16454 35012
rect 17497 35003 17555 35009
rect 17497 35000 17509 35003
rect 16448 34972 17509 35000
rect 16448 34960 16454 34972
rect 17497 34969 17509 34972
rect 17543 34969 17555 35003
rect 18892 35000 18920 35040
rect 18966 35028 18972 35080
rect 19024 35068 19030 35080
rect 19245 35071 19303 35077
rect 19245 35068 19257 35071
rect 19024 35040 19257 35068
rect 19024 35028 19030 35040
rect 19245 35037 19257 35040
rect 19291 35037 19303 35071
rect 21729 35071 21787 35077
rect 21729 35068 21741 35071
rect 19245 35031 19303 35037
rect 19352 35040 21741 35068
rect 19352 35000 19380 35040
rect 21729 35037 21741 35040
rect 21775 35037 21787 35071
rect 21729 35031 21787 35037
rect 21910 35028 21916 35080
rect 21968 35068 21974 35080
rect 22204 35077 22232 35108
rect 22738 35096 22744 35108
rect 22796 35096 22802 35148
rect 23017 35139 23075 35145
rect 23017 35105 23029 35139
rect 23063 35136 23075 35139
rect 24302 35136 24308 35148
rect 23063 35108 24308 35136
rect 23063 35105 23075 35108
rect 23017 35099 23075 35105
rect 24302 35096 24308 35108
rect 24360 35136 24366 35148
rect 24397 35139 24455 35145
rect 24397 35136 24409 35139
rect 24360 35108 24409 35136
rect 24360 35096 24366 35108
rect 24397 35105 24409 35108
rect 24443 35136 24455 35139
rect 24486 35136 24492 35148
rect 24443 35108 24492 35136
rect 24443 35105 24455 35108
rect 24397 35099 24455 35105
rect 24486 35096 24492 35108
rect 24544 35096 24550 35148
rect 24688 35145 24716 35176
rect 25700 35176 27988 35204
rect 24673 35139 24731 35145
rect 24673 35105 24685 35139
rect 24719 35136 24731 35139
rect 25498 35136 25504 35148
rect 24719 35108 25504 35136
rect 24719 35105 24731 35108
rect 24673 35099 24731 35105
rect 25498 35096 25504 35108
rect 25556 35096 25562 35148
rect 22078 35071 22136 35077
rect 21968 35040 22013 35068
rect 21968 35028 21974 35040
rect 22078 35037 22090 35071
rect 22124 35068 22136 35071
rect 22189 35071 22247 35077
rect 22124 35037 22140 35068
rect 22078 35031 22140 35037
rect 22189 35037 22201 35071
rect 22235 35037 22247 35071
rect 22189 35031 22247 35037
rect 22281 35071 22339 35077
rect 22281 35037 22293 35071
rect 22327 35068 22339 35071
rect 22646 35068 22652 35080
rect 22327 35040 22652 35068
rect 22327 35037 22339 35040
rect 22281 35031 22339 35037
rect 17497 34963 17555 34969
rect 17604 34972 18736 35000
rect 18892 34972 19380 35000
rect 13872 34904 14872 34932
rect 13872 34892 13878 34904
rect 14918 34892 14924 34944
rect 14976 34932 14982 34944
rect 17604 34932 17632 34972
rect 14976 34904 17632 34932
rect 17681 34935 17739 34941
rect 14976 34892 14982 34904
rect 17681 34901 17693 34935
rect 17727 34932 17739 34935
rect 17862 34932 17868 34944
rect 17727 34904 17868 34932
rect 17727 34901 17739 34904
rect 17681 34895 17739 34901
rect 17862 34892 17868 34904
rect 17920 34932 17926 34944
rect 18601 34935 18659 34941
rect 18601 34932 18613 34935
rect 17920 34904 18613 34932
rect 17920 34892 17926 34904
rect 18601 34901 18613 34904
rect 18647 34901 18659 34935
rect 18708 34932 18736 34972
rect 19610 34960 19616 35012
rect 19668 35000 19674 35012
rect 20134 35003 20192 35009
rect 20134 35000 20146 35003
rect 19668 34972 20146 35000
rect 19668 34960 19674 34972
rect 20134 34969 20146 34972
rect 20180 35000 20192 35003
rect 20990 35000 20996 35012
rect 20180 34972 20996 35000
rect 20180 34969 20192 34972
rect 20134 34963 20192 34969
rect 20990 34960 20996 34972
rect 21048 34960 21054 35012
rect 22112 35000 22140 35031
rect 22646 35028 22652 35040
rect 22704 35028 22710 35080
rect 22922 35068 22928 35080
rect 22883 35040 22928 35068
rect 22922 35028 22928 35040
rect 22980 35028 22986 35080
rect 24026 35028 24032 35080
rect 24084 35068 24090 35080
rect 24084 35040 24900 35068
rect 24084 35028 24090 35040
rect 22370 35000 22376 35012
rect 22112 34972 22376 35000
rect 22370 34960 22376 34972
rect 22428 34960 22434 35012
rect 24872 35000 24900 35040
rect 25406 35028 25412 35080
rect 25464 35068 25470 35080
rect 25700 35077 25728 35176
rect 27982 35164 27988 35176
rect 28040 35164 28046 35216
rect 26329 35139 26387 35145
rect 26329 35105 26341 35139
rect 26375 35136 26387 35139
rect 26602 35136 26608 35148
rect 26375 35108 26608 35136
rect 26375 35105 26387 35108
rect 26329 35099 26387 35105
rect 26602 35096 26608 35108
rect 26660 35096 26666 35148
rect 28166 35136 28172 35148
rect 28127 35108 28172 35136
rect 28166 35096 28172 35108
rect 28224 35096 28230 35148
rect 25685 35071 25743 35077
rect 25685 35068 25697 35071
rect 25464 35040 25697 35068
rect 25464 35028 25470 35040
rect 25685 35037 25697 35040
rect 25731 35037 25743 35071
rect 25685 35031 25743 35037
rect 26513 35003 26571 35009
rect 26513 35000 26525 35003
rect 24872 34972 26525 35000
rect 26513 34969 26525 34972
rect 26559 34969 26571 35003
rect 26513 34963 26571 34969
rect 20898 34932 20904 34944
rect 18708 34904 20904 34932
rect 18601 34895 18659 34901
rect 20898 34892 20904 34904
rect 20956 34892 20962 34944
rect 21266 34932 21272 34944
rect 21227 34904 21272 34932
rect 21266 34892 21272 34904
rect 21324 34892 21330 34944
rect 22830 34892 22836 34944
rect 22888 34932 22894 34944
rect 23293 34935 23351 34941
rect 23293 34932 23305 34935
rect 22888 34904 23305 34932
rect 22888 34892 22894 34904
rect 23293 34901 23305 34904
rect 23339 34901 23351 34935
rect 23293 34895 23351 34901
rect 23382 34892 23388 34944
rect 23440 34932 23446 34944
rect 24946 34932 24952 34944
rect 23440 34904 24952 34932
rect 23440 34892 23446 34904
rect 24946 34892 24952 34904
rect 25004 34892 25010 34944
rect 1104 34842 28888 34864
rect 1104 34790 10214 34842
rect 10266 34790 10278 34842
rect 10330 34790 10342 34842
rect 10394 34790 10406 34842
rect 10458 34790 10470 34842
rect 10522 34790 19478 34842
rect 19530 34790 19542 34842
rect 19594 34790 19606 34842
rect 19658 34790 19670 34842
rect 19722 34790 19734 34842
rect 19786 34790 28888 34842
rect 1104 34768 28888 34790
rect 3234 34728 3240 34740
rect 1688 34700 3240 34728
rect 1688 34601 1716 34700
rect 3234 34688 3240 34700
rect 3292 34688 3298 34740
rect 3786 34688 3792 34740
rect 3844 34728 3850 34740
rect 9030 34728 9036 34740
rect 3844 34700 9036 34728
rect 3844 34688 3850 34700
rect 9030 34688 9036 34700
rect 9088 34688 9094 34740
rect 9490 34728 9496 34740
rect 9451 34700 9496 34728
rect 9490 34688 9496 34700
rect 9548 34688 9554 34740
rect 10321 34731 10379 34737
rect 10321 34697 10333 34731
rect 10367 34728 10379 34731
rect 11238 34728 11244 34740
rect 10367 34700 11244 34728
rect 10367 34697 10379 34700
rect 10321 34691 10379 34697
rect 11238 34688 11244 34700
rect 11296 34688 11302 34740
rect 11974 34688 11980 34740
rect 12032 34728 12038 34740
rect 17037 34731 17095 34737
rect 17037 34728 17049 34731
rect 12032 34700 17049 34728
rect 12032 34688 12038 34700
rect 17037 34697 17049 34700
rect 17083 34697 17095 34731
rect 17037 34691 17095 34697
rect 17954 34688 17960 34740
rect 18012 34728 18018 34740
rect 20162 34728 20168 34740
rect 18012 34700 20168 34728
rect 18012 34688 18018 34700
rect 20162 34688 20168 34700
rect 20220 34688 20226 34740
rect 20272 34700 20576 34728
rect 1854 34660 1860 34672
rect 1815 34632 1860 34660
rect 1854 34620 1860 34632
rect 1912 34620 1918 34672
rect 8754 34660 8760 34672
rect 7760 34632 8760 34660
rect 7760 34601 7788 34632
rect 8754 34620 8760 34632
rect 8812 34620 8818 34672
rect 11762 34663 11820 34669
rect 11762 34660 11774 34663
rect 8864 34632 11774 34660
rect 1673 34595 1731 34601
rect 1673 34561 1685 34595
rect 1719 34561 1731 34595
rect 1673 34555 1731 34561
rect 7745 34595 7803 34601
rect 7745 34561 7757 34595
rect 7791 34561 7803 34595
rect 8386 34592 8392 34604
rect 8347 34564 8392 34592
rect 7745 34555 7803 34561
rect 8386 34552 8392 34564
rect 8444 34552 8450 34604
rect 2774 34484 2780 34536
rect 2832 34524 2838 34536
rect 2832 34496 2877 34524
rect 2832 34484 2838 34496
rect 7101 34459 7159 34465
rect 7101 34425 7113 34459
rect 7147 34456 7159 34459
rect 7466 34456 7472 34468
rect 7147 34428 7472 34456
rect 7147 34425 7159 34428
rect 7101 34419 7159 34425
rect 7466 34416 7472 34428
rect 7524 34416 7530 34468
rect 8864 34465 8892 34632
rect 11762 34629 11774 34632
rect 11808 34629 11820 34663
rect 11762 34623 11820 34629
rect 11882 34620 11888 34672
rect 11940 34660 11946 34672
rect 13078 34660 13084 34672
rect 11940 34632 13084 34660
rect 11940 34620 11946 34632
rect 13078 34620 13084 34632
rect 13136 34620 13142 34672
rect 13188 34632 16068 34660
rect 9033 34595 9091 34601
rect 9033 34561 9045 34595
rect 9079 34592 9091 34595
rect 9582 34592 9588 34604
rect 9079 34564 9588 34592
rect 9079 34561 9091 34564
rect 9033 34555 9091 34561
rect 9582 34552 9588 34564
rect 9640 34552 9646 34604
rect 9677 34595 9735 34601
rect 9677 34561 9689 34595
rect 9723 34561 9735 34595
rect 9677 34555 9735 34561
rect 9692 34524 9720 34555
rect 10042 34552 10048 34604
rect 10100 34592 10106 34604
rect 10137 34595 10195 34601
rect 10137 34592 10149 34595
rect 10100 34564 10149 34592
rect 10100 34552 10106 34564
rect 10137 34561 10149 34564
rect 10183 34561 10195 34595
rect 10137 34555 10195 34561
rect 10321 34595 10379 34601
rect 10321 34561 10333 34595
rect 10367 34592 10379 34595
rect 10781 34595 10839 34601
rect 10781 34592 10793 34595
rect 10367 34564 10793 34592
rect 10367 34561 10379 34564
rect 10321 34555 10379 34561
rect 10781 34561 10793 34564
rect 10827 34592 10839 34595
rect 11054 34592 11060 34604
rect 10827 34564 11060 34592
rect 10827 34561 10839 34564
rect 10781 34555 10839 34561
rect 11054 34552 11060 34564
rect 11112 34552 11118 34604
rect 13188 34592 13216 34632
rect 13613 34595 13671 34601
rect 13613 34592 13625 34595
rect 11440 34564 13216 34592
rect 13280 34564 13625 34592
rect 11440 34524 11468 34564
rect 9692 34496 11468 34524
rect 11517 34527 11575 34533
rect 11517 34493 11529 34527
rect 11563 34493 11575 34527
rect 11517 34487 11575 34493
rect 8849 34459 8907 34465
rect 8849 34425 8861 34459
rect 8895 34425 8907 34459
rect 8849 34419 8907 34425
rect 9508 34428 10827 34456
rect 1394 34348 1400 34400
rect 1452 34388 1458 34400
rect 4157 34391 4215 34397
rect 4157 34388 4169 34391
rect 1452 34360 4169 34388
rect 1452 34348 1458 34360
rect 4157 34357 4169 34360
rect 4203 34357 4215 34391
rect 7558 34388 7564 34400
rect 7519 34360 7564 34388
rect 4157 34351 4215 34357
rect 7558 34348 7564 34360
rect 7616 34348 7622 34400
rect 8205 34391 8263 34397
rect 8205 34357 8217 34391
rect 8251 34388 8263 34391
rect 9508 34388 9536 34428
rect 8251 34360 9536 34388
rect 8251 34357 8263 34360
rect 8205 34351 8263 34357
rect 9582 34348 9588 34400
rect 9640 34388 9646 34400
rect 10594 34388 10600 34400
rect 9640 34360 10600 34388
rect 9640 34348 9646 34360
rect 10594 34348 10600 34360
rect 10652 34348 10658 34400
rect 10799 34388 10827 34428
rect 10870 34416 10876 34468
rect 10928 34456 10934 34468
rect 10928 34428 10973 34456
rect 10928 34416 10934 34428
rect 11422 34416 11428 34468
rect 11480 34456 11486 34468
rect 11532 34456 11560 34487
rect 13280 34456 13308 34564
rect 13613 34561 13625 34564
rect 13659 34561 13671 34595
rect 13613 34555 13671 34561
rect 13906 34552 13912 34604
rect 13964 34592 13970 34604
rect 15930 34592 15936 34604
rect 13964 34564 15700 34592
rect 15891 34564 15936 34592
rect 13964 34552 13970 34564
rect 13354 34484 13360 34536
rect 13412 34524 13418 34536
rect 13412 34496 13457 34524
rect 13412 34484 13418 34496
rect 14550 34484 14556 34536
rect 14608 34524 14614 34536
rect 14608 34496 15608 34524
rect 14608 34484 14614 34496
rect 15470 34456 15476 34468
rect 11480 34428 11560 34456
rect 12443 34428 13308 34456
rect 14292 34428 15476 34456
rect 11480 34416 11486 34428
rect 12443 34388 12471 34428
rect 12894 34388 12900 34400
rect 10799 34360 12471 34388
rect 12855 34360 12900 34388
rect 12894 34348 12900 34360
rect 12952 34348 12958 34400
rect 12986 34348 12992 34400
rect 13044 34388 13050 34400
rect 14292 34388 14320 34428
rect 15470 34416 15476 34428
rect 15528 34416 15534 34468
rect 13044 34360 14320 34388
rect 13044 34348 13050 34360
rect 14642 34348 14648 34400
rect 14700 34388 14706 34400
rect 14737 34391 14795 34397
rect 14737 34388 14749 34391
rect 14700 34360 14749 34388
rect 14700 34348 14706 34360
rect 14737 34357 14749 34360
rect 14783 34357 14795 34391
rect 15580 34388 15608 34496
rect 15672 34456 15700 34564
rect 15930 34552 15936 34564
rect 15988 34552 15994 34604
rect 16040 34592 16068 34632
rect 16114 34620 16120 34672
rect 16172 34660 16178 34672
rect 18570 34663 18628 34669
rect 18570 34660 18582 34663
rect 16172 34632 18582 34660
rect 16172 34620 16178 34632
rect 18570 34629 18582 34632
rect 18616 34629 18628 34663
rect 18570 34623 18628 34629
rect 18690 34620 18696 34672
rect 18748 34660 18754 34672
rect 20272 34660 20300 34700
rect 18748 34632 20300 34660
rect 20442 34663 20500 34669
rect 18748 34620 18754 34632
rect 20442 34629 20454 34663
rect 20488 34629 20500 34663
rect 20548 34660 20576 34700
rect 20806 34688 20812 34740
rect 20864 34728 20870 34740
rect 22738 34728 22744 34740
rect 20864 34700 22744 34728
rect 20864 34688 20870 34700
rect 22738 34688 22744 34700
rect 22796 34688 22802 34740
rect 23658 34728 23664 34740
rect 22940 34700 23664 34728
rect 22940 34672 22968 34700
rect 23658 34688 23664 34700
rect 23716 34688 23722 34740
rect 24946 34728 24952 34740
rect 24907 34700 24952 34728
rect 24946 34688 24952 34700
rect 25004 34688 25010 34740
rect 25498 34688 25504 34740
rect 25556 34728 25562 34740
rect 26786 34728 26792 34740
rect 25556 34700 26792 34728
rect 25556 34688 25562 34700
rect 26786 34688 26792 34700
rect 26844 34728 26850 34740
rect 26844 34700 27108 34728
rect 26844 34688 26850 34700
rect 21913 34663 21971 34669
rect 21913 34660 21925 34663
rect 20548 34632 21925 34660
rect 20442 34623 20500 34629
rect 21913 34629 21925 34632
rect 21959 34629 21971 34663
rect 21913 34623 21971 34629
rect 22097 34663 22155 34669
rect 22097 34629 22109 34663
rect 22143 34660 22155 34663
rect 22922 34660 22928 34672
rect 22143 34632 22928 34660
rect 22143 34629 22155 34632
rect 22097 34623 22155 34629
rect 16482 34592 16488 34604
rect 16040 34564 16488 34592
rect 16482 34552 16488 34564
rect 16540 34552 16546 34604
rect 16666 34552 16672 34604
rect 16724 34592 16730 34604
rect 16853 34595 16911 34601
rect 16853 34592 16865 34595
rect 16724 34564 16769 34592
rect 16724 34552 16730 34564
rect 16837 34561 16865 34592
rect 16899 34561 16911 34595
rect 17494 34592 17500 34604
rect 17455 34564 17500 34592
rect 16837 34555 16911 34561
rect 15749 34527 15807 34533
rect 15749 34493 15761 34527
rect 15795 34524 15807 34527
rect 16574 34524 16580 34536
rect 15795 34496 16580 34524
rect 15795 34493 15807 34496
rect 15749 34487 15807 34493
rect 16574 34484 16580 34496
rect 16632 34484 16638 34536
rect 16117 34459 16175 34465
rect 16117 34456 16129 34459
rect 15672 34428 16129 34456
rect 16117 34425 16129 34428
rect 16163 34425 16175 34459
rect 16117 34419 16175 34425
rect 16206 34416 16212 34468
rect 16264 34456 16270 34468
rect 16837 34456 16865 34555
rect 17494 34552 17500 34564
rect 17552 34552 17558 34604
rect 17681 34595 17739 34601
rect 17681 34561 17693 34595
rect 17727 34592 17739 34595
rect 17770 34592 17776 34604
rect 17727 34564 17776 34592
rect 17727 34561 17739 34564
rect 17681 34555 17739 34561
rect 17770 34552 17776 34564
rect 17828 34552 17834 34604
rect 18322 34592 18328 34604
rect 18283 34564 18328 34592
rect 18322 34552 18328 34564
rect 18380 34552 18386 34604
rect 18432 34564 19564 34592
rect 18432 34524 18460 34564
rect 17972 34496 18460 34524
rect 19536 34524 19564 34564
rect 19978 34552 19984 34604
rect 20036 34592 20042 34604
rect 20349 34595 20407 34601
rect 20036 34590 20300 34592
rect 20349 34590 20361 34595
rect 20036 34564 20361 34590
rect 20036 34552 20042 34564
rect 20272 34562 20361 34564
rect 20349 34561 20361 34562
rect 20395 34561 20407 34595
rect 20349 34555 20407 34561
rect 20456 34536 20484 34623
rect 22922 34620 22928 34632
rect 22980 34620 22986 34672
rect 26973 34663 27031 34669
rect 26973 34660 26985 34663
rect 23032 34632 26985 34660
rect 20533 34595 20591 34601
rect 20533 34561 20545 34595
rect 20579 34561 20591 34595
rect 20533 34555 20591 34561
rect 20162 34524 20168 34536
rect 19536 34496 20168 34524
rect 16264 34428 16865 34456
rect 16264 34416 16270 34428
rect 17218 34416 17224 34468
rect 17276 34456 17282 34468
rect 17865 34459 17923 34465
rect 17865 34456 17877 34459
rect 17276 34428 17877 34456
rect 17276 34416 17282 34428
rect 17865 34425 17877 34428
rect 17911 34425 17923 34459
rect 17865 34419 17923 34425
rect 17972 34388 18000 34496
rect 20162 34484 20168 34496
rect 20220 34484 20226 34536
rect 20438 34484 20444 34536
rect 20496 34484 20502 34536
rect 19705 34459 19763 34465
rect 19705 34456 19717 34459
rect 19260 34428 19717 34456
rect 15580 34360 18000 34388
rect 14737 34351 14795 34357
rect 18506 34348 18512 34400
rect 18564 34388 18570 34400
rect 19260 34388 19288 34428
rect 19705 34425 19717 34428
rect 19751 34456 19763 34459
rect 20070 34456 20076 34468
rect 19751 34428 20076 34456
rect 19751 34425 19763 34428
rect 19705 34419 19763 34425
rect 20070 34416 20076 34428
rect 20128 34416 20134 34468
rect 20548 34400 20576 34555
rect 20622 34552 20628 34604
rect 20680 34601 20686 34604
rect 20680 34595 20709 34601
rect 20697 34561 20709 34595
rect 20680 34555 20709 34561
rect 20809 34595 20867 34601
rect 20809 34561 20821 34595
rect 20855 34592 20867 34595
rect 20990 34592 20996 34604
rect 20855 34564 20996 34592
rect 20855 34561 20867 34564
rect 20809 34555 20867 34561
rect 20680 34552 20686 34555
rect 20990 34552 20996 34564
rect 21048 34552 21054 34604
rect 21542 34552 21548 34604
rect 21600 34592 21606 34604
rect 21818 34592 21824 34604
rect 21600 34564 21824 34592
rect 21600 34552 21606 34564
rect 21818 34552 21824 34564
rect 21876 34552 21882 34604
rect 22002 34552 22008 34604
rect 22060 34592 22066 34604
rect 22830 34592 22836 34604
rect 22060 34564 22836 34592
rect 22060 34552 22066 34564
rect 22830 34552 22836 34564
rect 22888 34552 22894 34604
rect 23032 34601 23060 34632
rect 26973 34629 26985 34632
rect 27019 34629 27031 34663
rect 26973 34623 27031 34629
rect 23017 34595 23075 34601
rect 23017 34561 23029 34595
rect 23063 34561 23075 34595
rect 23017 34555 23075 34561
rect 23566 34552 23572 34604
rect 23624 34592 23630 34604
rect 23753 34595 23811 34601
rect 23753 34592 23765 34595
rect 23624 34564 23765 34592
rect 23624 34552 23630 34564
rect 23753 34561 23765 34564
rect 23799 34592 23811 34595
rect 23799 34564 24440 34592
rect 23799 34561 23811 34564
rect 23753 34555 23811 34561
rect 20898 34484 20904 34536
rect 20956 34524 20962 34536
rect 22741 34527 22799 34533
rect 22741 34524 22753 34527
rect 20956 34496 22753 34524
rect 20956 34484 20962 34496
rect 22741 34493 22753 34496
rect 22787 34493 22799 34527
rect 22741 34487 22799 34493
rect 22925 34527 22983 34533
rect 22925 34493 22937 34527
rect 22971 34524 22983 34527
rect 23106 34524 23112 34536
rect 22971 34496 23112 34524
rect 22971 34493 22983 34496
rect 22925 34487 22983 34493
rect 20990 34416 20996 34468
rect 21048 34456 21054 34468
rect 21174 34456 21180 34468
rect 21048 34428 21180 34456
rect 21048 34416 21054 34428
rect 21174 34416 21180 34428
rect 21232 34416 21238 34468
rect 22756 34456 22784 34487
rect 23106 34484 23112 34496
rect 23164 34484 23170 34536
rect 23845 34527 23903 34533
rect 23845 34493 23857 34527
rect 23891 34524 23903 34527
rect 24302 34524 24308 34536
rect 23891 34496 24308 34524
rect 23891 34493 23903 34496
rect 23845 34487 23903 34493
rect 24302 34484 24308 34496
rect 24360 34484 24366 34536
rect 24412 34524 24440 34564
rect 24486 34552 24492 34604
rect 24544 34592 24550 34604
rect 24581 34595 24639 34601
rect 24581 34592 24593 34595
rect 24544 34564 24593 34592
rect 24544 34552 24550 34564
rect 24581 34561 24593 34564
rect 24627 34561 24639 34595
rect 24762 34592 24768 34604
rect 24723 34564 24768 34592
rect 24581 34555 24639 34561
rect 24762 34552 24768 34564
rect 24820 34552 24826 34604
rect 25590 34592 25596 34604
rect 25551 34564 25596 34592
rect 25590 34552 25596 34564
rect 25648 34552 25654 34604
rect 27080 34592 27108 34700
rect 27157 34595 27215 34601
rect 27157 34592 27169 34595
rect 27080 34564 27169 34592
rect 27157 34561 27169 34564
rect 27203 34561 27215 34595
rect 27893 34595 27951 34601
rect 27893 34592 27905 34595
rect 27157 34555 27215 34561
rect 27264 34564 27905 34592
rect 24854 34524 24860 34536
rect 24412 34496 24860 34524
rect 24854 34484 24860 34496
rect 24912 34484 24918 34536
rect 25498 34524 25504 34536
rect 25459 34496 25504 34524
rect 25498 34484 25504 34496
rect 25556 34484 25562 34536
rect 27264 34524 27292 34564
rect 27893 34561 27905 34564
rect 27939 34561 27951 34595
rect 28074 34592 28080 34604
rect 28035 34564 28080 34592
rect 27893 34555 27951 34561
rect 28074 34552 28080 34564
rect 28132 34552 28138 34604
rect 28169 34595 28227 34601
rect 28169 34561 28181 34595
rect 28215 34592 28227 34595
rect 28258 34592 28264 34604
rect 28215 34564 28264 34592
rect 28215 34561 28227 34564
rect 28169 34555 28227 34561
rect 28258 34552 28264 34564
rect 28316 34552 28322 34604
rect 25608 34496 27292 34524
rect 27433 34527 27491 34533
rect 24121 34459 24179 34465
rect 24121 34456 24133 34459
rect 22756 34428 24133 34456
rect 24121 34425 24133 34428
rect 24167 34425 24179 34459
rect 24121 34419 24179 34425
rect 18564 34360 19288 34388
rect 18564 34348 18570 34360
rect 19886 34348 19892 34400
rect 19944 34388 19950 34400
rect 20165 34391 20223 34397
rect 20165 34388 20177 34391
rect 19944 34360 20177 34388
rect 19944 34348 19950 34360
rect 20165 34357 20177 34360
rect 20211 34357 20223 34391
rect 20165 34351 20223 34357
rect 20530 34348 20536 34400
rect 20588 34348 20594 34400
rect 20622 34348 20628 34400
rect 20680 34388 20686 34400
rect 22002 34388 22008 34400
rect 20680 34360 22008 34388
rect 20680 34348 20686 34360
rect 22002 34348 22008 34360
rect 22060 34348 22066 34400
rect 22554 34388 22560 34400
rect 22467 34360 22560 34388
rect 22554 34348 22560 34360
rect 22612 34388 22618 34400
rect 23106 34388 23112 34400
rect 22612 34360 23112 34388
rect 22612 34348 22618 34360
rect 23106 34348 23112 34360
rect 23164 34348 23170 34400
rect 24136 34388 24164 34419
rect 24210 34416 24216 34468
rect 24268 34456 24274 34468
rect 25608 34456 25636 34496
rect 27433 34493 27445 34527
rect 27479 34493 27491 34527
rect 28442 34524 28448 34536
rect 27433 34487 27491 34493
rect 27908 34496 28448 34524
rect 24268 34428 25636 34456
rect 25961 34459 26019 34465
rect 24268 34416 24274 34428
rect 25961 34425 25973 34459
rect 26007 34456 26019 34459
rect 26234 34456 26240 34468
rect 26007 34428 26240 34456
rect 26007 34425 26019 34428
rect 25961 34419 26019 34425
rect 26234 34416 26240 34428
rect 26292 34456 26298 34468
rect 27154 34456 27160 34468
rect 26292 34428 27160 34456
rect 26292 34416 26298 34428
rect 27154 34416 27160 34428
rect 27212 34416 27218 34468
rect 27338 34456 27344 34468
rect 27299 34428 27344 34456
rect 27338 34416 27344 34428
rect 27396 34416 27402 34468
rect 24486 34388 24492 34400
rect 24136 34360 24492 34388
rect 24486 34348 24492 34360
rect 24544 34348 24550 34400
rect 24854 34348 24860 34400
rect 24912 34388 24918 34400
rect 25130 34388 25136 34400
rect 24912 34360 25136 34388
rect 24912 34348 24918 34360
rect 25130 34348 25136 34360
rect 25188 34388 25194 34400
rect 27448 34388 27476 34487
rect 27908 34465 27936 34496
rect 28442 34484 28448 34496
rect 28500 34484 28506 34536
rect 27893 34459 27951 34465
rect 27893 34425 27905 34459
rect 27939 34425 27951 34459
rect 27893 34419 27951 34425
rect 25188 34360 27476 34388
rect 25188 34348 25194 34360
rect 1104 34298 28888 34320
rect 1104 34246 5582 34298
rect 5634 34246 5646 34298
rect 5698 34246 5710 34298
rect 5762 34246 5774 34298
rect 5826 34246 5838 34298
rect 5890 34246 14846 34298
rect 14898 34246 14910 34298
rect 14962 34246 14974 34298
rect 15026 34246 15038 34298
rect 15090 34246 15102 34298
rect 15154 34246 24110 34298
rect 24162 34246 24174 34298
rect 24226 34246 24238 34298
rect 24290 34246 24302 34298
rect 24354 34246 24366 34298
rect 24418 34246 28888 34298
rect 1104 34224 28888 34246
rect 7742 34144 7748 34196
rect 7800 34184 7806 34196
rect 11517 34187 11575 34193
rect 11517 34184 11529 34187
rect 7800 34156 11529 34184
rect 7800 34144 7806 34156
rect 11517 34153 11529 34156
rect 11563 34153 11575 34187
rect 12345 34187 12403 34193
rect 12345 34184 12357 34187
rect 11517 34147 11575 34153
rect 11624 34156 12357 34184
rect 6917 34119 6975 34125
rect 6917 34085 6929 34119
rect 6963 34085 6975 34119
rect 6917 34079 6975 34085
rect 8205 34119 8263 34125
rect 8205 34085 8217 34119
rect 8251 34116 8263 34119
rect 8846 34116 8852 34128
rect 8251 34088 8852 34116
rect 8251 34085 8263 34088
rect 8205 34079 8263 34085
rect 1394 34048 1400 34060
rect 1355 34020 1400 34048
rect 1394 34008 1400 34020
rect 1452 34008 1458 34060
rect 2774 34008 2780 34060
rect 2832 34048 2838 34060
rect 6932 34048 6960 34079
rect 8846 34076 8852 34088
rect 8904 34076 8910 34128
rect 9398 34076 9404 34128
rect 9456 34116 9462 34128
rect 9456 34088 10180 34116
rect 9456 34076 9462 34088
rect 9950 34048 9956 34060
rect 2832 34020 2877 34048
rect 6932 34020 9956 34048
rect 2832 34008 2838 34020
rect 9950 34008 9956 34020
rect 10008 34008 10014 34060
rect 7101 33983 7159 33989
rect 7101 33949 7113 33983
rect 7147 33980 7159 33983
rect 7650 33980 7656 33992
rect 7147 33952 7656 33980
rect 7147 33949 7159 33952
rect 7101 33943 7159 33949
rect 7650 33940 7656 33952
rect 7708 33940 7714 33992
rect 7742 33940 7748 33992
rect 7800 33980 7806 33992
rect 8389 33983 8447 33989
rect 7800 33952 7845 33980
rect 7800 33940 7806 33952
rect 8389 33949 8401 33983
rect 8435 33980 8447 33983
rect 8478 33980 8484 33992
rect 8435 33952 8484 33980
rect 8435 33949 8447 33952
rect 8389 33943 8447 33949
rect 8478 33940 8484 33952
rect 8536 33940 8542 33992
rect 9217 33983 9275 33989
rect 9217 33949 9229 33983
rect 9263 33980 9275 33983
rect 9306 33980 9312 33992
rect 9263 33952 9312 33980
rect 9263 33949 9275 33952
rect 9217 33943 9275 33949
rect 9306 33940 9312 33952
rect 9364 33940 9370 33992
rect 9398 33940 9404 33992
rect 9456 33980 9462 33992
rect 9665 33983 9723 33989
rect 9665 33980 9677 33983
rect 9456 33952 9677 33980
rect 9456 33940 9462 33952
rect 9665 33949 9677 33952
rect 9711 33949 9723 33983
rect 9665 33943 9723 33949
rect 9861 33983 9919 33989
rect 9861 33949 9873 33983
rect 9907 33949 9919 33983
rect 9861 33943 9919 33949
rect 1581 33915 1639 33921
rect 1581 33881 1593 33915
rect 1627 33912 1639 33915
rect 2222 33912 2228 33924
rect 1627 33884 2228 33912
rect 1627 33881 1639 33884
rect 1581 33875 1639 33881
rect 2222 33872 2228 33884
rect 2280 33872 2286 33924
rect 9490 33872 9496 33924
rect 9548 33912 9554 33924
rect 9769 33915 9827 33921
rect 9769 33912 9781 33915
rect 9548 33884 9781 33912
rect 9548 33872 9554 33884
rect 9769 33881 9781 33884
rect 9815 33881 9827 33915
rect 9876 33912 9904 33943
rect 10042 33940 10048 33992
rect 10100 33940 10106 33992
rect 10152 33980 10180 34088
rect 10226 34076 10232 34128
rect 10284 34116 10290 34128
rect 10962 34116 10968 34128
rect 10284 34088 10968 34116
rect 10284 34076 10290 34088
rect 10962 34076 10968 34088
rect 11020 34076 11026 34128
rect 11624 34116 11652 34156
rect 12345 34153 12357 34156
rect 12391 34153 12403 34187
rect 12345 34147 12403 34153
rect 12710 34144 12716 34196
rect 12768 34184 12774 34196
rect 12768 34156 12848 34184
rect 12768 34144 12774 34156
rect 11064 34088 11652 34116
rect 10336 34020 10732 34048
rect 10226 33980 10232 33992
rect 10152 33952 10232 33980
rect 10226 33940 10232 33952
rect 10284 33940 10290 33992
rect 10336 33989 10364 34020
rect 10321 33983 10379 33989
rect 10321 33949 10333 33983
rect 10367 33949 10379 33983
rect 10321 33943 10379 33949
rect 10410 33940 10416 33992
rect 10468 33980 10474 33992
rect 10505 33983 10563 33989
rect 10505 33980 10517 33983
rect 10468 33952 10517 33980
rect 10468 33940 10474 33952
rect 10505 33949 10517 33952
rect 10551 33949 10563 33983
rect 10704 33980 10732 34020
rect 10778 34008 10784 34060
rect 10836 34048 10842 34060
rect 11064 34048 11092 34088
rect 11698 34076 11704 34128
rect 11756 34116 11762 34128
rect 11882 34116 11888 34128
rect 11756 34088 11888 34116
rect 11756 34076 11762 34088
rect 11882 34076 11888 34088
rect 11940 34076 11946 34128
rect 12820 34116 12848 34156
rect 12894 34144 12900 34196
rect 12952 34184 12958 34196
rect 13357 34187 13415 34193
rect 13357 34184 13369 34187
rect 12952 34156 13369 34184
rect 12952 34144 12958 34156
rect 13357 34153 13369 34156
rect 13403 34184 13415 34187
rect 14182 34184 14188 34196
rect 13403 34156 14188 34184
rect 13403 34153 13415 34156
rect 13357 34147 13415 34153
rect 14182 34144 14188 34156
rect 14240 34144 14246 34196
rect 14458 34144 14464 34196
rect 14516 34184 14522 34196
rect 15930 34184 15936 34196
rect 14516 34156 15936 34184
rect 14516 34144 14522 34156
rect 15930 34144 15936 34156
rect 15988 34144 15994 34196
rect 16482 34144 16488 34196
rect 16540 34144 16546 34196
rect 16574 34144 16580 34196
rect 16632 34184 16638 34196
rect 16945 34187 17003 34193
rect 16945 34184 16957 34187
rect 16632 34156 16957 34184
rect 16632 34144 16638 34156
rect 16945 34153 16957 34156
rect 16991 34153 17003 34187
rect 16945 34147 17003 34153
rect 17494 34144 17500 34196
rect 17552 34184 17558 34196
rect 18598 34184 18604 34196
rect 17552 34156 18604 34184
rect 17552 34144 17558 34156
rect 18598 34144 18604 34156
rect 18656 34144 18662 34196
rect 18693 34187 18751 34193
rect 18693 34153 18705 34187
rect 18739 34184 18751 34187
rect 19978 34184 19984 34196
rect 18739 34156 19984 34184
rect 18739 34153 18751 34156
rect 18693 34147 18751 34153
rect 19978 34144 19984 34156
rect 20036 34144 20042 34196
rect 20162 34144 20168 34196
rect 20220 34184 20226 34196
rect 20622 34184 20628 34196
rect 20220 34156 20628 34184
rect 20220 34144 20226 34156
rect 20622 34144 20628 34156
rect 20680 34144 20686 34196
rect 21542 34144 21548 34196
rect 21600 34184 21606 34196
rect 21910 34184 21916 34196
rect 21600 34156 21916 34184
rect 21600 34144 21606 34156
rect 21910 34144 21916 34156
rect 21968 34144 21974 34196
rect 23658 34144 23664 34196
rect 23716 34184 23722 34196
rect 24581 34187 24639 34193
rect 24581 34184 24593 34187
rect 23716 34156 24593 34184
rect 23716 34144 23722 34156
rect 24581 34153 24593 34156
rect 24627 34153 24639 34187
rect 24581 34147 24639 34153
rect 13541 34119 13599 34125
rect 13541 34116 13553 34119
rect 11992 34088 12664 34116
rect 12820 34088 13553 34116
rect 11992 34048 12020 34088
rect 10836 34020 11092 34048
rect 11624 34020 12020 34048
rect 10836 34008 10842 34020
rect 11624 33996 11652 34020
rect 12066 34008 12072 34060
rect 12124 34048 12130 34060
rect 12434 34048 12440 34060
rect 12124 34020 12440 34048
rect 12124 34008 12130 34020
rect 12434 34008 12440 34020
rect 12492 34008 12498 34060
rect 12636 34048 12664 34088
rect 13541 34085 13553 34088
rect 13587 34085 13599 34119
rect 13541 34079 13599 34085
rect 13906 34076 13912 34128
rect 13964 34116 13970 34128
rect 14090 34116 14096 34128
rect 13964 34088 14096 34116
rect 13964 34076 13970 34088
rect 14090 34076 14096 34088
rect 14148 34076 14154 34128
rect 16500 34116 16528 34144
rect 17218 34116 17224 34128
rect 16500 34088 17224 34116
rect 17218 34076 17224 34088
rect 17276 34076 17282 34128
rect 18046 34076 18052 34128
rect 18104 34116 18110 34128
rect 18141 34119 18199 34125
rect 18141 34116 18153 34119
rect 18104 34088 18153 34116
rect 18104 34076 18110 34088
rect 18141 34085 18153 34088
rect 18187 34085 18199 34119
rect 18141 34079 18199 34085
rect 21082 34076 21088 34128
rect 21140 34116 21146 34128
rect 22281 34119 22339 34125
rect 22281 34116 22293 34119
rect 21140 34088 22293 34116
rect 21140 34076 21146 34088
rect 22281 34085 22293 34088
rect 22327 34085 22339 34119
rect 22462 34116 22468 34128
rect 22423 34088 22468 34116
rect 22281 34079 22339 34085
rect 22462 34076 22468 34088
rect 22520 34076 22526 34128
rect 23290 34116 23296 34128
rect 22572 34088 23296 34116
rect 12986 34048 12992 34060
rect 12636 34020 12992 34048
rect 12986 34008 12992 34020
rect 13044 34008 13050 34060
rect 13082 34020 15424 34048
rect 11146 33980 11152 33992
rect 10704 33952 11152 33980
rect 10505 33943 10563 33949
rect 11146 33940 11152 33952
rect 11204 33940 11210 33992
rect 11241 33983 11299 33989
rect 11241 33949 11253 33983
rect 11287 33949 11299 33983
rect 11241 33943 11299 33949
rect 11333 33983 11391 33989
rect 11333 33949 11345 33983
rect 11379 33980 11391 33983
rect 11440 33980 11652 33996
rect 11974 33980 11980 33992
rect 11379 33968 11652 33980
rect 11379 33952 11468 33968
rect 11935 33952 11980 33980
rect 11379 33949 11391 33952
rect 11333 33943 11391 33949
rect 9950 33912 9956 33924
rect 9876 33884 9956 33912
rect 9769 33875 9827 33881
rect 9950 33872 9956 33884
rect 10008 33872 10014 33924
rect 10060 33912 10088 33940
rect 10689 33915 10747 33921
rect 10689 33912 10701 33915
rect 10060 33884 10701 33912
rect 10689 33881 10701 33884
rect 10735 33881 10747 33915
rect 11256 33912 11284 33943
rect 11974 33940 11980 33952
rect 12032 33940 12038 33992
rect 12158 33940 12164 33992
rect 12216 33980 12222 33992
rect 12526 33980 12532 33992
rect 12216 33952 12532 33980
rect 12216 33940 12222 33952
rect 12526 33940 12532 33952
rect 12584 33940 12590 33992
rect 13082 33980 13110 34020
rect 12912 33952 13110 33980
rect 13265 33983 13323 33989
rect 12802 33912 12808 33924
rect 11256 33884 12808 33912
rect 10689 33875 10747 33881
rect 12802 33872 12808 33884
rect 12860 33872 12866 33924
rect 7558 33844 7564 33856
rect 7519 33816 7564 33844
rect 7558 33804 7564 33816
rect 7616 33804 7622 33856
rect 9033 33847 9091 33853
rect 9033 33813 9045 33847
rect 9079 33844 9091 33847
rect 12912 33844 12940 33952
rect 13265 33949 13277 33983
rect 13311 33949 13323 33983
rect 13265 33943 13323 33949
rect 13357 33983 13415 33989
rect 13357 33949 13369 33983
rect 13403 33980 13415 33983
rect 13906 33980 13912 33992
rect 13403 33952 13912 33980
rect 13403 33949 13415 33952
rect 13357 33943 13415 33949
rect 13081 33915 13139 33921
rect 13081 33881 13093 33915
rect 13127 33881 13139 33915
rect 13280 33912 13308 33943
rect 13906 33940 13912 33952
rect 13964 33980 13970 33992
rect 14093 33983 14151 33989
rect 14093 33980 14105 33983
rect 13964 33952 14105 33980
rect 13964 33940 13970 33952
rect 14093 33949 14105 33952
rect 14139 33949 14151 33983
rect 14093 33943 14151 33949
rect 14182 33940 14188 33992
rect 14240 33980 14246 33992
rect 14277 33983 14335 33989
rect 14277 33980 14289 33983
rect 14240 33952 14289 33980
rect 14240 33940 14246 33952
rect 14277 33949 14289 33952
rect 14323 33949 14335 33983
rect 14277 33943 14335 33949
rect 14366 33940 14372 33992
rect 14424 33980 14430 33992
rect 14642 33980 14648 33992
rect 14424 33952 14504 33980
rect 14603 33952 14648 33980
rect 14424 33940 14430 33952
rect 14476 33921 14504 33952
rect 14642 33940 14648 33952
rect 14700 33940 14706 33992
rect 14918 33980 14924 33992
rect 14752 33952 14924 33980
rect 14461 33915 14519 33921
rect 13280 33884 14412 33912
rect 13081 33875 13139 33881
rect 9079 33816 12940 33844
rect 13096 33844 13124 33875
rect 14274 33844 14280 33856
rect 13096 33816 14280 33844
rect 9079 33813 9091 33816
rect 9033 33807 9091 33813
rect 14274 33804 14280 33816
rect 14332 33804 14338 33856
rect 14384 33853 14412 33884
rect 14461 33881 14473 33915
rect 14507 33912 14519 33915
rect 14752 33912 14780 33952
rect 14918 33940 14924 33952
rect 14976 33940 14982 33992
rect 14507 33884 14780 33912
rect 14507 33881 14519 33884
rect 14461 33875 14519 33881
rect 14826 33872 14832 33924
rect 14884 33912 14890 33924
rect 15396 33912 15424 34020
rect 18322 34008 18328 34060
rect 18380 34048 18386 34060
rect 19242 34048 19248 34060
rect 18380 34020 19248 34048
rect 18380 34008 18386 34020
rect 19242 34008 19248 34020
rect 19300 34008 19306 34060
rect 20548 34020 21772 34048
rect 15565 33983 15623 33989
rect 15565 33949 15577 33983
rect 15611 33980 15623 33983
rect 15654 33980 15660 33992
rect 15611 33952 15660 33980
rect 15611 33949 15623 33952
rect 15565 33943 15623 33949
rect 15654 33940 15660 33952
rect 15712 33940 15718 33992
rect 16942 33940 16948 33992
rect 17000 33980 17006 33992
rect 17681 33983 17739 33989
rect 17000 33952 17612 33980
rect 17000 33940 17006 33952
rect 15810 33915 15868 33921
rect 15810 33912 15822 33915
rect 14884 33884 15332 33912
rect 15396 33884 15822 33912
rect 14884 33872 14890 33884
rect 14369 33847 14427 33853
rect 14369 33813 14381 33847
rect 14415 33844 14427 33847
rect 15194 33844 15200 33856
rect 14415 33816 15200 33844
rect 14415 33813 14427 33816
rect 14369 33807 14427 33813
rect 15194 33804 15200 33816
rect 15252 33804 15258 33856
rect 15304 33844 15332 33884
rect 15810 33881 15822 33884
rect 15856 33881 15868 33915
rect 15810 33875 15868 33881
rect 17126 33872 17132 33924
rect 17184 33912 17190 33924
rect 17497 33915 17555 33921
rect 17497 33912 17509 33915
rect 17184 33884 17509 33912
rect 17184 33872 17190 33884
rect 17497 33881 17509 33884
rect 17543 33881 17555 33915
rect 17584 33912 17612 33952
rect 17681 33949 17693 33983
rect 17727 33980 17739 33983
rect 20548 33980 20576 34020
rect 17727 33952 20576 33980
rect 17727 33949 17739 33952
rect 17681 33943 17739 33949
rect 20622 33940 20628 33992
rect 20680 33980 20686 33992
rect 21085 33983 21143 33989
rect 21085 33980 21097 33983
rect 20680 33952 21097 33980
rect 20680 33940 20686 33952
rect 21085 33949 21097 33952
rect 21131 33949 21143 33983
rect 21744 33980 21772 34020
rect 21818 34008 21824 34060
rect 21876 34048 21882 34060
rect 22005 34051 22063 34057
rect 22005 34048 22017 34051
rect 21876 34020 22017 34048
rect 21876 34008 21882 34020
rect 22005 34017 22017 34020
rect 22051 34017 22063 34051
rect 22572 34048 22600 34088
rect 23290 34076 23296 34088
rect 23348 34076 23354 34128
rect 23750 34076 23756 34128
rect 23808 34116 23814 34128
rect 24765 34119 24823 34125
rect 24765 34116 24777 34119
rect 23808 34088 24777 34116
rect 23808 34076 23814 34088
rect 24765 34085 24777 34088
rect 24811 34085 24823 34119
rect 26234 34116 26240 34128
rect 24765 34079 24823 34085
rect 25424 34088 26240 34116
rect 23382 34048 23388 34060
rect 22005 34011 22063 34017
rect 22204 34020 22600 34048
rect 23343 34020 23388 34048
rect 22204 33992 22232 34020
rect 23382 34008 23388 34020
rect 23440 34008 23446 34060
rect 23934 34008 23940 34060
rect 23992 34048 23998 34060
rect 24118 34048 24124 34060
rect 23992 34020 24124 34048
rect 23992 34008 23998 34020
rect 24118 34008 24124 34020
rect 24176 34008 24182 34060
rect 25424 34057 25452 34088
rect 26234 34076 26240 34088
rect 26292 34076 26298 34128
rect 25409 34051 25467 34057
rect 25409 34017 25421 34051
rect 25455 34017 25467 34051
rect 25682 34048 25688 34060
rect 25643 34020 25688 34048
rect 25409 34011 25467 34017
rect 25682 34008 25688 34020
rect 25740 34008 25746 34060
rect 26326 34048 26332 34060
rect 26287 34020 26332 34048
rect 26326 34008 26332 34020
rect 26384 34008 26390 34060
rect 28169 34051 28227 34057
rect 28169 34017 28181 34051
rect 28215 34048 28227 34051
rect 28902 34048 28908 34060
rect 28215 34020 28908 34048
rect 28215 34017 28227 34020
rect 28169 34011 28227 34017
rect 28902 34008 28908 34020
rect 28960 34008 28966 34060
rect 22186 33980 22192 33992
rect 21744 33952 22192 33980
rect 21085 33943 21143 33949
rect 22186 33940 22192 33952
rect 22244 33940 22250 33992
rect 22738 33940 22744 33992
rect 22796 33980 22802 33992
rect 23109 33983 23167 33989
rect 23109 33980 23121 33983
rect 22796 33952 23121 33980
rect 22796 33940 22802 33952
rect 23109 33949 23121 33952
rect 23155 33949 23167 33983
rect 23109 33943 23167 33949
rect 25038 33940 25044 33992
rect 25096 33980 25102 33992
rect 25501 33983 25559 33989
rect 25501 33980 25513 33983
rect 25096 33952 25513 33980
rect 25096 33940 25102 33952
rect 25501 33949 25513 33952
rect 25547 33949 25559 33983
rect 25501 33943 25559 33949
rect 25593 33983 25651 33989
rect 25593 33949 25605 33983
rect 25639 33949 25651 33983
rect 25593 33943 25651 33949
rect 18230 33912 18236 33924
rect 17584 33884 18236 33912
rect 17497 33875 17555 33881
rect 18230 33872 18236 33884
rect 18288 33912 18294 33924
rect 18325 33915 18383 33921
rect 18325 33912 18337 33915
rect 18288 33884 18337 33912
rect 18288 33872 18294 33884
rect 18325 33881 18337 33884
rect 18371 33912 18383 33915
rect 18966 33912 18972 33924
rect 18371 33884 18972 33912
rect 18371 33881 18383 33884
rect 18325 33875 18383 33881
rect 18966 33872 18972 33884
rect 19024 33872 19030 33924
rect 19334 33872 19340 33924
rect 19392 33912 19398 33924
rect 19490 33915 19548 33921
rect 19490 33912 19502 33915
rect 19392 33884 19502 33912
rect 19392 33872 19398 33884
rect 19490 33881 19502 33884
rect 19536 33881 19548 33915
rect 21361 33915 21419 33921
rect 21361 33912 21373 33915
rect 19490 33875 19548 33881
rect 19628 33884 21373 33912
rect 18138 33844 18144 33856
rect 15304 33816 18144 33844
rect 18138 33804 18144 33816
rect 18196 33804 18202 33856
rect 18414 33844 18420 33856
rect 18375 33816 18420 33844
rect 18414 33804 18420 33816
rect 18472 33804 18478 33856
rect 18506 33804 18512 33856
rect 18564 33844 18570 33856
rect 18564 33816 18609 33844
rect 18564 33804 18570 33816
rect 18782 33804 18788 33856
rect 18840 33844 18846 33856
rect 19628 33844 19656 33884
rect 21361 33881 21373 33884
rect 21407 33881 21419 33915
rect 24397 33915 24455 33921
rect 24397 33912 24409 33915
rect 21361 33875 21419 33881
rect 22066 33884 24409 33912
rect 18840 33816 19656 33844
rect 18840 33804 18846 33816
rect 20162 33804 20168 33856
rect 20220 33844 20226 33856
rect 20625 33847 20683 33853
rect 20625 33844 20637 33847
rect 20220 33816 20637 33844
rect 20220 33804 20226 33816
rect 20625 33813 20637 33816
rect 20671 33813 20683 33847
rect 20625 33807 20683 33813
rect 20806 33804 20812 33856
rect 20864 33844 20870 33856
rect 22066 33844 22094 33884
rect 24397 33881 24409 33884
rect 24443 33881 24455 33915
rect 24397 33875 24455 33881
rect 24486 33872 24492 33924
rect 24544 33912 24550 33924
rect 24597 33915 24655 33921
rect 24597 33912 24609 33915
rect 24544 33884 24609 33912
rect 24544 33872 24550 33884
rect 24597 33881 24609 33884
rect 24643 33881 24655 33915
rect 25608 33912 25636 33943
rect 26510 33912 26516 33924
rect 24597 33875 24655 33881
rect 24688 33884 25636 33912
rect 26471 33884 26516 33912
rect 22922 33844 22928 33856
rect 20864 33816 22094 33844
rect 22883 33816 22928 33844
rect 20864 33804 20870 33816
rect 22922 33804 22928 33816
rect 22980 33804 22986 33856
rect 23106 33804 23112 33856
rect 23164 33844 23170 33856
rect 24688 33844 24716 33884
rect 26510 33872 26516 33884
rect 26568 33872 26574 33924
rect 25222 33844 25228 33856
rect 23164 33816 24716 33844
rect 25183 33816 25228 33844
rect 23164 33804 23170 33816
rect 25222 33804 25228 33816
rect 25280 33804 25286 33856
rect 1104 33754 28888 33776
rect 1104 33702 10214 33754
rect 10266 33702 10278 33754
rect 10330 33702 10342 33754
rect 10394 33702 10406 33754
rect 10458 33702 10470 33754
rect 10522 33702 19478 33754
rect 19530 33702 19542 33754
rect 19594 33702 19606 33754
rect 19658 33702 19670 33754
rect 19722 33702 19734 33754
rect 19786 33702 28888 33754
rect 1104 33680 28888 33702
rect 1581 33643 1639 33649
rect 1581 33609 1593 33643
rect 1627 33640 1639 33643
rect 2038 33640 2044 33652
rect 1627 33612 2044 33640
rect 1627 33609 1639 33612
rect 1581 33603 1639 33609
rect 2038 33600 2044 33612
rect 2096 33600 2102 33652
rect 2222 33640 2228 33652
rect 2183 33612 2228 33640
rect 2222 33600 2228 33612
rect 2280 33600 2286 33652
rect 9585 33643 9643 33649
rect 9585 33609 9597 33643
rect 9631 33640 9643 33643
rect 9950 33640 9956 33652
rect 9631 33612 9956 33640
rect 9631 33609 9643 33612
rect 9585 33603 9643 33609
rect 9950 33600 9956 33612
rect 10008 33600 10014 33652
rect 11422 33640 11428 33652
rect 10152 33612 11428 33640
rect 10152 33572 10180 33612
rect 11422 33600 11428 33612
rect 11480 33600 11486 33652
rect 11882 33600 11888 33652
rect 11940 33640 11946 33652
rect 12066 33640 12072 33652
rect 11940 33612 12072 33640
rect 11940 33600 11946 33612
rect 12066 33600 12072 33612
rect 12124 33600 12130 33652
rect 15562 33640 15568 33652
rect 12406 33612 15568 33640
rect 12406 33572 12434 33612
rect 15562 33600 15568 33612
rect 15620 33600 15626 33652
rect 18414 33600 18420 33652
rect 18472 33640 18478 33652
rect 20162 33640 20168 33652
rect 18472 33612 20168 33640
rect 18472 33600 18478 33612
rect 20162 33600 20168 33612
rect 20220 33600 20226 33652
rect 21082 33600 21088 33652
rect 21140 33640 21146 33652
rect 21177 33643 21235 33649
rect 21177 33640 21189 33643
rect 21140 33612 21189 33640
rect 21140 33600 21146 33612
rect 21177 33609 21189 33612
rect 21223 33609 21235 33643
rect 21177 33603 21235 33609
rect 25958 33600 25964 33652
rect 26016 33640 26022 33652
rect 28077 33643 28135 33649
rect 28077 33640 28089 33643
rect 26016 33612 28089 33640
rect 26016 33600 26022 33612
rect 28077 33609 28089 33612
rect 28123 33609 28135 33643
rect 28077 33603 28135 33609
rect 9048 33544 10180 33572
rect 10244 33544 12434 33572
rect 1394 33504 1400 33516
rect 1355 33476 1400 33504
rect 1394 33464 1400 33476
rect 1452 33464 1458 33516
rect 1946 33464 1952 33516
rect 2004 33504 2010 33516
rect 2133 33507 2191 33513
rect 2133 33504 2145 33507
rect 2004 33476 2145 33504
rect 2004 33464 2010 33476
rect 2133 33473 2145 33476
rect 2179 33504 2191 33507
rect 7834 33504 7840 33516
rect 2179 33476 7840 33504
rect 2179 33473 2191 33476
rect 2133 33467 2191 33473
rect 7834 33464 7840 33476
rect 7892 33464 7898 33516
rect 8389 33507 8447 33513
rect 8389 33473 8401 33507
rect 8435 33504 8447 33507
rect 8478 33504 8484 33516
rect 8435 33476 8484 33504
rect 8435 33473 8447 33476
rect 8389 33467 8447 33473
rect 8478 33464 8484 33476
rect 8536 33464 8542 33516
rect 9048 33513 9076 33544
rect 9033 33507 9091 33513
rect 9033 33473 9045 33507
rect 9079 33473 9091 33507
rect 9033 33467 9091 33473
rect 9398 33464 9404 33516
rect 9456 33504 9462 33516
rect 9493 33507 9551 33513
rect 9493 33504 9505 33507
rect 9456 33476 9505 33504
rect 9456 33464 9462 33476
rect 9493 33473 9505 33476
rect 9539 33473 9551 33507
rect 9493 33467 9551 33473
rect 9582 33464 9588 33516
rect 9640 33504 9646 33516
rect 9677 33507 9735 33513
rect 9677 33504 9689 33507
rect 9640 33476 9689 33504
rect 9640 33464 9646 33476
rect 9677 33473 9689 33476
rect 9723 33473 9735 33507
rect 9677 33467 9735 33473
rect 10042 33464 10048 33516
rect 10100 33504 10106 33516
rect 10137 33507 10195 33513
rect 10137 33504 10149 33507
rect 10100 33476 10149 33504
rect 10100 33464 10106 33476
rect 10137 33473 10149 33476
rect 10183 33473 10195 33507
rect 10137 33467 10195 33473
rect 7745 33439 7803 33445
rect 7745 33405 7757 33439
rect 7791 33436 7803 33439
rect 10244 33436 10272 33544
rect 12986 33532 12992 33584
rect 13044 33572 13050 33584
rect 17466 33575 17524 33581
rect 17466 33572 17478 33575
rect 13044 33544 17478 33572
rect 13044 33532 13050 33544
rect 17466 33541 17478 33544
rect 17512 33541 17524 33575
rect 17466 33535 17524 33541
rect 18046 33532 18052 33584
rect 18104 33572 18110 33584
rect 18598 33572 18604 33584
rect 18104 33544 18604 33572
rect 18104 33532 18110 33544
rect 18598 33532 18604 33544
rect 18656 33532 18662 33584
rect 19426 33572 19432 33584
rect 18708 33544 19432 33572
rect 10321 33507 10379 33513
rect 10321 33473 10333 33507
rect 10367 33504 10379 33507
rect 10594 33504 10600 33516
rect 10367 33476 10600 33504
rect 10367 33473 10379 33476
rect 10321 33467 10379 33473
rect 10594 33464 10600 33476
rect 10652 33464 10658 33516
rect 10781 33507 10839 33513
rect 10781 33473 10793 33507
rect 10827 33504 10839 33507
rect 10870 33504 10876 33516
rect 10827 33476 10876 33504
rect 10827 33473 10839 33476
rect 10781 33467 10839 33473
rect 10870 33464 10876 33476
rect 10928 33464 10934 33516
rect 10965 33507 11023 33513
rect 10965 33473 10977 33507
rect 11011 33504 11023 33507
rect 11054 33504 11060 33516
rect 11011 33476 11060 33504
rect 11011 33473 11023 33476
rect 10965 33467 11023 33473
rect 11054 33464 11060 33476
rect 11112 33464 11118 33516
rect 11882 33464 11888 33516
rect 11940 33504 11946 33516
rect 11977 33507 12035 33513
rect 11977 33504 11989 33507
rect 11940 33476 11989 33504
rect 11940 33464 11946 33476
rect 11977 33473 11989 33476
rect 12023 33473 12035 33507
rect 12158 33504 12164 33516
rect 12119 33476 12164 33504
rect 11977 33467 12035 33473
rect 12158 33464 12164 33476
rect 12216 33464 12222 33516
rect 12618 33464 12624 33516
rect 12676 33504 12682 33516
rect 12805 33507 12863 33513
rect 12805 33504 12817 33507
rect 12676 33476 12817 33504
rect 12676 33464 12682 33476
rect 12805 33473 12817 33476
rect 12851 33473 12863 33507
rect 12805 33467 12863 33473
rect 13354 33464 13360 33516
rect 13412 33504 13418 33516
rect 13449 33507 13507 33513
rect 13449 33504 13461 33507
rect 13412 33476 13461 33504
rect 13412 33464 13418 33476
rect 13449 33473 13461 33476
rect 13495 33473 13507 33507
rect 13705 33507 13763 33513
rect 13705 33504 13717 33507
rect 13449 33467 13507 33473
rect 13556 33476 13717 33504
rect 7791 33408 10272 33436
rect 7791 33405 7803 33408
rect 7745 33399 7803 33405
rect 10410 33396 10416 33448
rect 10468 33436 10474 33448
rect 12345 33439 12403 33445
rect 12345 33436 12357 33439
rect 10468 33408 10916 33436
rect 10468 33396 10474 33408
rect 8849 33371 8907 33377
rect 8849 33337 8861 33371
rect 8895 33368 8907 33371
rect 10502 33368 10508 33380
rect 8895 33340 10508 33368
rect 8895 33337 8907 33340
rect 8849 33331 8907 33337
rect 10502 33328 10508 33340
rect 10560 33328 10566 33380
rect 10594 33328 10600 33380
rect 10652 33368 10658 33380
rect 10781 33371 10839 33377
rect 10781 33368 10793 33371
rect 10652 33340 10793 33368
rect 10652 33328 10658 33340
rect 10781 33337 10793 33340
rect 10827 33337 10839 33371
rect 10888 33368 10916 33408
rect 11064 33408 12357 33436
rect 11064 33368 11092 33408
rect 12345 33405 12357 33408
rect 12391 33405 12403 33439
rect 12345 33399 12403 33405
rect 12434 33396 12440 33448
rect 12492 33436 12498 33448
rect 12710 33436 12716 33448
rect 12492 33408 12716 33436
rect 12492 33396 12498 33408
rect 12710 33396 12716 33408
rect 12768 33396 12774 33448
rect 12894 33436 12900 33448
rect 12855 33408 12900 33436
rect 12894 33396 12900 33408
rect 12952 33396 12958 33448
rect 12986 33396 12992 33448
rect 13044 33436 13050 33448
rect 13556 33436 13584 33476
rect 13705 33473 13717 33476
rect 13751 33473 13763 33507
rect 13705 33467 13763 33473
rect 13998 33464 14004 33516
rect 14056 33504 14062 33516
rect 15194 33504 15200 33516
rect 14056 33476 15200 33504
rect 14056 33464 14062 33476
rect 15194 33464 15200 33476
rect 15252 33464 15258 33516
rect 15654 33464 15660 33516
rect 15712 33504 15718 33516
rect 17221 33507 17279 33513
rect 17221 33504 17233 33507
rect 15712 33476 17233 33504
rect 15712 33464 15718 33476
rect 17221 33473 17233 33476
rect 17267 33473 17279 33507
rect 18708 33504 18736 33544
rect 19426 33532 19432 33544
rect 19484 33532 19490 33584
rect 19886 33532 19892 33584
rect 19944 33572 19950 33584
rect 20042 33575 20100 33581
rect 20042 33572 20054 33575
rect 19944 33544 20054 33572
rect 19944 33532 19950 33544
rect 20042 33541 20054 33544
rect 20088 33541 20100 33575
rect 20042 33535 20100 33541
rect 23290 33532 23296 33584
rect 23348 33572 23354 33584
rect 23348 33544 23796 33572
rect 23348 33532 23354 33544
rect 17221 33467 17279 33473
rect 17328 33476 18736 33504
rect 13044 33408 13584 33436
rect 13044 33396 13050 33408
rect 14458 33396 14464 33448
rect 14516 33436 14522 33448
rect 14516 33408 14964 33436
rect 14516 33396 14522 33408
rect 13354 33368 13360 33380
rect 10888 33340 11092 33368
rect 11164 33340 13360 33368
rect 10781 33331 10839 33337
rect 8205 33303 8263 33309
rect 8205 33269 8217 33303
rect 8251 33300 8263 33303
rect 10042 33300 10048 33312
rect 8251 33272 10048 33300
rect 8251 33269 8263 33272
rect 8205 33263 8263 33269
rect 10042 33260 10048 33272
rect 10100 33260 10106 33312
rect 10137 33303 10195 33309
rect 10137 33269 10149 33303
rect 10183 33300 10195 33303
rect 11164 33300 11192 33340
rect 13354 33328 13360 33340
rect 13412 33328 13418 33380
rect 14826 33368 14832 33380
rect 14787 33340 14832 33368
rect 14826 33328 14832 33340
rect 14884 33328 14890 33380
rect 14936 33368 14964 33408
rect 15102 33396 15108 33448
rect 15160 33436 15166 33448
rect 15289 33439 15347 33445
rect 15289 33436 15301 33439
rect 15160 33408 15301 33436
rect 15160 33396 15166 33408
rect 15289 33405 15301 33408
rect 15335 33405 15347 33439
rect 17328 33436 17356 33476
rect 19150 33464 19156 33516
rect 19208 33504 19214 33516
rect 19208 33476 19253 33504
rect 19208 33464 19214 33476
rect 19334 33464 19340 33516
rect 19392 33504 19398 33516
rect 19610 33504 19616 33516
rect 19392 33476 19616 33504
rect 19392 33464 19398 33476
rect 19610 33464 19616 33476
rect 19668 33504 19674 33516
rect 19797 33507 19855 33513
rect 19797 33504 19809 33507
rect 19668 33476 19809 33504
rect 19668 33464 19674 33476
rect 19797 33473 19809 33476
rect 19843 33473 19855 33507
rect 22002 33504 22008 33516
rect 19797 33467 19855 33473
rect 19904 33476 22008 33504
rect 19904 33436 19932 33476
rect 22002 33464 22008 33476
rect 22060 33513 22066 33516
rect 22060 33507 22109 33513
rect 22060 33473 22063 33507
rect 22097 33473 22109 33507
rect 22186 33504 22192 33516
rect 22147 33476 22192 33504
rect 22060 33467 22109 33473
rect 22060 33464 22066 33467
rect 22186 33464 22192 33476
rect 22244 33464 22250 33516
rect 22302 33507 22360 33513
rect 22302 33473 22314 33507
rect 22348 33504 22360 33507
rect 22348 33476 22416 33504
rect 22348 33473 22360 33476
rect 22302 33467 22360 33473
rect 15289 33399 15347 33405
rect 15396 33408 17356 33436
rect 19260 33408 19932 33436
rect 22388 33436 22416 33476
rect 22462 33464 22468 33516
rect 22520 33504 22526 33516
rect 23638 33504 23644 33516
rect 22520 33476 22565 33504
rect 23599 33476 23644 33504
rect 22520 33464 22526 33476
rect 23638 33464 23644 33476
rect 23696 33464 23702 33516
rect 23768 33513 23796 33544
rect 24762 33532 24768 33584
rect 24820 33572 24826 33584
rect 27614 33572 27620 33584
rect 24820 33544 27620 33572
rect 24820 33532 24826 33544
rect 27614 33532 27620 33544
rect 27672 33532 27678 33584
rect 23753 33507 23811 33513
rect 23753 33473 23765 33507
rect 23799 33473 23811 33507
rect 23753 33467 23811 33473
rect 23842 33464 23848 33516
rect 23900 33507 23906 33516
rect 24029 33507 24087 33513
rect 23900 33479 23942 33507
rect 23900 33464 23906 33479
rect 24029 33473 24041 33507
rect 24075 33473 24087 33507
rect 24029 33467 24087 33473
rect 22554 33436 22560 33448
rect 22388 33408 22560 33436
rect 15396 33368 15424 33408
rect 14936 33340 15424 33368
rect 15470 33328 15476 33380
rect 15528 33377 15534 33380
rect 15528 33371 15577 33377
rect 15528 33337 15531 33371
rect 15565 33368 15577 33371
rect 16298 33368 16304 33380
rect 15565 33340 16304 33368
rect 15565 33337 15577 33340
rect 15528 33331 15577 33337
rect 15528 33328 15534 33331
rect 16298 33328 16304 33340
rect 16356 33328 16362 33380
rect 18598 33368 18604 33380
rect 18559 33340 18604 33368
rect 18598 33328 18604 33340
rect 18656 33328 18662 33380
rect 10183 33272 11192 33300
rect 10183 33269 10195 33272
rect 10137 33263 10195 33269
rect 11238 33260 11244 33312
rect 11296 33300 11302 33312
rect 14734 33300 14740 33312
rect 11296 33272 14740 33300
rect 11296 33260 11302 33272
rect 14734 33260 14740 33272
rect 14792 33260 14798 33312
rect 15194 33260 15200 33312
rect 15252 33300 15258 33312
rect 19260 33300 19288 33408
rect 22554 33396 22560 33408
rect 22612 33396 22618 33448
rect 22830 33396 22836 33448
rect 22888 33436 22894 33448
rect 24044 33436 24072 33467
rect 26970 33464 26976 33516
rect 27028 33504 27034 33516
rect 27157 33507 27215 33513
rect 27157 33504 27169 33507
rect 27028 33476 27169 33504
rect 27028 33464 27034 33476
rect 27157 33473 27169 33476
rect 27203 33473 27215 33507
rect 27157 33467 27215 33473
rect 27985 33507 28043 33513
rect 27985 33473 27997 33507
rect 28031 33504 28043 33507
rect 28166 33504 28172 33516
rect 28031 33476 28172 33504
rect 28031 33473 28043 33476
rect 27985 33467 28043 33473
rect 22888 33408 24072 33436
rect 22888 33396 22894 33408
rect 19337 33371 19395 33377
rect 19337 33337 19349 33371
rect 19383 33368 19395 33371
rect 19794 33368 19800 33380
rect 19383 33340 19800 33368
rect 19383 33337 19395 33340
rect 19337 33331 19395 33337
rect 19794 33328 19800 33340
rect 19852 33328 19858 33380
rect 24044 33368 24072 33408
rect 24118 33396 24124 33448
rect 24176 33436 24182 33448
rect 24581 33439 24639 33445
rect 24581 33436 24593 33439
rect 24176 33408 24593 33436
rect 24176 33396 24182 33408
rect 24581 33405 24593 33408
rect 24627 33405 24639 33439
rect 24581 33399 24639 33405
rect 24765 33439 24823 33445
rect 24765 33405 24777 33439
rect 24811 33436 24823 33439
rect 24946 33436 24952 33448
rect 24811 33408 24952 33436
rect 24811 33405 24823 33408
rect 24765 33399 24823 33405
rect 24946 33396 24952 33408
rect 25004 33396 25010 33448
rect 25314 33436 25320 33448
rect 25148 33408 25320 33436
rect 25148 33368 25176 33408
rect 25314 33396 25320 33408
rect 25372 33396 25378 33448
rect 26142 33436 26148 33448
rect 26103 33408 26148 33436
rect 26142 33396 26148 33408
rect 26200 33396 26206 33448
rect 27249 33439 27307 33445
rect 27249 33405 27261 33439
rect 27295 33436 27307 33439
rect 27706 33436 27712 33448
rect 27295 33408 27712 33436
rect 27295 33405 27307 33408
rect 27249 33399 27307 33405
rect 27264 33368 27292 33399
rect 27706 33396 27712 33408
rect 27764 33396 27770 33448
rect 20732 33340 23980 33368
rect 24044 33340 25176 33368
rect 25240 33340 27292 33368
rect 15252 33272 19288 33300
rect 15252 33260 15258 33272
rect 19426 33260 19432 33312
rect 19484 33300 19490 33312
rect 20732 33300 20760 33340
rect 21818 33300 21824 33312
rect 19484 33272 20760 33300
rect 21779 33272 21824 33300
rect 19484 33260 19490 33272
rect 21818 33260 21824 33272
rect 21876 33260 21882 33312
rect 22002 33260 22008 33312
rect 22060 33300 22066 33312
rect 22646 33300 22652 33312
rect 22060 33272 22652 33300
rect 22060 33260 22066 33272
rect 22646 33260 22652 33272
rect 22704 33260 22710 33312
rect 23385 33303 23443 33309
rect 23385 33269 23397 33303
rect 23431 33300 23443 33303
rect 23750 33300 23756 33312
rect 23431 33272 23756 33300
rect 23431 33269 23443 33272
rect 23385 33263 23443 33269
rect 23750 33260 23756 33272
rect 23808 33260 23814 33312
rect 23952 33300 23980 33340
rect 25240 33300 25268 33340
rect 23952 33272 25268 33300
rect 27246 33260 27252 33312
rect 27304 33300 27310 33312
rect 27433 33303 27491 33309
rect 27433 33300 27445 33303
rect 27304 33272 27445 33300
rect 27304 33260 27310 33272
rect 27433 33269 27445 33272
rect 27479 33269 27491 33303
rect 27433 33263 27491 33269
rect 27706 33260 27712 33312
rect 27764 33300 27770 33312
rect 28000 33300 28028 33467
rect 28166 33464 28172 33476
rect 28224 33464 28230 33516
rect 27764 33272 28028 33300
rect 27764 33260 27770 33272
rect 1104 33210 28888 33232
rect 1104 33158 5582 33210
rect 5634 33158 5646 33210
rect 5698 33158 5710 33210
rect 5762 33158 5774 33210
rect 5826 33158 5838 33210
rect 5890 33158 14846 33210
rect 14898 33158 14910 33210
rect 14962 33158 14974 33210
rect 15026 33158 15038 33210
rect 15090 33158 15102 33210
rect 15154 33158 24110 33210
rect 24162 33158 24174 33210
rect 24226 33158 24238 33210
rect 24290 33158 24302 33210
rect 24354 33158 24366 33210
rect 24418 33158 28888 33210
rect 1104 33136 28888 33158
rect 1397 33099 1455 33105
rect 1397 33065 1409 33099
rect 1443 33096 1455 33099
rect 3418 33096 3424 33108
rect 1443 33068 3424 33096
rect 1443 33065 1455 33068
rect 1397 33059 1455 33065
rect 3418 33056 3424 33068
rect 3476 33056 3482 33108
rect 8205 33099 8263 33105
rect 8205 33065 8217 33099
rect 8251 33096 8263 33099
rect 10594 33096 10600 33108
rect 8251 33068 10600 33096
rect 8251 33065 8263 33068
rect 8205 33059 8263 33065
rect 10594 33056 10600 33068
rect 10652 33056 10658 33108
rect 10686 33056 10692 33108
rect 10744 33096 10750 33108
rect 11606 33096 11612 33108
rect 10744 33068 11612 33096
rect 10744 33056 10750 33068
rect 11606 33056 11612 33068
rect 11664 33056 11670 33108
rect 12066 33056 12072 33108
rect 12124 33096 12130 33108
rect 12345 33099 12403 33105
rect 12345 33096 12357 33099
rect 12124 33068 12357 33096
rect 12124 33056 12130 33068
rect 12345 33065 12357 33068
rect 12391 33065 12403 33099
rect 13262 33096 13268 33108
rect 12345 33059 12403 33065
rect 12547 33068 13268 33096
rect 9030 32988 9036 33040
rect 9088 33028 9094 33040
rect 9490 33028 9496 33040
rect 9088 33000 9496 33028
rect 9088 32988 9094 33000
rect 9490 32988 9496 33000
rect 9548 32988 9554 33040
rect 9585 33031 9643 33037
rect 9585 32997 9597 33031
rect 9631 33028 9643 33031
rect 10778 33028 10784 33040
rect 9631 33000 10784 33028
rect 9631 32997 9643 33000
rect 9585 32991 9643 32997
rect 10778 32988 10784 33000
rect 10836 32988 10842 33040
rect 11974 32988 11980 33040
rect 12032 33028 12038 33040
rect 12547 33028 12575 33068
rect 13262 33056 13268 33068
rect 13320 33056 13326 33108
rect 13354 33056 13360 33108
rect 13412 33096 13418 33108
rect 17681 33099 17739 33105
rect 13412 33068 17632 33096
rect 13412 33056 13418 33068
rect 12032 33000 12575 33028
rect 12032 32988 12038 33000
rect 13078 32988 13084 33040
rect 13136 33028 13142 33040
rect 17604 33028 17632 33068
rect 17681 33065 17693 33099
rect 17727 33096 17739 33099
rect 18046 33096 18052 33108
rect 17727 33068 18052 33096
rect 17727 33065 17739 33068
rect 17681 33059 17739 33065
rect 18046 33056 18052 33068
rect 18104 33056 18110 33108
rect 18230 33096 18236 33108
rect 18191 33068 18236 33096
rect 18230 33056 18236 33068
rect 18288 33056 18294 33108
rect 18340 33068 23244 33096
rect 18340 33028 18368 33068
rect 21082 33028 21088 33040
rect 13136 33000 15516 33028
rect 17604 33000 18368 33028
rect 18432 33000 21088 33028
rect 13136 32988 13142 33000
rect 10870 32960 10876 32972
rect 9508 32932 10876 32960
rect 1486 32852 1492 32904
rect 1544 32892 1550 32904
rect 1581 32895 1639 32901
rect 1581 32892 1593 32895
rect 1544 32864 1593 32892
rect 1544 32852 1550 32864
rect 1581 32861 1593 32864
rect 1627 32861 1639 32895
rect 1581 32855 1639 32861
rect 7745 32895 7803 32901
rect 7745 32861 7757 32895
rect 7791 32892 7803 32895
rect 7834 32892 7840 32904
rect 7791 32864 7840 32892
rect 7791 32861 7803 32864
rect 7745 32855 7803 32861
rect 7834 32852 7840 32864
rect 7892 32852 7898 32904
rect 8389 32895 8447 32901
rect 8389 32861 8401 32895
rect 8435 32892 8447 32895
rect 8938 32892 8944 32904
rect 8435 32864 8944 32892
rect 8435 32861 8447 32864
rect 8389 32855 8447 32861
rect 8938 32852 8944 32864
rect 8996 32852 9002 32904
rect 9508 32901 9536 32932
rect 10870 32920 10876 32932
rect 10928 32920 10934 32972
rect 12066 32920 12072 32972
rect 12124 32960 12130 32972
rect 12124 32932 13124 32960
rect 12124 32920 12130 32932
rect 13096 32904 13124 32932
rect 14182 32920 14188 32972
rect 14240 32960 14246 32972
rect 14737 32963 14795 32969
rect 14240 32932 14504 32960
rect 14240 32920 14246 32932
rect 9493 32895 9551 32901
rect 9493 32861 9505 32895
rect 9539 32861 9551 32895
rect 9493 32855 9551 32861
rect 9677 32895 9735 32901
rect 9677 32861 9689 32895
rect 9723 32892 9735 32895
rect 9766 32892 9772 32904
rect 9723 32864 9772 32892
rect 9723 32861 9735 32864
rect 9677 32855 9735 32861
rect 8754 32784 8760 32836
rect 8812 32824 8818 32836
rect 9692 32824 9720 32855
rect 9766 32852 9772 32864
rect 9824 32852 9830 32904
rect 9858 32852 9864 32904
rect 9916 32892 9922 32904
rect 10134 32892 10140 32904
rect 9916 32864 10140 32892
rect 9916 32852 9922 32864
rect 10134 32852 10140 32864
rect 10192 32852 10198 32904
rect 10229 32895 10287 32901
rect 10229 32861 10241 32895
rect 10275 32861 10287 32895
rect 10229 32855 10287 32861
rect 8812 32796 9720 32824
rect 10244 32824 10272 32855
rect 10318 32852 10324 32904
rect 10376 32892 10382 32904
rect 10376 32864 10421 32892
rect 10376 32852 10382 32864
rect 10594 32852 10600 32904
rect 10652 32892 10658 32904
rect 10965 32895 11023 32901
rect 10652 32864 10732 32892
rect 10652 32852 10658 32864
rect 10704 32824 10732 32864
rect 10965 32861 10977 32895
rect 11011 32892 11023 32895
rect 11514 32892 11520 32904
rect 11011 32864 11520 32892
rect 11011 32861 11023 32864
rect 10965 32855 11023 32861
rect 11514 32852 11520 32864
rect 11572 32852 11578 32904
rect 11624 32864 12575 32892
rect 11210 32827 11268 32833
rect 11210 32824 11222 32827
rect 10244 32796 10640 32824
rect 10704 32796 11222 32824
rect 8812 32784 8818 32796
rect 9490 32716 9496 32768
rect 9548 32756 9554 32768
rect 10505 32759 10563 32765
rect 10505 32756 10517 32759
rect 9548 32728 10517 32756
rect 9548 32716 9554 32728
rect 10505 32725 10517 32728
rect 10551 32725 10563 32759
rect 10612 32756 10640 32796
rect 11210 32793 11222 32796
rect 11256 32793 11268 32827
rect 11210 32787 11268 32793
rect 11330 32784 11336 32836
rect 11388 32824 11394 32836
rect 11624 32824 11652 32864
rect 11388 32796 11652 32824
rect 11388 32784 11394 32796
rect 11698 32784 11704 32836
rect 11756 32824 11762 32836
rect 12434 32824 12440 32836
rect 11756 32796 12440 32824
rect 11756 32784 11762 32796
rect 12434 32784 12440 32796
rect 12492 32784 12498 32836
rect 12547 32824 12575 32864
rect 12618 32852 12624 32904
rect 12676 32892 12682 32904
rect 12676 32864 13032 32892
rect 12676 32852 12682 32864
rect 12802 32824 12808 32836
rect 12547 32796 12808 32824
rect 12802 32784 12808 32796
rect 12860 32784 12866 32836
rect 13004 32833 13032 32864
rect 13078 32852 13084 32904
rect 13136 32892 13142 32904
rect 14476 32901 14504 32932
rect 14737 32929 14749 32963
rect 14783 32960 14795 32963
rect 14826 32960 14832 32972
rect 14783 32932 14832 32960
rect 14783 32929 14795 32932
rect 14737 32923 14795 32929
rect 14826 32920 14832 32932
rect 14884 32920 14890 32972
rect 13357 32895 13415 32901
rect 13136 32864 13229 32892
rect 13136 32852 13142 32864
rect 13357 32861 13369 32895
rect 13403 32892 13415 32895
rect 14277 32895 14335 32901
rect 14277 32892 14289 32895
rect 13403 32864 14289 32892
rect 13403 32861 13415 32864
rect 13357 32855 13415 32861
rect 14277 32861 14289 32864
rect 14323 32861 14335 32895
rect 14277 32855 14335 32861
rect 14461 32895 14519 32901
rect 14461 32861 14473 32895
rect 14507 32892 14519 32895
rect 15378 32892 15384 32904
rect 14507 32864 15384 32892
rect 14507 32861 14519 32864
rect 14461 32855 14519 32861
rect 15378 32852 15384 32864
rect 15436 32852 15442 32904
rect 15488 32892 15516 33000
rect 15654 32960 15660 32972
rect 15615 32932 15660 32960
rect 15654 32920 15660 32932
rect 15712 32920 15718 32972
rect 18432 32960 18460 33000
rect 21082 32988 21088 33000
rect 21140 32988 21146 33040
rect 22646 33028 22652 33040
rect 22607 33000 22652 33028
rect 22646 32988 22652 33000
rect 22704 32988 22710 33040
rect 17420 32932 18460 32960
rect 17420 32892 17448 32932
rect 19610 32920 19616 32972
rect 19668 32960 19674 32972
rect 23216 32969 23244 33068
rect 23934 33056 23940 33108
rect 23992 33096 23998 33108
rect 27430 33096 27436 33108
rect 23992 33068 27436 33096
rect 23992 33056 23998 33068
rect 23201 32963 23259 32969
rect 19668 32932 21312 32960
rect 19668 32920 19674 32932
rect 21284 32904 21312 32932
rect 23201 32929 23213 32963
rect 23247 32929 23259 32963
rect 24670 32960 24676 32972
rect 23201 32923 23259 32929
rect 23308 32932 24676 32960
rect 15488 32864 17448 32892
rect 17494 32852 17500 32904
rect 17552 32892 17558 32904
rect 17552 32864 17597 32892
rect 17552 32852 17558 32864
rect 18230 32852 18236 32904
rect 18288 32892 18294 32904
rect 18414 32892 18420 32904
rect 18288 32864 18333 32892
rect 18375 32864 18420 32892
rect 18288 32852 18294 32864
rect 18414 32852 18420 32864
rect 18472 32852 18478 32904
rect 18509 32895 18567 32901
rect 18509 32861 18521 32895
rect 18555 32892 18567 32895
rect 18598 32892 18604 32904
rect 18555 32864 18604 32892
rect 18555 32861 18567 32864
rect 18509 32855 18567 32861
rect 18598 32852 18604 32864
rect 18656 32852 18662 32904
rect 19242 32892 19248 32904
rect 19203 32864 19248 32892
rect 19242 32852 19248 32864
rect 19300 32852 19306 32904
rect 19426 32892 19432 32904
rect 19387 32864 19432 32892
rect 19426 32852 19432 32864
rect 19484 32892 19490 32904
rect 19702 32892 19708 32904
rect 19484 32864 19708 32892
rect 19484 32852 19490 32864
rect 19702 32852 19708 32864
rect 19760 32852 19766 32904
rect 19794 32852 19800 32904
rect 19852 32892 19858 32904
rect 20165 32895 20223 32901
rect 20165 32892 20177 32895
rect 19852 32864 20177 32892
rect 19852 32852 19858 32864
rect 20165 32861 20177 32864
rect 20211 32892 20223 32895
rect 20622 32892 20628 32904
rect 20211 32864 20628 32892
rect 20211 32861 20223 32864
rect 20165 32855 20223 32861
rect 20622 32852 20628 32864
rect 20680 32852 20686 32904
rect 21266 32892 21272 32904
rect 21227 32864 21272 32892
rect 21266 32852 21272 32864
rect 21324 32852 21330 32904
rect 21536 32895 21594 32901
rect 21536 32861 21548 32895
rect 21582 32892 21594 32895
rect 21818 32892 21824 32904
rect 21582 32864 21824 32892
rect 21582 32861 21594 32864
rect 21536 32855 21594 32861
rect 21818 32852 21824 32864
rect 21876 32852 21882 32904
rect 21910 32852 21916 32904
rect 21968 32892 21974 32904
rect 23308 32892 23336 32932
rect 24670 32920 24676 32932
rect 24728 32960 24734 32972
rect 24728 32932 24799 32960
rect 24728 32920 24734 32932
rect 21968 32864 23336 32892
rect 23371 32895 23429 32901
rect 21968 32852 21974 32864
rect 23371 32861 23383 32895
rect 23417 32892 23429 32895
rect 23474 32892 23480 32904
rect 23417 32864 23480 32892
rect 23417 32861 23429 32864
rect 23371 32855 23429 32861
rect 23474 32852 23480 32864
rect 23532 32852 23538 32904
rect 24771 32901 24799 32932
rect 24872 32901 24900 33068
rect 27430 33056 27436 33068
rect 27488 33056 27494 33108
rect 28350 33028 28356 33040
rect 25884 33000 28356 33028
rect 25038 32960 25044 32972
rect 24964 32932 25044 32960
rect 24964 32901 24992 32932
rect 25038 32920 25044 32932
rect 25096 32920 25102 32972
rect 25406 32920 25412 32972
rect 25464 32960 25470 32972
rect 25685 32963 25743 32969
rect 25685 32960 25697 32963
rect 25464 32932 25697 32960
rect 25464 32920 25470 32932
rect 25685 32929 25697 32932
rect 25731 32929 25743 32963
rect 25685 32923 25743 32929
rect 25774 32920 25780 32972
rect 25832 32960 25838 32972
rect 25884 32969 25912 33000
rect 28350 32988 28356 33000
rect 28408 32988 28414 33040
rect 25869 32963 25927 32969
rect 25869 32960 25881 32963
rect 25832 32932 25881 32960
rect 25832 32920 25838 32932
rect 25869 32929 25881 32932
rect 25915 32929 25927 32963
rect 26326 32960 26332 32972
rect 26287 32932 26332 32960
rect 25869 32923 25927 32929
rect 26326 32920 26332 32932
rect 26384 32920 26390 32972
rect 28166 32960 28172 32972
rect 28127 32932 28172 32960
rect 28166 32920 28172 32932
rect 28224 32920 28230 32972
rect 24765 32895 24823 32901
rect 24765 32861 24777 32895
rect 24811 32861 24823 32895
rect 24765 32855 24823 32861
rect 24854 32895 24912 32901
rect 24854 32861 24866 32895
rect 24900 32861 24912 32895
rect 24854 32855 24912 32861
rect 24954 32895 25012 32901
rect 24954 32861 24966 32895
rect 25000 32861 25012 32895
rect 24954 32855 25012 32861
rect 25133 32895 25191 32901
rect 25133 32861 25145 32895
rect 25179 32892 25191 32895
rect 25314 32892 25320 32904
rect 25179 32864 25320 32892
rect 25179 32861 25191 32864
rect 25133 32855 25191 32861
rect 25314 32852 25320 32864
rect 25372 32852 25378 32904
rect 25498 32852 25504 32904
rect 25556 32892 25562 32904
rect 25593 32895 25651 32901
rect 25593 32892 25605 32895
rect 25556 32864 25605 32892
rect 25556 32852 25562 32864
rect 25593 32861 25605 32864
rect 25639 32861 25651 32895
rect 25593 32855 25651 32861
rect 12989 32827 13047 32833
rect 12989 32793 13001 32827
rect 13035 32824 13047 32827
rect 13446 32824 13452 32836
rect 13035 32796 13452 32824
rect 13035 32793 13047 32796
rect 12989 32787 13047 32793
rect 13446 32784 13452 32796
rect 13504 32784 13510 32836
rect 13538 32784 13544 32836
rect 13596 32824 13602 32836
rect 14366 32824 14372 32836
rect 13596 32796 14289 32824
rect 14327 32796 14372 32824
rect 13596 32784 13602 32796
rect 12710 32756 12716 32768
rect 10612 32728 12716 32756
rect 10505 32719 10563 32725
rect 12710 32716 12716 32728
rect 12768 32716 12774 32768
rect 13170 32756 13176 32768
rect 13131 32728 13176 32756
rect 13170 32716 13176 32728
rect 13228 32716 13234 32768
rect 14090 32756 14096 32768
rect 14051 32728 14096 32756
rect 14090 32716 14096 32728
rect 14148 32716 14154 32768
rect 14261 32756 14289 32796
rect 14366 32784 14372 32796
rect 14424 32784 14430 32836
rect 14550 32784 14556 32836
rect 14608 32833 14614 32836
rect 14608 32827 14637 32833
rect 14625 32793 14637 32827
rect 14608 32787 14637 32793
rect 14608 32784 14614 32787
rect 14734 32784 14740 32836
rect 14792 32824 14798 32836
rect 15902 32827 15960 32833
rect 15902 32824 15914 32827
rect 14792 32796 15914 32824
rect 14792 32784 14798 32796
rect 15902 32793 15914 32796
rect 15948 32793 15960 32827
rect 15902 32787 15960 32793
rect 15988 32796 20024 32824
rect 15988 32756 16016 32796
rect 14261 32728 16016 32756
rect 16298 32716 16304 32768
rect 16356 32756 16362 32768
rect 17037 32759 17095 32765
rect 17037 32756 17049 32759
rect 16356 32728 17049 32756
rect 16356 32716 16362 32728
rect 17037 32725 17049 32728
rect 17083 32756 17095 32759
rect 17126 32756 17132 32768
rect 17083 32728 17132 32756
rect 17083 32725 17095 32728
rect 17037 32719 17095 32725
rect 17126 32716 17132 32728
rect 17184 32716 17190 32768
rect 18230 32716 18236 32768
rect 18288 32756 18294 32768
rect 18506 32756 18512 32768
rect 18288 32728 18512 32756
rect 18288 32716 18294 32728
rect 18506 32716 18512 32728
rect 18564 32716 18570 32768
rect 18690 32756 18696 32768
rect 18651 32728 18696 32756
rect 18690 32716 18696 32728
rect 18748 32716 18754 32768
rect 19334 32716 19340 32768
rect 19392 32756 19398 32768
rect 19613 32759 19671 32765
rect 19613 32756 19625 32759
rect 19392 32728 19625 32756
rect 19392 32716 19398 32728
rect 19613 32725 19625 32728
rect 19659 32725 19671 32759
rect 19886 32756 19892 32768
rect 19847 32728 19892 32756
rect 19613 32719 19671 32725
rect 19886 32716 19892 32728
rect 19944 32716 19950 32768
rect 19996 32756 20024 32796
rect 20346 32784 20352 32836
rect 20404 32824 20410 32836
rect 20533 32827 20591 32833
rect 20533 32824 20545 32827
rect 20404 32796 20545 32824
rect 20404 32784 20410 32796
rect 20533 32793 20545 32796
rect 20579 32793 20591 32827
rect 20533 32787 20591 32793
rect 21082 32784 21088 32836
rect 21140 32824 21146 32836
rect 26513 32827 26571 32833
rect 26513 32824 26525 32827
rect 21140 32796 26525 32824
rect 21140 32784 21146 32796
rect 26513 32793 26525 32796
rect 26559 32793 26571 32827
rect 26513 32787 26571 32793
rect 23661 32759 23719 32765
rect 23661 32756 23673 32759
rect 19996 32728 23673 32756
rect 23661 32725 23673 32728
rect 23707 32725 23719 32759
rect 23661 32719 23719 32725
rect 24489 32759 24547 32765
rect 24489 32725 24501 32759
rect 24535 32756 24547 32759
rect 24578 32756 24584 32768
rect 24535 32728 24584 32756
rect 24535 32725 24547 32728
rect 24489 32719 24547 32725
rect 24578 32716 24584 32728
rect 24636 32716 24642 32768
rect 24946 32716 24952 32768
rect 25004 32756 25010 32768
rect 25869 32759 25927 32765
rect 25869 32756 25881 32759
rect 25004 32728 25881 32756
rect 25004 32716 25010 32728
rect 25869 32725 25881 32728
rect 25915 32725 25927 32759
rect 25869 32719 25927 32725
rect 1104 32666 28888 32688
rect 1104 32614 10214 32666
rect 10266 32614 10278 32666
rect 10330 32614 10342 32666
rect 10394 32614 10406 32666
rect 10458 32614 10470 32666
rect 10522 32614 19478 32666
rect 19530 32614 19542 32666
rect 19594 32614 19606 32666
rect 19658 32614 19670 32666
rect 19722 32614 19734 32666
rect 19786 32614 28888 32666
rect 1104 32592 28888 32614
rect 7929 32555 7987 32561
rect 7929 32521 7941 32555
rect 7975 32552 7987 32555
rect 12894 32552 12900 32564
rect 7975 32524 10364 32552
rect 7975 32521 7987 32524
rect 7929 32515 7987 32521
rect 10336 32496 10364 32524
rect 10428 32524 12900 32552
rect 9490 32484 9496 32496
rect 7484 32456 9496 32484
rect 7484 32425 7512 32456
rect 9490 32444 9496 32456
rect 9548 32444 9554 32496
rect 9858 32484 9864 32496
rect 9646 32456 9864 32484
rect 7469 32419 7527 32425
rect 7469 32385 7481 32419
rect 7515 32385 7527 32419
rect 8110 32416 8116 32428
rect 8071 32388 8116 32416
rect 7469 32379 7527 32385
rect 8110 32376 8116 32388
rect 8168 32376 8174 32428
rect 8573 32419 8631 32425
rect 8573 32385 8585 32419
rect 8619 32385 8631 32419
rect 8754 32416 8760 32428
rect 8715 32388 8760 32416
rect 8573 32379 8631 32385
rect 1486 32348 1492 32360
rect 1447 32320 1492 32348
rect 1486 32308 1492 32320
rect 1544 32308 1550 32360
rect 1673 32351 1731 32357
rect 1673 32317 1685 32351
rect 1719 32348 1731 32351
rect 1762 32348 1768 32360
rect 1719 32320 1768 32348
rect 1719 32317 1731 32320
rect 1673 32311 1731 32317
rect 1762 32308 1768 32320
rect 1820 32308 1826 32360
rect 2866 32348 2872 32360
rect 2827 32320 2872 32348
rect 2866 32308 2872 32320
rect 2924 32308 2930 32360
rect 8588 32348 8616 32379
rect 8754 32376 8760 32388
rect 8812 32376 8818 32428
rect 9401 32419 9459 32425
rect 9401 32385 9413 32419
rect 9447 32416 9459 32419
rect 9646 32416 9674 32456
rect 9858 32444 9864 32456
rect 9916 32444 9922 32496
rect 9953 32487 10011 32493
rect 9953 32453 9965 32487
rect 9999 32484 10011 32487
rect 10042 32484 10048 32496
rect 9999 32456 10048 32484
rect 9999 32453 10011 32456
rect 9953 32447 10011 32453
rect 10042 32444 10048 32456
rect 10100 32444 10106 32496
rect 10318 32444 10324 32496
rect 10376 32444 10382 32496
rect 10428 32416 10456 32524
rect 12894 32512 12900 32524
rect 12952 32512 12958 32564
rect 13354 32512 13360 32564
rect 13412 32552 13418 32564
rect 13412 32524 25728 32552
rect 13412 32512 13418 32524
rect 12158 32484 12164 32496
rect 11164 32456 12164 32484
rect 10686 32416 10692 32428
rect 9447 32388 9674 32416
rect 10066 32388 10456 32416
rect 10520 32388 10692 32416
rect 9447 32385 9459 32388
rect 9401 32379 9459 32385
rect 10066 32348 10094 32388
rect 8588 32320 9812 32348
rect 8662 32280 8668 32292
rect 8623 32252 8668 32280
rect 8662 32240 8668 32252
rect 8720 32240 8726 32292
rect 9674 32280 9680 32292
rect 9048 32252 9680 32280
rect 7285 32215 7343 32221
rect 7285 32181 7297 32215
rect 7331 32212 7343 32215
rect 9048 32212 9076 32252
rect 9674 32240 9680 32252
rect 9732 32240 9738 32292
rect 9784 32280 9812 32320
rect 9876 32320 10094 32348
rect 10137 32351 10195 32357
rect 9876 32280 9904 32320
rect 10137 32317 10149 32351
rect 10183 32348 10195 32351
rect 10410 32348 10416 32360
rect 10183 32320 10416 32348
rect 10183 32317 10195 32320
rect 10137 32311 10195 32317
rect 10410 32308 10416 32320
rect 10468 32348 10474 32360
rect 10520 32348 10548 32388
rect 10686 32376 10692 32388
rect 10744 32376 10750 32428
rect 10778 32376 10784 32428
rect 10836 32416 10842 32428
rect 11164 32416 11192 32456
rect 12158 32444 12164 32456
rect 12216 32444 12222 32496
rect 12802 32444 12808 32496
rect 12860 32484 12866 32496
rect 12860 32456 13676 32484
rect 12860 32444 12866 32456
rect 11773 32419 11831 32425
rect 11773 32416 11785 32419
rect 10836 32388 11192 32416
rect 11245 32388 11785 32416
rect 10836 32376 10842 32388
rect 10468 32320 10548 32348
rect 10597 32351 10655 32357
rect 10468 32308 10474 32320
rect 10597 32317 10609 32351
rect 10643 32348 10655 32351
rect 11146 32348 11152 32360
rect 10643 32320 11152 32348
rect 10643 32317 10655 32320
rect 10597 32311 10655 32317
rect 11146 32308 11152 32320
rect 11204 32308 11210 32360
rect 9784 32252 9904 32280
rect 10318 32240 10324 32292
rect 10376 32280 10382 32292
rect 11245 32280 11273 32388
rect 11773 32385 11785 32388
rect 11819 32385 11831 32419
rect 11773 32379 11831 32385
rect 13170 32376 13176 32428
rect 13228 32416 13234 32428
rect 13648 32425 13676 32456
rect 13722 32444 13728 32496
rect 13780 32484 13786 32496
rect 14182 32484 14188 32496
rect 13780 32456 14188 32484
rect 13780 32444 13786 32456
rect 14182 32444 14188 32456
rect 14240 32444 14246 32496
rect 14366 32444 14372 32496
rect 14424 32484 14430 32496
rect 17037 32487 17095 32493
rect 14424 32456 15332 32484
rect 14424 32444 14430 32456
rect 13357 32419 13415 32425
rect 13228 32414 13308 32416
rect 13357 32414 13369 32419
rect 13228 32388 13369 32414
rect 13228 32376 13234 32388
rect 13280 32386 13369 32388
rect 13357 32385 13369 32386
rect 13403 32385 13415 32419
rect 13357 32379 13415 32385
rect 13633 32419 13691 32425
rect 13633 32385 13645 32419
rect 13679 32385 13691 32419
rect 13633 32379 13691 32385
rect 13814 32376 13820 32428
rect 13872 32416 13878 32428
rect 14277 32419 14335 32425
rect 14277 32416 14289 32419
rect 13872 32388 14289 32416
rect 13872 32376 13878 32388
rect 14277 32385 14289 32388
rect 14323 32385 14335 32419
rect 14533 32419 14591 32425
rect 14533 32416 14545 32419
rect 14277 32379 14335 32385
rect 14384 32388 14545 32416
rect 11514 32348 11520 32360
rect 11475 32320 11520 32348
rect 11514 32308 11520 32320
rect 11572 32308 11578 32360
rect 13078 32308 13084 32360
rect 13136 32348 13142 32360
rect 13449 32351 13507 32357
rect 13449 32348 13461 32351
rect 13136 32320 13461 32348
rect 13136 32308 13142 32320
rect 13449 32317 13461 32320
rect 13495 32317 13507 32351
rect 14384 32348 14412 32388
rect 14533 32385 14545 32388
rect 14579 32385 14591 32419
rect 14533 32379 14591 32385
rect 13449 32311 13507 32317
rect 13556 32320 14412 32348
rect 15304 32348 15332 32456
rect 17037 32453 17049 32487
rect 17083 32484 17095 32487
rect 17218 32484 17224 32496
rect 17083 32456 17224 32484
rect 17083 32453 17095 32456
rect 17037 32447 17095 32453
rect 17218 32444 17224 32456
rect 17276 32444 17282 32496
rect 17494 32444 17500 32496
rect 17552 32484 17558 32496
rect 18478 32487 18536 32493
rect 18478 32484 18490 32487
rect 17552 32456 18490 32484
rect 17552 32444 17558 32456
rect 18478 32453 18490 32456
rect 18524 32453 18536 32487
rect 18478 32447 18536 32453
rect 18690 32444 18696 32496
rect 18748 32484 18754 32496
rect 20714 32484 20720 32496
rect 18748 32456 20720 32484
rect 18748 32444 18754 32456
rect 20714 32444 20720 32456
rect 20772 32444 20778 32496
rect 21177 32487 21235 32493
rect 21177 32453 21189 32487
rect 21223 32484 21235 32487
rect 21634 32484 21640 32496
rect 21223 32456 21640 32484
rect 21223 32453 21235 32456
rect 21177 32447 21235 32453
rect 21634 32444 21640 32456
rect 21692 32444 21698 32496
rect 25700 32484 25728 32524
rect 27338 32484 27344 32496
rect 21836 32456 23704 32484
rect 16574 32376 16580 32428
rect 16632 32416 16638 32428
rect 16761 32419 16819 32425
rect 16761 32416 16773 32419
rect 16632 32388 16773 32416
rect 16632 32376 16638 32388
rect 16761 32385 16773 32388
rect 16807 32385 16819 32419
rect 16942 32416 16948 32428
rect 16903 32388 16948 32416
rect 16761 32379 16819 32385
rect 16942 32376 16948 32388
rect 17000 32376 17006 32428
rect 17126 32416 17132 32428
rect 17087 32388 17132 32416
rect 17126 32376 17132 32388
rect 17184 32376 17190 32428
rect 18230 32416 18236 32428
rect 18191 32388 18236 32416
rect 18230 32376 18236 32388
rect 18288 32376 18294 32428
rect 19978 32416 19984 32428
rect 18340 32388 19984 32416
rect 18340 32348 18368 32388
rect 19978 32376 19984 32388
rect 20036 32376 20042 32428
rect 20622 32416 20628 32428
rect 20583 32388 20628 32416
rect 20622 32376 20628 32388
rect 20680 32376 20686 32428
rect 21266 32376 21272 32428
rect 21324 32416 21330 32428
rect 21836 32425 21864 32456
rect 21821 32419 21879 32425
rect 21821 32416 21833 32419
rect 21324 32388 21833 32416
rect 21324 32376 21330 32388
rect 21821 32385 21833 32388
rect 21867 32385 21879 32419
rect 21821 32379 21879 32385
rect 21910 32376 21916 32428
rect 21968 32376 21974 32428
rect 22088 32419 22146 32425
rect 22088 32385 22100 32419
rect 22134 32416 22146 32419
rect 22922 32416 22928 32428
rect 22134 32388 22928 32416
rect 22134 32385 22146 32388
rect 22088 32379 22146 32385
rect 22922 32376 22928 32388
rect 22980 32376 22986 32428
rect 23676 32425 23704 32456
rect 25700 32456 27344 32484
rect 23661 32419 23719 32425
rect 23661 32385 23673 32419
rect 23707 32385 23719 32419
rect 23661 32379 23719 32385
rect 23750 32376 23756 32428
rect 23808 32416 23814 32428
rect 23917 32419 23975 32425
rect 23917 32416 23929 32419
rect 23808 32388 23929 32416
rect 23808 32376 23814 32388
rect 23917 32385 23929 32388
rect 23963 32385 23975 32419
rect 23917 32379 23975 32385
rect 24670 32376 24676 32428
rect 24728 32416 24734 32428
rect 25314 32416 25320 32428
rect 24728 32388 25320 32416
rect 24728 32376 24734 32388
rect 25314 32376 25320 32388
rect 25372 32376 25378 32428
rect 25700 32425 25728 32456
rect 27338 32444 27344 32456
rect 27396 32444 27402 32496
rect 25685 32419 25743 32425
rect 25685 32385 25697 32419
rect 25731 32385 25743 32419
rect 27154 32416 27160 32428
rect 27115 32388 27160 32416
rect 25685 32379 25743 32385
rect 27154 32376 27160 32388
rect 27212 32376 27218 32428
rect 27982 32416 27988 32428
rect 27943 32388 27988 32416
rect 27982 32376 27988 32388
rect 28040 32376 28046 32428
rect 15304 32320 18368 32348
rect 10376 32252 11273 32280
rect 10376 32240 10382 32252
rect 12526 32240 12532 32292
rect 12584 32280 12590 32292
rect 13556 32280 13584 32320
rect 19242 32308 19248 32360
rect 19300 32348 19306 32360
rect 21928 32348 21956 32376
rect 19300 32320 21956 32348
rect 19300 32308 19306 32320
rect 25222 32308 25228 32360
rect 25280 32348 25286 32360
rect 25590 32348 25596 32360
rect 25280 32320 25596 32348
rect 25280 32308 25286 32320
rect 25590 32308 25596 32320
rect 25648 32308 25654 32360
rect 27246 32348 27252 32360
rect 27207 32320 27252 32348
rect 27246 32308 27252 32320
rect 27304 32308 27310 32360
rect 12584 32252 13584 32280
rect 12584 32240 12590 32252
rect 13722 32240 13728 32292
rect 13780 32280 13786 32292
rect 14274 32280 14280 32292
rect 13780 32252 14280 32280
rect 13780 32240 13786 32252
rect 14274 32240 14280 32252
rect 14332 32240 14338 32292
rect 16206 32280 16212 32292
rect 15212 32252 16212 32280
rect 7331 32184 9076 32212
rect 7331 32181 7343 32184
rect 7285 32175 7343 32181
rect 9122 32172 9128 32224
rect 9180 32212 9186 32224
rect 9217 32215 9275 32221
rect 9217 32212 9229 32215
rect 9180 32184 9229 32212
rect 9180 32172 9186 32184
rect 9217 32181 9229 32184
rect 9263 32181 9275 32215
rect 9217 32175 9275 32181
rect 9306 32172 9312 32224
rect 9364 32212 9370 32224
rect 10965 32215 11023 32221
rect 10965 32212 10977 32215
rect 9364 32184 10977 32212
rect 9364 32172 9370 32184
rect 10965 32181 10977 32184
rect 11011 32181 11023 32215
rect 10965 32175 11023 32181
rect 11054 32172 11060 32224
rect 11112 32212 11118 32224
rect 12710 32212 12716 32224
rect 11112 32184 12716 32212
rect 11112 32172 11118 32184
rect 12710 32172 12716 32184
rect 12768 32172 12774 32224
rect 12802 32172 12808 32224
rect 12860 32212 12866 32224
rect 12897 32215 12955 32221
rect 12897 32212 12909 32215
rect 12860 32184 12909 32212
rect 12860 32172 12866 32184
rect 12897 32181 12909 32184
rect 12943 32181 12955 32215
rect 13446 32212 13452 32224
rect 13407 32184 13452 32212
rect 12897 32175 12955 32181
rect 13446 32172 13452 32184
rect 13504 32172 13510 32224
rect 13814 32212 13820 32224
rect 13775 32184 13820 32212
rect 13814 32172 13820 32184
rect 13872 32172 13878 32224
rect 13998 32172 14004 32224
rect 14056 32212 14062 32224
rect 15212 32212 15240 32252
rect 16206 32240 16212 32252
rect 16264 32240 16270 32292
rect 23201 32283 23259 32289
rect 16546 32252 18276 32280
rect 14056 32184 15240 32212
rect 14056 32172 14062 32184
rect 15286 32172 15292 32224
rect 15344 32212 15350 32224
rect 15657 32215 15715 32221
rect 15657 32212 15669 32215
rect 15344 32184 15669 32212
rect 15344 32172 15350 32184
rect 15657 32181 15669 32184
rect 15703 32181 15715 32215
rect 15657 32175 15715 32181
rect 15930 32172 15936 32224
rect 15988 32212 15994 32224
rect 16546 32212 16574 32252
rect 15988 32184 16574 32212
rect 15988 32172 15994 32184
rect 17034 32172 17040 32224
rect 17092 32212 17098 32224
rect 17313 32215 17371 32221
rect 17313 32212 17325 32215
rect 17092 32184 17325 32212
rect 17092 32172 17098 32184
rect 17313 32181 17325 32184
rect 17359 32181 17371 32215
rect 18248 32212 18276 32252
rect 19306 32252 21036 32280
rect 19306 32212 19334 32252
rect 18248 32184 19334 32212
rect 19613 32215 19671 32221
rect 17313 32175 17371 32181
rect 19613 32181 19625 32215
rect 19659 32212 19671 32215
rect 19978 32212 19984 32224
rect 19659 32184 19984 32212
rect 19659 32181 19671 32184
rect 19613 32175 19671 32181
rect 19978 32172 19984 32184
rect 20036 32172 20042 32224
rect 21008 32212 21036 32252
rect 23201 32249 23213 32283
rect 23247 32280 23259 32283
rect 23474 32280 23480 32292
rect 23247 32252 23480 32280
rect 23247 32249 23259 32252
rect 23201 32243 23259 32249
rect 23474 32240 23480 32252
rect 23532 32240 23538 32292
rect 24670 32240 24676 32292
rect 24728 32280 24734 32292
rect 24854 32280 24860 32292
rect 24728 32252 24860 32280
rect 24728 32240 24734 32252
rect 24854 32240 24860 32252
rect 24912 32240 24918 32292
rect 25041 32283 25099 32289
rect 25041 32249 25053 32283
rect 25087 32280 25099 32283
rect 25130 32280 25136 32292
rect 25087 32252 25136 32280
rect 25087 32249 25099 32252
rect 25041 32243 25099 32249
rect 25130 32240 25136 32252
rect 25188 32240 25194 32292
rect 24946 32212 24952 32224
rect 21008 32184 24952 32212
rect 24946 32172 24952 32184
rect 25004 32172 25010 32224
rect 25958 32212 25964 32224
rect 25919 32184 25964 32212
rect 25958 32172 25964 32184
rect 26016 32172 26022 32224
rect 26050 32172 26056 32224
rect 26108 32212 26114 32224
rect 27433 32215 27491 32221
rect 27433 32212 27445 32215
rect 26108 32184 27445 32212
rect 26108 32172 26114 32184
rect 27433 32181 27445 32184
rect 27479 32181 27491 32215
rect 27433 32175 27491 32181
rect 27522 32172 27528 32224
rect 27580 32212 27586 32224
rect 28077 32215 28135 32221
rect 28077 32212 28089 32215
rect 27580 32184 28089 32212
rect 27580 32172 27586 32184
rect 28077 32181 28089 32184
rect 28123 32181 28135 32215
rect 28077 32175 28135 32181
rect 1104 32122 28888 32144
rect 1104 32070 5582 32122
rect 5634 32070 5646 32122
rect 5698 32070 5710 32122
rect 5762 32070 5774 32122
rect 5826 32070 5838 32122
rect 5890 32070 14846 32122
rect 14898 32070 14910 32122
rect 14962 32070 14974 32122
rect 15026 32070 15038 32122
rect 15090 32070 15102 32122
rect 15154 32070 24110 32122
rect 24162 32070 24174 32122
rect 24226 32070 24238 32122
rect 24290 32070 24302 32122
rect 24354 32070 24366 32122
rect 24418 32070 28888 32122
rect 1104 32048 28888 32070
rect 1486 31968 1492 32020
rect 1544 32008 1550 32020
rect 1765 32011 1823 32017
rect 1765 32008 1777 32011
rect 1544 31980 1777 32008
rect 1544 31968 1550 31980
rect 1765 31977 1777 31980
rect 1811 31977 1823 32011
rect 1765 31971 1823 31977
rect 7561 32011 7619 32017
rect 7561 31977 7573 32011
rect 7607 32008 7619 32011
rect 10226 32008 10232 32020
rect 7607 31980 10232 32008
rect 7607 31977 7619 31980
rect 7561 31971 7619 31977
rect 10226 31968 10232 31980
rect 10284 31968 10290 32020
rect 10318 31968 10324 32020
rect 10376 32008 10382 32020
rect 10962 32008 10968 32020
rect 10376 31980 10968 32008
rect 10376 31968 10382 31980
rect 10962 31968 10968 31980
rect 11020 31968 11026 32020
rect 11514 31968 11520 32020
rect 11572 32008 11578 32020
rect 13814 32008 13820 32020
rect 11572 31980 13820 32008
rect 11572 31968 11578 31980
rect 13814 31968 13820 31980
rect 13872 31968 13878 32020
rect 13924 31980 15056 32008
rect 9398 31940 9404 31952
rect 6932 31912 9404 31940
rect 1670 31764 1676 31816
rect 1728 31804 1734 31816
rect 2409 31807 2467 31813
rect 2409 31804 2421 31807
rect 1728 31776 2421 31804
rect 1728 31764 1734 31776
rect 2409 31773 2421 31776
rect 2455 31773 2467 31807
rect 6270 31804 6276 31816
rect 6231 31776 6276 31804
rect 2409 31767 2467 31773
rect 6270 31764 6276 31776
rect 6328 31764 6334 31816
rect 6932 31813 6960 31912
rect 9398 31900 9404 31912
rect 9456 31900 9462 31952
rect 9493 31943 9551 31949
rect 9493 31909 9505 31943
rect 9539 31940 9551 31943
rect 11698 31940 11704 31952
rect 9539 31912 11704 31940
rect 9539 31909 9551 31912
rect 9493 31903 9551 31909
rect 11698 31900 11704 31912
rect 11756 31900 11762 31952
rect 12710 31900 12716 31952
rect 12768 31940 12774 31952
rect 13538 31940 13544 31952
rect 12768 31912 13544 31940
rect 12768 31900 12774 31912
rect 13538 31900 13544 31912
rect 13596 31900 13602 31952
rect 9306 31872 9312 31884
rect 7760 31844 9312 31872
rect 7760 31813 7788 31844
rect 9306 31832 9312 31844
rect 9364 31832 9370 31884
rect 10045 31875 10103 31881
rect 10045 31841 10057 31875
rect 10091 31872 10103 31875
rect 13722 31872 13728 31884
rect 10091 31844 11836 31872
rect 10091 31841 10103 31844
rect 10045 31835 10103 31841
rect 6917 31807 6975 31813
rect 6917 31773 6929 31807
rect 6963 31773 6975 31807
rect 6917 31767 6975 31773
rect 7745 31807 7803 31813
rect 7745 31773 7757 31807
rect 7791 31773 7803 31807
rect 7745 31767 7803 31773
rect 7926 31764 7932 31816
rect 7984 31804 7990 31816
rect 8205 31807 8263 31813
rect 8205 31804 8217 31807
rect 7984 31776 8217 31804
rect 7984 31764 7990 31776
rect 8205 31773 8217 31776
rect 8251 31773 8263 31807
rect 8205 31767 8263 31773
rect 8389 31807 8447 31813
rect 8389 31773 8401 31807
rect 8435 31804 8447 31807
rect 9398 31804 9404 31816
rect 8435 31776 9404 31804
rect 8435 31773 8447 31776
rect 8389 31767 8447 31773
rect 9398 31764 9404 31776
rect 9456 31764 9462 31816
rect 9582 31764 9588 31816
rect 9640 31804 9646 31816
rect 10134 31804 10140 31816
rect 9640 31776 10140 31804
rect 9640 31764 9646 31776
rect 10134 31764 10140 31776
rect 10192 31804 10198 31816
rect 10229 31807 10287 31813
rect 10229 31804 10241 31807
rect 10192 31776 10241 31804
rect 10192 31764 10198 31776
rect 10229 31773 10241 31776
rect 10275 31773 10287 31807
rect 10229 31767 10287 31773
rect 10318 31764 10324 31816
rect 10376 31804 10382 31816
rect 11057 31807 11115 31813
rect 10376 31776 11008 31804
rect 10376 31764 10382 31776
rect 2222 31696 2228 31748
rect 2280 31736 2286 31748
rect 8297 31739 8355 31745
rect 2280 31708 6868 31736
rect 2280 31696 2286 31708
rect 6730 31668 6736 31680
rect 6691 31640 6736 31668
rect 6730 31628 6736 31640
rect 6788 31628 6794 31680
rect 6840 31668 6868 31708
rect 8297 31705 8309 31739
rect 8343 31736 8355 31739
rect 9122 31736 9128 31748
rect 8343 31708 9128 31736
rect 8343 31705 8355 31708
rect 8297 31699 8355 31705
rect 9122 31696 9128 31708
rect 9180 31696 9186 31748
rect 9306 31696 9312 31748
rect 9364 31736 9370 31748
rect 9950 31736 9956 31748
rect 9364 31708 9956 31736
rect 9364 31696 9370 31708
rect 9950 31696 9956 31708
rect 10008 31696 10014 31748
rect 10042 31696 10048 31748
rect 10100 31736 10106 31748
rect 10778 31736 10784 31748
rect 10100 31708 10784 31736
rect 10100 31696 10106 31708
rect 10778 31696 10784 31708
rect 10836 31696 10842 31748
rect 10873 31739 10931 31745
rect 10873 31705 10885 31739
rect 10919 31705 10931 31739
rect 10980 31736 11008 31776
rect 11057 31773 11069 31807
rect 11103 31804 11115 31807
rect 11514 31804 11520 31816
rect 11103 31776 11520 31804
rect 11103 31773 11115 31776
rect 11057 31767 11115 31773
rect 11514 31764 11520 31776
rect 11572 31764 11578 31816
rect 11698 31804 11704 31816
rect 11659 31776 11704 31804
rect 11698 31764 11704 31776
rect 11756 31764 11762 31816
rect 11808 31804 11836 31844
rect 12728 31844 13728 31872
rect 12728 31804 12756 31844
rect 13722 31832 13728 31844
rect 13780 31832 13786 31884
rect 11808 31776 12756 31804
rect 12894 31764 12900 31816
rect 12952 31804 12958 31816
rect 13924 31804 13952 31980
rect 14090 31900 14096 31952
rect 14148 31900 14154 31952
rect 15028 31940 15056 31980
rect 15194 31968 15200 32020
rect 15252 32008 15258 32020
rect 15473 32011 15531 32017
rect 15473 32008 15485 32011
rect 15252 31980 15485 32008
rect 15252 31968 15258 31980
rect 15473 31977 15485 31980
rect 15519 31977 15531 32011
rect 18509 32011 18567 32017
rect 15473 31971 15531 31977
rect 15580 31980 17172 32008
rect 15580 31940 15608 31980
rect 15028 31912 15608 31940
rect 17144 31940 17172 31980
rect 18509 31977 18521 32011
rect 18555 32008 18567 32011
rect 18598 32008 18604 32020
rect 18555 31980 18604 32008
rect 18555 31977 18567 31980
rect 18509 31971 18567 31977
rect 18598 31968 18604 31980
rect 18656 31968 18662 32020
rect 19702 31968 19708 32020
rect 19760 32008 19766 32020
rect 20254 32008 20260 32020
rect 19760 31980 20260 32008
rect 19760 31968 19766 31980
rect 20254 31968 20260 31980
rect 20312 31968 20318 32020
rect 20349 32011 20407 32017
rect 20349 31977 20361 32011
rect 20395 32008 20407 32011
rect 20438 32008 20444 32020
rect 20395 31980 20444 32008
rect 20395 31977 20407 31980
rect 20349 31971 20407 31977
rect 20438 31968 20444 31980
rect 20496 31968 20502 32020
rect 22833 32011 22891 32017
rect 22833 31977 22845 32011
rect 22879 32008 22891 32011
rect 23106 32008 23112 32020
rect 22879 31980 23112 32008
rect 22879 31977 22891 31980
rect 22833 31971 22891 31977
rect 23106 31968 23112 31980
rect 23164 31968 23170 32020
rect 23474 32008 23480 32020
rect 23435 31980 23480 32008
rect 23474 31968 23480 31980
rect 23532 31968 23538 32020
rect 25958 32008 25964 32020
rect 23584 31980 25964 32008
rect 23584 31940 23612 31980
rect 25958 31968 25964 31980
rect 26016 31968 26022 32020
rect 17144 31912 23612 31940
rect 14108 31872 14136 31900
rect 14108 31844 14228 31872
rect 14090 31804 14096 31816
rect 12952 31776 13952 31804
rect 14051 31776 14096 31804
rect 12952 31764 12958 31776
rect 14090 31764 14096 31776
rect 14148 31764 14154 31816
rect 14200 31804 14228 31844
rect 15654 31832 15660 31884
rect 15712 31872 15718 31884
rect 16209 31875 16267 31881
rect 16209 31872 16221 31875
rect 15712 31844 16221 31872
rect 15712 31832 15718 31844
rect 16209 31841 16221 31844
rect 16255 31841 16267 31875
rect 16209 31835 16267 31841
rect 17310 31832 17316 31884
rect 17368 31872 17374 31884
rect 19518 31872 19524 31884
rect 17368 31844 19524 31872
rect 17368 31832 17374 31844
rect 19518 31832 19524 31844
rect 19576 31832 19582 31884
rect 19886 31832 19892 31884
rect 19944 31872 19950 31884
rect 19944 31844 20208 31872
rect 19944 31832 19950 31844
rect 14349 31807 14407 31813
rect 14349 31804 14361 31807
rect 14200 31776 14361 31804
rect 14349 31773 14361 31776
rect 14395 31773 14407 31807
rect 14349 31767 14407 31773
rect 14734 31764 14740 31816
rect 14792 31804 14798 31816
rect 15672 31804 15700 31832
rect 14792 31776 15700 31804
rect 16316 31776 16703 31804
rect 14792 31764 14798 31776
rect 11946 31739 12004 31745
rect 11946 31736 11958 31739
rect 10980 31708 11958 31736
rect 10873 31699 10931 31705
rect 11946 31705 11958 31708
rect 11992 31705 12004 31739
rect 14550 31736 14556 31748
rect 11946 31699 12004 31705
rect 12268 31708 14556 31736
rect 8386 31668 8392 31680
rect 6840 31640 8392 31668
rect 8386 31628 8392 31640
rect 8444 31628 8450 31680
rect 9674 31628 9680 31680
rect 9732 31668 9738 31680
rect 10413 31671 10471 31677
rect 10413 31668 10425 31671
rect 9732 31640 10425 31668
rect 9732 31628 9738 31640
rect 10413 31637 10425 31640
rect 10459 31637 10471 31671
rect 10888 31668 10916 31699
rect 11146 31668 11152 31680
rect 10888 31640 11152 31668
rect 10413 31631 10471 31637
rect 11146 31628 11152 31640
rect 11204 31628 11210 31680
rect 11241 31671 11299 31677
rect 11241 31637 11253 31671
rect 11287 31668 11299 31671
rect 12268 31668 12296 31708
rect 14550 31696 14556 31708
rect 14608 31696 14614 31748
rect 14826 31696 14832 31748
rect 14884 31736 14890 31748
rect 16316 31736 16344 31776
rect 16482 31745 16488 31748
rect 14884 31708 16344 31736
rect 14884 31696 14890 31708
rect 16476 31699 16488 31745
rect 16540 31736 16546 31748
rect 16675 31736 16703 31776
rect 17494 31764 17500 31816
rect 17552 31804 17558 31816
rect 19702 31804 19708 31816
rect 17552 31776 19708 31804
rect 17552 31764 17558 31776
rect 19702 31764 19708 31776
rect 19760 31764 19766 31816
rect 20070 31804 20076 31816
rect 20031 31776 20076 31804
rect 20070 31764 20076 31776
rect 20128 31764 20134 31816
rect 20180 31813 20208 31844
rect 20254 31832 20260 31884
rect 20312 31872 20318 31884
rect 26326 31872 26332 31884
rect 20312 31844 24072 31872
rect 26287 31844 26332 31872
rect 20312 31832 20318 31844
rect 20165 31807 20223 31813
rect 20165 31773 20177 31807
rect 20211 31773 20223 31807
rect 20806 31804 20812 31816
rect 20767 31776 20812 31804
rect 20165 31767 20223 31773
rect 20806 31764 20812 31776
rect 20864 31804 20870 31816
rect 21729 31807 21787 31813
rect 21729 31804 21741 31807
rect 20864 31776 21741 31804
rect 20864 31764 20870 31776
rect 21729 31773 21741 31776
rect 21775 31773 21787 31807
rect 21729 31767 21787 31773
rect 22554 31764 22560 31816
rect 22612 31804 22618 31816
rect 23106 31804 23112 31816
rect 22612 31776 23112 31804
rect 22612 31764 22618 31776
rect 23106 31764 23112 31776
rect 23164 31764 23170 31816
rect 23382 31804 23388 31816
rect 23343 31776 23388 31804
rect 23382 31764 23388 31776
rect 23440 31764 23446 31816
rect 17402 31736 17408 31748
rect 16540 31708 16576 31736
rect 16675 31708 17408 31736
rect 16482 31696 16488 31699
rect 16540 31696 16546 31708
rect 17402 31696 17408 31708
rect 17460 31736 17466 31748
rect 18230 31736 18236 31748
rect 17460 31708 18236 31736
rect 17460 31696 17466 31708
rect 18230 31696 18236 31708
rect 18288 31696 18294 31748
rect 18325 31739 18383 31745
rect 18325 31705 18337 31739
rect 18371 31736 18383 31739
rect 18371 31708 19288 31736
rect 18371 31705 18383 31708
rect 18325 31699 18383 31705
rect 11287 31640 12296 31668
rect 11287 31637 11299 31640
rect 11241 31631 11299 31637
rect 12342 31628 12348 31680
rect 12400 31668 12406 31680
rect 13081 31671 13139 31677
rect 13081 31668 13093 31671
rect 12400 31640 13093 31668
rect 12400 31628 12406 31640
rect 13081 31637 13093 31640
rect 13127 31668 13139 31671
rect 13170 31668 13176 31680
rect 13127 31640 13176 31668
rect 13127 31637 13139 31640
rect 13081 31631 13139 31637
rect 13170 31628 13176 31640
rect 13228 31628 13234 31680
rect 13906 31628 13912 31680
rect 13964 31668 13970 31680
rect 16298 31668 16304 31680
rect 13964 31640 16304 31668
rect 13964 31628 13970 31640
rect 16298 31628 16304 31640
rect 16356 31628 16362 31680
rect 16758 31628 16764 31680
rect 16816 31668 16822 31680
rect 17218 31668 17224 31680
rect 16816 31640 17224 31668
rect 16816 31628 16822 31640
rect 17218 31628 17224 31640
rect 17276 31668 17282 31680
rect 17589 31671 17647 31677
rect 17589 31668 17601 31671
rect 17276 31640 17601 31668
rect 17276 31628 17282 31640
rect 17589 31637 17601 31640
rect 17635 31637 17647 31671
rect 17589 31631 17647 31637
rect 18506 31628 18512 31680
rect 18564 31677 18570 31680
rect 18564 31671 18583 31677
rect 18571 31637 18583 31671
rect 18690 31668 18696 31680
rect 18651 31640 18696 31668
rect 18564 31631 18583 31637
rect 18564 31628 18570 31631
rect 18690 31628 18696 31640
rect 18748 31628 18754 31680
rect 19260 31668 19288 31708
rect 19334 31696 19340 31748
rect 19392 31736 19398 31748
rect 19797 31739 19855 31745
rect 19797 31736 19809 31739
rect 19392 31708 19809 31736
rect 19392 31696 19398 31708
rect 19797 31705 19809 31708
rect 19843 31705 19855 31739
rect 19978 31736 19984 31748
rect 19939 31708 19984 31736
rect 19797 31699 19855 31705
rect 19978 31696 19984 31708
rect 20036 31696 20042 31748
rect 20990 31696 20996 31748
rect 21048 31736 21054 31748
rect 21085 31739 21143 31745
rect 21085 31736 21097 31739
rect 21048 31708 21097 31736
rect 21048 31696 21054 31708
rect 21085 31705 21097 31708
rect 21131 31705 21143 31739
rect 21085 31699 21143 31705
rect 21910 31696 21916 31748
rect 21968 31736 21974 31748
rect 22005 31739 22063 31745
rect 22005 31736 22017 31739
rect 21968 31708 22017 31736
rect 21968 31696 21974 31708
rect 22005 31705 22017 31708
rect 22051 31705 22063 31739
rect 22005 31699 22063 31705
rect 22741 31739 22799 31745
rect 22741 31705 22753 31739
rect 22787 31705 22799 31739
rect 22741 31699 22799 31705
rect 20346 31668 20352 31680
rect 19260 31640 20352 31668
rect 20346 31628 20352 31640
rect 20404 31628 20410 31680
rect 20806 31628 20812 31680
rect 20864 31668 20870 31680
rect 22756 31668 22784 31699
rect 22922 31696 22928 31748
rect 22980 31736 22986 31748
rect 23400 31736 23428 31764
rect 22980 31708 23428 31736
rect 22980 31696 22986 31708
rect 23474 31696 23480 31748
rect 23532 31736 23538 31748
rect 24044 31736 24072 31844
rect 26326 31832 26332 31844
rect 26384 31832 26390 31884
rect 28166 31872 28172 31884
rect 28127 31844 28172 31872
rect 28166 31832 28172 31844
rect 28224 31832 28230 31884
rect 24486 31804 24492 31816
rect 24447 31776 24492 31804
rect 24486 31764 24492 31776
rect 24544 31764 24550 31816
rect 24578 31764 24584 31816
rect 24636 31804 24642 31816
rect 24745 31807 24803 31813
rect 24745 31804 24757 31807
rect 24636 31776 24757 31804
rect 24636 31764 24642 31776
rect 24745 31773 24757 31776
rect 24791 31773 24803 31807
rect 24745 31767 24803 31773
rect 26513 31739 26571 31745
rect 26513 31736 26525 31739
rect 23532 31708 23980 31736
rect 24044 31708 26525 31736
rect 23532 31696 23538 31708
rect 23842 31668 23848 31680
rect 20864 31640 22784 31668
rect 23803 31640 23848 31668
rect 20864 31628 20870 31640
rect 23842 31628 23848 31640
rect 23900 31628 23906 31680
rect 23952 31668 23980 31708
rect 26513 31705 26525 31708
rect 26559 31705 26571 31739
rect 26513 31699 26571 31705
rect 24854 31668 24860 31680
rect 23952 31640 24860 31668
rect 24854 31628 24860 31640
rect 24912 31628 24918 31680
rect 25314 31628 25320 31680
rect 25372 31668 25378 31680
rect 25869 31671 25927 31677
rect 25869 31668 25881 31671
rect 25372 31640 25881 31668
rect 25372 31628 25378 31640
rect 25869 31637 25881 31640
rect 25915 31637 25927 31671
rect 25869 31631 25927 31637
rect 1104 31578 28888 31600
rect 1104 31526 10214 31578
rect 10266 31526 10278 31578
rect 10330 31526 10342 31578
rect 10394 31526 10406 31578
rect 10458 31526 10470 31578
rect 10522 31526 19478 31578
rect 19530 31526 19542 31578
rect 19594 31526 19606 31578
rect 19658 31526 19670 31578
rect 19722 31526 19734 31578
rect 19786 31526 28888 31578
rect 1104 31504 28888 31526
rect 7837 31467 7895 31473
rect 7837 31433 7849 31467
rect 7883 31464 7895 31467
rect 9950 31464 9956 31476
rect 7883 31436 9956 31464
rect 7883 31433 7895 31436
rect 7837 31427 7895 31433
rect 9950 31424 9956 31436
rect 10008 31424 10014 31476
rect 10042 31424 10048 31476
rect 10100 31464 10106 31476
rect 10137 31467 10195 31473
rect 10137 31464 10149 31467
rect 10100 31436 10149 31464
rect 10100 31424 10106 31436
rect 10137 31433 10149 31436
rect 10183 31433 10195 31467
rect 14277 31467 14335 31473
rect 14277 31464 14289 31467
rect 10137 31427 10195 31433
rect 10244 31436 14289 31464
rect 10244 31408 10272 31436
rect 14277 31433 14289 31436
rect 14323 31433 14335 31467
rect 14277 31427 14335 31433
rect 14458 31424 14464 31476
rect 14516 31464 14522 31476
rect 14516 31436 15148 31464
rect 14516 31424 14522 31436
rect 9674 31396 9680 31408
rect 6748 31368 9680 31396
rect 1670 31328 1676 31340
rect 1631 31300 1676 31328
rect 1670 31288 1676 31300
rect 1728 31288 1734 31340
rect 6748 31337 6776 31368
rect 9674 31356 9680 31368
rect 9732 31356 9738 31408
rect 9876 31368 10180 31396
rect 6733 31331 6791 31337
rect 6733 31297 6745 31331
rect 6779 31297 6791 31331
rect 6733 31291 6791 31297
rect 7377 31331 7435 31337
rect 7377 31297 7389 31331
rect 7423 31297 7435 31331
rect 7377 31291 7435 31297
rect 8021 31331 8079 31337
rect 8021 31297 8033 31331
rect 8067 31328 8079 31331
rect 8294 31328 8300 31340
rect 8067 31300 8300 31328
rect 8067 31297 8079 31300
rect 8021 31291 8079 31297
rect 1857 31263 1915 31269
rect 1857 31229 1869 31263
rect 1903 31260 1915 31263
rect 2314 31260 2320 31272
rect 1903 31232 2320 31260
rect 1903 31229 1915 31232
rect 1857 31223 1915 31229
rect 2314 31220 2320 31232
rect 2372 31220 2378 31272
rect 2774 31220 2780 31272
rect 2832 31260 2838 31272
rect 7392 31260 7420 31291
rect 8294 31288 8300 31300
rect 8352 31288 8358 31340
rect 8481 31331 8539 31337
rect 8481 31297 8493 31331
rect 8527 31328 8539 31331
rect 8938 31328 8944 31340
rect 8527 31300 8944 31328
rect 8527 31297 8539 31300
rect 8481 31291 8539 31297
rect 8938 31288 8944 31300
rect 8996 31288 9002 31340
rect 9122 31328 9128 31340
rect 9083 31300 9128 31328
rect 9122 31288 9128 31300
rect 9180 31288 9186 31340
rect 9876 31337 9904 31368
rect 9861 31331 9919 31337
rect 9861 31297 9873 31331
rect 9907 31297 9919 31331
rect 9861 31291 9919 31297
rect 9953 31331 10011 31337
rect 9953 31297 9965 31331
rect 9999 31297 10011 31331
rect 10152 31328 10180 31368
rect 10226 31356 10232 31408
rect 10284 31356 10290 31408
rect 12250 31396 12256 31408
rect 10612 31368 12256 31396
rect 10612 31328 10640 31368
rect 12250 31356 12256 31368
rect 12308 31356 12314 31408
rect 12342 31356 12348 31408
rect 12400 31396 12406 31408
rect 12400 31368 13676 31396
rect 12400 31356 12406 31368
rect 10152 31300 10640 31328
rect 9953 31291 10011 31297
rect 8202 31260 8208 31272
rect 2832 31232 2877 31260
rect 7392 31232 8208 31260
rect 2832 31220 2838 31232
rect 8202 31220 8208 31232
rect 8260 31220 8266 31272
rect 9582 31260 9588 31272
rect 8404 31232 9588 31260
rect 6549 31195 6607 31201
rect 6549 31161 6561 31195
rect 6595 31192 6607 31195
rect 8110 31192 8116 31204
rect 6595 31164 8116 31192
rect 6595 31161 6607 31164
rect 6549 31155 6607 31161
rect 8110 31152 8116 31164
rect 8168 31152 8174 31204
rect 7193 31127 7251 31133
rect 7193 31093 7205 31127
rect 7239 31124 7251 31127
rect 8404 31124 8432 31232
rect 9582 31220 9588 31232
rect 9640 31260 9646 31272
rect 9968 31260 9996 31291
rect 10686 31288 10692 31340
rect 10744 31328 10750 31340
rect 10781 31331 10839 31337
rect 10781 31328 10793 31331
rect 10744 31300 10793 31328
rect 10744 31288 10750 31300
rect 10781 31297 10793 31300
rect 10827 31297 10839 31331
rect 10781 31291 10839 31297
rect 10962 31288 10968 31340
rect 11020 31328 11026 31340
rect 11609 31331 11667 31337
rect 11609 31328 11621 31331
rect 11020 31300 11621 31328
rect 11020 31288 11026 31300
rect 11609 31297 11621 31300
rect 11655 31297 11667 31331
rect 11609 31291 11667 31297
rect 11698 31288 11704 31340
rect 11756 31328 11762 31340
rect 11793 31331 11851 31337
rect 11793 31328 11805 31331
rect 11756 31300 11805 31328
rect 11756 31288 11762 31300
rect 11793 31297 11805 31300
rect 11839 31328 11851 31331
rect 12066 31328 12072 31340
rect 11839 31300 12072 31328
rect 11839 31297 11851 31300
rect 11793 31291 11851 31297
rect 12066 31288 12072 31300
rect 12124 31288 12130 31340
rect 12437 31331 12495 31337
rect 12437 31297 12449 31331
rect 12483 31328 12495 31331
rect 13170 31328 13176 31340
rect 12483 31300 13176 31328
rect 12483 31297 12495 31300
rect 12437 31291 12495 31297
rect 13170 31288 13176 31300
rect 13228 31328 13234 31340
rect 13265 31331 13323 31337
rect 13265 31328 13277 31331
rect 13228 31300 13277 31328
rect 13228 31288 13234 31300
rect 13265 31297 13277 31300
rect 13311 31297 13323 31331
rect 13446 31328 13452 31340
rect 13407 31300 13452 31328
rect 13265 31291 13323 31297
rect 13446 31288 13452 31300
rect 13504 31288 13510 31340
rect 13648 31328 13676 31368
rect 13722 31356 13728 31408
rect 13780 31396 13786 31408
rect 14982 31399 15040 31405
rect 14982 31396 14994 31399
rect 13780 31368 14994 31396
rect 13780 31356 13786 31368
rect 14982 31365 14994 31368
rect 15028 31365 15040 31399
rect 15120 31396 15148 31436
rect 15194 31424 15200 31476
rect 15252 31464 15258 31476
rect 15252 31436 17080 31464
rect 15252 31424 15258 31436
rect 15120 31368 16436 31396
rect 14982 31359 15040 31365
rect 14093 31331 14151 31337
rect 14093 31328 14105 31331
rect 13648 31300 14105 31328
rect 14093 31297 14105 31300
rect 14139 31328 14151 31331
rect 14366 31328 14372 31340
rect 14139 31300 14372 31328
rect 14139 31297 14151 31300
rect 14093 31291 14151 31297
rect 14366 31288 14372 31300
rect 14424 31288 14430 31340
rect 14734 31328 14740 31340
rect 14695 31300 14740 31328
rect 14734 31288 14740 31300
rect 14792 31288 14798 31340
rect 15838 31328 15844 31340
rect 14844 31300 15844 31328
rect 9640 31232 9996 31260
rect 9640 31220 9646 31232
rect 10042 31220 10048 31272
rect 10100 31260 10106 31272
rect 10410 31260 10416 31272
rect 10100 31232 10416 31260
rect 10100 31220 10106 31232
rect 10410 31220 10416 31232
rect 10468 31220 10474 31272
rect 10597 31263 10655 31269
rect 10597 31229 10609 31263
rect 10643 31260 10655 31263
rect 12158 31260 12164 31272
rect 10643 31232 12164 31260
rect 10643 31229 10655 31232
rect 10597 31223 10655 31229
rect 12158 31220 12164 31232
rect 12216 31220 12222 31272
rect 12253 31263 12311 31269
rect 12253 31229 12265 31263
rect 12299 31260 12311 31263
rect 12802 31260 12808 31272
rect 12299 31232 12808 31260
rect 12299 31229 12311 31232
rect 12253 31223 12311 31229
rect 12802 31220 12808 31232
rect 12860 31220 12866 31272
rect 13081 31263 13139 31269
rect 13081 31229 13093 31263
rect 13127 31260 13139 31263
rect 13127 31232 13860 31260
rect 13127 31229 13139 31232
rect 13081 31223 13139 31229
rect 9217 31195 9275 31201
rect 9217 31161 9229 31195
rect 9263 31192 9275 31195
rect 10318 31192 10324 31204
rect 9263 31164 10324 31192
rect 9263 31161 9275 31164
rect 9217 31155 9275 31161
rect 10318 31152 10324 31164
rect 10376 31152 10382 31204
rect 10502 31152 10508 31204
rect 10560 31192 10566 31204
rect 13832 31192 13860 31232
rect 13906 31220 13912 31272
rect 13964 31260 13970 31272
rect 13964 31232 14009 31260
rect 13964 31220 13970 31232
rect 14182 31220 14188 31272
rect 14240 31260 14246 31272
rect 14458 31260 14464 31272
rect 14240 31232 14464 31260
rect 14240 31220 14246 31232
rect 14458 31220 14464 31232
rect 14516 31220 14522 31272
rect 14844 31260 14872 31300
rect 15838 31288 15844 31300
rect 15896 31288 15902 31340
rect 14752 31232 14872 31260
rect 16408 31260 16436 31368
rect 16574 31356 16580 31408
rect 16632 31396 16638 31408
rect 17052 31396 17080 31436
rect 20070 31424 20076 31476
rect 20128 31464 20134 31476
rect 21269 31467 21327 31473
rect 21269 31464 21281 31467
rect 20128 31436 21281 31464
rect 20128 31424 20134 31436
rect 21269 31433 21281 31436
rect 21315 31433 21327 31467
rect 21269 31427 21327 31433
rect 22278 31424 22284 31476
rect 22336 31464 22342 31476
rect 22336 31436 23336 31464
rect 22336 31424 22342 31436
rect 17926 31399 17984 31405
rect 17926 31396 17938 31399
rect 16632 31368 16988 31396
rect 17052 31368 17938 31396
rect 16632 31356 16638 31368
rect 16482 31288 16488 31340
rect 16540 31328 16546 31340
rect 16960 31337 16988 31368
rect 17926 31365 17938 31368
rect 17972 31365 17984 31399
rect 17926 31359 17984 31365
rect 21913 31399 21971 31405
rect 21913 31365 21925 31399
rect 21959 31396 21971 31399
rect 22922 31396 22928 31408
rect 21959 31368 22928 31396
rect 21959 31365 21971 31368
rect 21913 31359 21971 31365
rect 22922 31356 22928 31368
rect 22980 31356 22986 31408
rect 23198 31396 23204 31408
rect 23032 31368 23204 31396
rect 16669 31331 16727 31337
rect 16669 31328 16681 31331
rect 16540 31300 16681 31328
rect 16540 31288 16546 31300
rect 16669 31297 16681 31300
rect 16715 31297 16727 31331
rect 16669 31291 16727 31297
rect 16945 31331 17003 31337
rect 16945 31297 16957 31331
rect 16991 31297 17003 31331
rect 16945 31291 17003 31297
rect 17126 31288 17132 31340
rect 17184 31328 17190 31340
rect 23032 31337 23060 31368
rect 23198 31356 23204 31368
rect 23256 31356 23262 31408
rect 20145 31331 20203 31337
rect 20145 31328 20157 31331
rect 17184 31300 20157 31328
rect 17184 31288 17190 31300
rect 20145 31297 20157 31300
rect 20191 31297 20203 31331
rect 20145 31291 20203 31297
rect 23017 31331 23075 31337
rect 23017 31297 23029 31331
rect 23063 31297 23075 31331
rect 23017 31291 23075 31297
rect 23106 31288 23112 31340
rect 23164 31328 23170 31340
rect 23308 31328 23336 31436
rect 23750 31424 23756 31476
rect 23808 31464 23814 31476
rect 23808 31436 24348 31464
rect 23808 31424 23814 31436
rect 23842 31356 23848 31408
rect 23900 31396 23906 31408
rect 24320 31405 24348 31436
rect 24854 31424 24860 31476
rect 24912 31464 24918 31476
rect 25498 31464 25504 31476
rect 24912 31436 25504 31464
rect 24912 31424 24918 31436
rect 25498 31424 25504 31436
rect 25556 31424 25562 31476
rect 26418 31464 26424 31476
rect 26379 31436 26424 31464
rect 26418 31424 26424 31436
rect 26476 31424 26482 31476
rect 26973 31467 27031 31473
rect 26973 31433 26985 31467
rect 27019 31464 27031 31467
rect 27154 31464 27160 31476
rect 27019 31436 27160 31464
rect 27019 31433 27031 31436
rect 26973 31427 27031 31433
rect 27154 31424 27160 31436
rect 27212 31424 27218 31476
rect 27338 31464 27344 31476
rect 27299 31436 27344 31464
rect 27338 31424 27344 31436
rect 27396 31424 27402 31476
rect 28074 31464 28080 31476
rect 28035 31436 28080 31464
rect 28074 31424 28080 31436
rect 28132 31424 28138 31476
rect 24213 31399 24271 31405
rect 24213 31396 24225 31399
rect 23900 31368 24225 31396
rect 23900 31356 23906 31368
rect 24213 31365 24225 31368
rect 24259 31365 24271 31399
rect 24213 31359 24271 31365
rect 24305 31399 24363 31405
rect 24305 31365 24317 31399
rect 24351 31365 24363 31399
rect 24946 31396 24952 31408
rect 24305 31359 24363 31365
rect 24412 31368 24952 31396
rect 23382 31328 23388 31340
rect 23164 31300 23209 31328
rect 23295 31300 23388 31328
rect 23164 31288 23170 31300
rect 23382 31288 23388 31300
rect 23440 31288 23446 31340
rect 24026 31328 24032 31340
rect 23987 31300 24032 31328
rect 24026 31288 24032 31300
rect 24084 31288 24090 31340
rect 24412 31337 24440 31368
rect 24946 31356 24952 31368
rect 25004 31356 25010 31408
rect 25406 31396 25412 31408
rect 25148 31368 25412 31396
rect 24397 31331 24455 31337
rect 24397 31297 24409 31331
rect 24443 31297 24455 31331
rect 24397 31291 24455 31297
rect 24486 31288 24492 31340
rect 24544 31328 24550 31340
rect 25041 31331 25099 31337
rect 25041 31328 25053 31331
rect 24544 31300 25053 31328
rect 24544 31288 24550 31300
rect 25041 31297 25053 31300
rect 25087 31297 25099 31331
rect 25041 31291 25099 31297
rect 16758 31260 16764 31272
rect 16408 31232 16764 31260
rect 14752 31192 14780 31232
rect 16758 31220 16764 31232
rect 16816 31220 16822 31272
rect 17678 31260 17684 31272
rect 17639 31232 17684 31260
rect 17678 31220 17684 31232
rect 17736 31220 17742 31272
rect 19886 31260 19892 31272
rect 19847 31232 19892 31260
rect 19886 31220 19892 31232
rect 19944 31220 19950 31272
rect 24670 31220 24676 31272
rect 24728 31260 24734 31272
rect 25148 31260 25176 31368
rect 25406 31356 25412 31368
rect 25464 31356 25470 31408
rect 25314 31337 25320 31340
rect 25308 31291 25320 31337
rect 25372 31328 25378 31340
rect 25372 31300 25408 31328
rect 25314 31288 25320 31291
rect 25372 31288 25378 31300
rect 25590 31288 25596 31340
rect 25648 31328 25654 31340
rect 25648 31300 26096 31328
rect 25648 31288 25654 31300
rect 24728 31232 25176 31260
rect 26068 31260 26096 31300
rect 26142 31288 26148 31340
rect 26200 31328 26206 31340
rect 27157 31331 27215 31337
rect 27157 31328 27169 31331
rect 26200 31300 27169 31328
rect 26200 31288 26206 31300
rect 27157 31297 27169 31300
rect 27203 31297 27215 31331
rect 27157 31291 27215 31297
rect 27433 31331 27491 31337
rect 27433 31297 27445 31331
rect 27479 31297 27491 31331
rect 27433 31291 27491 31297
rect 27448 31260 27476 31291
rect 27614 31288 27620 31340
rect 27672 31328 27678 31340
rect 27893 31331 27951 31337
rect 27893 31328 27905 31331
rect 27672 31300 27905 31328
rect 27672 31288 27678 31300
rect 27893 31297 27905 31300
rect 27939 31297 27951 31331
rect 27893 31291 27951 31297
rect 28169 31331 28227 31337
rect 28169 31297 28181 31331
rect 28215 31328 28227 31331
rect 28258 31328 28264 31340
rect 28215 31300 28264 31328
rect 28215 31297 28227 31300
rect 28169 31291 28227 31297
rect 28258 31288 28264 31300
rect 28316 31288 28322 31340
rect 26068 31232 27476 31260
rect 24728 31220 24734 31232
rect 10560 31164 13584 31192
rect 13832 31164 14780 31192
rect 15948 31164 17264 31192
rect 10560 31152 10566 31164
rect 8570 31124 8576 31136
rect 7239 31096 8432 31124
rect 8531 31096 8576 31124
rect 7239 31093 7251 31096
rect 7193 31087 7251 31093
rect 8570 31084 8576 31096
rect 8628 31084 8634 31136
rect 8662 31084 8668 31136
rect 8720 31124 8726 31136
rect 10226 31124 10232 31136
rect 8720 31096 10232 31124
rect 8720 31084 8726 31096
rect 10226 31084 10232 31096
rect 10284 31084 10290 31136
rect 10410 31084 10416 31136
rect 10468 31124 10474 31136
rect 10965 31127 11023 31133
rect 10965 31124 10977 31127
rect 10468 31096 10977 31124
rect 10468 31084 10474 31096
rect 10965 31093 10977 31096
rect 11011 31093 11023 31127
rect 10965 31087 11023 31093
rect 11330 31084 11336 31136
rect 11388 31124 11394 31136
rect 11974 31124 11980 31136
rect 11388 31096 11980 31124
rect 11388 31084 11394 31096
rect 11974 31084 11980 31096
rect 12032 31084 12038 31136
rect 12618 31084 12624 31136
rect 12676 31124 12682 31136
rect 13556 31124 13584 31164
rect 15948 31124 15976 31164
rect 12676 31096 12721 31124
rect 13556 31096 15976 31124
rect 12676 31084 12682 31096
rect 16022 31084 16028 31136
rect 16080 31124 16086 31136
rect 16117 31127 16175 31133
rect 16117 31124 16129 31127
rect 16080 31096 16129 31124
rect 16080 31084 16086 31096
rect 16117 31093 16129 31096
rect 16163 31093 16175 31127
rect 16850 31124 16856 31136
rect 16811 31096 16856 31124
rect 16117 31087 16175 31093
rect 16850 31084 16856 31096
rect 16908 31084 16914 31136
rect 16942 31084 16948 31136
rect 17000 31124 17006 31136
rect 17129 31127 17187 31133
rect 17129 31124 17141 31127
rect 17000 31096 17141 31124
rect 17000 31084 17006 31096
rect 17129 31093 17141 31096
rect 17175 31093 17187 31127
rect 17236 31124 17264 31164
rect 18616 31164 19334 31192
rect 18616 31124 18644 31164
rect 19058 31124 19064 31136
rect 17236 31096 18644 31124
rect 19019 31096 19064 31124
rect 17129 31087 17187 31093
rect 19058 31084 19064 31096
rect 19116 31084 19122 31136
rect 19306 31124 19334 31164
rect 21082 31152 21088 31204
rect 21140 31192 21146 31204
rect 21910 31192 21916 31204
rect 21140 31164 21916 31192
rect 21140 31152 21146 31164
rect 21910 31152 21916 31164
rect 21968 31152 21974 31204
rect 22281 31195 22339 31201
rect 22281 31161 22293 31195
rect 22327 31192 22339 31195
rect 23293 31195 23351 31201
rect 22327 31164 23244 31192
rect 22327 31161 22339 31164
rect 22281 31155 22339 31161
rect 20254 31124 20260 31136
rect 19306 31096 20260 31124
rect 20254 31084 20260 31096
rect 20312 31084 20318 31136
rect 20622 31084 20628 31136
rect 20680 31124 20686 31136
rect 21358 31124 21364 31136
rect 20680 31096 21364 31124
rect 20680 31084 20686 31096
rect 21358 31084 21364 31096
rect 21416 31084 21422 31136
rect 22370 31124 22376 31136
rect 22331 31096 22376 31124
rect 22370 31084 22376 31096
rect 22428 31084 22434 31136
rect 22830 31124 22836 31136
rect 22791 31096 22836 31124
rect 22830 31084 22836 31096
rect 22888 31084 22894 31136
rect 23216 31124 23244 31164
rect 23293 31161 23305 31195
rect 23339 31192 23351 31195
rect 23934 31192 23940 31204
rect 23339 31164 23940 31192
rect 23339 31161 23351 31164
rect 23293 31155 23351 31161
rect 23934 31152 23940 31164
rect 23992 31152 23998 31204
rect 23474 31124 23480 31136
rect 23216 31096 23480 31124
rect 23474 31084 23480 31096
rect 23532 31084 23538 31136
rect 24581 31127 24639 31133
rect 24581 31093 24593 31127
rect 24627 31124 24639 31127
rect 25222 31124 25228 31136
rect 24627 31096 25228 31124
rect 24627 31093 24639 31096
rect 24581 31087 24639 31093
rect 25222 31084 25228 31096
rect 25280 31084 25286 31136
rect 25774 31084 25780 31136
rect 25832 31124 25838 31136
rect 27893 31127 27951 31133
rect 27893 31124 27905 31127
rect 25832 31096 27905 31124
rect 25832 31084 25838 31096
rect 27893 31093 27905 31096
rect 27939 31093 27951 31127
rect 27893 31087 27951 31093
rect 1104 31034 28888 31056
rect 1104 30982 5582 31034
rect 5634 30982 5646 31034
rect 5698 30982 5710 31034
rect 5762 30982 5774 31034
rect 5826 30982 5838 31034
rect 5890 30982 14846 31034
rect 14898 30982 14910 31034
rect 14962 30982 14974 31034
rect 15026 30982 15038 31034
rect 15090 30982 15102 31034
rect 15154 30982 24110 31034
rect 24162 30982 24174 31034
rect 24226 30982 24238 31034
rect 24290 30982 24302 31034
rect 24354 30982 24366 31034
rect 24418 30982 28888 31034
rect 1104 30960 28888 30982
rect 2314 30920 2320 30932
rect 2275 30892 2320 30920
rect 2314 30880 2320 30892
rect 2372 30880 2378 30932
rect 6917 30923 6975 30929
rect 6917 30889 6929 30923
rect 6963 30920 6975 30923
rect 7006 30920 7012 30932
rect 6963 30892 7012 30920
rect 6963 30889 6975 30892
rect 6917 30883 6975 30889
rect 7006 30880 7012 30892
rect 7064 30880 7070 30932
rect 7561 30923 7619 30929
rect 7561 30889 7573 30923
rect 7607 30920 7619 30923
rect 11606 30920 11612 30932
rect 7607 30892 11612 30920
rect 7607 30889 7619 30892
rect 7561 30883 7619 30889
rect 11606 30880 11612 30892
rect 11664 30880 11670 30932
rect 11974 30880 11980 30932
rect 12032 30920 12038 30932
rect 12618 30920 12624 30932
rect 12032 30892 12624 30920
rect 12032 30880 12038 30892
rect 12618 30880 12624 30892
rect 12676 30880 12682 30932
rect 12710 30880 12716 30932
rect 12768 30920 12774 30932
rect 15289 30923 15347 30929
rect 15289 30920 15301 30923
rect 12768 30892 15301 30920
rect 12768 30880 12774 30892
rect 15289 30889 15301 30892
rect 15335 30889 15347 30923
rect 15289 30883 15347 30889
rect 15378 30880 15384 30932
rect 15436 30920 15442 30932
rect 17218 30920 17224 30932
rect 15436 30892 17224 30920
rect 15436 30880 15442 30892
rect 17218 30880 17224 30892
rect 17276 30880 17282 30932
rect 19978 30920 19984 30932
rect 19939 30892 19984 30920
rect 19978 30880 19984 30892
rect 20036 30880 20042 30932
rect 20162 30920 20168 30932
rect 20123 30892 20168 30920
rect 20162 30880 20168 30892
rect 20220 30880 20226 30932
rect 20254 30880 20260 30932
rect 20312 30920 20318 30932
rect 20312 30892 22094 30920
rect 20312 30880 20318 30892
rect 8205 30855 8263 30861
rect 8205 30821 8217 30855
rect 8251 30852 8263 30855
rect 9306 30852 9312 30864
rect 8251 30824 9312 30852
rect 8251 30821 8263 30824
rect 8205 30815 8263 30821
rect 9306 30812 9312 30824
rect 9364 30812 9370 30864
rect 12158 30852 12164 30864
rect 9876 30824 12164 30852
rect 8294 30744 8300 30796
rect 8352 30784 8358 30796
rect 9876 30793 9904 30824
rect 12158 30812 12164 30824
rect 12216 30812 12222 30864
rect 12250 30812 12256 30864
rect 12308 30852 12314 30864
rect 16942 30852 16948 30864
rect 12308 30824 16948 30852
rect 12308 30812 12314 30824
rect 16942 30812 16948 30824
rect 17000 30812 17006 30864
rect 17402 30812 17408 30864
rect 17460 30852 17466 30864
rect 22066 30852 22094 30892
rect 22646 30880 22652 30932
rect 22704 30920 22710 30932
rect 23198 30920 23204 30932
rect 22704 30892 23204 30920
rect 22704 30880 22710 30892
rect 23198 30880 23204 30892
rect 23256 30920 23262 30932
rect 24765 30923 24823 30929
rect 23256 30892 23336 30920
rect 23256 30880 23262 30892
rect 23308 30852 23336 30892
rect 24765 30889 24777 30923
rect 24811 30920 24823 30923
rect 25038 30920 25044 30932
rect 24811 30892 25044 30920
rect 24811 30889 24823 30892
rect 24765 30883 24823 30889
rect 25038 30880 25044 30892
rect 25096 30880 25102 30932
rect 28074 30920 28080 30932
rect 25148 30892 28080 30920
rect 23842 30852 23848 30864
rect 17460 30824 19012 30852
rect 22066 30824 23244 30852
rect 23308 30824 23848 30852
rect 17460 30812 17466 30824
rect 9861 30787 9919 30793
rect 8352 30756 9812 30784
rect 8352 30744 8358 30756
rect 2222 30716 2228 30728
rect 2183 30688 2228 30716
rect 2222 30676 2228 30688
rect 2280 30676 2286 30728
rect 7101 30719 7159 30725
rect 7101 30685 7113 30719
rect 7147 30685 7159 30719
rect 7101 30679 7159 30685
rect 7745 30719 7803 30725
rect 7745 30685 7757 30719
rect 7791 30716 7803 30719
rect 8018 30716 8024 30728
rect 7791 30688 8024 30716
rect 7791 30685 7803 30688
rect 7745 30679 7803 30685
rect 7116 30648 7144 30679
rect 8018 30676 8024 30688
rect 8076 30676 8082 30728
rect 8389 30719 8447 30725
rect 8389 30685 8401 30719
rect 8435 30716 8447 30719
rect 8662 30716 8668 30728
rect 8435 30688 8668 30716
rect 8435 30685 8447 30688
rect 8389 30679 8447 30685
rect 8662 30676 8668 30688
rect 8720 30676 8726 30728
rect 9217 30719 9275 30725
rect 9217 30685 9229 30719
rect 9263 30716 9275 30719
rect 9398 30716 9404 30728
rect 9263 30688 9404 30716
rect 9263 30685 9275 30688
rect 9217 30679 9275 30685
rect 9398 30676 9404 30688
rect 9456 30676 9462 30728
rect 9784 30716 9812 30756
rect 9861 30753 9873 30787
rect 9907 30753 9919 30787
rect 10502 30784 10508 30796
rect 9861 30747 9919 30753
rect 9968 30756 10508 30784
rect 9968 30716 9996 30756
rect 10502 30744 10508 30756
rect 10560 30744 10566 30796
rect 10686 30744 10692 30796
rect 10744 30744 10750 30796
rect 11330 30784 11336 30796
rect 10796 30756 11336 30784
rect 9784 30688 9996 30716
rect 10045 30719 10103 30725
rect 10045 30685 10057 30719
rect 10091 30716 10103 30719
rect 10704 30716 10732 30744
rect 10796 30725 10824 30756
rect 11330 30744 11336 30756
rect 11388 30744 11394 30796
rect 12710 30744 12716 30796
rect 12768 30784 12774 30796
rect 14461 30787 14519 30793
rect 14461 30784 14473 30787
rect 12768 30756 14473 30784
rect 12768 30744 12774 30756
rect 14461 30753 14473 30756
rect 14507 30753 14519 30787
rect 14461 30747 14519 30753
rect 14550 30744 14556 30796
rect 14608 30784 14614 30796
rect 14608 30756 14964 30784
rect 14608 30744 14614 30756
rect 10091 30688 10732 30716
rect 10781 30719 10839 30725
rect 10091 30685 10103 30688
rect 10045 30679 10103 30685
rect 10781 30685 10793 30719
rect 10827 30685 10839 30719
rect 10781 30679 10839 30685
rect 10870 30676 10876 30728
rect 10928 30716 10934 30728
rect 12250 30716 12256 30728
rect 10928 30688 10973 30716
rect 11716 30688 12256 30716
rect 10928 30676 10934 30688
rect 11716 30657 11744 30688
rect 12250 30676 12256 30688
rect 12308 30676 12314 30728
rect 12342 30676 12348 30728
rect 12400 30716 12406 30728
rect 12529 30719 12587 30725
rect 12400 30688 12445 30716
rect 12400 30676 12406 30688
rect 12529 30685 12541 30719
rect 12575 30716 12587 30719
rect 12618 30716 12624 30728
rect 12575 30688 12624 30716
rect 12575 30685 12587 30688
rect 12529 30679 12587 30685
rect 12618 30676 12624 30688
rect 12676 30716 12682 30728
rect 13170 30716 13176 30728
rect 12676 30688 13176 30716
rect 12676 30676 12682 30688
rect 13170 30676 13176 30688
rect 13228 30676 13234 30728
rect 13265 30719 13323 30725
rect 13265 30685 13277 30719
rect 13311 30685 13323 30719
rect 13265 30679 13323 30685
rect 13357 30719 13415 30725
rect 13357 30685 13369 30719
rect 13403 30716 13415 30719
rect 13446 30716 13452 30728
rect 13403 30688 13452 30716
rect 13403 30685 13415 30688
rect 13357 30679 13415 30685
rect 11057 30651 11115 30657
rect 7116 30620 10732 30648
rect 9030 30540 9036 30592
rect 9088 30580 9094 30592
rect 9309 30583 9367 30589
rect 9309 30580 9321 30583
rect 9088 30552 9321 30580
rect 9088 30540 9094 30552
rect 9309 30549 9321 30552
rect 9355 30549 9367 30583
rect 9309 30543 9367 30549
rect 9398 30540 9404 30592
rect 9456 30580 9462 30592
rect 10229 30583 10287 30589
rect 10229 30580 10241 30583
rect 9456 30552 10241 30580
rect 9456 30540 9462 30552
rect 10229 30549 10241 30552
rect 10275 30549 10287 30583
rect 10704 30580 10732 30620
rect 11057 30617 11069 30651
rect 11103 30617 11115 30651
rect 11057 30611 11115 30617
rect 11517 30651 11575 30657
rect 11517 30617 11529 30651
rect 11563 30617 11575 30651
rect 11517 30611 11575 30617
rect 11701 30651 11759 30657
rect 11701 30617 11713 30651
rect 11747 30617 11759 30651
rect 11701 30611 11759 30617
rect 11885 30651 11943 30657
rect 11885 30617 11897 30651
rect 11931 30648 11943 30651
rect 12986 30648 12992 30660
rect 11931 30620 12992 30648
rect 11931 30617 11943 30620
rect 11885 30611 11943 30617
rect 11072 30580 11100 30611
rect 10704 30552 11100 30580
rect 11532 30580 11560 30611
rect 12986 30608 12992 30620
rect 13044 30608 13050 30660
rect 13280 30648 13308 30679
rect 13446 30676 13452 30688
rect 13504 30676 13510 30728
rect 13630 30676 13636 30728
rect 13688 30716 13694 30728
rect 14182 30716 14188 30728
rect 13688 30688 14044 30716
rect 14143 30688 14188 30716
rect 13688 30676 13694 30688
rect 14016 30648 14044 30688
rect 14182 30676 14188 30688
rect 14240 30676 14246 30728
rect 14277 30719 14335 30725
rect 14277 30685 14289 30719
rect 14323 30716 14335 30719
rect 14366 30716 14372 30728
rect 14323 30688 14372 30716
rect 14323 30685 14335 30688
rect 14277 30679 14335 30685
rect 14366 30676 14372 30688
rect 14424 30716 14430 30728
rect 14734 30716 14740 30728
rect 14424 30688 14740 30716
rect 14424 30676 14430 30688
rect 14734 30676 14740 30688
rect 14792 30676 14798 30728
rect 14936 30725 14964 30756
rect 15028 30756 17382 30784
rect 14921 30719 14979 30725
rect 14921 30685 14933 30719
rect 14967 30685 14979 30719
rect 14921 30679 14979 30685
rect 15028 30648 15056 30756
rect 15105 30719 15163 30725
rect 15105 30685 15117 30719
rect 15151 30716 15163 30719
rect 15194 30716 15200 30728
rect 15151 30688 15200 30716
rect 15151 30685 15163 30688
rect 15105 30679 15163 30685
rect 15194 30676 15200 30688
rect 15252 30716 15258 30728
rect 15470 30716 15476 30728
rect 15252 30688 15476 30716
rect 15252 30676 15258 30688
rect 15470 30676 15476 30688
rect 15528 30676 15534 30728
rect 15838 30716 15844 30728
rect 15799 30688 15844 30716
rect 15838 30676 15844 30688
rect 15896 30676 15902 30728
rect 17034 30716 17040 30728
rect 16995 30688 17040 30716
rect 17034 30676 17040 30688
rect 17092 30676 17098 30728
rect 17218 30716 17224 30728
rect 17179 30688 17224 30716
rect 17218 30676 17224 30688
rect 17276 30676 17282 30728
rect 17354 30725 17382 30756
rect 17770 30744 17776 30796
rect 17828 30784 17834 30796
rect 18414 30784 18420 30796
rect 17828 30756 18420 30784
rect 17828 30744 17834 30756
rect 18414 30744 18420 30756
rect 18472 30784 18478 30796
rect 18472 30756 18552 30784
rect 18472 30744 18478 30756
rect 17339 30719 17397 30725
rect 17339 30685 17351 30719
rect 17385 30685 17397 30719
rect 17494 30716 17500 30728
rect 17455 30688 17500 30716
rect 17339 30679 17397 30685
rect 17494 30676 17500 30688
rect 17552 30676 17558 30728
rect 18524 30725 18552 30756
rect 18325 30719 18383 30725
rect 18325 30685 18337 30719
rect 18371 30685 18383 30719
rect 18325 30679 18383 30685
rect 18509 30719 18567 30725
rect 18509 30685 18521 30719
rect 18555 30685 18567 30719
rect 18984 30716 19012 30824
rect 19058 30744 19064 30796
rect 19116 30784 19122 30796
rect 19334 30784 19340 30796
rect 19116 30756 19340 30784
rect 19116 30744 19122 30756
rect 19334 30744 19340 30756
rect 19392 30784 19398 30796
rect 19889 30787 19947 30793
rect 19392 30756 19840 30784
rect 19392 30744 19398 30756
rect 19610 30716 19616 30728
rect 18984 30688 19616 30716
rect 18509 30679 18567 30685
rect 13280 30620 13952 30648
rect 14016 30620 15056 30648
rect 12342 30580 12348 30592
rect 11532 30552 12348 30580
rect 10229 30543 10287 30549
rect 12342 30540 12348 30552
rect 12400 30540 12406 30592
rect 12434 30540 12440 30592
rect 12492 30580 12498 30592
rect 12713 30583 12771 30589
rect 12713 30580 12725 30583
rect 12492 30552 12725 30580
rect 12492 30540 12498 30552
rect 12713 30549 12725 30552
rect 12759 30549 12771 30583
rect 12713 30543 12771 30549
rect 12810 30540 12816 30592
rect 12868 30580 12874 30592
rect 13541 30583 13599 30589
rect 13541 30580 13553 30583
rect 12868 30552 13553 30580
rect 12868 30540 12874 30552
rect 13541 30549 13553 30552
rect 13587 30549 13599 30583
rect 13924 30580 13952 30620
rect 15286 30608 15292 30660
rect 15344 30648 15350 30660
rect 16206 30648 16212 30660
rect 15344 30620 16212 30648
rect 15344 30608 15350 30620
rect 16206 30608 16212 30620
rect 16264 30608 16270 30660
rect 16393 30651 16451 30657
rect 16393 30617 16405 30651
rect 16439 30648 16451 30651
rect 17129 30651 17187 30657
rect 17129 30648 17141 30651
rect 16439 30620 17141 30648
rect 16439 30617 16451 30620
rect 16393 30611 16451 30617
rect 17129 30617 17141 30620
rect 17175 30617 17187 30651
rect 18340 30648 18368 30679
rect 19610 30676 19616 30688
rect 19668 30676 19674 30728
rect 19812 30716 19840 30756
rect 19889 30753 19901 30787
rect 19935 30784 19947 30787
rect 20070 30784 20076 30796
rect 19935 30756 20076 30784
rect 19935 30753 19947 30756
rect 19889 30747 19947 30753
rect 20070 30744 20076 30756
rect 20128 30744 20134 30796
rect 23216 30784 23244 30824
rect 23842 30812 23848 30824
rect 23900 30852 23906 30864
rect 25148 30852 25176 30892
rect 28074 30880 28080 30892
rect 28132 30880 28138 30932
rect 23900 30824 25176 30852
rect 23900 30812 23906 30824
rect 25682 30812 25688 30864
rect 25740 30812 25746 30864
rect 27062 30852 27068 30864
rect 26160 30824 27068 30852
rect 25700 30784 25728 30812
rect 23216 30756 24992 30784
rect 19981 30719 20039 30725
rect 19981 30716 19993 30719
rect 19812 30688 19993 30716
rect 19981 30685 19993 30688
rect 20027 30685 20039 30719
rect 19981 30679 20039 30685
rect 20162 30676 20168 30728
rect 20220 30716 20226 30728
rect 20717 30719 20775 30725
rect 20717 30716 20729 30719
rect 20220 30688 20729 30716
rect 20220 30676 20226 30688
rect 20717 30685 20729 30688
rect 20763 30685 20775 30719
rect 20717 30679 20775 30685
rect 20984 30719 21042 30725
rect 20984 30685 20996 30719
rect 21030 30716 21042 30719
rect 21542 30716 21548 30728
rect 21030 30688 21548 30716
rect 21030 30685 21042 30688
rect 20984 30679 21042 30685
rect 21542 30676 21548 30688
rect 21600 30676 21606 30728
rect 22922 30716 22928 30728
rect 22883 30688 22928 30716
rect 22922 30676 22928 30688
rect 22980 30676 22986 30728
rect 23017 30719 23075 30725
rect 23017 30685 23029 30719
rect 23063 30685 23075 30719
rect 23198 30716 23204 30728
rect 23159 30688 23204 30716
rect 23017 30679 23075 30685
rect 18782 30648 18788 30660
rect 18340 30620 18788 30648
rect 17129 30611 17187 30617
rect 18782 30608 18788 30620
rect 18840 30608 18846 30660
rect 18874 30608 18880 30660
rect 18932 30648 18938 30660
rect 19705 30651 19763 30657
rect 19705 30648 19717 30651
rect 18932 30620 19717 30648
rect 18932 30608 18938 30620
rect 19705 30617 19717 30620
rect 19751 30648 19763 30651
rect 19794 30648 19800 30660
rect 19751 30620 19800 30648
rect 19751 30617 19763 30620
rect 19705 30611 19763 30617
rect 19794 30608 19800 30620
rect 19852 30648 19858 30660
rect 20254 30648 20260 30660
rect 19852 30620 20260 30648
rect 19852 30608 19858 30620
rect 20254 30608 20260 30620
rect 20312 30608 20318 30660
rect 22462 30608 22468 30660
rect 22520 30648 22526 30660
rect 23032 30648 23060 30679
rect 23198 30676 23204 30688
rect 23256 30676 23262 30728
rect 23290 30676 23296 30728
rect 23348 30716 23354 30728
rect 24489 30719 24547 30725
rect 23348 30688 23393 30716
rect 23348 30676 23354 30688
rect 24489 30685 24501 30719
rect 24535 30685 24547 30719
rect 24489 30679 24547 30685
rect 24581 30719 24639 30725
rect 24581 30685 24593 30719
rect 24627 30716 24639 30719
rect 24670 30716 24676 30728
rect 24627 30688 24676 30716
rect 24627 30685 24639 30688
rect 24581 30679 24639 30685
rect 23106 30648 23112 30660
rect 22520 30620 23112 30648
rect 22520 30608 22526 30620
rect 23106 30608 23112 30620
rect 23164 30608 23170 30660
rect 24504 30648 24532 30679
rect 24670 30676 24676 30688
rect 24728 30676 24734 30728
rect 24854 30648 24860 30660
rect 24504 30620 24860 30648
rect 24854 30608 24860 30620
rect 24912 30608 24918 30660
rect 16022 30580 16028 30592
rect 13924 30552 16028 30580
rect 13541 30543 13599 30549
rect 16022 30540 16028 30552
rect 16080 30540 16086 30592
rect 16114 30540 16120 30592
rect 16172 30580 16178 30592
rect 16850 30580 16856 30592
rect 16172 30552 16217 30580
rect 16811 30552 16856 30580
rect 16172 30540 16178 30552
rect 16850 30540 16856 30552
rect 16908 30540 16914 30592
rect 16942 30540 16948 30592
rect 17000 30580 17006 30592
rect 18693 30583 18751 30589
rect 18693 30580 18705 30583
rect 17000 30552 18705 30580
rect 17000 30540 17006 30552
rect 18693 30549 18705 30552
rect 18739 30549 18751 30583
rect 18693 30543 18751 30549
rect 18966 30540 18972 30592
rect 19024 30580 19030 30592
rect 22097 30583 22155 30589
rect 22097 30580 22109 30583
rect 19024 30552 22109 30580
rect 19024 30540 19030 30552
rect 22097 30549 22109 30552
rect 22143 30549 22155 30583
rect 22097 30543 22155 30549
rect 22741 30583 22799 30589
rect 22741 30549 22753 30583
rect 22787 30580 22799 30583
rect 23474 30580 23480 30592
rect 22787 30552 23480 30580
rect 22787 30549 22799 30552
rect 22741 30543 22799 30549
rect 23474 30540 23480 30552
rect 23532 30540 23538 30592
rect 24964 30580 24992 30756
rect 25388 30756 25728 30784
rect 25130 30676 25136 30728
rect 25188 30716 25194 30728
rect 25388 30725 25416 30756
rect 25225 30719 25283 30725
rect 25225 30716 25237 30719
rect 25188 30688 25237 30716
rect 25188 30676 25194 30688
rect 25225 30685 25237 30688
rect 25271 30685 25283 30719
rect 25225 30679 25283 30685
rect 25373 30719 25431 30725
rect 25373 30685 25385 30719
rect 25419 30685 25431 30719
rect 25373 30679 25431 30685
rect 25731 30719 25789 30725
rect 25731 30685 25743 30719
rect 25777 30716 25789 30719
rect 26160 30716 26188 30824
rect 27062 30812 27068 30824
rect 27120 30812 27126 30864
rect 26513 30787 26571 30793
rect 26513 30753 26525 30787
rect 26559 30784 26571 30787
rect 27522 30784 27528 30796
rect 26559 30756 27528 30784
rect 26559 30753 26571 30756
rect 26513 30747 26571 30753
rect 27522 30744 27528 30756
rect 27580 30744 27586 30796
rect 28169 30787 28227 30793
rect 28169 30753 28181 30787
rect 28215 30784 28227 30787
rect 28718 30784 28724 30796
rect 28215 30756 28724 30784
rect 28215 30753 28227 30756
rect 28169 30747 28227 30753
rect 28718 30744 28724 30756
rect 28776 30744 28782 30796
rect 26326 30716 26332 30728
rect 25777 30688 26188 30716
rect 26287 30688 26332 30716
rect 25777 30685 25789 30688
rect 25731 30679 25789 30685
rect 26326 30676 26332 30688
rect 26384 30676 26390 30728
rect 25498 30648 25504 30660
rect 25459 30620 25504 30648
rect 25498 30608 25504 30620
rect 25556 30608 25562 30660
rect 25593 30651 25651 30657
rect 25593 30617 25605 30651
rect 25639 30648 25651 30651
rect 27246 30648 27252 30660
rect 25639 30620 27252 30648
rect 25639 30617 25651 30620
rect 25593 30611 25651 30617
rect 25608 30580 25636 30611
rect 27246 30608 27252 30620
rect 27304 30608 27310 30660
rect 24964 30552 25636 30580
rect 25869 30583 25927 30589
rect 25869 30549 25881 30583
rect 25915 30580 25927 30583
rect 26970 30580 26976 30592
rect 25915 30552 26976 30580
rect 25915 30549 25927 30552
rect 25869 30543 25927 30549
rect 26970 30540 26976 30552
rect 27028 30540 27034 30592
rect 1104 30490 28888 30512
rect 1104 30438 10214 30490
rect 10266 30438 10278 30490
rect 10330 30438 10342 30490
rect 10394 30438 10406 30490
rect 10458 30438 10470 30490
rect 10522 30438 19478 30490
rect 19530 30438 19542 30490
rect 19594 30438 19606 30490
rect 19658 30438 19670 30490
rect 19722 30438 19734 30490
rect 19786 30438 28888 30490
rect 1104 30416 28888 30438
rect 8021 30379 8079 30385
rect 8021 30345 8033 30379
rect 8067 30376 8079 30379
rect 8067 30348 9628 30376
rect 8067 30345 8079 30348
rect 8021 30339 8079 30345
rect 9398 30308 9404 30320
rect 7944 30280 9404 30308
rect 7944 30249 7972 30280
rect 9398 30268 9404 30280
rect 9456 30268 9462 30320
rect 9600 30308 9628 30348
rect 9674 30336 9680 30388
rect 9732 30376 9738 30388
rect 10594 30376 10600 30388
rect 9732 30348 10600 30376
rect 9732 30336 9738 30348
rect 10594 30336 10600 30348
rect 10652 30336 10658 30388
rect 12342 30376 12348 30388
rect 10704 30348 12348 30376
rect 10045 30311 10103 30317
rect 9600 30280 9720 30308
rect 6917 30243 6975 30249
rect 6917 30209 6929 30243
rect 6963 30240 6975 30243
rect 7929 30243 7987 30249
rect 6963 30212 7328 30240
rect 6963 30209 6975 30212
rect 6917 30203 6975 30209
rect 6730 30036 6736 30048
rect 6691 30008 6736 30036
rect 6730 29996 6736 30008
rect 6788 29996 6794 30048
rect 7300 30045 7328 30212
rect 7929 30209 7941 30243
rect 7975 30209 7987 30243
rect 7929 30203 7987 30209
rect 8205 30243 8263 30249
rect 8205 30209 8217 30243
rect 8251 30209 8263 30243
rect 8205 30203 8263 30209
rect 8220 30172 8248 30203
rect 8478 30200 8484 30252
rect 8536 30240 8542 30252
rect 8754 30240 8760 30252
rect 8536 30212 8760 30240
rect 8536 30200 8542 30212
rect 8754 30200 8760 30212
rect 8812 30240 8818 30252
rect 8849 30243 8907 30249
rect 8849 30240 8861 30243
rect 8812 30212 8861 30240
rect 8812 30200 8818 30212
rect 8849 30209 8861 30212
rect 8895 30209 8907 30243
rect 8849 30203 8907 30209
rect 9493 30243 9551 30249
rect 9493 30209 9505 30243
rect 9539 30240 9551 30243
rect 9582 30240 9588 30252
rect 9539 30212 9588 30240
rect 9539 30209 9551 30212
rect 9493 30203 9551 30209
rect 9582 30200 9588 30212
rect 9640 30200 9646 30252
rect 9692 30240 9720 30280
rect 10045 30277 10057 30311
rect 10091 30308 10103 30311
rect 10134 30308 10140 30320
rect 10091 30280 10140 30308
rect 10091 30277 10103 30280
rect 10045 30271 10103 30277
rect 10134 30268 10140 30280
rect 10192 30268 10198 30320
rect 10229 30311 10287 30317
rect 10229 30277 10241 30311
rect 10275 30308 10287 30311
rect 10502 30308 10508 30320
rect 10275 30280 10508 30308
rect 10275 30277 10287 30280
rect 10229 30271 10287 30277
rect 10502 30268 10508 30280
rect 10560 30268 10566 30320
rect 10704 30240 10732 30348
rect 12342 30336 12348 30348
rect 12400 30336 12406 30388
rect 12526 30336 12532 30388
rect 12584 30376 12590 30388
rect 15286 30376 15292 30388
rect 12584 30348 15292 30376
rect 12584 30336 12590 30348
rect 15286 30336 15292 30348
rect 15344 30336 15350 30388
rect 15381 30379 15439 30385
rect 15381 30345 15393 30379
rect 15427 30376 15439 30379
rect 15838 30376 15844 30388
rect 15427 30348 15844 30376
rect 15427 30345 15439 30348
rect 15381 30339 15439 30345
rect 15838 30336 15844 30348
rect 15896 30376 15902 30388
rect 16298 30376 16304 30388
rect 15896 30348 16304 30376
rect 15896 30336 15902 30348
rect 16298 30336 16304 30348
rect 16356 30336 16362 30388
rect 18046 30336 18052 30388
rect 18104 30376 18110 30388
rect 18966 30376 18972 30388
rect 18104 30348 18972 30376
rect 18104 30336 18110 30348
rect 18966 30336 18972 30348
rect 19024 30336 19030 30388
rect 19886 30376 19892 30388
rect 19076 30348 19892 30376
rect 10781 30311 10839 30317
rect 10781 30277 10793 30311
rect 10827 30308 10839 30311
rect 11514 30308 11520 30320
rect 10827 30280 11520 30308
rect 10827 30277 10839 30280
rect 10781 30271 10839 30277
rect 11514 30268 11520 30280
rect 11572 30268 11578 30320
rect 11606 30268 11612 30320
rect 11664 30308 11670 30320
rect 11762 30311 11820 30317
rect 11762 30308 11774 30311
rect 11664 30280 11774 30308
rect 11664 30268 11670 30280
rect 11762 30277 11774 30280
rect 11808 30277 11820 30311
rect 12710 30308 12716 30320
rect 11762 30271 11820 30277
rect 11900 30280 12716 30308
rect 11900 30240 11928 30280
rect 12710 30268 12716 30280
rect 12768 30268 12774 30320
rect 14246 30311 14304 30317
rect 14246 30308 14258 30311
rect 13188 30280 14258 30308
rect 9692 30212 10732 30240
rect 10888 30212 11928 30240
rect 10888 30172 10916 30212
rect 12342 30200 12348 30252
rect 12400 30240 12406 30252
rect 13188 30240 13216 30280
rect 14246 30277 14258 30280
rect 14292 30277 14304 30311
rect 14246 30271 14304 30277
rect 14366 30268 14372 30320
rect 14424 30308 14430 30320
rect 16025 30311 16083 30317
rect 14424 30280 15332 30308
rect 14424 30268 14430 30280
rect 15304 30252 15332 30280
rect 15396 30280 15976 30308
rect 15396 30252 15424 30280
rect 12400 30212 13216 30240
rect 13357 30243 13415 30249
rect 12400 30200 12406 30212
rect 13357 30209 13369 30243
rect 13403 30240 13415 30243
rect 13446 30240 13452 30252
rect 13403 30212 13452 30240
rect 13403 30209 13415 30212
rect 13357 30203 13415 30209
rect 13446 30200 13452 30212
rect 13504 30200 13510 30252
rect 13998 30240 14004 30252
rect 13959 30212 14004 30240
rect 13998 30200 14004 30212
rect 14056 30200 14062 30252
rect 14108 30212 15056 30240
rect 8220 30144 10916 30172
rect 10965 30175 11023 30181
rect 10965 30141 10977 30175
rect 11011 30172 11023 30175
rect 11238 30172 11244 30184
rect 11011 30144 11244 30172
rect 11011 30141 11023 30144
rect 10965 30135 11023 30141
rect 11238 30132 11244 30144
rect 11296 30172 11302 30184
rect 11517 30175 11575 30181
rect 11517 30172 11529 30175
rect 11296 30144 11529 30172
rect 11296 30132 11302 30144
rect 11517 30141 11529 30144
rect 11563 30141 11575 30175
rect 11517 30135 11575 30141
rect 12986 30132 12992 30184
rect 13044 30172 13050 30184
rect 14108 30172 14136 30212
rect 13044 30144 14136 30172
rect 15028 30172 15056 30212
rect 15286 30200 15292 30252
rect 15344 30200 15350 30252
rect 15378 30200 15384 30252
rect 15436 30200 15442 30252
rect 15838 30240 15844 30252
rect 15799 30212 15844 30240
rect 15838 30200 15844 30212
rect 15896 30200 15902 30252
rect 15948 30240 15976 30280
rect 16025 30277 16037 30311
rect 16071 30308 16083 30311
rect 16071 30280 16804 30308
rect 16071 30277 16083 30280
rect 16025 30271 16083 30277
rect 16117 30243 16175 30249
rect 16117 30240 16129 30243
rect 15948 30212 16129 30240
rect 16117 30209 16129 30212
rect 16163 30209 16175 30243
rect 16776 30240 16804 30280
rect 16850 30268 16856 30320
rect 16908 30308 16914 30320
rect 17374 30311 17432 30317
rect 17374 30308 17386 30311
rect 16908 30280 17386 30308
rect 16908 30268 16914 30280
rect 17374 30277 17386 30280
rect 17420 30277 17432 30311
rect 18874 30308 18880 30320
rect 17374 30271 17432 30277
rect 17604 30280 18880 30308
rect 17604 30240 17632 30280
rect 18874 30268 18880 30280
rect 18932 30268 18938 30320
rect 19076 30308 19104 30348
rect 19886 30336 19892 30348
rect 19944 30336 19950 30388
rect 20070 30336 20076 30388
rect 20128 30376 20134 30388
rect 20990 30376 20996 30388
rect 20128 30348 20996 30376
rect 20128 30336 20134 30348
rect 20990 30336 20996 30348
rect 21048 30336 21054 30388
rect 22922 30336 22928 30388
rect 22980 30376 22986 30388
rect 23201 30379 23259 30385
rect 23201 30376 23213 30379
rect 22980 30348 23213 30376
rect 22980 30336 22986 30348
rect 23201 30345 23213 30348
rect 23247 30345 23259 30379
rect 23201 30339 23259 30345
rect 25130 30336 25136 30388
rect 25188 30376 25194 30388
rect 25961 30379 26019 30385
rect 25961 30376 25973 30379
rect 25188 30348 25973 30376
rect 25188 30336 25194 30348
rect 25961 30345 25973 30348
rect 26007 30345 26019 30379
rect 25961 30339 26019 30345
rect 19242 30317 19248 30320
rect 18984 30280 19104 30308
rect 16776 30212 17632 30240
rect 16117 30203 16175 30209
rect 17678 30200 17684 30252
rect 17736 30240 17742 30252
rect 18984 30249 19012 30280
rect 19236 30271 19248 30317
rect 19300 30308 19306 30320
rect 19904 30308 19932 30336
rect 23566 30308 23572 30320
rect 19300 30280 19336 30308
rect 19904 30280 23572 30308
rect 19242 30268 19248 30271
rect 19300 30268 19306 30280
rect 18969 30243 19027 30249
rect 18969 30240 18981 30243
rect 17736 30212 18981 30240
rect 17736 30200 17742 30212
rect 18969 30209 18981 30212
rect 19015 30209 19027 30243
rect 18969 30203 19027 30209
rect 19058 30200 19064 30252
rect 19116 30240 19122 30252
rect 20714 30240 20720 30252
rect 19116 30212 20720 30240
rect 19116 30200 19122 30212
rect 20714 30200 20720 30212
rect 20772 30200 20778 30252
rect 20809 30243 20867 30249
rect 20809 30209 20821 30243
rect 20855 30209 20867 30243
rect 20809 30203 20867 30209
rect 16850 30172 16856 30184
rect 15028 30144 16856 30172
rect 13044 30132 13050 30144
rect 16850 30132 16856 30144
rect 16908 30132 16914 30184
rect 17034 30132 17040 30184
rect 17092 30172 17098 30184
rect 17129 30175 17187 30181
rect 17129 30172 17141 30175
rect 17092 30144 17141 30172
rect 17092 30132 17098 30144
rect 17129 30141 17141 30144
rect 17175 30141 17187 30175
rect 19076 30172 19104 30200
rect 17129 30135 17187 30141
rect 18524 30144 19104 30172
rect 7745 30107 7803 30113
rect 7745 30073 7757 30107
rect 7791 30104 7803 30107
rect 7791 30076 10272 30104
rect 7791 30073 7803 30076
rect 7745 30067 7803 30073
rect 7285 30039 7343 30045
rect 7285 30005 7297 30039
rect 7331 30036 7343 30039
rect 7653 30039 7711 30045
rect 7653 30036 7665 30039
rect 7331 30008 7665 30036
rect 7331 30005 7343 30008
rect 7285 29999 7343 30005
rect 7653 30005 7665 30008
rect 7699 30036 7711 30039
rect 8570 30036 8576 30048
rect 7699 30008 8576 30036
rect 7699 30005 7711 30008
rect 7653 29999 7711 30005
rect 8570 29996 8576 30008
rect 8628 29996 8634 30048
rect 8662 29996 8668 30048
rect 8720 30036 8726 30048
rect 9309 30039 9367 30045
rect 8720 30008 8765 30036
rect 8720 29996 8726 30008
rect 9309 30005 9321 30039
rect 9355 30036 9367 30039
rect 9950 30036 9956 30048
rect 9355 30008 9956 30036
rect 9355 30005 9367 30008
rect 9309 29999 9367 30005
rect 9950 29996 9956 30008
rect 10008 29996 10014 30048
rect 10244 30036 10272 30076
rect 10318 30064 10324 30116
rect 10376 30104 10382 30116
rect 11330 30104 11336 30116
rect 10376 30076 11336 30104
rect 10376 30064 10382 30076
rect 11330 30064 11336 30076
rect 11388 30064 11394 30116
rect 12710 30104 12716 30116
rect 12452 30076 12716 30104
rect 12452 30036 12480 30076
rect 12710 30064 12716 30076
rect 12768 30064 12774 30116
rect 13449 30107 13507 30113
rect 13449 30073 13461 30107
rect 13495 30104 13507 30107
rect 13906 30104 13912 30116
rect 13495 30076 13912 30104
rect 13495 30073 13507 30076
rect 13449 30067 13507 30073
rect 13906 30064 13912 30076
rect 13964 30064 13970 30116
rect 16942 30104 16948 30116
rect 14936 30076 16948 30104
rect 10244 30008 12480 30036
rect 12802 29996 12808 30048
rect 12860 30036 12866 30048
rect 12897 30039 12955 30045
rect 12897 30036 12909 30039
rect 12860 30008 12909 30036
rect 12860 29996 12866 30008
rect 12897 30005 12909 30008
rect 12943 30005 12955 30039
rect 12897 29999 12955 30005
rect 13722 29996 13728 30048
rect 13780 30036 13786 30048
rect 14936 30036 14964 30076
rect 16942 30064 16948 30076
rect 17000 30064 17006 30116
rect 13780 30008 14964 30036
rect 15841 30039 15899 30045
rect 13780 29996 13786 30008
rect 15841 30005 15853 30039
rect 15887 30036 15899 30039
rect 18414 30036 18420 30048
rect 15887 30008 18420 30036
rect 15887 30005 15899 30008
rect 15841 29999 15899 30005
rect 18414 29996 18420 30008
rect 18472 29996 18478 30048
rect 18524 30045 18552 30144
rect 20162 30132 20168 30184
rect 20220 30172 20226 30184
rect 20622 30172 20628 30184
rect 20220 30144 20628 30172
rect 20220 30132 20226 30144
rect 20622 30132 20628 30144
rect 20680 30132 20686 30184
rect 20824 30172 20852 30203
rect 20898 30200 20904 30252
rect 20956 30240 20962 30252
rect 21836 30249 21864 30280
rect 23566 30268 23572 30280
rect 23624 30268 23630 30320
rect 24946 30268 24952 30320
rect 25004 30308 25010 30320
rect 25004 30280 25452 30308
rect 25004 30268 25010 30280
rect 25424 30252 25452 30280
rect 25498 30268 25504 30320
rect 25556 30308 25562 30320
rect 25556 30280 25636 30308
rect 25556 30268 25562 30280
rect 22094 30249 22100 30252
rect 21821 30243 21879 30249
rect 20956 30212 21001 30240
rect 20956 30200 20962 30212
rect 21821 30209 21833 30243
rect 21867 30209 21879 30243
rect 21821 30203 21879 30209
rect 22088 30203 22100 30249
rect 22152 30240 22158 30252
rect 22152 30212 22188 30240
rect 22094 30200 22100 30203
rect 22152 30200 22158 30212
rect 22922 30200 22928 30252
rect 22980 30240 22986 30252
rect 23661 30243 23719 30249
rect 23661 30240 23673 30243
rect 22980 30212 23673 30240
rect 22980 30200 22986 30212
rect 23661 30209 23673 30212
rect 23707 30209 23719 30243
rect 25222 30240 25228 30252
rect 25183 30212 25228 30240
rect 23661 30203 23719 30209
rect 25222 30200 25228 30212
rect 25280 30200 25286 30252
rect 25406 30200 25412 30252
rect 25464 30240 25470 30252
rect 25608 30249 25636 30280
rect 26878 30268 26884 30320
rect 26936 30308 26942 30320
rect 26936 30280 27568 30308
rect 26936 30268 26942 30280
rect 25593 30243 25651 30249
rect 25464 30212 25557 30240
rect 25464 30200 25470 30212
rect 25593 30209 25605 30243
rect 25639 30209 25651 30243
rect 25593 30203 25651 30209
rect 25682 30200 25688 30252
rect 25740 30240 25746 30252
rect 25777 30243 25835 30249
rect 25777 30240 25789 30243
rect 25740 30212 25789 30240
rect 25740 30200 25746 30212
rect 25777 30209 25789 30212
rect 25823 30209 25835 30243
rect 26970 30240 26976 30252
rect 26931 30212 26976 30240
rect 25777 30203 25835 30209
rect 26970 30200 26976 30212
rect 27028 30200 27034 30252
rect 27062 30200 27068 30252
rect 27120 30240 27126 30252
rect 27157 30243 27215 30249
rect 27157 30240 27169 30243
rect 27120 30212 27169 30240
rect 27120 30200 27126 30212
rect 27157 30209 27169 30212
rect 27203 30209 27215 30243
rect 27157 30203 27215 30209
rect 27246 30200 27252 30252
rect 27304 30240 27310 30252
rect 27540 30249 27568 30280
rect 27525 30243 27583 30249
rect 27304 30212 27349 30240
rect 27304 30200 27310 30212
rect 27525 30209 27537 30243
rect 27571 30209 27583 30243
rect 27525 30203 27583 30209
rect 21174 30172 21180 30184
rect 20824 30144 20944 30172
rect 21135 30144 21180 30172
rect 20916 30104 20944 30144
rect 21174 30132 21180 30144
rect 21232 30132 21238 30184
rect 23842 30132 23848 30184
rect 23900 30172 23906 30184
rect 23937 30175 23995 30181
rect 23937 30172 23949 30175
rect 23900 30144 23949 30172
rect 23900 30132 23906 30144
rect 23937 30141 23949 30144
rect 23983 30141 23995 30175
rect 23937 30135 23995 30141
rect 25501 30175 25559 30181
rect 25501 30141 25513 30175
rect 25547 30141 25559 30175
rect 25501 30135 25559 30141
rect 21358 30104 21364 30116
rect 19904 30076 20484 30104
rect 20916 30076 21364 30104
rect 18509 30039 18567 30045
rect 18509 30005 18521 30039
rect 18555 30005 18567 30039
rect 18509 29999 18567 30005
rect 19150 29996 19156 30048
rect 19208 30036 19214 30048
rect 19904 30036 19932 30076
rect 19208 30008 19932 30036
rect 19208 29996 19214 30008
rect 20254 29996 20260 30048
rect 20312 30036 20318 30048
rect 20349 30039 20407 30045
rect 20349 30036 20361 30039
rect 20312 30008 20361 30036
rect 20312 29996 20318 30008
rect 20349 30005 20361 30008
rect 20395 30005 20407 30039
rect 20456 30036 20484 30076
rect 21358 30064 21364 30076
rect 21416 30064 21422 30116
rect 23750 30064 23756 30116
rect 23808 30104 23814 30116
rect 25516 30104 25544 30135
rect 25958 30132 25964 30184
rect 26016 30172 26022 30184
rect 26878 30172 26884 30184
rect 26016 30144 26884 30172
rect 26016 30132 26022 30144
rect 26878 30132 26884 30144
rect 26936 30172 26942 30184
rect 27341 30175 27399 30181
rect 27341 30172 27353 30175
rect 26936 30144 27353 30172
rect 26936 30132 26942 30144
rect 27341 30141 27353 30144
rect 27387 30141 27399 30175
rect 27341 30135 27399 30141
rect 23808 30076 25544 30104
rect 23808 30064 23814 30076
rect 21085 30039 21143 30045
rect 21085 30036 21097 30039
rect 20456 30008 21097 30036
rect 20349 29999 20407 30005
rect 21085 30005 21097 30008
rect 21131 30005 21143 30039
rect 21085 29999 21143 30005
rect 21269 30039 21327 30045
rect 21269 30005 21281 30039
rect 21315 30036 21327 30039
rect 25314 30036 25320 30048
rect 21315 30008 25320 30036
rect 21315 30005 21327 30008
rect 21269 29999 21327 30005
rect 25314 29996 25320 30008
rect 25372 29996 25378 30048
rect 27246 29996 27252 30048
rect 27304 30036 27310 30048
rect 27709 30039 27767 30045
rect 27709 30036 27721 30039
rect 27304 30008 27721 30036
rect 27304 29996 27310 30008
rect 27709 30005 27721 30008
rect 27755 30005 27767 30039
rect 27709 29999 27767 30005
rect 1104 29946 28888 29968
rect 1104 29894 5582 29946
rect 5634 29894 5646 29946
rect 5698 29894 5710 29946
rect 5762 29894 5774 29946
rect 5826 29894 5838 29946
rect 5890 29894 14846 29946
rect 14898 29894 14910 29946
rect 14962 29894 14974 29946
rect 15026 29894 15038 29946
rect 15090 29894 15102 29946
rect 15154 29894 24110 29946
rect 24162 29894 24174 29946
rect 24226 29894 24238 29946
rect 24290 29894 24302 29946
rect 24354 29894 24366 29946
rect 24418 29894 28888 29946
rect 1104 29872 28888 29894
rect 9217 29835 9275 29841
rect 9217 29801 9229 29835
rect 9263 29832 9275 29835
rect 9306 29832 9312 29844
rect 9263 29804 9312 29832
rect 9263 29801 9275 29804
rect 9217 29795 9275 29801
rect 9306 29792 9312 29804
rect 9364 29792 9370 29844
rect 9398 29792 9404 29844
rect 9456 29832 9462 29844
rect 10410 29832 10416 29844
rect 9456 29804 10416 29832
rect 9456 29792 9462 29804
rect 10410 29792 10416 29804
rect 10468 29792 10474 29844
rect 10502 29792 10508 29844
rect 10560 29832 10566 29844
rect 17678 29832 17684 29844
rect 10560 29804 17684 29832
rect 10560 29792 10566 29804
rect 8205 29767 8263 29773
rect 8205 29733 8217 29767
rect 8251 29764 8263 29767
rect 12158 29764 12164 29776
rect 8251 29736 12164 29764
rect 8251 29733 8263 29736
rect 8205 29727 8263 29733
rect 12158 29724 12164 29736
rect 12216 29724 12222 29776
rect 13446 29724 13452 29776
rect 13504 29764 13510 29776
rect 13541 29767 13599 29773
rect 13541 29764 13553 29767
rect 13504 29736 13553 29764
rect 13504 29724 13510 29736
rect 13541 29733 13553 29736
rect 13587 29733 13599 29767
rect 14642 29764 14648 29776
rect 13541 29727 13599 29733
rect 13740 29736 14648 29764
rect 6730 29656 6736 29708
rect 6788 29696 6794 29708
rect 6788 29668 9352 29696
rect 6788 29656 6794 29668
rect 1394 29588 1400 29640
rect 1452 29628 1458 29640
rect 1581 29631 1639 29637
rect 1581 29628 1593 29631
rect 1452 29600 1593 29628
rect 1452 29588 1458 29600
rect 1581 29597 1593 29600
rect 1627 29597 1639 29631
rect 1581 29591 1639 29597
rect 3878 29588 3884 29640
rect 3936 29628 3942 29640
rect 7558 29628 7564 29640
rect 3936 29600 7564 29628
rect 3936 29588 3942 29600
rect 7558 29588 7564 29600
rect 7616 29588 7622 29640
rect 7745 29631 7803 29637
rect 7745 29597 7757 29631
rect 7791 29597 7803 29631
rect 8386 29628 8392 29640
rect 8347 29600 8392 29628
rect 7745 29591 7803 29597
rect 7760 29560 7788 29591
rect 8386 29588 8392 29600
rect 8444 29588 8450 29640
rect 9214 29560 9220 29572
rect 7760 29532 9220 29560
rect 9214 29520 9220 29532
rect 9272 29520 9278 29572
rect 9324 29560 9352 29668
rect 9416 29668 12296 29696
rect 9416 29637 9444 29668
rect 9401 29631 9459 29637
rect 9401 29597 9413 29631
rect 9447 29597 9459 29631
rect 9401 29591 9459 29597
rect 10045 29631 10103 29637
rect 10045 29597 10057 29631
rect 10091 29628 10103 29631
rect 10134 29628 10140 29640
rect 10091 29600 10140 29628
rect 10091 29597 10103 29600
rect 10045 29591 10103 29597
rect 10134 29588 10140 29600
rect 10192 29588 10198 29640
rect 10229 29631 10287 29637
rect 10229 29597 10241 29631
rect 10275 29597 10287 29631
rect 10229 29591 10287 29597
rect 9674 29560 9680 29572
rect 9324 29532 9680 29560
rect 9674 29520 9680 29532
rect 9732 29520 9738 29572
rect 9769 29563 9827 29569
rect 9769 29529 9781 29563
rect 9815 29560 9827 29563
rect 10244 29560 10272 29591
rect 10410 29588 10416 29640
rect 10468 29628 10474 29640
rect 10689 29631 10747 29637
rect 10689 29628 10701 29631
rect 10468 29600 10701 29628
rect 10468 29588 10474 29600
rect 10689 29597 10701 29600
rect 10735 29597 10747 29631
rect 10689 29591 10747 29597
rect 10778 29588 10784 29640
rect 10836 29628 10842 29640
rect 11146 29628 11152 29640
rect 10836 29600 11152 29628
rect 10836 29588 10842 29600
rect 11146 29588 11152 29600
rect 11204 29588 11210 29640
rect 11425 29631 11483 29637
rect 11425 29597 11437 29631
rect 11471 29597 11483 29631
rect 11425 29591 11483 29597
rect 11440 29560 11468 29591
rect 11514 29588 11520 29640
rect 11572 29628 11578 29640
rect 11698 29628 11704 29640
rect 11572 29600 11617 29628
rect 11659 29600 11704 29628
rect 11572 29588 11578 29600
rect 11698 29588 11704 29600
rect 11756 29588 11762 29640
rect 11790 29588 11796 29640
rect 11848 29628 11854 29640
rect 12158 29628 12164 29640
rect 11848 29600 12164 29628
rect 11848 29588 11854 29600
rect 12158 29588 12164 29600
rect 12216 29588 12222 29640
rect 12268 29630 12296 29668
rect 13170 29656 13176 29708
rect 13228 29696 13234 29708
rect 13740 29696 13768 29736
rect 14642 29724 14648 29736
rect 14700 29724 14706 29776
rect 15746 29724 15752 29776
rect 15804 29764 15810 29776
rect 16117 29767 16175 29773
rect 16117 29764 16129 29767
rect 15804 29736 16129 29764
rect 15804 29724 15810 29736
rect 16117 29733 16129 29736
rect 16163 29764 16175 29767
rect 16206 29764 16212 29776
rect 16163 29736 16212 29764
rect 16163 29733 16175 29736
rect 16117 29727 16175 29733
rect 16206 29724 16212 29736
rect 16264 29724 16270 29776
rect 13228 29668 13768 29696
rect 13228 29656 13234 29668
rect 13998 29656 14004 29708
rect 14056 29696 14062 29708
rect 16592 29705 16620 29804
rect 17678 29792 17684 29804
rect 17736 29792 17742 29844
rect 18601 29835 18659 29841
rect 18601 29832 18613 29835
rect 17926 29804 18613 29832
rect 17586 29724 17592 29776
rect 17644 29764 17650 29776
rect 17926 29764 17954 29804
rect 18601 29801 18613 29804
rect 18647 29801 18659 29835
rect 18601 29795 18659 29801
rect 18874 29792 18880 29844
rect 18932 29832 18938 29844
rect 19978 29832 19984 29844
rect 18932 29804 19984 29832
rect 18932 29792 18938 29804
rect 19978 29792 19984 29804
rect 20036 29792 20042 29844
rect 20714 29792 20720 29844
rect 20772 29832 20778 29844
rect 20898 29832 20904 29844
rect 20772 29804 20904 29832
rect 20772 29792 20778 29804
rect 20898 29792 20904 29804
rect 20956 29792 20962 29844
rect 21174 29792 21180 29844
rect 21232 29832 21238 29844
rect 22094 29832 22100 29844
rect 21232 29804 22100 29832
rect 21232 29792 21238 29804
rect 22094 29792 22100 29804
rect 22152 29792 22158 29844
rect 23845 29835 23903 29841
rect 23845 29801 23857 29835
rect 23891 29832 23903 29835
rect 24026 29832 24032 29844
rect 23891 29804 24032 29832
rect 23891 29801 23903 29804
rect 23845 29795 23903 29801
rect 24026 29792 24032 29804
rect 24084 29792 24090 29844
rect 25774 29832 25780 29844
rect 24136 29804 25780 29832
rect 17644 29736 17954 29764
rect 17644 29724 17650 29736
rect 18414 29724 18420 29776
rect 18472 29764 18478 29776
rect 21542 29764 21548 29776
rect 18472 29736 21548 29764
rect 18472 29724 18478 29736
rect 21542 29724 21548 29736
rect 21600 29724 21606 29776
rect 22278 29724 22284 29776
rect 22336 29764 22342 29776
rect 24136 29764 24164 29804
rect 25774 29792 25780 29804
rect 25832 29792 25838 29844
rect 25869 29835 25927 29841
rect 25869 29801 25881 29835
rect 25915 29832 25927 29835
rect 25958 29832 25964 29844
rect 25915 29804 25964 29832
rect 25915 29801 25927 29804
rect 25869 29795 25927 29801
rect 25958 29792 25964 29804
rect 26016 29792 26022 29844
rect 22336 29736 24164 29764
rect 22336 29724 22342 29736
rect 25590 29724 25596 29776
rect 25648 29764 25654 29776
rect 28258 29764 28264 29776
rect 25648 29736 28264 29764
rect 25648 29724 25654 29736
rect 28258 29724 28264 29736
rect 28316 29724 28322 29776
rect 14737 29699 14795 29705
rect 14737 29696 14749 29699
rect 14056 29668 14749 29696
rect 14056 29656 14062 29668
rect 14737 29665 14749 29668
rect 14783 29665 14795 29699
rect 14737 29659 14795 29665
rect 16577 29699 16635 29705
rect 16577 29665 16589 29699
rect 16623 29665 16635 29699
rect 16577 29659 16635 29665
rect 17862 29656 17868 29708
rect 17920 29696 17926 29708
rect 21726 29696 21732 29708
rect 17920 29668 21732 29696
rect 17920 29656 17926 29668
rect 21726 29656 21732 29668
rect 21784 29656 21790 29708
rect 21910 29696 21916 29708
rect 21871 29668 21916 29696
rect 21910 29656 21916 29668
rect 21968 29656 21974 29708
rect 22830 29656 22836 29708
rect 22888 29696 22894 29708
rect 22888 29668 23336 29696
rect 22888 29656 22894 29668
rect 12268 29628 12388 29630
rect 12452 29628 12572 29630
rect 13814 29628 13820 29640
rect 12268 29602 13820 29628
rect 12360 29600 12480 29602
rect 12544 29600 13820 29602
rect 13814 29588 13820 29600
rect 13872 29588 13878 29640
rect 14090 29628 14096 29640
rect 14051 29600 14096 29628
rect 14090 29588 14096 29600
rect 14148 29588 14154 29640
rect 14185 29631 14243 29637
rect 14185 29597 14197 29631
rect 14231 29628 14243 29631
rect 14231 29600 18644 29628
rect 14231 29597 14243 29600
rect 14185 29591 14243 29597
rect 12250 29560 12256 29572
rect 9815 29532 10916 29560
rect 11440 29532 12256 29560
rect 9815 29529 9827 29532
rect 9769 29523 9827 29529
rect 7561 29495 7619 29501
rect 7561 29461 7573 29495
rect 7607 29492 7619 29495
rect 9122 29492 9128 29504
rect 7607 29464 9128 29492
rect 7607 29461 7619 29464
rect 7561 29455 7619 29461
rect 9122 29452 9128 29464
rect 9180 29452 9186 29504
rect 9398 29452 9404 29504
rect 9456 29492 9462 29504
rect 10137 29495 10195 29501
rect 10137 29492 10149 29495
rect 9456 29464 10149 29492
rect 9456 29452 9462 29464
rect 10137 29461 10149 29464
rect 10183 29461 10195 29495
rect 10778 29492 10784 29504
rect 10739 29464 10784 29492
rect 10137 29455 10195 29461
rect 10778 29452 10784 29464
rect 10836 29452 10842 29504
rect 10888 29492 10916 29532
rect 12250 29520 12256 29532
rect 12308 29520 12314 29572
rect 12428 29563 12486 29569
rect 12428 29529 12440 29563
rect 12474 29560 12486 29563
rect 12526 29560 12532 29572
rect 12474 29532 12532 29560
rect 12474 29529 12486 29532
rect 12428 29523 12486 29529
rect 12526 29520 12532 29532
rect 12584 29520 12590 29572
rect 12618 29520 12624 29572
rect 12676 29560 12682 29572
rect 14982 29563 15040 29569
rect 14982 29560 14994 29563
rect 12676 29532 14994 29560
rect 12676 29520 12682 29532
rect 14982 29529 14994 29532
rect 15028 29529 15040 29563
rect 14982 29523 15040 29529
rect 15654 29520 15660 29572
rect 15712 29560 15718 29572
rect 16822 29563 16880 29569
rect 16822 29560 16834 29563
rect 15712 29532 16834 29560
rect 15712 29520 15718 29532
rect 16822 29529 16834 29532
rect 16868 29529 16880 29563
rect 17862 29560 17868 29572
rect 16822 29523 16880 29529
rect 16929 29532 17868 29560
rect 16929 29492 16957 29532
rect 17862 29520 17868 29532
rect 17920 29520 17926 29572
rect 18509 29563 18567 29569
rect 18509 29529 18521 29563
rect 18555 29529 18567 29563
rect 18616 29560 18644 29600
rect 19242 29588 19248 29640
rect 19300 29628 19306 29640
rect 19300 29600 19345 29628
rect 19300 29588 19306 29600
rect 19426 29588 19432 29640
rect 19484 29628 19490 29640
rect 20346 29628 20352 29640
rect 19484 29600 19529 29628
rect 20307 29600 20352 29628
rect 19484 29588 19490 29600
rect 20346 29588 20352 29600
rect 20404 29588 20410 29640
rect 22370 29588 22376 29640
rect 22428 29628 22434 29640
rect 23308 29637 23336 29668
rect 24394 29656 24400 29708
rect 24452 29696 24458 29708
rect 24489 29699 24547 29705
rect 24489 29696 24501 29699
rect 24452 29668 24501 29696
rect 24452 29656 24458 29668
rect 24489 29665 24501 29668
rect 24535 29665 24547 29699
rect 24489 29659 24547 29665
rect 25866 29656 25872 29708
rect 25924 29696 25930 29708
rect 26789 29699 26847 29705
rect 26789 29696 26801 29699
rect 25924 29668 26801 29696
rect 25924 29656 25930 29668
rect 26789 29665 26801 29668
rect 26835 29665 26847 29699
rect 26789 29659 26847 29665
rect 23201 29631 23259 29637
rect 23201 29628 23213 29631
rect 22428 29600 23213 29628
rect 22428 29588 22434 29600
rect 23201 29597 23213 29600
rect 23247 29597 23259 29631
rect 23201 29591 23259 29597
rect 23294 29631 23352 29637
rect 23294 29597 23306 29631
rect 23340 29597 23352 29631
rect 23294 29591 23352 29597
rect 23474 29588 23480 29640
rect 23532 29628 23538 29640
rect 23707 29631 23765 29637
rect 23532 29600 23577 29628
rect 23532 29588 23538 29600
rect 23707 29597 23719 29631
rect 23753 29628 23765 29631
rect 23934 29628 23940 29640
rect 23753 29600 23940 29628
rect 23753 29597 23765 29600
rect 23707 29591 23765 29597
rect 23934 29588 23940 29600
rect 23992 29588 23998 29640
rect 24756 29631 24814 29637
rect 24756 29597 24768 29631
rect 24802 29628 24814 29631
rect 25038 29628 25044 29640
rect 24802 29600 25044 29628
rect 24802 29597 24814 29600
rect 24756 29591 24814 29597
rect 25038 29588 25044 29600
rect 25096 29588 25102 29640
rect 26326 29628 26332 29640
rect 26287 29600 26332 29628
rect 26326 29588 26332 29600
rect 26384 29588 26390 29640
rect 18616 29532 19932 29560
rect 18509 29523 18567 29529
rect 17954 29492 17960 29504
rect 10888 29464 16957 29492
rect 17915 29464 17960 29492
rect 17954 29452 17960 29464
rect 18012 29452 18018 29504
rect 18322 29452 18328 29504
rect 18380 29492 18386 29504
rect 18524 29492 18552 29523
rect 18380 29464 18552 29492
rect 18380 29452 18386 29464
rect 18874 29452 18880 29504
rect 18932 29492 18938 29504
rect 19613 29495 19671 29501
rect 19613 29492 19625 29495
rect 18932 29464 19625 29492
rect 18932 29452 18938 29464
rect 19613 29461 19625 29464
rect 19659 29461 19671 29495
rect 19904 29492 19932 29532
rect 19978 29520 19984 29572
rect 20036 29560 20042 29572
rect 20533 29563 20591 29569
rect 20533 29560 20545 29563
rect 20036 29532 20545 29560
rect 20036 29520 20042 29532
rect 20533 29529 20545 29532
rect 20579 29529 20591 29563
rect 20533 29523 20591 29529
rect 23382 29520 23388 29572
rect 23440 29560 23446 29572
rect 23569 29563 23627 29569
rect 23569 29560 23581 29563
rect 23440 29532 23581 29560
rect 23440 29520 23446 29532
rect 23569 29529 23581 29532
rect 23615 29529 23627 29563
rect 26513 29563 26571 29569
rect 26513 29560 26525 29563
rect 23569 29523 23627 29529
rect 23676 29532 26525 29560
rect 23676 29492 23704 29532
rect 26513 29529 26525 29532
rect 26559 29529 26571 29563
rect 26513 29523 26571 29529
rect 19904 29464 23704 29492
rect 19613 29455 19671 29461
rect 1104 29402 28888 29424
rect 1104 29350 10214 29402
rect 10266 29350 10278 29402
rect 10330 29350 10342 29402
rect 10394 29350 10406 29402
rect 10458 29350 10470 29402
rect 10522 29350 19478 29402
rect 19530 29350 19542 29402
rect 19594 29350 19606 29402
rect 19658 29350 19670 29402
rect 19722 29350 19734 29402
rect 19786 29350 28888 29402
rect 1104 29328 28888 29350
rect 9214 29248 9220 29300
rect 9272 29288 9278 29300
rect 10686 29288 10692 29300
rect 9272 29260 10692 29288
rect 9272 29248 9278 29260
rect 10686 29248 10692 29260
rect 10744 29248 10750 29300
rect 10778 29248 10784 29300
rect 10836 29288 10842 29300
rect 13722 29288 13728 29300
rect 10836 29260 13728 29288
rect 10836 29248 10842 29260
rect 13722 29248 13728 29260
rect 13780 29248 13786 29300
rect 13814 29248 13820 29300
rect 13872 29288 13878 29300
rect 18874 29288 18880 29300
rect 13872 29260 18880 29288
rect 13872 29248 13878 29260
rect 18874 29248 18880 29260
rect 18932 29248 18938 29300
rect 19058 29248 19064 29300
rect 19116 29288 19122 29300
rect 21542 29288 21548 29300
rect 19116 29260 21548 29288
rect 19116 29248 19122 29260
rect 21542 29248 21548 29260
rect 21600 29248 21606 29300
rect 21726 29248 21732 29300
rect 21784 29288 21790 29300
rect 24946 29288 24952 29300
rect 21784 29260 24952 29288
rect 21784 29248 21790 29260
rect 24946 29248 24952 29260
rect 25004 29248 25010 29300
rect 26786 29248 26792 29300
rect 26844 29288 26850 29300
rect 27065 29291 27123 29297
rect 27065 29288 27077 29291
rect 26844 29260 27077 29288
rect 26844 29248 26850 29260
rect 27065 29257 27077 29260
rect 27111 29257 27123 29291
rect 27065 29251 27123 29257
rect 10870 29220 10876 29232
rect 9048 29192 10876 29220
rect 1394 29152 1400 29164
rect 1355 29124 1400 29152
rect 1394 29112 1400 29124
rect 1452 29112 1458 29164
rect 9048 29161 9076 29192
rect 10870 29180 10876 29192
rect 10928 29180 10934 29232
rect 11790 29220 11796 29232
rect 11348 29192 11796 29220
rect 8389 29155 8447 29161
rect 8389 29121 8401 29155
rect 8435 29121 8447 29155
rect 8389 29115 8447 29121
rect 9033 29155 9091 29161
rect 9033 29121 9045 29155
rect 9079 29121 9091 29155
rect 9033 29115 9091 29121
rect 9677 29155 9735 29161
rect 9677 29121 9689 29155
rect 9723 29152 9735 29155
rect 10042 29152 10048 29164
rect 9723 29124 10048 29152
rect 9723 29121 9735 29124
rect 9677 29115 9735 29121
rect 1578 29084 1584 29096
rect 1539 29056 1584 29084
rect 1578 29044 1584 29056
rect 1636 29044 1642 29096
rect 2774 29044 2780 29096
rect 2832 29084 2838 29096
rect 8404 29084 8432 29115
rect 10042 29112 10048 29124
rect 10100 29112 10106 29164
rect 10137 29155 10195 29161
rect 10137 29121 10149 29155
rect 10183 29152 10195 29155
rect 10226 29152 10232 29164
rect 10183 29124 10232 29152
rect 10183 29121 10195 29124
rect 10137 29115 10195 29121
rect 10226 29112 10232 29124
rect 10284 29112 10290 29164
rect 10321 29155 10379 29161
rect 10321 29121 10333 29155
rect 10367 29152 10379 29155
rect 10410 29152 10416 29164
rect 10367 29124 10416 29152
rect 10367 29121 10379 29124
rect 10321 29115 10379 29121
rect 10410 29112 10416 29124
rect 10468 29112 10474 29164
rect 10502 29112 10508 29164
rect 10560 29152 10566 29164
rect 10781 29155 10839 29161
rect 10781 29152 10793 29155
rect 10560 29124 10793 29152
rect 10560 29112 10566 29124
rect 10781 29121 10793 29124
rect 10827 29121 10839 29155
rect 11348 29152 11376 29192
rect 11790 29180 11796 29192
rect 11848 29180 11854 29232
rect 11885 29223 11943 29229
rect 11885 29189 11897 29223
rect 11931 29220 11943 29223
rect 12250 29220 12256 29232
rect 11931 29192 12256 29220
rect 11931 29189 11943 29192
rect 11885 29183 11943 29189
rect 10781 29115 10839 29121
rect 10980 29124 11376 29152
rect 10980 29084 11008 29124
rect 11422 29112 11428 29164
rect 11480 29152 11486 29164
rect 11900 29152 11928 29183
rect 12250 29180 12256 29192
rect 12308 29180 12314 29232
rect 14090 29220 14096 29232
rect 12544 29192 14096 29220
rect 11480 29124 11928 29152
rect 11480 29112 11486 29124
rect 12158 29112 12164 29164
rect 12216 29152 12222 29164
rect 12544 29161 12572 29192
rect 14090 29180 14096 29192
rect 14148 29180 14154 29232
rect 14182 29180 14188 29232
rect 14240 29220 14246 29232
rect 15562 29220 15568 29232
rect 14240 29192 15568 29220
rect 14240 29180 14246 29192
rect 15562 29180 15568 29192
rect 15620 29180 15626 29232
rect 15657 29223 15715 29229
rect 15657 29189 15669 29223
rect 15703 29220 15715 29223
rect 15746 29220 15752 29232
rect 15703 29192 15752 29220
rect 15703 29189 15715 29192
rect 15657 29183 15715 29189
rect 15746 29180 15752 29192
rect 15804 29180 15810 29232
rect 16114 29220 16120 29232
rect 15856 29192 16120 29220
rect 12529 29155 12587 29161
rect 12529 29152 12541 29155
rect 12216 29124 12541 29152
rect 12216 29112 12222 29124
rect 12529 29121 12541 29124
rect 12575 29121 12587 29155
rect 12785 29155 12843 29161
rect 12785 29152 12797 29155
rect 12529 29115 12587 29121
rect 12636 29124 12797 29152
rect 11514 29084 11520 29096
rect 2832 29056 2877 29084
rect 8404 29056 11008 29084
rect 11064 29056 11520 29084
rect 2832 29044 2838 29056
rect 7742 29016 7748 29028
rect 7703 28988 7748 29016
rect 7742 28976 7748 28988
rect 7800 28976 7806 29028
rect 8205 29019 8263 29025
rect 8205 28985 8217 29019
rect 8251 29016 8263 29019
rect 11064 29016 11092 29056
rect 11514 29044 11520 29056
rect 11572 29044 11578 29096
rect 11606 29044 11612 29096
rect 11664 29084 11670 29096
rect 12636 29084 12664 29124
rect 12785 29121 12797 29124
rect 12831 29121 12843 29155
rect 12785 29115 12843 29121
rect 13078 29112 13084 29164
rect 13136 29152 13142 29164
rect 14921 29155 14979 29161
rect 13136 29124 13584 29152
rect 13136 29112 13142 29124
rect 11664 29056 12664 29084
rect 13556 29084 13584 29124
rect 14921 29121 14933 29155
rect 14967 29121 14979 29155
rect 14921 29115 14979 29121
rect 14936 29084 14964 29115
rect 15010 29112 15016 29164
rect 15068 29152 15074 29164
rect 15856 29161 15884 29192
rect 16114 29180 16120 29192
rect 16172 29220 16178 29232
rect 17954 29220 17960 29232
rect 16172 29192 17960 29220
rect 16172 29180 16178 29192
rect 17954 29180 17960 29192
rect 18012 29180 18018 29232
rect 18046 29180 18052 29232
rect 18104 29220 18110 29232
rect 22094 29220 22100 29232
rect 18104 29192 22100 29220
rect 18104 29180 18110 29192
rect 22094 29180 22100 29192
rect 22152 29180 22158 29232
rect 23474 29180 23480 29232
rect 23532 29220 23538 29232
rect 23532 29192 25360 29220
rect 23532 29180 23538 29192
rect 15841 29155 15899 29161
rect 15068 29124 15113 29152
rect 15068 29112 15074 29124
rect 15841 29121 15853 29155
rect 15887 29121 15899 29155
rect 15841 29115 15899 29121
rect 15933 29155 15991 29161
rect 15933 29121 15945 29155
rect 15979 29152 15991 29155
rect 16298 29152 16304 29164
rect 15979 29124 16304 29152
rect 15979 29121 15991 29124
rect 15933 29115 15991 29121
rect 16298 29112 16304 29124
rect 16356 29112 16362 29164
rect 16669 29155 16727 29161
rect 16669 29121 16681 29155
rect 16715 29121 16727 29155
rect 16669 29115 16727 29121
rect 16684 29084 16712 29115
rect 16758 29112 16764 29164
rect 16816 29152 16822 29164
rect 17661 29155 17719 29161
rect 17661 29152 17673 29155
rect 16816 29124 17673 29152
rect 16816 29112 16822 29124
rect 17661 29121 17673 29124
rect 17707 29121 17719 29155
rect 17661 29115 17719 29121
rect 18138 29112 18144 29164
rect 18196 29152 18202 29164
rect 19961 29155 20019 29161
rect 19961 29152 19973 29155
rect 18196 29124 19973 29152
rect 18196 29112 18202 29124
rect 19961 29121 19973 29124
rect 20007 29121 20019 29155
rect 19961 29115 20019 29121
rect 22002 29112 22008 29164
rect 22060 29112 22066 29164
rect 22189 29155 22247 29161
rect 22189 29121 22201 29155
rect 22235 29152 22247 29155
rect 22278 29152 22284 29164
rect 22235 29124 22284 29152
rect 22235 29121 22247 29124
rect 22189 29115 22247 29121
rect 22278 29112 22284 29124
rect 22336 29112 22342 29164
rect 22646 29152 22652 29164
rect 22572 29124 22652 29152
rect 16850 29084 16856 29096
rect 13556 29056 14841 29084
rect 14936 29056 16620 29084
rect 16684 29056 16856 29084
rect 11664 29044 11670 29056
rect 8251 28988 11092 29016
rect 8251 28985 8263 28988
rect 8205 28979 8263 28985
rect 11330 28976 11336 29028
rect 11388 29016 11394 29028
rect 12069 29019 12127 29025
rect 12069 29016 12081 29019
rect 11388 28988 12081 29016
rect 11388 28976 11394 28988
rect 12069 28985 12081 28988
rect 12115 29016 12127 29019
rect 12526 29016 12532 29028
rect 12115 28988 12532 29016
rect 12115 28985 12127 28988
rect 12069 28979 12127 28985
rect 12526 28976 12532 28988
rect 12584 28976 12590 29028
rect 13630 28976 13636 29028
rect 13688 29016 13694 29028
rect 14813 29016 14841 29056
rect 15654 29016 15660 29028
rect 13688 28988 14136 29016
rect 14813 28988 15660 29016
rect 13688 28976 13694 28988
rect 8849 28951 8907 28957
rect 8849 28917 8861 28951
rect 8895 28948 8907 28951
rect 9122 28948 9128 28960
rect 8895 28920 9128 28948
rect 8895 28917 8907 28920
rect 8849 28911 8907 28917
rect 9122 28908 9128 28920
rect 9180 28908 9186 28960
rect 9490 28948 9496 28960
rect 9451 28920 9496 28948
rect 9490 28908 9496 28920
rect 9548 28908 9554 28960
rect 10134 28948 10140 28960
rect 10095 28920 10140 28948
rect 10134 28908 10140 28920
rect 10192 28908 10198 28960
rect 10873 28951 10931 28957
rect 10873 28917 10885 28951
rect 10919 28948 10931 28951
rect 11422 28948 11428 28960
rect 10919 28920 11428 28948
rect 10919 28917 10931 28920
rect 10873 28911 10931 28917
rect 11422 28908 11428 28920
rect 11480 28908 11486 28960
rect 13906 28908 13912 28960
rect 13964 28948 13970 28960
rect 14108 28948 14136 28988
rect 15654 28976 15660 28988
rect 15712 28976 15718 29028
rect 16117 29019 16175 29025
rect 16117 29016 16129 29019
rect 15764 28988 16129 29016
rect 15197 28951 15255 28957
rect 15197 28948 15209 28951
rect 13964 28920 14009 28948
rect 14108 28920 15209 28948
rect 13964 28908 13970 28920
rect 15197 28917 15209 28920
rect 15243 28917 15255 28951
rect 15197 28911 15255 28917
rect 15562 28908 15568 28960
rect 15620 28948 15626 28960
rect 15764 28948 15792 28988
rect 16117 28985 16129 28988
rect 16163 28985 16175 29019
rect 16592 29016 16620 29056
rect 16850 29044 16856 29056
rect 16908 29044 16914 29096
rect 17034 29044 17040 29096
rect 17092 29084 17098 29096
rect 17405 29087 17463 29093
rect 17405 29084 17417 29087
rect 17092 29056 17417 29084
rect 17092 29044 17098 29056
rect 17405 29053 17417 29056
rect 17451 29053 17463 29087
rect 17405 29047 17463 29053
rect 18414 29044 18420 29096
rect 18472 29084 18478 29096
rect 18472 29056 19656 29084
rect 18472 29044 18478 29056
rect 17218 29016 17224 29028
rect 16592 28988 17224 29016
rect 16117 28979 16175 28985
rect 17218 28976 17224 28988
rect 17276 28976 17282 29028
rect 18782 29016 18788 29028
rect 18743 28988 18788 29016
rect 18782 28976 18788 28988
rect 18840 28976 18846 29028
rect 15620 28920 15792 28948
rect 15933 28951 15991 28957
rect 15620 28908 15626 28920
rect 15933 28917 15945 28951
rect 15979 28948 15991 28951
rect 16022 28948 16028 28960
rect 15979 28920 16028 28948
rect 15979 28917 15991 28920
rect 15933 28911 15991 28917
rect 16022 28908 16028 28920
rect 16080 28908 16086 28960
rect 16853 28951 16911 28957
rect 16853 28917 16865 28951
rect 16899 28948 16911 28951
rect 16942 28948 16948 28960
rect 16899 28920 16948 28948
rect 16899 28917 16911 28920
rect 16853 28911 16911 28917
rect 16942 28908 16948 28920
rect 17000 28908 17006 28960
rect 17126 28908 17132 28960
rect 17184 28948 17190 28960
rect 18322 28948 18328 28960
rect 17184 28920 18328 28948
rect 17184 28908 17190 28920
rect 18322 28908 18328 28920
rect 18380 28908 18386 28960
rect 19628 28948 19656 29056
rect 19702 29044 19708 29096
rect 19760 29084 19766 29096
rect 21726 29084 21732 29096
rect 19760 29056 19805 29084
rect 20732 29056 21732 29084
rect 19760 29044 19766 29056
rect 20732 29016 20760 29056
rect 21726 29044 21732 29056
rect 21784 29044 21790 29096
rect 20640 28988 20760 29016
rect 20640 28948 20668 28988
rect 19628 28920 20668 28948
rect 21085 28951 21143 28957
rect 21085 28917 21097 28951
rect 21131 28948 21143 28951
rect 21174 28948 21180 28960
rect 21131 28920 21180 28948
rect 21131 28917 21143 28920
rect 21085 28911 21143 28917
rect 21174 28908 21180 28920
rect 21232 28908 21238 28960
rect 21358 28908 21364 28960
rect 21416 28948 21422 28960
rect 21910 28948 21916 28960
rect 21416 28920 21916 28948
rect 21416 28908 21422 28920
rect 21910 28908 21916 28920
rect 21968 28908 21974 28960
rect 22020 28957 22048 29112
rect 22465 29087 22523 29093
rect 22465 29053 22477 29087
rect 22511 29084 22523 29087
rect 22572 29084 22600 29124
rect 22646 29112 22652 29124
rect 22704 29152 22710 29164
rect 22922 29152 22928 29164
rect 22704 29124 22928 29152
rect 22704 29112 22710 29124
rect 22922 29112 22928 29124
rect 22980 29112 22986 29164
rect 23017 29155 23075 29161
rect 23017 29121 23029 29155
rect 23063 29152 23075 29155
rect 23198 29152 23204 29164
rect 23063 29124 23204 29152
rect 23063 29121 23075 29124
rect 23017 29115 23075 29121
rect 23198 29112 23204 29124
rect 23256 29112 23262 29164
rect 23290 29112 23296 29164
rect 23348 29152 23354 29164
rect 23348 29124 23393 29152
rect 23348 29112 23354 29124
rect 23566 29112 23572 29164
rect 23624 29152 23630 29164
rect 24305 29155 24363 29161
rect 24305 29152 24317 29155
rect 23624 29124 24317 29152
rect 23624 29112 23630 29124
rect 24305 29121 24317 29124
rect 24351 29152 24363 29155
rect 24394 29152 24400 29164
rect 24351 29124 24400 29152
rect 24351 29121 24363 29124
rect 24305 29115 24363 29121
rect 24394 29112 24400 29124
rect 24452 29112 24458 29164
rect 24578 29161 24584 29164
rect 24572 29115 24584 29161
rect 24636 29152 24642 29164
rect 24636 29124 24672 29152
rect 24578 29112 24584 29115
rect 24636 29112 24642 29124
rect 22511 29056 22600 29084
rect 22511 29053 22523 29056
rect 22465 29047 22523 29053
rect 22830 29044 22836 29096
rect 22888 29084 22894 29096
rect 23308 29084 23336 29112
rect 22888 29056 23336 29084
rect 22888 29044 22894 29056
rect 23382 29044 23388 29096
rect 23440 29084 23446 29096
rect 25332 29084 25360 29192
rect 26326 29180 26332 29232
rect 26384 29220 26390 29232
rect 27433 29223 27491 29229
rect 27433 29220 27445 29223
rect 26384 29192 27445 29220
rect 26384 29180 26390 29192
rect 27433 29189 27445 29192
rect 27479 29189 27491 29223
rect 27433 29183 27491 29189
rect 26050 29112 26056 29164
rect 26108 29152 26114 29164
rect 26145 29155 26203 29161
rect 26145 29152 26157 29155
rect 26108 29124 26157 29152
rect 26108 29112 26114 29124
rect 26145 29121 26157 29124
rect 26191 29121 26203 29155
rect 26145 29115 26203 29121
rect 26878 29112 26884 29164
rect 26936 29152 26942 29164
rect 26973 29155 27031 29161
rect 26973 29152 26985 29155
rect 26936 29124 26985 29152
rect 26936 29112 26942 29124
rect 26973 29121 26985 29124
rect 27019 29121 27031 29155
rect 27246 29152 27252 29164
rect 27207 29124 27252 29152
rect 26973 29115 27031 29121
rect 27246 29112 27252 29124
rect 27304 29112 27310 29164
rect 27893 29155 27951 29161
rect 27893 29121 27905 29155
rect 27939 29121 27951 29155
rect 27893 29115 27951 29121
rect 27341 29087 27399 29093
rect 27341 29084 27353 29087
rect 23440 29056 24348 29084
rect 25332 29056 27353 29084
rect 23440 29044 23446 29056
rect 22005 28951 22063 28957
rect 22005 28917 22017 28951
rect 22051 28917 22063 28951
rect 22005 28911 22063 28917
rect 22278 28908 22284 28960
rect 22336 28948 22342 28960
rect 22373 28951 22431 28957
rect 22373 28948 22385 28951
rect 22336 28920 22385 28948
rect 22336 28908 22342 28920
rect 22373 28917 22385 28920
rect 22419 28948 22431 28951
rect 22830 28948 22836 28960
rect 22419 28920 22836 28948
rect 22419 28917 22431 28920
rect 22373 28911 22431 28917
rect 22830 28908 22836 28920
rect 22888 28908 22894 28960
rect 22922 28908 22928 28960
rect 22980 28948 22986 28960
rect 23290 28948 23296 28960
rect 22980 28920 23296 28948
rect 22980 28908 22986 28920
rect 23290 28908 23296 28920
rect 23348 28908 23354 28960
rect 24320 28948 24348 29056
rect 27341 29053 27353 29056
rect 27387 29053 27399 29087
rect 27341 29047 27399 29053
rect 25406 28976 25412 29028
rect 25464 29016 25470 29028
rect 25685 29019 25743 29025
rect 25685 29016 25697 29019
rect 25464 28988 25697 29016
rect 25464 28976 25470 28988
rect 25685 28985 25697 28988
rect 25731 29016 25743 29019
rect 25866 29016 25872 29028
rect 25731 28988 25872 29016
rect 25731 28985 25743 28988
rect 25685 28979 25743 28985
rect 25866 28976 25872 28988
rect 25924 28976 25930 29028
rect 26050 28976 26056 29028
rect 26108 29016 26114 29028
rect 27908 29016 27936 29115
rect 26108 28988 27936 29016
rect 28077 29019 28135 29025
rect 26108 28976 26114 28988
rect 28077 28985 28089 29019
rect 28123 29016 28135 29019
rect 28626 29016 28632 29028
rect 28123 28988 28632 29016
rect 28123 28985 28135 28988
rect 28077 28979 28135 28985
rect 28626 28976 28632 28988
rect 28684 28976 28690 29028
rect 26329 28951 26387 28957
rect 26329 28948 26341 28951
rect 24320 28920 26341 28948
rect 26329 28917 26341 28920
rect 26375 28948 26387 28951
rect 27614 28948 27620 28960
rect 26375 28920 27620 28948
rect 26375 28917 26387 28920
rect 26329 28911 26387 28917
rect 27614 28908 27620 28920
rect 27672 28908 27678 28960
rect 1104 28858 28888 28880
rect 1104 28806 5582 28858
rect 5634 28806 5646 28858
rect 5698 28806 5710 28858
rect 5762 28806 5774 28858
rect 5826 28806 5838 28858
rect 5890 28806 14846 28858
rect 14898 28806 14910 28858
rect 14962 28806 14974 28858
rect 15026 28806 15038 28858
rect 15090 28806 15102 28858
rect 15154 28806 24110 28858
rect 24162 28806 24174 28858
rect 24226 28806 24238 28858
rect 24290 28806 24302 28858
rect 24354 28806 24366 28858
rect 24418 28806 28888 28858
rect 1104 28784 28888 28806
rect 1578 28704 1584 28756
rect 1636 28744 1642 28756
rect 1673 28747 1731 28753
rect 1673 28744 1685 28747
rect 1636 28716 1685 28744
rect 1636 28704 1642 28716
rect 1673 28713 1685 28716
rect 1719 28713 1731 28747
rect 10594 28744 10600 28756
rect 1673 28707 1731 28713
rect 9416 28716 10600 28744
rect 8846 28608 8852 28620
rect 2746 28580 8852 28608
rect 1581 28543 1639 28549
rect 1581 28509 1593 28543
rect 1627 28540 1639 28543
rect 1670 28540 1676 28552
rect 1627 28512 1676 28540
rect 1627 28509 1639 28512
rect 1581 28503 1639 28509
rect 1670 28500 1676 28512
rect 1728 28540 1734 28552
rect 2746 28540 2774 28580
rect 8846 28568 8852 28580
rect 8904 28568 8910 28620
rect 1728 28512 2774 28540
rect 8389 28543 8447 28549
rect 1728 28500 1734 28512
rect 8389 28509 8401 28543
rect 8435 28540 8447 28543
rect 8754 28540 8760 28552
rect 8435 28512 8760 28540
rect 8435 28509 8447 28512
rect 8389 28503 8447 28509
rect 8754 28500 8760 28512
rect 8812 28500 8818 28552
rect 9416 28549 9444 28716
rect 10594 28704 10600 28716
rect 10652 28704 10658 28756
rect 10689 28747 10747 28753
rect 10689 28713 10701 28747
rect 10735 28713 10747 28747
rect 10689 28707 10747 28713
rect 10704 28676 10732 28707
rect 10870 28704 10876 28756
rect 10928 28744 10934 28756
rect 10928 28716 12296 28744
rect 10928 28704 10934 28716
rect 11054 28676 11060 28688
rect 10704 28648 11060 28676
rect 11054 28636 11060 28648
rect 11112 28636 11118 28688
rect 10226 28568 10232 28620
rect 10284 28608 10290 28620
rect 10594 28608 10600 28620
rect 10284 28580 10600 28608
rect 10284 28568 10290 28580
rect 10594 28568 10600 28580
rect 10652 28568 10658 28620
rect 11238 28617 11244 28620
rect 11230 28611 11244 28617
rect 11230 28608 11242 28611
rect 11199 28580 11242 28608
rect 11230 28577 11242 28580
rect 11230 28571 11244 28577
rect 11238 28568 11244 28571
rect 11296 28568 11302 28620
rect 12268 28608 12296 28716
rect 12342 28704 12348 28756
rect 12400 28744 12406 28756
rect 12400 28716 16574 28744
rect 12400 28704 12406 28716
rect 12434 28636 12440 28688
rect 12492 28676 12498 28688
rect 16209 28679 16267 28685
rect 16209 28676 16221 28679
rect 12492 28648 16221 28676
rect 12492 28636 12498 28648
rect 16209 28645 16221 28648
rect 16255 28645 16267 28679
rect 16546 28676 16574 28716
rect 17862 28704 17868 28756
rect 17920 28744 17926 28756
rect 17957 28747 18015 28753
rect 17957 28744 17969 28747
rect 17920 28716 17969 28744
rect 17920 28704 17926 28716
rect 17957 28713 17969 28716
rect 18003 28713 18015 28747
rect 17957 28707 18015 28713
rect 18322 28704 18328 28756
rect 18380 28744 18386 28756
rect 18380 28716 20300 28744
rect 18380 28704 18386 28716
rect 19886 28676 19892 28688
rect 16546 28648 19892 28676
rect 16209 28639 16267 28645
rect 19886 28636 19892 28648
rect 19944 28636 19950 28688
rect 20272 28624 20300 28716
rect 22002 28704 22008 28756
rect 22060 28744 22066 28756
rect 23109 28747 23167 28753
rect 22060 28716 22692 28744
rect 22060 28704 22066 28716
rect 21542 28636 21548 28688
rect 21600 28676 21606 28688
rect 21726 28676 21732 28688
rect 21600 28648 21732 28676
rect 21600 28636 21606 28648
rect 21726 28636 21732 28648
rect 21784 28636 21790 28688
rect 22664 28676 22692 28716
rect 23109 28713 23121 28747
rect 23155 28744 23167 28747
rect 23198 28744 23204 28756
rect 23155 28716 23204 28744
rect 23155 28713 23167 28716
rect 23109 28707 23167 28713
rect 23198 28704 23204 28716
rect 23256 28704 23262 28756
rect 27614 28744 27620 28756
rect 24412 28716 27620 28744
rect 24412 28676 24440 28716
rect 27614 28704 27620 28716
rect 27672 28704 27678 28756
rect 22664 28648 24440 28676
rect 13354 28608 13360 28620
rect 12268 28580 13360 28608
rect 13354 28568 13360 28580
rect 13412 28568 13418 28620
rect 13449 28611 13507 28617
rect 13449 28577 13461 28611
rect 13495 28608 13507 28611
rect 13722 28608 13728 28620
rect 13495 28580 13728 28608
rect 13495 28577 13507 28580
rect 13449 28571 13507 28577
rect 13722 28568 13728 28580
rect 13780 28568 13786 28620
rect 14182 28568 14188 28620
rect 14240 28608 14246 28620
rect 15841 28611 15899 28617
rect 15841 28608 15853 28611
rect 14240 28580 15853 28608
rect 14240 28568 14246 28580
rect 15841 28577 15853 28580
rect 15887 28577 15899 28611
rect 16669 28611 16727 28617
rect 16669 28608 16681 28611
rect 15841 28571 15899 28577
rect 15948 28580 16681 28608
rect 9401 28543 9459 28549
rect 9401 28509 9413 28543
rect 9447 28509 9459 28543
rect 9401 28503 9459 28509
rect 9861 28543 9919 28549
rect 9861 28509 9873 28543
rect 9907 28509 9919 28543
rect 10042 28540 10048 28552
rect 10003 28512 10048 28540
rect 9861 28503 9919 28509
rect 8202 28404 8208 28416
rect 8163 28376 8208 28404
rect 8202 28364 8208 28376
rect 8260 28364 8266 28416
rect 9214 28404 9220 28416
rect 9175 28376 9220 28404
rect 9214 28364 9220 28376
rect 9272 28364 9278 28416
rect 9876 28404 9904 28503
rect 10042 28500 10048 28512
rect 10100 28500 10106 28552
rect 10520 28512 11275 28540
rect 9953 28475 10011 28481
rect 9953 28441 9965 28475
rect 9999 28472 10011 28475
rect 10520 28472 10548 28512
rect 9999 28444 10548 28472
rect 10597 28475 10655 28481
rect 9999 28441 10011 28444
rect 9953 28435 10011 28441
rect 10597 28441 10609 28475
rect 10643 28472 10655 28475
rect 10686 28472 10692 28484
rect 10643 28444 10692 28472
rect 10643 28441 10655 28444
rect 10597 28435 10655 28441
rect 10686 28432 10692 28444
rect 10744 28432 10750 28484
rect 11247 28472 11275 28512
rect 11330 28500 11336 28552
rect 11388 28540 11394 28552
rect 11497 28543 11555 28549
rect 11497 28540 11509 28543
rect 11388 28512 11509 28540
rect 11388 28500 11394 28512
rect 11497 28509 11509 28512
rect 11543 28509 11555 28543
rect 12894 28540 12900 28552
rect 11497 28503 11555 28509
rect 11624 28512 12900 28540
rect 11624 28484 11652 28512
rect 12894 28500 12900 28512
rect 12952 28500 12958 28552
rect 13078 28500 13084 28552
rect 13136 28540 13142 28552
rect 13265 28543 13323 28549
rect 13265 28540 13277 28543
rect 13136 28512 13277 28540
rect 13136 28500 13142 28512
rect 13265 28509 13277 28512
rect 13311 28509 13323 28543
rect 13538 28540 13544 28552
rect 13499 28512 13544 28540
rect 13265 28503 13323 28509
rect 13538 28500 13544 28512
rect 13596 28500 13602 28552
rect 14093 28543 14151 28549
rect 14093 28509 14105 28543
rect 14139 28540 14151 28543
rect 14366 28540 14372 28552
rect 14139 28512 14372 28540
rect 14139 28509 14151 28512
rect 14093 28503 14151 28509
rect 14366 28500 14372 28512
rect 14424 28540 14430 28552
rect 14642 28540 14648 28552
rect 14424 28512 14648 28540
rect 14424 28500 14430 28512
rect 14642 28500 14648 28512
rect 14700 28500 14706 28552
rect 14734 28500 14740 28552
rect 14792 28540 14798 28552
rect 14921 28543 14979 28549
rect 14792 28512 14837 28540
rect 14792 28500 14798 28512
rect 14921 28509 14933 28543
rect 14967 28540 14979 28543
rect 15948 28540 15976 28580
rect 16669 28577 16681 28580
rect 16715 28608 16727 28611
rect 17126 28608 17132 28620
rect 16715 28580 17132 28608
rect 16715 28577 16727 28580
rect 16669 28571 16727 28577
rect 17126 28568 17132 28580
rect 17184 28568 17190 28620
rect 17494 28568 17500 28620
rect 17552 28608 17558 28620
rect 17552 28580 18276 28608
rect 17552 28568 17558 28580
rect 14967 28512 15976 28540
rect 16025 28543 16083 28549
rect 14967 28509 14979 28512
rect 14921 28503 14979 28509
rect 16025 28509 16037 28543
rect 16071 28540 16083 28543
rect 16298 28540 16304 28552
rect 16071 28512 16304 28540
rect 16071 28509 16083 28512
rect 16025 28503 16083 28509
rect 16298 28500 16304 28512
rect 16356 28500 16362 28552
rect 16991 28543 17049 28549
rect 16991 28509 17003 28543
rect 17037 28540 17049 28543
rect 17037 28512 17172 28540
rect 17037 28509 17049 28512
rect 16991 28503 17049 28509
rect 17144 28484 17172 28512
rect 17218 28500 17224 28552
rect 17276 28540 17282 28552
rect 17957 28543 18015 28549
rect 17957 28540 17969 28543
rect 17276 28512 17969 28540
rect 17276 28500 17282 28512
rect 17957 28509 17969 28512
rect 18003 28509 18015 28543
rect 17957 28503 18015 28509
rect 18046 28500 18052 28552
rect 18104 28540 18110 28552
rect 18248 28549 18276 28580
rect 18322 28568 18328 28620
rect 18380 28608 18386 28620
rect 19150 28608 19156 28620
rect 18380 28580 19156 28608
rect 18380 28568 18386 28580
rect 19150 28568 19156 28580
rect 19208 28608 19214 28620
rect 19702 28608 19708 28620
rect 19208 28580 19708 28608
rect 19208 28568 19214 28580
rect 19702 28568 19708 28580
rect 19760 28568 19766 28620
rect 20272 28608 20484 28624
rect 20272 28596 21864 28608
rect 20456 28580 21864 28596
rect 18141 28543 18199 28549
rect 18141 28540 18153 28543
rect 18104 28512 18153 28540
rect 18104 28500 18110 28512
rect 18141 28509 18153 28512
rect 18187 28509 18199 28543
rect 18141 28503 18199 28509
rect 18233 28543 18291 28549
rect 18233 28509 18245 28543
rect 18279 28509 18291 28543
rect 20441 28543 20499 28549
rect 20441 28540 20453 28543
rect 18233 28503 18291 28509
rect 19168 28512 20453 28540
rect 11247 28444 11567 28472
rect 11054 28404 11060 28416
rect 9876 28376 11060 28404
rect 11054 28364 11060 28376
rect 11112 28364 11118 28416
rect 11539 28404 11567 28444
rect 11606 28432 11612 28484
rect 11664 28432 11670 28484
rect 11698 28432 11704 28484
rect 11756 28472 11762 28484
rect 15105 28475 15163 28481
rect 15105 28472 15117 28475
rect 11756 28444 15117 28472
rect 11756 28432 11762 28444
rect 15105 28441 15117 28444
rect 15151 28441 15163 28475
rect 17126 28472 17132 28484
rect 17039 28444 17132 28472
rect 15105 28435 15163 28441
rect 17126 28432 17132 28444
rect 17184 28472 17190 28484
rect 19168 28472 19196 28512
rect 20441 28509 20453 28512
rect 20487 28540 20499 28543
rect 20622 28540 20628 28552
rect 20487 28512 20628 28540
rect 20487 28509 20499 28512
rect 20441 28503 20499 28509
rect 20622 28500 20628 28512
rect 20680 28500 20686 28552
rect 20714 28500 20720 28552
rect 20772 28540 20778 28552
rect 21726 28540 21732 28552
rect 20772 28512 20817 28540
rect 21687 28512 21732 28540
rect 20772 28500 20778 28512
rect 21726 28500 21732 28512
rect 21784 28500 21790 28552
rect 21836 28540 21864 28580
rect 23106 28568 23112 28620
rect 23164 28608 23170 28620
rect 28166 28608 28172 28620
rect 23164 28580 24256 28608
rect 28127 28580 28172 28608
rect 23164 28568 23170 28580
rect 23845 28543 23903 28549
rect 23845 28540 23857 28543
rect 21836 28512 23857 28540
rect 23845 28509 23857 28512
rect 23891 28509 23903 28543
rect 23845 28503 23903 28509
rect 17184 28444 19196 28472
rect 17184 28432 17190 28444
rect 19334 28432 19340 28484
rect 19392 28472 19398 28484
rect 19613 28475 19671 28481
rect 19613 28472 19625 28475
rect 19392 28444 19625 28472
rect 19392 28432 19398 28444
rect 19613 28441 19625 28444
rect 19659 28441 19671 28475
rect 19794 28472 19800 28484
rect 19755 28444 19800 28472
rect 19613 28435 19671 28441
rect 19794 28432 19800 28444
rect 19852 28432 19858 28484
rect 20806 28432 20812 28484
rect 20864 28472 20870 28484
rect 21974 28475 22032 28481
rect 21974 28472 21986 28475
rect 20864 28444 21986 28472
rect 20864 28432 20870 28444
rect 21974 28441 21986 28444
rect 22020 28441 22032 28475
rect 22922 28472 22928 28484
rect 21974 28435 22032 28441
rect 22066 28444 22928 28472
rect 12342 28404 12348 28416
rect 11539 28376 12348 28404
rect 12342 28364 12348 28376
rect 12400 28364 12406 28416
rect 12434 28364 12440 28416
rect 12492 28404 12498 28416
rect 12621 28407 12679 28413
rect 12621 28404 12633 28407
rect 12492 28376 12633 28404
rect 12492 28364 12498 28376
rect 12621 28373 12633 28376
rect 12667 28373 12679 28407
rect 12621 28367 12679 28373
rect 13081 28407 13139 28413
rect 13081 28373 13093 28407
rect 13127 28404 13139 28407
rect 13170 28404 13176 28416
rect 13127 28376 13176 28404
rect 13127 28373 13139 28376
rect 13081 28367 13139 28373
rect 13170 28364 13176 28376
rect 13228 28364 13234 28416
rect 14185 28407 14243 28413
rect 14185 28373 14197 28407
rect 14231 28404 14243 28407
rect 16114 28404 16120 28416
rect 14231 28376 16120 28404
rect 14231 28373 14243 28376
rect 14185 28367 14243 28373
rect 16114 28364 16120 28376
rect 16172 28364 16178 28416
rect 16482 28364 16488 28416
rect 16540 28404 16546 28416
rect 18230 28404 18236 28416
rect 16540 28376 18236 28404
rect 16540 28364 16546 28376
rect 18230 28364 18236 28376
rect 18288 28364 18294 28416
rect 18417 28407 18475 28413
rect 18417 28373 18429 28407
rect 18463 28404 18475 28407
rect 19886 28404 19892 28416
rect 18463 28376 19892 28404
rect 18463 28373 18475 28376
rect 18417 28367 18475 28373
rect 19886 28364 19892 28376
rect 19944 28364 19950 28416
rect 19981 28407 20039 28413
rect 19981 28373 19993 28407
rect 20027 28404 20039 28407
rect 22066 28404 22094 28444
rect 22922 28432 22928 28444
rect 22980 28432 22986 28484
rect 23658 28472 23664 28484
rect 23619 28444 23664 28472
rect 23658 28432 23664 28444
rect 23716 28432 23722 28484
rect 23750 28432 23756 28484
rect 23808 28472 23814 28484
rect 24118 28472 24124 28484
rect 23808 28444 24124 28472
rect 23808 28432 23814 28444
rect 24118 28432 24124 28444
rect 24176 28432 24182 28484
rect 24228 28472 24256 28580
rect 28166 28568 28172 28580
rect 28224 28568 28230 28620
rect 24397 28543 24455 28549
rect 24397 28509 24409 28543
rect 24443 28540 24455 28543
rect 24486 28540 24492 28552
rect 24443 28512 24492 28540
rect 24443 28509 24455 28512
rect 24397 28503 24455 28509
rect 24486 28500 24492 28512
rect 24544 28500 24550 28552
rect 24946 28500 24952 28552
rect 25004 28540 25010 28552
rect 25682 28540 25688 28552
rect 25004 28512 25688 28540
rect 25004 28500 25010 28512
rect 25682 28500 25688 28512
rect 25740 28500 25746 28552
rect 26326 28540 26332 28552
rect 26287 28512 26332 28540
rect 26326 28500 26332 28512
rect 26384 28500 26390 28552
rect 24642 28475 24700 28481
rect 24642 28472 24654 28475
rect 24228 28444 24654 28472
rect 24642 28441 24654 28444
rect 24688 28472 24700 28475
rect 26053 28475 26111 28481
rect 26053 28472 26065 28475
rect 24688 28444 26065 28472
rect 24688 28441 24700 28444
rect 24642 28435 24700 28441
rect 26053 28441 26065 28444
rect 26099 28441 26111 28475
rect 26510 28472 26516 28484
rect 26471 28444 26516 28472
rect 26053 28435 26111 28441
rect 26510 28432 26516 28444
rect 26568 28432 26574 28484
rect 20027 28376 22094 28404
rect 20027 28373 20039 28376
rect 19981 28367 20039 28373
rect 22186 28364 22192 28416
rect 22244 28404 22250 28416
rect 25590 28404 25596 28416
rect 22244 28376 25596 28404
rect 22244 28364 22250 28376
rect 25590 28364 25596 28376
rect 25648 28364 25654 28416
rect 25682 28364 25688 28416
rect 25740 28404 25746 28416
rect 25777 28407 25835 28413
rect 25777 28404 25789 28407
rect 25740 28376 25789 28404
rect 25740 28364 25746 28376
rect 25777 28373 25789 28376
rect 25823 28373 25835 28407
rect 25777 28367 25835 28373
rect 1104 28314 28888 28336
rect 1104 28262 10214 28314
rect 10266 28262 10278 28314
rect 10330 28262 10342 28314
rect 10394 28262 10406 28314
rect 10458 28262 10470 28314
rect 10522 28262 19478 28314
rect 19530 28262 19542 28314
rect 19594 28262 19606 28314
rect 19658 28262 19670 28314
rect 19722 28262 19734 28314
rect 19786 28262 28888 28314
rect 1104 28240 28888 28262
rect 8205 28203 8263 28209
rect 8205 28169 8217 28203
rect 8251 28200 8263 28203
rect 8294 28200 8300 28212
rect 8251 28172 8300 28200
rect 8251 28169 8263 28172
rect 8205 28163 8263 28169
rect 8294 28160 8300 28172
rect 8352 28160 8358 28212
rect 12345 28203 12403 28209
rect 12345 28200 12357 28203
rect 8404 28172 12357 28200
rect 8404 28073 8432 28172
rect 12345 28169 12357 28172
rect 12391 28169 12403 28203
rect 12345 28163 12403 28169
rect 12618 28160 12624 28212
rect 12676 28160 12682 28212
rect 12802 28160 12808 28212
rect 12860 28200 12866 28212
rect 13170 28200 13176 28212
rect 12860 28172 13176 28200
rect 12860 28160 12866 28172
rect 13170 28160 13176 28172
rect 13228 28200 13234 28212
rect 13541 28203 13599 28209
rect 13541 28200 13553 28203
rect 13228 28172 13553 28200
rect 13228 28160 13234 28172
rect 13541 28169 13553 28172
rect 13587 28200 13599 28203
rect 13906 28200 13912 28212
rect 13587 28172 13912 28200
rect 13587 28169 13599 28172
rect 13541 28163 13599 28169
rect 13906 28160 13912 28172
rect 13964 28160 13970 28212
rect 13998 28160 14004 28212
rect 14056 28200 14062 28212
rect 14056 28172 14596 28200
rect 14056 28160 14062 28172
rect 9674 28092 9680 28144
rect 9732 28132 9738 28144
rect 10965 28135 11023 28141
rect 10965 28132 10977 28135
rect 9732 28104 10977 28132
rect 9732 28092 9738 28104
rect 10965 28101 10977 28104
rect 11011 28101 11023 28135
rect 10965 28095 11023 28101
rect 11238 28092 11244 28144
rect 11296 28132 11302 28144
rect 11974 28132 11980 28144
rect 11296 28104 11980 28132
rect 11296 28092 11302 28104
rect 11974 28092 11980 28104
rect 12032 28092 12038 28144
rect 12636 28132 12664 28160
rect 12084 28104 12296 28132
rect 12636 28104 14044 28132
rect 8389 28067 8447 28073
rect 8389 28033 8401 28067
rect 8435 28033 8447 28067
rect 9490 28064 9496 28076
rect 9451 28036 9496 28064
rect 8389 28027 8447 28033
rect 9490 28024 9496 28036
rect 9548 28024 9554 28076
rect 9950 28024 9956 28076
rect 10008 28064 10014 28076
rect 10137 28067 10195 28073
rect 10137 28064 10149 28067
rect 10008 28036 10149 28064
rect 10008 28024 10014 28036
rect 10137 28033 10149 28036
rect 10183 28033 10195 28067
rect 10781 28067 10839 28073
rect 10781 28064 10793 28067
rect 10137 28027 10195 28033
rect 10520 28036 10793 28064
rect 8202 27956 8208 28008
rect 8260 27996 8266 28008
rect 10520 27996 10548 28036
rect 10781 28033 10793 28036
rect 10827 28064 10839 28067
rect 11514 28064 11520 28076
rect 10827 28036 11520 28064
rect 10827 28033 10839 28036
rect 10781 28027 10839 28033
rect 11514 28024 11520 28036
rect 11572 28064 11578 28076
rect 12084 28073 12112 28104
rect 12069 28067 12127 28073
rect 11572 28036 12020 28064
rect 11572 28024 11578 28036
rect 8260 27968 10548 27996
rect 10597 27999 10655 28005
rect 8260 27956 8266 27968
rect 10597 27965 10609 27999
rect 10643 27996 10655 27999
rect 11790 27996 11796 28008
rect 10643 27968 11796 27996
rect 10643 27965 10655 27968
rect 10597 27959 10655 27965
rect 11790 27956 11796 27968
rect 11848 27956 11854 28008
rect 11992 27996 12020 28036
rect 12069 28033 12081 28067
rect 12115 28033 12127 28067
rect 12069 28027 12127 28033
rect 12161 28067 12219 28073
rect 12161 28033 12173 28067
rect 12207 28033 12219 28067
rect 12268 28064 12296 28104
rect 12802 28064 12808 28076
rect 12268 28036 12808 28064
rect 12161 28027 12219 28033
rect 12176 27996 12204 28027
rect 12802 28024 12808 28036
rect 12860 28024 12866 28076
rect 13262 28064 13268 28076
rect 13223 28036 13268 28064
rect 13262 28024 13268 28036
rect 13320 28024 13326 28076
rect 13446 28024 13452 28076
rect 13504 28064 13510 28076
rect 13633 28067 13691 28073
rect 13633 28064 13645 28067
rect 13504 28036 13645 28064
rect 13504 28024 13510 28036
rect 13633 28033 13645 28036
rect 13679 28033 13691 28067
rect 13633 28027 13691 28033
rect 13725 28067 13783 28073
rect 13725 28033 13737 28067
rect 13771 28064 13783 28067
rect 13771 28036 13952 28064
rect 13771 28033 13783 28036
rect 13725 28027 13783 28033
rect 11992 27968 12204 27996
rect 12986 27956 12992 28008
rect 13044 27996 13050 28008
rect 13357 27999 13415 28005
rect 13357 27996 13369 27999
rect 13044 27968 13369 27996
rect 13044 27956 13050 27968
rect 13357 27965 13369 27968
rect 13403 27996 13415 27999
rect 13814 27996 13820 28008
rect 13403 27968 13820 27996
rect 13403 27965 13415 27968
rect 13357 27959 13415 27965
rect 13814 27956 13820 27968
rect 13872 27956 13878 28008
rect 9309 27931 9367 27937
rect 9309 27897 9321 27931
rect 9355 27928 9367 27931
rect 11882 27928 11888 27940
rect 9355 27900 11888 27928
rect 9355 27897 9367 27900
rect 9309 27891 9367 27897
rect 11882 27888 11888 27900
rect 11940 27888 11946 27940
rect 12618 27928 12624 27940
rect 12084 27900 12624 27928
rect 9953 27863 10011 27869
rect 9953 27829 9965 27863
rect 9999 27860 10011 27863
rect 12084 27860 12112 27900
rect 12618 27888 12624 27900
rect 12676 27888 12682 27940
rect 13924 27928 13952 28036
rect 12728 27900 13952 27928
rect 14016 27928 14044 28104
rect 14274 28092 14280 28144
rect 14332 28132 14338 28144
rect 14430 28135 14488 28141
rect 14430 28132 14442 28135
rect 14332 28104 14442 28132
rect 14332 28092 14338 28104
rect 14430 28101 14442 28104
rect 14476 28101 14488 28135
rect 14430 28095 14488 28101
rect 14568 28064 14596 28172
rect 14642 28160 14648 28212
rect 14700 28200 14706 28212
rect 15470 28200 15476 28212
rect 14700 28172 15476 28200
rect 14700 28160 14706 28172
rect 15470 28160 15476 28172
rect 15528 28160 15534 28212
rect 15565 28203 15623 28209
rect 15565 28169 15577 28203
rect 15611 28200 15623 28203
rect 15838 28200 15844 28212
rect 15611 28172 15844 28200
rect 15611 28169 15623 28172
rect 15565 28163 15623 28169
rect 15838 28160 15844 28172
rect 15896 28160 15902 28212
rect 16114 28160 16120 28212
rect 16172 28200 16178 28212
rect 26510 28200 26516 28212
rect 16172 28172 26516 28200
rect 16172 28160 16178 28172
rect 26510 28160 26516 28172
rect 26568 28160 26574 28212
rect 28074 28200 28080 28212
rect 28035 28172 28080 28200
rect 28074 28160 28080 28172
rect 28132 28160 28138 28212
rect 15286 28092 15292 28144
rect 15344 28132 15350 28144
rect 17374 28135 17432 28141
rect 17374 28132 17386 28135
rect 15344 28104 17386 28132
rect 15344 28092 15350 28104
rect 17374 28101 17386 28104
rect 17420 28101 17432 28135
rect 17374 28095 17432 28101
rect 18230 28092 18236 28144
rect 18288 28132 18294 28144
rect 21358 28132 21364 28144
rect 18288 28104 21364 28132
rect 18288 28092 18294 28104
rect 21358 28092 21364 28104
rect 21416 28092 21422 28144
rect 21913 28135 21971 28141
rect 21913 28101 21925 28135
rect 21959 28132 21971 28135
rect 22370 28132 22376 28144
rect 21959 28104 22376 28132
rect 21959 28101 21971 28104
rect 21913 28095 21971 28101
rect 22370 28092 22376 28104
rect 22428 28092 22434 28144
rect 25038 28092 25044 28144
rect 25096 28132 25102 28144
rect 26973 28135 27031 28141
rect 26973 28132 26985 28135
rect 25096 28104 26985 28132
rect 25096 28092 25102 28104
rect 26973 28101 26985 28104
rect 27019 28101 27031 28135
rect 26973 28095 27031 28101
rect 27430 28092 27436 28144
rect 27488 28132 27494 28144
rect 27488 28104 27936 28132
rect 27488 28092 27494 28104
rect 17218 28064 17224 28076
rect 14568 28036 17224 28064
rect 17218 28024 17224 28036
rect 17276 28024 17282 28076
rect 17678 28024 17684 28076
rect 17736 28064 17742 28076
rect 18969 28067 19027 28073
rect 18969 28064 18981 28067
rect 17736 28036 18981 28064
rect 17736 28024 17742 28036
rect 18969 28033 18981 28036
rect 19015 28033 19027 28067
rect 18969 28027 19027 28033
rect 19058 28024 19064 28076
rect 19116 28064 19122 28076
rect 19225 28067 19283 28073
rect 19225 28064 19237 28067
rect 19116 28036 19237 28064
rect 19116 28024 19122 28036
rect 19225 28033 19237 28036
rect 19271 28033 19283 28067
rect 19225 28027 19283 28033
rect 21085 28067 21143 28073
rect 21085 28033 21097 28067
rect 21131 28064 21143 28067
rect 21174 28064 21180 28076
rect 21131 28036 21180 28064
rect 21131 28033 21143 28036
rect 21085 28027 21143 28033
rect 21174 28024 21180 28036
rect 21232 28024 21238 28076
rect 21542 28024 21548 28076
rect 21600 28064 21606 28076
rect 21829 28065 21887 28071
rect 21600 28062 21772 28064
rect 21829 28062 21841 28065
rect 21600 28036 21841 28062
rect 21600 28024 21606 28036
rect 21744 28034 21841 28036
rect 21829 28031 21841 28034
rect 21875 28031 21887 28065
rect 21829 28025 21887 28031
rect 22732 28067 22790 28073
rect 22732 28033 22744 28067
rect 22778 28064 22790 28067
rect 23842 28064 23848 28076
rect 22778 28036 23848 28064
rect 22778 28033 22790 28036
rect 22732 28027 22790 28033
rect 23842 28024 23848 28036
rect 23900 28024 23906 28076
rect 24305 28067 24363 28073
rect 24305 28033 24317 28067
rect 24351 28033 24363 28067
rect 24305 28027 24363 28033
rect 14090 27956 14096 28008
rect 14148 27996 14154 28008
rect 14185 27999 14243 28005
rect 14185 27996 14197 27999
rect 14148 27968 14197 27996
rect 14148 27956 14154 27968
rect 14185 27965 14197 27968
rect 14231 27965 14243 27999
rect 14185 27959 14243 27965
rect 17034 27956 17040 28008
rect 17092 27996 17098 28008
rect 17129 27999 17187 28005
rect 17129 27996 17141 27999
rect 17092 27968 17141 27996
rect 17092 27956 17098 27968
rect 17129 27965 17141 27968
rect 17175 27965 17187 27999
rect 17129 27959 17187 27965
rect 18230 27956 18236 28008
rect 18288 27996 18294 28008
rect 18690 27996 18696 28008
rect 18288 27968 18696 27996
rect 18288 27956 18294 27968
rect 18690 27956 18696 27968
rect 18748 27956 18754 28008
rect 20806 27956 20812 28008
rect 20864 27996 20870 28008
rect 20901 27999 20959 28005
rect 20901 27996 20913 27999
rect 20864 27968 20913 27996
rect 20864 27956 20870 27968
rect 20901 27965 20913 27968
rect 20947 27965 20959 27999
rect 20901 27959 20959 27965
rect 22465 27999 22523 28005
rect 22465 27965 22477 27999
rect 22511 27965 22523 27999
rect 22465 27959 22523 27965
rect 14016 27900 14136 27928
rect 9999 27832 12112 27860
rect 9999 27829 10011 27832
rect 9953 27823 10011 27829
rect 12158 27820 12164 27872
rect 12216 27860 12222 27872
rect 12728 27860 12756 27900
rect 12216 27832 12756 27860
rect 13081 27863 13139 27869
rect 12216 27820 12222 27832
rect 13081 27829 13093 27863
rect 13127 27860 13139 27863
rect 13998 27860 14004 27872
rect 13127 27832 14004 27860
rect 13127 27829 13139 27832
rect 13081 27823 13139 27829
rect 13998 27820 14004 27832
rect 14056 27820 14062 27872
rect 14108 27860 14136 27900
rect 15378 27888 15384 27940
rect 15436 27928 15442 27940
rect 16482 27928 16488 27940
rect 15436 27900 16488 27928
rect 15436 27888 15442 27900
rect 16482 27888 16488 27900
rect 16540 27888 16546 27940
rect 18322 27888 18328 27940
rect 18380 27928 18386 27940
rect 18509 27931 18567 27937
rect 18509 27928 18521 27931
rect 18380 27900 18521 27928
rect 18380 27888 18386 27900
rect 18509 27897 18521 27900
rect 18555 27928 18567 27931
rect 18598 27928 18604 27940
rect 18555 27900 18604 27928
rect 18555 27897 18567 27900
rect 18509 27891 18567 27897
rect 18598 27888 18604 27900
rect 18656 27888 18662 27940
rect 20254 27888 20260 27940
rect 20312 27928 20318 27940
rect 20349 27931 20407 27937
rect 20349 27928 20361 27931
rect 20312 27900 20361 27928
rect 20312 27888 20318 27900
rect 20349 27897 20361 27900
rect 20395 27897 20407 27931
rect 20349 27891 20407 27897
rect 20622 27888 20628 27940
rect 20680 27928 20686 27940
rect 21726 27928 21732 27940
rect 20680 27900 21732 27928
rect 20680 27888 20686 27900
rect 21726 27888 21732 27900
rect 21784 27928 21790 27940
rect 22480 27928 22508 27959
rect 23474 27956 23480 28008
rect 23532 27996 23538 28008
rect 24320 27996 24348 28027
rect 24486 28024 24492 28076
rect 24544 28064 24550 28076
rect 25297 28067 25355 28073
rect 25297 28064 25309 28067
rect 24544 28036 25309 28064
rect 24544 28024 24550 28036
rect 25297 28033 25309 28036
rect 25343 28033 25355 28067
rect 25297 28027 25355 28033
rect 25590 28024 25596 28076
rect 25648 28064 25654 28076
rect 27157 28067 27215 28073
rect 27157 28064 27169 28067
rect 25648 28036 27169 28064
rect 25648 28024 25654 28036
rect 27157 28033 27169 28036
rect 27203 28033 27215 28067
rect 27157 28027 27215 28033
rect 27341 28067 27399 28073
rect 27341 28033 27353 28067
rect 27387 28064 27399 28067
rect 27614 28064 27620 28076
rect 27387 28036 27620 28064
rect 27387 28033 27399 28036
rect 27341 28027 27399 28033
rect 27614 28024 27620 28036
rect 27672 28024 27678 28076
rect 27908 28073 27936 28104
rect 27893 28067 27951 28073
rect 27893 28033 27905 28067
rect 27939 28033 27951 28067
rect 27893 28027 27951 28033
rect 25038 27996 25044 28008
rect 23532 27968 24348 27996
rect 24999 27968 25044 27996
rect 23532 27956 23538 27968
rect 21784 27900 22508 27928
rect 21784 27888 21790 27900
rect 23934 27888 23940 27940
rect 23992 27888 23998 27940
rect 24118 27888 24124 27940
rect 24176 27888 24182 27940
rect 24320 27928 24348 27968
rect 25038 27956 25044 27968
rect 25096 27956 25102 28008
rect 26970 27956 26976 28008
rect 27028 27996 27034 28008
rect 27433 27999 27491 28005
rect 27433 27996 27445 27999
rect 27028 27968 27445 27996
rect 27028 27956 27034 27968
rect 27433 27965 27445 27968
rect 27479 27965 27491 27999
rect 27433 27959 27491 27965
rect 24320 27900 25084 27928
rect 20714 27860 20720 27872
rect 14108 27832 20720 27860
rect 20714 27820 20720 27832
rect 20772 27820 20778 27872
rect 21269 27863 21327 27869
rect 21269 27829 21281 27863
rect 21315 27860 21327 27863
rect 21818 27860 21824 27872
rect 21315 27832 21824 27860
rect 21315 27829 21327 27832
rect 21269 27823 21327 27829
rect 21818 27820 21824 27832
rect 21876 27820 21882 27872
rect 22370 27820 22376 27872
rect 22428 27860 22434 27872
rect 23750 27860 23756 27872
rect 22428 27832 23756 27860
rect 22428 27820 22434 27832
rect 23750 27820 23756 27832
rect 23808 27820 23814 27872
rect 23845 27863 23903 27869
rect 23845 27829 23857 27863
rect 23891 27860 23903 27863
rect 23952 27860 23980 27888
rect 23891 27832 23980 27860
rect 24136 27860 24164 27888
rect 24489 27863 24547 27869
rect 24489 27860 24501 27863
rect 24136 27832 24501 27860
rect 23891 27829 23903 27832
rect 23845 27823 23903 27829
rect 24489 27829 24501 27832
rect 24535 27829 24547 27863
rect 25056 27860 25084 27900
rect 26050 27860 26056 27872
rect 25056 27832 26056 27860
rect 24489 27823 24547 27829
rect 26050 27820 26056 27832
rect 26108 27820 26114 27872
rect 26421 27863 26479 27869
rect 26421 27829 26433 27863
rect 26467 27860 26479 27863
rect 27062 27860 27068 27872
rect 26467 27832 27068 27860
rect 26467 27829 26479 27832
rect 26421 27823 26479 27829
rect 27062 27820 27068 27832
rect 27120 27820 27126 27872
rect 1104 27770 28888 27792
rect 1104 27718 5582 27770
rect 5634 27718 5646 27770
rect 5698 27718 5710 27770
rect 5762 27718 5774 27770
rect 5826 27718 5838 27770
rect 5890 27718 14846 27770
rect 14898 27718 14910 27770
rect 14962 27718 14974 27770
rect 15026 27718 15038 27770
rect 15090 27718 15102 27770
rect 15154 27718 24110 27770
rect 24162 27718 24174 27770
rect 24226 27718 24238 27770
rect 24290 27718 24302 27770
rect 24354 27718 24366 27770
rect 24418 27718 28888 27770
rect 1104 27696 28888 27718
rect 9490 27616 9496 27668
rect 9548 27656 9554 27668
rect 10870 27656 10876 27668
rect 9548 27628 10876 27656
rect 9548 27616 9554 27628
rect 10870 27616 10876 27628
rect 10928 27616 10934 27668
rect 11256 27628 12204 27656
rect 8205 27591 8263 27597
rect 8205 27557 8217 27591
rect 8251 27557 8263 27591
rect 8205 27551 8263 27557
rect 9309 27591 9367 27597
rect 9309 27557 9321 27591
rect 9355 27588 9367 27591
rect 11256 27588 11284 27628
rect 9355 27560 11284 27588
rect 12176 27588 12204 27628
rect 12710 27616 12716 27668
rect 12768 27656 12774 27668
rect 13081 27659 13139 27665
rect 13081 27656 13093 27659
rect 12768 27628 13093 27656
rect 12768 27616 12774 27628
rect 13081 27625 13093 27628
rect 13127 27625 13139 27659
rect 13081 27619 13139 27625
rect 13446 27616 13452 27668
rect 13504 27656 13510 27668
rect 13541 27659 13599 27665
rect 13541 27656 13553 27659
rect 13504 27628 13553 27656
rect 13504 27616 13510 27628
rect 13541 27625 13553 27628
rect 13587 27625 13599 27659
rect 15930 27656 15936 27668
rect 13541 27619 13599 27625
rect 14108 27628 15936 27656
rect 14108 27588 14136 27628
rect 15930 27616 15936 27628
rect 15988 27616 15994 27668
rect 17034 27656 17040 27668
rect 16316 27628 17040 27656
rect 12176 27560 12664 27588
rect 9355 27557 9367 27560
rect 9309 27551 9367 27557
rect 8220 27520 8248 27551
rect 12636 27520 12664 27560
rect 13096 27560 14136 27588
rect 13096 27520 13124 27560
rect 15102 27548 15108 27600
rect 15160 27588 15166 27600
rect 16206 27588 16212 27600
rect 15160 27560 16212 27588
rect 15160 27548 15166 27560
rect 16206 27548 16212 27560
rect 16264 27548 16270 27600
rect 8220 27492 11376 27520
rect 12636 27492 13124 27520
rect 13173 27523 13231 27529
rect 8389 27455 8447 27461
rect 8389 27421 8401 27455
rect 8435 27421 8447 27455
rect 9490 27452 9496 27464
rect 9451 27424 9496 27452
rect 8389 27415 8447 27421
rect 8404 27384 8432 27415
rect 9490 27412 9496 27424
rect 9548 27412 9554 27464
rect 10134 27412 10140 27464
rect 10192 27452 10198 27464
rect 10597 27455 10655 27461
rect 10192 27424 10237 27452
rect 10192 27412 10198 27424
rect 10597 27421 10609 27455
rect 10643 27452 10655 27455
rect 10686 27452 10692 27464
rect 10643 27424 10692 27452
rect 10643 27421 10655 27424
rect 10597 27415 10655 27421
rect 10686 27412 10692 27424
rect 10744 27412 10750 27464
rect 10778 27412 10784 27464
rect 10836 27452 10842 27464
rect 11238 27452 11244 27464
rect 10836 27424 10881 27452
rect 11199 27424 11244 27452
rect 10836 27412 10842 27424
rect 11238 27412 11244 27424
rect 11296 27412 11302 27464
rect 11348 27452 11376 27492
rect 13173 27489 13185 27523
rect 13219 27489 13231 27523
rect 13173 27483 13231 27489
rect 11348 27424 11468 27452
rect 9674 27384 9680 27396
rect 8404 27356 9680 27384
rect 9674 27344 9680 27356
rect 9732 27344 9738 27396
rect 11054 27384 11060 27396
rect 9968 27356 11060 27384
rect 6822 27276 6828 27328
rect 6880 27316 6886 27328
rect 9582 27316 9588 27328
rect 6880 27288 9588 27316
rect 6880 27276 6886 27288
rect 9582 27276 9588 27288
rect 9640 27276 9646 27328
rect 9968 27325 9996 27356
rect 11054 27344 11060 27356
rect 11112 27344 11118 27396
rect 11440 27384 11468 27424
rect 11974 27412 11980 27464
rect 12032 27452 12038 27464
rect 12434 27452 12440 27464
rect 12032 27424 12440 27452
rect 12032 27412 12038 27424
rect 12434 27412 12440 27424
rect 12492 27452 12498 27464
rect 13188 27452 13216 27483
rect 15746 27480 15752 27532
rect 15804 27520 15810 27532
rect 16316 27529 16344 27628
rect 17034 27616 17040 27628
rect 17092 27616 17098 27668
rect 17402 27616 17408 27668
rect 17460 27656 17466 27668
rect 21726 27656 21732 27668
rect 17460 27628 21732 27656
rect 17460 27616 17466 27628
rect 21726 27616 21732 27628
rect 21784 27616 21790 27668
rect 22002 27616 22008 27668
rect 22060 27656 22066 27668
rect 23198 27656 23204 27668
rect 22060 27628 23204 27656
rect 22060 27616 22066 27628
rect 23198 27616 23204 27628
rect 23256 27616 23262 27668
rect 23290 27616 23296 27668
rect 23348 27656 23354 27668
rect 23348 27628 23393 27656
rect 23348 27616 23354 27628
rect 23750 27616 23756 27668
rect 23808 27656 23814 27668
rect 23808 27628 26556 27656
rect 23808 27616 23814 27628
rect 17681 27591 17739 27597
rect 17681 27557 17693 27591
rect 17727 27588 17739 27591
rect 17862 27588 17868 27600
rect 17727 27560 17868 27588
rect 17727 27557 17739 27560
rect 17681 27551 17739 27557
rect 17862 27548 17868 27560
rect 17920 27588 17926 27600
rect 18046 27588 18052 27600
rect 17920 27560 18052 27588
rect 17920 27548 17926 27560
rect 18046 27548 18052 27560
rect 18104 27548 18110 27600
rect 18156 27560 18635 27588
rect 16301 27523 16359 27529
rect 16301 27520 16313 27523
rect 15804 27492 16313 27520
rect 15804 27480 15810 27492
rect 16301 27489 16313 27492
rect 16347 27489 16359 27523
rect 18156 27520 18184 27560
rect 16301 27483 16359 27489
rect 17926 27492 18184 27520
rect 12492 27424 13216 27452
rect 13357 27455 13415 27461
rect 12492 27412 12498 27424
rect 13357 27421 13369 27455
rect 13403 27452 13415 27455
rect 13814 27452 13820 27464
rect 13403 27424 13820 27452
rect 13403 27421 13415 27424
rect 13357 27415 13415 27421
rect 13814 27412 13820 27424
rect 13872 27412 13878 27464
rect 14090 27452 14096 27464
rect 14003 27424 14096 27452
rect 14090 27412 14096 27424
rect 14148 27452 14154 27464
rect 15764 27452 15792 27480
rect 17926 27452 17954 27492
rect 18230 27480 18236 27532
rect 18288 27520 18294 27532
rect 18325 27523 18383 27529
rect 18325 27520 18337 27523
rect 18288 27492 18337 27520
rect 18288 27480 18294 27492
rect 18325 27489 18337 27492
rect 18371 27489 18383 27523
rect 18325 27483 18383 27489
rect 18414 27480 18420 27532
rect 18472 27520 18478 27532
rect 18607 27520 18635 27560
rect 18874 27548 18880 27600
rect 18932 27588 18938 27600
rect 23106 27588 23112 27600
rect 18932 27560 23112 27588
rect 18932 27548 18938 27560
rect 23106 27548 23112 27560
rect 23164 27548 23170 27600
rect 25498 27548 25504 27600
rect 25556 27588 25562 27600
rect 25869 27591 25927 27597
rect 25869 27588 25881 27591
rect 25556 27560 25881 27588
rect 25556 27548 25562 27560
rect 25869 27557 25881 27560
rect 25915 27588 25927 27591
rect 25958 27588 25964 27600
rect 25915 27560 25964 27588
rect 25915 27557 25927 27560
rect 25869 27551 25927 27557
rect 25958 27548 25964 27560
rect 26016 27548 26022 27600
rect 21910 27520 21916 27532
rect 18472 27492 18517 27520
rect 18607 27492 21916 27520
rect 18472 27480 18478 27492
rect 21910 27480 21916 27492
rect 21968 27480 21974 27532
rect 24118 27520 24124 27532
rect 22112 27492 24124 27520
rect 14148 27424 15792 27452
rect 15825 27424 17954 27452
rect 14148 27412 14154 27424
rect 11497 27387 11555 27393
rect 11497 27384 11509 27387
rect 11440 27356 11509 27384
rect 11497 27353 11509 27356
rect 11543 27353 11555 27387
rect 11497 27347 11555 27353
rect 11606 27344 11612 27396
rect 11664 27384 11670 27396
rect 11664 27356 12856 27384
rect 11664 27344 11670 27356
rect 9953 27319 10011 27325
rect 9953 27285 9965 27319
rect 9999 27285 10011 27319
rect 9953 27279 10011 27285
rect 10689 27319 10747 27325
rect 10689 27285 10701 27319
rect 10735 27316 10747 27319
rect 12434 27316 12440 27328
rect 10735 27288 12440 27316
rect 10735 27285 10747 27288
rect 10689 27279 10747 27285
rect 12434 27276 12440 27288
rect 12492 27276 12498 27328
rect 12621 27319 12679 27325
rect 12621 27285 12633 27319
rect 12667 27316 12679 27319
rect 12710 27316 12716 27328
rect 12667 27288 12716 27316
rect 12667 27285 12679 27288
rect 12621 27279 12679 27285
rect 12710 27276 12716 27288
rect 12768 27276 12774 27328
rect 12828 27316 12856 27356
rect 12894 27344 12900 27396
rect 12952 27384 12958 27396
rect 13081 27387 13139 27393
rect 13081 27384 13093 27387
rect 12952 27356 13093 27384
rect 12952 27344 12958 27356
rect 13081 27353 13093 27356
rect 13127 27353 13139 27387
rect 13081 27347 13139 27353
rect 13998 27344 14004 27396
rect 14056 27384 14062 27396
rect 14338 27387 14396 27393
rect 14338 27384 14350 27387
rect 14056 27356 14350 27384
rect 14056 27344 14062 27356
rect 14338 27353 14350 27356
rect 14384 27353 14396 27387
rect 15825 27384 15853 27424
rect 18046 27412 18052 27464
rect 18104 27452 18110 27464
rect 18509 27455 18567 27461
rect 18509 27452 18521 27455
rect 18104 27424 18521 27452
rect 18104 27412 18110 27424
rect 18509 27421 18521 27424
rect 18555 27421 18567 27455
rect 18509 27415 18567 27421
rect 18598 27412 18604 27464
rect 18656 27452 18662 27464
rect 22112 27452 22140 27492
rect 24118 27480 24124 27492
rect 24176 27480 24182 27532
rect 26528 27529 26556 27628
rect 26513 27523 26571 27529
rect 26513 27489 26525 27523
rect 26559 27489 26571 27523
rect 26513 27483 26571 27489
rect 22278 27452 22284 27464
rect 18656 27424 18701 27452
rect 18769 27424 22140 27452
rect 22239 27424 22284 27452
rect 18656 27412 18662 27424
rect 14338 27347 14396 27353
rect 14660 27356 15853 27384
rect 14660 27316 14688 27356
rect 15930 27344 15936 27396
rect 15988 27384 15994 27396
rect 16546 27387 16604 27393
rect 16546 27384 16558 27387
rect 15988 27356 16558 27384
rect 15988 27344 15994 27356
rect 16546 27353 16558 27356
rect 16592 27353 16604 27387
rect 16546 27347 16604 27353
rect 16850 27344 16856 27396
rect 16908 27384 16914 27396
rect 18769 27384 18797 27424
rect 22278 27412 22284 27424
rect 22336 27412 22342 27464
rect 22370 27412 22376 27464
rect 22428 27452 22434 27464
rect 22557 27455 22615 27461
rect 22557 27452 22569 27455
rect 22428 27424 22569 27452
rect 22428 27412 22434 27424
rect 22557 27421 22569 27424
rect 22603 27421 22615 27455
rect 22557 27415 22615 27421
rect 23566 27412 23572 27464
rect 23624 27452 23630 27464
rect 24489 27455 24547 27461
rect 24489 27452 24501 27455
rect 23624 27424 24501 27452
rect 23624 27412 23630 27424
rect 24489 27421 24501 27424
rect 24535 27452 24547 27455
rect 25038 27452 25044 27464
rect 24535 27424 25044 27452
rect 24535 27421 24547 27424
rect 24489 27415 24547 27421
rect 25038 27412 25044 27424
rect 25096 27412 25102 27464
rect 26326 27452 26332 27464
rect 26287 27424 26332 27452
rect 26326 27412 26332 27424
rect 26384 27412 26390 27464
rect 16908 27356 18797 27384
rect 16908 27344 16914 27356
rect 19058 27344 19064 27396
rect 19116 27384 19122 27396
rect 19242 27384 19248 27396
rect 19116 27356 19248 27384
rect 19116 27344 19122 27356
rect 19242 27344 19248 27356
rect 19300 27384 19306 27396
rect 19334 27384 19340 27396
rect 19300 27356 19340 27384
rect 19300 27344 19306 27356
rect 19334 27344 19340 27356
rect 19392 27344 19398 27396
rect 19613 27387 19671 27393
rect 19613 27353 19625 27387
rect 19659 27384 19671 27387
rect 20714 27384 20720 27396
rect 19659 27356 20720 27384
rect 19659 27353 19671 27356
rect 19613 27347 19671 27353
rect 20714 27344 20720 27356
rect 20772 27344 20778 27396
rect 20806 27344 20812 27396
rect 20864 27384 20870 27396
rect 21082 27384 21088 27396
rect 20864 27356 21088 27384
rect 20864 27344 20870 27356
rect 21082 27344 21088 27356
rect 21140 27344 21146 27396
rect 22097 27387 22155 27393
rect 22097 27353 22109 27387
rect 22143 27384 22155 27387
rect 22646 27384 22652 27396
rect 22143 27356 22652 27384
rect 22143 27353 22155 27356
rect 22097 27347 22155 27353
rect 22646 27344 22652 27356
rect 22704 27344 22710 27396
rect 23109 27387 23167 27393
rect 23109 27353 23121 27387
rect 23155 27384 23167 27387
rect 23934 27384 23940 27396
rect 23155 27356 23940 27384
rect 23155 27353 23167 27356
rect 23109 27347 23167 27353
rect 23934 27344 23940 27356
rect 23992 27344 23998 27396
rect 24756 27387 24814 27393
rect 24756 27353 24768 27387
rect 24802 27384 24814 27387
rect 25406 27384 25412 27396
rect 24802 27356 25412 27384
rect 24802 27353 24814 27356
rect 24756 27347 24814 27353
rect 25406 27344 25412 27356
rect 25464 27344 25470 27396
rect 28166 27384 28172 27396
rect 28127 27356 28172 27384
rect 28166 27344 28172 27356
rect 28224 27344 28230 27396
rect 12828 27288 14688 27316
rect 14734 27276 14740 27328
rect 14792 27316 14798 27328
rect 15194 27316 15200 27328
rect 14792 27288 15200 27316
rect 14792 27276 14798 27288
rect 15194 27276 15200 27288
rect 15252 27316 15258 27328
rect 15473 27319 15531 27325
rect 15473 27316 15485 27319
rect 15252 27288 15485 27316
rect 15252 27276 15258 27288
rect 15473 27285 15485 27288
rect 15519 27285 15531 27319
rect 15473 27279 15531 27285
rect 17954 27276 17960 27328
rect 18012 27316 18018 27328
rect 18141 27319 18199 27325
rect 18141 27316 18153 27319
rect 18012 27288 18153 27316
rect 18012 27276 18018 27288
rect 18141 27285 18153 27288
rect 18187 27285 18199 27319
rect 18141 27279 18199 27285
rect 18230 27276 18236 27328
rect 18288 27316 18294 27328
rect 20901 27319 20959 27325
rect 20901 27316 20913 27319
rect 18288 27288 20913 27316
rect 18288 27276 18294 27288
rect 20901 27285 20913 27288
rect 20947 27285 20959 27319
rect 20901 27279 20959 27285
rect 22186 27276 22192 27328
rect 22244 27316 22250 27328
rect 22465 27319 22523 27325
rect 22465 27316 22477 27319
rect 22244 27288 22477 27316
rect 22244 27276 22250 27288
rect 22465 27285 22477 27288
rect 22511 27285 22523 27319
rect 22465 27279 22523 27285
rect 22554 27276 22560 27328
rect 22612 27316 22618 27328
rect 23309 27319 23367 27325
rect 23309 27316 23321 27319
rect 22612 27288 23321 27316
rect 22612 27276 22618 27288
rect 23309 27285 23321 27288
rect 23355 27285 23367 27319
rect 23309 27279 23367 27285
rect 23477 27319 23535 27325
rect 23477 27285 23489 27319
rect 23523 27316 23535 27319
rect 24670 27316 24676 27328
rect 23523 27288 24676 27316
rect 23523 27285 23535 27288
rect 23477 27279 23535 27285
rect 24670 27276 24676 27288
rect 24728 27316 24734 27328
rect 24854 27316 24860 27328
rect 24728 27288 24860 27316
rect 24728 27276 24734 27288
rect 24854 27276 24860 27288
rect 24912 27276 24918 27328
rect 1104 27226 28888 27248
rect 1104 27174 10214 27226
rect 10266 27174 10278 27226
rect 10330 27174 10342 27226
rect 10394 27174 10406 27226
rect 10458 27174 10470 27226
rect 10522 27174 19478 27226
rect 19530 27174 19542 27226
rect 19594 27174 19606 27226
rect 19658 27174 19670 27226
rect 19722 27174 19734 27226
rect 19786 27174 28888 27226
rect 1104 27152 28888 27174
rect 9214 27072 9220 27124
rect 9272 27112 9278 27124
rect 11422 27112 11428 27124
rect 9272 27084 11428 27112
rect 9272 27072 9278 27084
rect 11422 27072 11428 27084
rect 11480 27072 11486 27124
rect 12250 27072 12256 27124
rect 12308 27112 12314 27124
rect 13446 27112 13452 27124
rect 12308 27084 13452 27112
rect 12308 27072 12314 27084
rect 13446 27072 13452 27084
rect 13504 27112 13510 27124
rect 18230 27112 18236 27124
rect 13504 27084 18236 27112
rect 13504 27072 13510 27084
rect 18230 27072 18236 27084
rect 18288 27072 18294 27124
rect 18506 27112 18512 27124
rect 18340 27084 18512 27112
rect 10134 27004 10140 27056
rect 10192 27044 10198 27056
rect 11606 27044 11612 27056
rect 10192 27016 11612 27044
rect 10192 27004 10198 27016
rect 11606 27004 11612 27016
rect 11664 27004 11670 27056
rect 11793 27047 11851 27053
rect 11793 27013 11805 27047
rect 11839 27013 11851 27047
rect 11793 27007 11851 27013
rect 12009 27047 12067 27053
rect 12009 27013 12021 27047
rect 12055 27044 12067 27047
rect 12055 27016 12664 27044
rect 12055 27013 12067 27016
rect 12009 27007 12067 27013
rect 10321 26979 10379 26985
rect 10321 26945 10333 26979
rect 10367 26976 10379 26979
rect 10778 26976 10784 26988
rect 10367 26948 10640 26976
rect 10739 26948 10784 26976
rect 10367 26945 10379 26948
rect 10321 26939 10379 26945
rect 9766 26868 9772 26920
rect 9824 26908 9830 26920
rect 9950 26908 9956 26920
rect 9824 26880 9956 26908
rect 9824 26868 9830 26880
rect 9950 26868 9956 26880
rect 10008 26868 10014 26920
rect 9674 26840 9680 26852
rect 9635 26812 9680 26840
rect 9674 26800 9680 26812
rect 9732 26800 9738 26852
rect 10612 26840 10640 26948
rect 10778 26936 10784 26948
rect 10836 26936 10842 26988
rect 10965 26979 11023 26985
rect 10965 26945 10977 26979
rect 11011 26976 11023 26979
rect 11698 26976 11704 26988
rect 11011 26948 11704 26976
rect 11011 26945 11023 26948
rect 10965 26939 11023 26945
rect 11698 26936 11704 26948
rect 11756 26936 11762 26988
rect 11808 26976 11836 27007
rect 12526 26976 12532 26988
rect 11808 26948 12532 26976
rect 12526 26936 12532 26948
rect 12584 26936 12590 26988
rect 10873 26911 10931 26917
rect 10873 26877 10885 26911
rect 10919 26908 10931 26911
rect 11790 26908 11796 26920
rect 10919 26880 11796 26908
rect 10919 26877 10931 26880
rect 10873 26871 10931 26877
rect 11790 26868 11796 26880
rect 11848 26868 11854 26920
rect 12342 26908 12348 26920
rect 11900 26880 12348 26908
rect 11900 26840 11928 26880
rect 12342 26868 12348 26880
rect 12400 26868 12406 26920
rect 12636 26908 12664 27016
rect 14182 27004 14188 27056
rect 14240 27044 14246 27056
rect 16850 27044 16856 27056
rect 14240 27016 16856 27044
rect 14240 27004 14246 27016
rect 16850 27004 16856 27016
rect 16908 27004 16914 27056
rect 17954 27004 17960 27056
rect 18012 27044 18018 27056
rect 18012 27016 18057 27044
rect 18012 27004 18018 27016
rect 18138 27004 18144 27056
rect 18196 27004 18202 27056
rect 12710 26936 12716 26988
rect 12768 26976 12774 26988
rect 12805 26979 12863 26985
rect 12805 26976 12817 26979
rect 12768 26948 12817 26976
rect 12768 26936 12774 26948
rect 12805 26945 12817 26948
rect 12851 26945 12863 26979
rect 12805 26939 12863 26945
rect 12897 26979 12955 26985
rect 12897 26945 12909 26979
rect 12943 26945 12955 26979
rect 12897 26939 12955 26945
rect 12912 26908 12940 26939
rect 12986 26936 12992 26988
rect 13044 26976 13050 26988
rect 13633 26979 13691 26985
rect 13633 26976 13645 26979
rect 13044 26948 13645 26976
rect 13044 26946 13124 26948
rect 13044 26936 13050 26946
rect 13633 26945 13645 26948
rect 13679 26945 13691 26979
rect 13633 26939 13691 26945
rect 13814 26936 13820 26988
rect 13872 26976 13878 26988
rect 13909 26979 13967 26985
rect 13909 26976 13921 26979
rect 13872 26948 13921 26976
rect 13872 26936 13878 26948
rect 13909 26945 13921 26948
rect 13955 26945 13967 26979
rect 13909 26939 13967 26945
rect 14090 26936 14096 26988
rect 14148 26976 14154 26988
rect 14642 26976 14648 26988
rect 14148 26948 14648 26976
rect 14148 26936 14154 26948
rect 14642 26936 14648 26948
rect 14700 26936 14706 26988
rect 14734 26936 14740 26988
rect 14792 26976 14798 26988
rect 14829 26979 14887 26985
rect 14829 26976 14841 26979
rect 14792 26948 14841 26976
rect 14792 26936 14798 26948
rect 14829 26945 14841 26948
rect 14875 26945 14887 26979
rect 14829 26939 14887 26945
rect 15010 26936 15016 26988
rect 15068 26976 15074 26988
rect 15654 26976 15660 26988
rect 15068 26948 15660 26976
rect 15068 26936 15074 26948
rect 15654 26936 15660 26948
rect 15712 26936 15718 26988
rect 15838 26936 15844 26988
rect 15896 26976 15902 26988
rect 15933 26979 15991 26985
rect 15933 26976 15945 26979
rect 15896 26948 15945 26976
rect 15896 26936 15902 26948
rect 15933 26945 15945 26948
rect 15979 26945 15991 26979
rect 16942 26976 16948 26988
rect 16903 26948 16948 26976
rect 15933 26939 15991 26945
rect 16942 26936 16948 26948
rect 17000 26936 17006 26988
rect 17037 26979 17095 26985
rect 17037 26945 17049 26979
rect 17083 26976 17095 26979
rect 17678 26976 17684 26988
rect 17083 26948 17684 26976
rect 17083 26945 17095 26948
rect 17037 26939 17095 26945
rect 13538 26908 13544 26920
rect 12636 26880 12756 26908
rect 12912 26880 13544 26908
rect 12158 26840 12164 26852
rect 10612 26812 11928 26840
rect 12119 26812 12164 26840
rect 12158 26800 12164 26812
rect 12216 26800 12222 26852
rect 12618 26840 12624 26852
rect 12579 26812 12624 26840
rect 12618 26800 12624 26812
rect 12676 26800 12682 26852
rect 12728 26840 12756 26880
rect 13538 26868 13544 26880
rect 13596 26908 13602 26920
rect 13725 26911 13783 26917
rect 13725 26908 13737 26911
rect 13596 26880 13737 26908
rect 13596 26868 13602 26880
rect 13725 26877 13737 26880
rect 13771 26877 13783 26911
rect 13725 26871 13783 26877
rect 13812 26880 15240 26908
rect 13173 26843 13231 26849
rect 13173 26840 13185 26843
rect 12728 26812 13185 26840
rect 13173 26809 13185 26812
rect 13219 26809 13231 26843
rect 13173 26803 13231 26809
rect 13262 26800 13268 26852
rect 13320 26840 13326 26852
rect 13812 26840 13840 26880
rect 13320 26812 13840 26840
rect 13320 26800 13326 26812
rect 13998 26800 14004 26852
rect 14056 26840 14062 26852
rect 15010 26840 15016 26852
rect 14056 26812 15016 26840
rect 14056 26800 14062 26812
rect 15010 26800 15016 26812
rect 15068 26800 15074 26852
rect 15105 26843 15163 26849
rect 15105 26809 15117 26843
rect 15151 26809 15163 26843
rect 15212 26840 15240 26880
rect 15562 26868 15568 26920
rect 15620 26908 15626 26920
rect 15749 26911 15807 26917
rect 15749 26908 15761 26911
rect 15620 26880 15761 26908
rect 15620 26868 15626 26880
rect 15749 26877 15761 26880
rect 15795 26877 15807 26911
rect 15749 26871 15807 26877
rect 16758 26868 16764 26920
rect 16816 26908 16822 26920
rect 17052 26908 17080 26939
rect 17678 26936 17684 26948
rect 17736 26936 17742 26988
rect 17770 26936 17776 26988
rect 17828 26966 17834 26988
rect 17865 26979 17923 26985
rect 17865 26966 17877 26979
rect 17828 26945 17877 26966
rect 17911 26945 17923 26979
rect 17828 26939 17923 26945
rect 18049 26979 18107 26985
rect 18049 26945 18061 26979
rect 18095 26976 18107 26979
rect 18156 26976 18184 27004
rect 18095 26948 18184 26976
rect 18233 26979 18291 26985
rect 18095 26945 18107 26948
rect 18049 26939 18107 26945
rect 18233 26945 18245 26979
rect 18279 26976 18291 26979
rect 18340 26976 18368 27084
rect 18506 27072 18512 27084
rect 18564 27072 18570 27124
rect 18785 27115 18843 27121
rect 18785 27081 18797 27115
rect 18831 27112 18843 27115
rect 19978 27112 19984 27124
rect 18831 27084 19984 27112
rect 18831 27081 18843 27084
rect 18785 27075 18843 27081
rect 19978 27072 19984 27084
rect 20036 27072 20042 27124
rect 22370 27112 22376 27124
rect 22112 27084 22376 27112
rect 18414 27004 18420 27056
rect 18472 27044 18478 27056
rect 19582 27047 19640 27053
rect 19582 27044 19594 27047
rect 18472 27016 19594 27044
rect 18472 27004 18478 27016
rect 19582 27013 19594 27016
rect 19628 27013 19640 27047
rect 19582 27007 19640 27013
rect 22112 26988 22140 27084
rect 22370 27072 22376 27084
rect 22428 27072 22434 27124
rect 24578 27072 24584 27124
rect 24636 27112 24642 27124
rect 25409 27115 25467 27121
rect 25409 27112 25421 27115
rect 24636 27084 25421 27112
rect 24636 27072 24642 27084
rect 25409 27081 25421 27084
rect 25455 27081 25467 27115
rect 25409 27075 25467 27081
rect 27338 27072 27344 27124
rect 27396 27112 27402 27124
rect 27890 27112 27896 27124
rect 27396 27084 27896 27112
rect 27396 27072 27402 27084
rect 27890 27072 27896 27084
rect 27948 27072 27954 27124
rect 22186 27004 22192 27056
rect 22244 27044 22250 27056
rect 27798 27044 27804 27056
rect 22244 27016 22416 27044
rect 27759 27016 27804 27044
rect 22244 27004 22250 27016
rect 22388 26988 22416 27016
rect 27798 27004 27804 27016
rect 27856 27004 27862 27056
rect 18693 26979 18751 26985
rect 18693 26976 18705 26979
rect 18279 26948 18368 26976
rect 18432 26948 18705 26976
rect 18279 26945 18291 26948
rect 18233 26939 18291 26945
rect 17828 26938 17908 26939
rect 17828 26936 17834 26938
rect 16816 26880 17080 26908
rect 16816 26868 16822 26880
rect 17402 26868 17408 26920
rect 17460 26908 17466 26920
rect 18432 26908 18460 26948
rect 18693 26945 18705 26948
rect 18739 26945 18751 26979
rect 18693 26939 18751 26945
rect 18874 26936 18880 26988
rect 18932 26976 18938 26988
rect 21726 26976 21732 26988
rect 18932 26948 21732 26976
rect 18932 26936 18938 26948
rect 21726 26936 21732 26948
rect 21784 26936 21790 26988
rect 21818 26936 21824 26988
rect 21876 26976 21882 26988
rect 22005 26979 22063 26985
rect 22005 26976 22017 26979
rect 21876 26948 22017 26976
rect 21876 26936 21882 26948
rect 22005 26945 22017 26948
rect 22051 26945 22063 26979
rect 22005 26939 22063 26945
rect 22094 26936 22100 26988
rect 22152 26976 22158 26988
rect 22370 26976 22376 26988
rect 22152 26948 22197 26976
rect 22331 26948 22376 26976
rect 22152 26936 22158 26948
rect 22370 26936 22376 26948
rect 22428 26936 22434 26988
rect 22554 26936 22560 26988
rect 22612 26976 22618 26988
rect 23842 26985 23848 26988
rect 22925 26979 22983 26985
rect 22925 26976 22937 26979
rect 22612 26948 22937 26976
rect 22612 26936 22618 26948
rect 22925 26945 22937 26948
rect 22971 26945 22983 26979
rect 22925 26939 22983 26945
rect 23836 26939 23848 26985
rect 23900 26976 23906 26988
rect 23900 26948 23936 26976
rect 23842 26936 23848 26939
rect 23900 26936 23906 26948
rect 24118 26936 24124 26988
rect 24176 26976 24182 26988
rect 25593 26979 25651 26985
rect 25593 26976 25605 26979
rect 24176 26948 25605 26976
rect 24176 26936 24182 26948
rect 25593 26945 25605 26948
rect 25639 26945 25651 26979
rect 25866 26976 25872 26988
rect 25827 26948 25872 26976
rect 25593 26939 25651 26945
rect 25866 26936 25872 26948
rect 25924 26936 25930 26988
rect 27430 26976 27436 26988
rect 27391 26948 27436 26976
rect 27430 26936 27436 26948
rect 27488 26936 27494 26988
rect 17460 26880 18460 26908
rect 17460 26868 17466 26880
rect 17221 26843 17279 26849
rect 17221 26840 17233 26843
rect 15212 26812 17233 26840
rect 15105 26803 15163 26809
rect 17221 26809 17233 26812
rect 17267 26809 17279 26843
rect 17221 26803 17279 26809
rect 9030 26772 9036 26784
rect 8991 26744 9036 26772
rect 9030 26732 9036 26744
rect 9088 26732 9094 26784
rect 10137 26775 10195 26781
rect 10137 26741 10149 26775
rect 10183 26772 10195 26775
rect 10226 26772 10232 26784
rect 10183 26744 10232 26772
rect 10183 26741 10195 26744
rect 10137 26735 10195 26741
rect 10226 26732 10232 26744
rect 10284 26732 10290 26784
rect 11974 26772 11980 26784
rect 11935 26744 11980 26772
rect 11974 26732 11980 26744
rect 12032 26732 12038 26784
rect 12250 26732 12256 26784
rect 12308 26772 12314 26784
rect 12710 26772 12716 26784
rect 12308 26744 12716 26772
rect 12308 26732 12314 26744
rect 12710 26732 12716 26744
rect 12768 26772 12774 26784
rect 13633 26775 13691 26781
rect 13633 26772 13645 26775
rect 12768 26744 13645 26772
rect 12768 26732 12774 26744
rect 13633 26741 13645 26744
rect 13679 26741 13691 26775
rect 13633 26735 13691 26741
rect 13722 26732 13728 26784
rect 13780 26772 13786 26784
rect 14093 26775 14151 26781
rect 14093 26772 14105 26775
rect 13780 26744 14105 26772
rect 13780 26732 13786 26744
rect 14093 26741 14105 26744
rect 14139 26741 14151 26775
rect 14093 26735 14151 26741
rect 14550 26732 14556 26784
rect 14608 26772 14614 26784
rect 15120 26772 15148 26803
rect 17494 26800 17500 26852
rect 17552 26840 17558 26852
rect 17681 26843 17739 26849
rect 17681 26840 17693 26843
rect 17552 26812 17693 26840
rect 17552 26800 17558 26812
rect 17681 26809 17693 26812
rect 17727 26809 17739 26843
rect 18432 26840 18460 26880
rect 18506 26868 18512 26920
rect 18564 26908 18570 26920
rect 19337 26911 19395 26917
rect 19337 26908 19349 26911
rect 18564 26880 19349 26908
rect 18564 26868 18570 26880
rect 19337 26877 19349 26880
rect 19383 26877 19395 26911
rect 19337 26871 19395 26877
rect 20622 26868 20628 26920
rect 20680 26908 20686 26920
rect 23566 26908 23572 26920
rect 20680 26880 23572 26908
rect 20680 26868 20686 26880
rect 23566 26868 23572 26880
rect 23624 26868 23630 26920
rect 24578 26868 24584 26920
rect 24636 26908 24642 26920
rect 25884 26908 25912 26936
rect 24636 26880 25912 26908
rect 24636 26868 24642 26880
rect 19242 26840 19248 26852
rect 18432 26812 19248 26840
rect 17681 26803 17739 26809
rect 14608 26744 15148 26772
rect 15289 26775 15347 26781
rect 14608 26732 14614 26744
rect 15289 26741 15301 26775
rect 15335 26772 15347 26775
rect 15470 26772 15476 26784
rect 15335 26744 15476 26772
rect 15335 26741 15347 26744
rect 15289 26735 15347 26741
rect 15470 26732 15476 26744
rect 15528 26732 15534 26784
rect 16114 26772 16120 26784
rect 16075 26744 16120 26772
rect 16114 26732 16120 26744
rect 16172 26732 16178 26784
rect 17696 26772 17724 26803
rect 19242 26800 19248 26812
rect 19300 26800 19306 26852
rect 22002 26800 22008 26852
rect 22060 26840 22066 26852
rect 23109 26843 23167 26849
rect 23109 26840 23121 26843
rect 22060 26812 23121 26840
rect 22060 26800 22066 26812
rect 23109 26809 23121 26812
rect 23155 26809 23167 26843
rect 23109 26803 23167 26809
rect 24762 26800 24768 26852
rect 24820 26840 24826 26852
rect 24820 26812 25084 26840
rect 24820 26800 24826 26812
rect 18046 26772 18052 26784
rect 17696 26744 18052 26772
rect 18046 26732 18052 26744
rect 18104 26732 18110 26784
rect 18138 26732 18144 26784
rect 18196 26772 18202 26784
rect 20070 26772 20076 26784
rect 18196 26744 20076 26772
rect 18196 26732 18202 26744
rect 20070 26732 20076 26744
rect 20128 26732 20134 26784
rect 20717 26775 20775 26781
rect 20717 26741 20729 26775
rect 20763 26772 20775 26775
rect 20806 26772 20812 26784
rect 20763 26744 20812 26772
rect 20763 26741 20775 26744
rect 20717 26735 20775 26741
rect 20806 26732 20812 26744
rect 20864 26732 20870 26784
rect 21266 26732 21272 26784
rect 21324 26772 21330 26784
rect 21542 26772 21548 26784
rect 21324 26744 21548 26772
rect 21324 26732 21330 26744
rect 21542 26732 21548 26744
rect 21600 26732 21606 26784
rect 21634 26732 21640 26784
rect 21692 26772 21698 26784
rect 21821 26775 21879 26781
rect 21821 26772 21833 26775
rect 21692 26744 21833 26772
rect 21692 26732 21698 26744
rect 21821 26741 21833 26744
rect 21867 26741 21879 26775
rect 21821 26735 21879 26741
rect 22186 26732 22192 26784
rect 22244 26772 22250 26784
rect 22281 26775 22339 26781
rect 22281 26772 22293 26775
rect 22244 26744 22293 26772
rect 22244 26732 22250 26744
rect 22281 26741 22293 26744
rect 22327 26741 22339 26775
rect 22281 26735 22339 26741
rect 23566 26732 23572 26784
rect 23624 26772 23630 26784
rect 24949 26775 25007 26781
rect 24949 26772 24961 26775
rect 23624 26744 24961 26772
rect 23624 26732 23630 26744
rect 24949 26741 24961 26744
rect 24995 26741 25007 26775
rect 25056 26772 25084 26812
rect 25130 26800 25136 26852
rect 25188 26840 25194 26852
rect 25777 26843 25835 26849
rect 25777 26840 25789 26843
rect 25188 26812 25789 26840
rect 25188 26800 25194 26812
rect 25777 26809 25789 26812
rect 25823 26809 25835 26843
rect 25777 26803 25835 26809
rect 25682 26772 25688 26784
rect 25056 26744 25688 26772
rect 24949 26735 25007 26741
rect 25682 26732 25688 26744
rect 25740 26732 25746 26784
rect 1104 26682 28888 26704
rect 1104 26630 5582 26682
rect 5634 26630 5646 26682
rect 5698 26630 5710 26682
rect 5762 26630 5774 26682
rect 5826 26630 5838 26682
rect 5890 26630 14846 26682
rect 14898 26630 14910 26682
rect 14962 26630 14974 26682
rect 15026 26630 15038 26682
rect 15090 26630 15102 26682
rect 15154 26630 24110 26682
rect 24162 26630 24174 26682
rect 24226 26630 24238 26682
rect 24290 26630 24302 26682
rect 24354 26630 24366 26682
rect 24418 26630 28888 26682
rect 1104 26608 28888 26630
rect 10045 26571 10103 26577
rect 10045 26537 10057 26571
rect 10091 26568 10103 26571
rect 13538 26568 13544 26580
rect 10091 26540 13400 26568
rect 13499 26540 13544 26568
rect 10091 26537 10103 26540
rect 10045 26531 10103 26537
rect 12066 26500 12072 26512
rect 10888 26472 12072 26500
rect 9582 26364 9588 26376
rect 9543 26336 9588 26364
rect 9582 26324 9588 26336
rect 9640 26324 9646 26376
rect 9858 26324 9864 26376
rect 9916 26364 9922 26376
rect 10888 26373 10916 26472
rect 12066 26460 12072 26472
rect 12124 26460 12130 26512
rect 13372 26500 13400 26540
rect 13538 26528 13544 26540
rect 13596 26528 13602 26580
rect 14093 26571 14151 26577
rect 14093 26537 14105 26571
rect 14139 26568 14151 26571
rect 18414 26568 18420 26580
rect 14139 26540 18092 26568
rect 18375 26540 18420 26568
rect 14139 26537 14151 26540
rect 14093 26531 14151 26537
rect 15194 26500 15200 26512
rect 13372 26472 14504 26500
rect 15155 26472 15200 26500
rect 12158 26432 12164 26444
rect 12119 26404 12164 26432
rect 12158 26392 12164 26404
rect 12216 26392 12222 26444
rect 13354 26392 13360 26444
rect 13412 26432 13418 26444
rect 13906 26432 13912 26444
rect 13412 26404 13912 26432
rect 13412 26392 13418 26404
rect 13906 26392 13912 26404
rect 13964 26392 13970 26444
rect 10229 26367 10287 26373
rect 10229 26364 10241 26367
rect 9916 26336 10241 26364
rect 9916 26324 9922 26336
rect 10229 26333 10241 26336
rect 10275 26333 10287 26367
rect 10229 26327 10287 26333
rect 10873 26367 10931 26373
rect 10873 26333 10885 26367
rect 10919 26333 10931 26367
rect 11330 26364 11336 26376
rect 11291 26336 11336 26364
rect 10873 26327 10931 26333
rect 11330 26324 11336 26336
rect 11388 26324 11394 26376
rect 11514 26364 11520 26376
rect 11475 26336 11520 26364
rect 11514 26324 11520 26336
rect 11572 26324 11578 26376
rect 11882 26324 11888 26376
rect 11940 26364 11946 26376
rect 11940 26336 14228 26364
rect 11940 26324 11946 26336
rect 11606 26296 11612 26308
rect 10704 26268 11612 26296
rect 10704 26237 10732 26268
rect 11606 26256 11612 26268
rect 11664 26256 11670 26308
rect 11974 26256 11980 26308
rect 12032 26296 12038 26308
rect 12250 26296 12256 26308
rect 12032 26268 12256 26296
rect 12032 26256 12038 26268
rect 12250 26256 12256 26268
rect 12308 26256 12314 26308
rect 12428 26299 12486 26305
rect 12428 26265 12440 26299
rect 12474 26296 12486 26299
rect 12526 26296 12532 26308
rect 12474 26268 12532 26296
rect 12474 26265 12486 26268
rect 12428 26259 12486 26265
rect 12526 26256 12532 26268
rect 12584 26256 12590 26308
rect 12618 26256 12624 26308
rect 12676 26296 12682 26308
rect 13814 26296 13820 26308
rect 12676 26268 13820 26296
rect 12676 26256 12682 26268
rect 13814 26256 13820 26268
rect 13872 26256 13878 26308
rect 13998 26256 14004 26308
rect 14056 26296 14062 26308
rect 14093 26299 14151 26305
rect 14093 26296 14105 26299
rect 14056 26268 14105 26296
rect 14056 26256 14062 26268
rect 14093 26265 14105 26268
rect 14139 26265 14151 26299
rect 14200 26296 14228 26336
rect 14274 26324 14280 26376
rect 14332 26364 14338 26376
rect 14369 26367 14427 26373
rect 14369 26364 14381 26367
rect 14332 26336 14381 26364
rect 14332 26324 14338 26336
rect 14369 26333 14381 26336
rect 14415 26333 14427 26367
rect 14476 26364 14504 26472
rect 15194 26460 15200 26472
rect 15252 26460 15258 26512
rect 17129 26503 17187 26509
rect 17129 26469 17141 26503
rect 17175 26500 17187 26503
rect 17310 26500 17316 26512
rect 17175 26472 17316 26500
rect 17175 26469 17187 26472
rect 17129 26463 17187 26469
rect 17310 26460 17316 26472
rect 17368 26460 17374 26512
rect 17586 26460 17592 26512
rect 17644 26500 17650 26512
rect 17862 26500 17868 26512
rect 17644 26472 17868 26500
rect 17644 26460 17650 26472
rect 17862 26460 17868 26472
rect 17920 26460 17926 26512
rect 18064 26500 18092 26540
rect 18414 26528 18420 26540
rect 18472 26528 18478 26580
rect 18598 26528 18604 26580
rect 18656 26568 18662 26580
rect 19521 26571 19579 26577
rect 19521 26568 19533 26571
rect 18656 26540 19533 26568
rect 18656 26528 18662 26540
rect 19521 26537 19533 26540
rect 19567 26537 19579 26571
rect 19521 26531 19579 26537
rect 19610 26528 19616 26580
rect 19668 26568 19674 26580
rect 20162 26568 20168 26580
rect 19668 26540 20168 26568
rect 19668 26528 19674 26540
rect 20162 26528 20168 26540
rect 20220 26528 20226 26580
rect 21729 26571 21787 26577
rect 21729 26537 21741 26571
rect 21775 26568 21787 26571
rect 22278 26568 22284 26580
rect 21775 26540 22284 26568
rect 21775 26537 21787 26540
rect 21729 26531 21787 26537
rect 22278 26528 22284 26540
rect 22336 26528 22342 26580
rect 23842 26568 23848 26580
rect 22388 26540 23244 26568
rect 23803 26540 23848 26568
rect 22388 26500 22416 26540
rect 18064 26472 22416 26500
rect 22465 26503 22523 26509
rect 22465 26469 22477 26503
rect 22511 26469 22523 26503
rect 22465 26463 22523 26469
rect 14550 26392 14556 26444
rect 14608 26432 14614 26444
rect 14734 26432 14740 26444
rect 14608 26404 14740 26432
rect 14608 26392 14614 26404
rect 14734 26392 14740 26404
rect 14792 26432 14798 26444
rect 14829 26435 14887 26441
rect 14829 26432 14841 26435
rect 14792 26404 14841 26432
rect 14792 26392 14798 26404
rect 14829 26401 14841 26404
rect 14875 26401 14887 26435
rect 14829 26395 14887 26401
rect 14918 26392 14924 26444
rect 14976 26432 14982 26444
rect 15562 26432 15568 26444
rect 14976 26404 15568 26432
rect 14976 26392 14982 26404
rect 15562 26392 15568 26404
rect 15620 26392 15626 26444
rect 15746 26432 15752 26444
rect 15707 26404 15752 26432
rect 15746 26392 15752 26404
rect 15804 26392 15810 26444
rect 18138 26392 18144 26444
rect 18196 26432 18202 26444
rect 18322 26432 18328 26444
rect 18196 26404 18328 26432
rect 18196 26392 18202 26404
rect 18322 26392 18328 26404
rect 18380 26392 18386 26444
rect 18782 26432 18788 26444
rect 18524 26404 18788 26432
rect 16005 26367 16063 26373
rect 16005 26364 16017 26367
rect 14476 26336 16017 26364
rect 14369 26327 14427 26333
rect 16005 26333 16017 26336
rect 16051 26333 16063 26367
rect 17586 26364 17592 26376
rect 17547 26336 17592 26364
rect 16005 26327 16063 26333
rect 17586 26324 17592 26336
rect 17644 26324 17650 26376
rect 18524 26373 18552 26404
rect 18782 26392 18788 26404
rect 18840 26392 18846 26444
rect 19996 26404 20852 26432
rect 17681 26367 17739 26373
rect 17681 26333 17693 26367
rect 17727 26364 17739 26367
rect 18509 26367 18567 26373
rect 17727 26336 18460 26364
rect 17727 26333 17739 26336
rect 17681 26327 17739 26333
rect 18230 26296 18236 26308
rect 14200 26268 18092 26296
rect 18191 26268 18236 26296
rect 14093 26259 14151 26265
rect 10689 26231 10747 26237
rect 10689 26197 10701 26231
rect 10735 26197 10747 26231
rect 10689 26191 10747 26197
rect 10962 26188 10968 26240
rect 11020 26228 11026 26240
rect 11701 26231 11759 26237
rect 11701 26228 11713 26231
rect 11020 26200 11713 26228
rect 11020 26188 11026 26200
rect 11701 26197 11713 26200
rect 11747 26197 11759 26231
rect 11701 26191 11759 26197
rect 12342 26188 12348 26240
rect 12400 26228 12406 26240
rect 13078 26228 13084 26240
rect 12400 26200 13084 26228
rect 12400 26188 12406 26200
rect 13078 26188 13084 26200
rect 13136 26188 13142 26240
rect 13262 26188 13268 26240
rect 13320 26228 13326 26240
rect 14277 26231 14335 26237
rect 14277 26228 14289 26231
rect 13320 26200 14289 26228
rect 13320 26188 13326 26200
rect 14277 26197 14289 26200
rect 14323 26228 14335 26231
rect 15194 26228 15200 26240
rect 14323 26200 15200 26228
rect 14323 26197 14335 26200
rect 14277 26191 14335 26197
rect 15194 26188 15200 26200
rect 15252 26188 15258 26240
rect 15289 26231 15347 26237
rect 15289 26197 15301 26231
rect 15335 26228 15347 26231
rect 15930 26228 15936 26240
rect 15335 26200 15936 26228
rect 15335 26197 15347 26200
rect 15289 26191 15347 26197
rect 15930 26188 15936 26200
rect 15988 26188 15994 26240
rect 18064 26228 18092 26268
rect 18230 26256 18236 26268
rect 18288 26256 18294 26308
rect 18432 26296 18460 26336
rect 18509 26333 18521 26367
rect 18555 26333 18567 26367
rect 18509 26327 18567 26333
rect 18874 26324 18880 26376
rect 18932 26364 18938 26376
rect 19996 26373 20024 26404
rect 20824 26376 20852 26404
rect 21174 26392 21180 26444
rect 21232 26432 21238 26444
rect 21453 26435 21511 26441
rect 21453 26432 21465 26435
rect 21232 26404 21465 26432
rect 21232 26392 21238 26404
rect 21453 26401 21465 26404
rect 21499 26401 21511 26435
rect 21453 26395 21511 26401
rect 19797 26367 19855 26373
rect 19981 26367 20039 26373
rect 19797 26364 19809 26367
rect 18932 26336 19809 26364
rect 18932 26324 18938 26336
rect 19797 26333 19809 26336
rect 19843 26333 19855 26367
rect 19797 26327 19855 26333
rect 19886 26361 19944 26367
rect 19886 26327 19898 26361
rect 19932 26327 19944 26361
rect 19981 26333 19993 26367
rect 20027 26333 20039 26367
rect 20162 26364 20168 26376
rect 20123 26336 20168 26364
rect 19981 26327 20039 26333
rect 19886 26321 19944 26327
rect 20162 26324 20168 26336
rect 20220 26324 20226 26376
rect 20806 26324 20812 26376
rect 20864 26364 20870 26376
rect 21085 26367 21143 26373
rect 21085 26364 21097 26367
rect 20864 26336 21097 26364
rect 20864 26324 20870 26336
rect 21085 26333 21097 26336
rect 21131 26364 21143 26367
rect 22480 26364 22508 26463
rect 21131 26362 21496 26364
rect 21652 26362 22508 26364
rect 21131 26336 22508 26362
rect 21131 26333 21143 26336
rect 21468 26334 21680 26336
rect 21085 26327 21143 26333
rect 22738 26324 22744 26376
rect 22796 26364 22802 26376
rect 23109 26367 23167 26373
rect 23109 26364 23121 26367
rect 22796 26336 23121 26364
rect 22796 26324 22802 26336
rect 23109 26333 23121 26336
rect 23155 26333 23167 26367
rect 23216 26364 23244 26540
rect 23842 26528 23848 26540
rect 23900 26528 23906 26580
rect 24762 26568 24768 26580
rect 24723 26540 24768 26568
rect 24762 26528 24768 26540
rect 24820 26528 24826 26580
rect 24946 26568 24952 26580
rect 24907 26540 24952 26568
rect 24946 26528 24952 26540
rect 25004 26568 25010 26580
rect 25774 26568 25780 26580
rect 25004 26540 25780 26568
rect 25004 26528 25010 26540
rect 25774 26528 25780 26540
rect 25832 26528 25838 26580
rect 23290 26460 23296 26512
rect 23348 26500 23354 26512
rect 23348 26472 23520 26500
rect 23348 26460 23354 26472
rect 23382 26432 23388 26444
rect 23343 26404 23388 26432
rect 23382 26392 23388 26404
rect 23440 26392 23446 26444
rect 23492 26441 23520 26472
rect 23477 26435 23535 26441
rect 23477 26401 23489 26435
rect 23523 26401 23535 26435
rect 23477 26395 23535 26401
rect 23566 26392 23572 26444
rect 23624 26432 23630 26444
rect 26513 26435 26571 26441
rect 26513 26432 26525 26435
rect 23624 26404 26525 26432
rect 23624 26392 23630 26404
rect 26513 26401 26525 26404
rect 26559 26401 26571 26435
rect 28166 26432 28172 26444
rect 28127 26404 28172 26432
rect 26513 26395 26571 26401
rect 28166 26392 28172 26404
rect 28224 26392 28230 26444
rect 23293 26367 23351 26373
rect 23293 26364 23305 26367
rect 23216 26336 23305 26364
rect 23109 26327 23167 26333
rect 23293 26333 23305 26336
rect 23339 26333 23351 26367
rect 23658 26364 23664 26376
rect 23619 26336 23664 26364
rect 23293 26327 23351 26333
rect 23658 26324 23664 26336
rect 23716 26324 23722 26376
rect 25590 26364 25596 26376
rect 24811 26333 24869 26339
rect 25551 26336 25596 26364
rect 24811 26330 24823 26333
rect 19702 26296 19708 26308
rect 18432 26268 19708 26296
rect 19702 26256 19708 26268
rect 19760 26256 19766 26308
rect 19904 26240 19932 26321
rect 20990 26256 20996 26308
rect 21048 26296 21054 26308
rect 21570 26299 21628 26305
rect 21570 26296 21582 26299
rect 21048 26268 21582 26296
rect 21048 26256 21054 26268
rect 21570 26265 21582 26268
rect 21616 26296 21628 26299
rect 22189 26299 22247 26305
rect 22189 26296 22201 26299
rect 21616 26268 22201 26296
rect 21616 26265 21628 26268
rect 21570 26259 21628 26265
rect 22189 26265 22201 26268
rect 22235 26265 22247 26299
rect 24578 26296 24584 26308
rect 24539 26268 24584 26296
rect 22189 26259 22247 26265
rect 24578 26256 24584 26268
rect 24636 26256 24642 26308
rect 24796 26299 24823 26330
rect 24857 26308 24869 26333
rect 25590 26324 25596 26336
rect 25648 26324 25654 26376
rect 25869 26367 25927 26373
rect 25869 26333 25881 26367
rect 25915 26364 25927 26367
rect 25958 26364 25964 26376
rect 25915 26336 25964 26364
rect 25915 26333 25927 26336
rect 25869 26327 25927 26333
rect 25958 26324 25964 26336
rect 26016 26324 26022 26376
rect 26050 26324 26056 26376
rect 26108 26364 26114 26376
rect 26329 26367 26387 26373
rect 26329 26364 26341 26367
rect 26108 26336 26341 26364
rect 26108 26324 26114 26336
rect 26329 26333 26341 26336
rect 26375 26333 26387 26367
rect 26329 26327 26387 26333
rect 24857 26299 24860 26308
rect 24796 26268 24860 26299
rect 24854 26256 24860 26268
rect 24912 26256 24918 26308
rect 18598 26228 18604 26240
rect 18064 26200 18604 26228
rect 18598 26188 18604 26200
rect 18656 26188 18662 26240
rect 18693 26231 18751 26237
rect 18693 26197 18705 26231
rect 18739 26228 18751 26231
rect 18874 26228 18880 26240
rect 18739 26200 18880 26228
rect 18739 26197 18751 26200
rect 18693 26191 18751 26197
rect 18874 26188 18880 26200
rect 18932 26188 18938 26240
rect 19886 26188 19892 26240
rect 19944 26188 19950 26240
rect 21082 26188 21088 26240
rect 21140 26228 21146 26240
rect 21361 26231 21419 26237
rect 21361 26228 21373 26231
rect 21140 26200 21373 26228
rect 21140 26188 21146 26200
rect 21361 26197 21373 26200
rect 21407 26197 21419 26231
rect 21361 26191 21419 26197
rect 22370 26188 22376 26240
rect 22428 26228 22434 26240
rect 22649 26231 22707 26237
rect 22649 26228 22661 26231
rect 22428 26200 22661 26228
rect 22428 26188 22434 26200
rect 22649 26197 22661 26200
rect 22695 26197 22707 26231
rect 22649 26191 22707 26197
rect 25409 26231 25467 26237
rect 25409 26197 25421 26231
rect 25455 26228 25467 26231
rect 25498 26228 25504 26240
rect 25455 26200 25504 26228
rect 25455 26197 25467 26200
rect 25409 26191 25467 26197
rect 25498 26188 25504 26200
rect 25556 26188 25562 26240
rect 1104 26138 28888 26160
rect 1104 26086 10214 26138
rect 10266 26086 10278 26138
rect 10330 26086 10342 26138
rect 10394 26086 10406 26138
rect 10458 26086 10470 26138
rect 10522 26086 19478 26138
rect 19530 26086 19542 26138
rect 19594 26086 19606 26138
rect 19658 26086 19670 26138
rect 19722 26086 19734 26138
rect 19786 26086 28888 26138
rect 1104 26064 28888 26086
rect 9493 26027 9551 26033
rect 9493 25993 9505 26027
rect 9539 25993 9551 26027
rect 9493 25987 9551 25993
rect 10137 26027 10195 26033
rect 10137 25993 10149 26027
rect 10183 26024 10195 26027
rect 10183 25996 16048 26024
rect 10183 25993 10195 25996
rect 10137 25987 10195 25993
rect 9508 25956 9536 25987
rect 13538 25956 13544 25968
rect 9508 25928 10640 25956
rect 9677 25891 9735 25897
rect 9677 25857 9689 25891
rect 9723 25857 9735 25891
rect 9677 25851 9735 25857
rect 10321 25891 10379 25897
rect 10321 25857 10333 25891
rect 10367 25857 10379 25891
rect 10321 25851 10379 25857
rect 9692 25684 9720 25851
rect 10336 25752 10364 25851
rect 10612 25820 10640 25928
rect 11532 25928 13544 25956
rect 10778 25888 10784 25900
rect 10739 25860 10784 25888
rect 10778 25848 10784 25860
rect 10836 25848 10842 25900
rect 10873 25891 10931 25897
rect 10873 25857 10885 25891
rect 10919 25888 10931 25891
rect 11330 25888 11336 25900
rect 10919 25860 11336 25888
rect 10919 25857 10931 25860
rect 10873 25851 10931 25857
rect 11330 25848 11336 25860
rect 11388 25848 11394 25900
rect 11422 25848 11428 25900
rect 11480 25888 11486 25900
rect 11532 25897 11560 25928
rect 13538 25916 13544 25928
rect 13596 25916 13602 25968
rect 15866 25959 15924 25965
rect 15866 25956 15878 25959
rect 13740 25928 14964 25956
rect 11517 25891 11575 25897
rect 11517 25888 11529 25891
rect 11480 25860 11529 25888
rect 11480 25848 11486 25860
rect 11517 25857 11529 25860
rect 11563 25857 11575 25891
rect 11773 25891 11831 25897
rect 11773 25888 11785 25891
rect 11517 25851 11575 25857
rect 11624 25860 11785 25888
rect 11624 25820 11652 25860
rect 11773 25857 11785 25860
rect 11819 25857 11831 25891
rect 11773 25851 11831 25857
rect 12158 25848 12164 25900
rect 12216 25888 12222 25900
rect 13262 25888 13268 25900
rect 12216 25860 13268 25888
rect 12216 25848 12222 25860
rect 13262 25848 13268 25860
rect 13320 25848 13326 25900
rect 13740 25888 13768 25928
rect 13814 25897 13820 25900
rect 13378 25860 13768 25888
rect 10612 25792 11652 25820
rect 10336 25724 11563 25752
rect 11238 25684 11244 25696
rect 9692 25656 11244 25684
rect 11238 25644 11244 25656
rect 11296 25644 11302 25696
rect 11535 25684 11563 25724
rect 12618 25712 12624 25764
rect 12676 25752 12682 25764
rect 12897 25755 12955 25761
rect 12897 25752 12909 25755
rect 12676 25724 12909 25752
rect 12676 25712 12682 25724
rect 12897 25721 12909 25724
rect 12943 25721 12955 25755
rect 12897 25715 12955 25721
rect 13378 25684 13406 25860
rect 13808 25851 13820 25897
rect 13872 25888 13878 25900
rect 13872 25860 13908 25888
rect 13814 25848 13820 25851
rect 13872 25848 13878 25860
rect 14826 25848 14832 25900
rect 14884 25848 14890 25900
rect 13538 25820 13544 25832
rect 13451 25792 13544 25820
rect 13538 25780 13544 25792
rect 13596 25780 13602 25832
rect 11535 25656 13406 25684
rect 13556 25684 13584 25780
rect 14844 25752 14872 25848
rect 14936 25820 14964 25928
rect 15028 25928 15878 25956
rect 15028 25900 15056 25928
rect 15866 25925 15878 25928
rect 15912 25925 15924 25959
rect 16020 25956 16048 25996
rect 16574 25984 16580 26036
rect 16632 26024 16638 26036
rect 21269 26027 21327 26033
rect 16632 25996 19334 26024
rect 16632 25984 16638 25996
rect 16020 25928 16344 25956
rect 15866 25919 15924 25925
rect 15010 25848 15016 25900
rect 15068 25848 15074 25900
rect 15102 25848 15108 25900
rect 15160 25888 15166 25900
rect 15381 25891 15439 25897
rect 15381 25888 15393 25891
rect 15160 25860 15393 25888
rect 15160 25848 15166 25860
rect 15381 25857 15393 25860
rect 15427 25857 15439 25891
rect 16206 25888 16212 25900
rect 15381 25851 15439 25857
rect 15488 25860 16212 25888
rect 15488 25820 15516 25860
rect 16206 25848 16212 25860
rect 16264 25848 16270 25900
rect 14936 25792 15516 25820
rect 15657 25823 15715 25829
rect 15657 25789 15669 25823
rect 15703 25789 15715 25823
rect 15657 25783 15715 25789
rect 14476 25724 14872 25752
rect 13722 25684 13728 25696
rect 13556 25656 13728 25684
rect 13722 25644 13728 25656
rect 13780 25684 13786 25696
rect 14476 25684 14504 25724
rect 15672 25696 15700 25783
rect 15746 25780 15752 25832
rect 15804 25820 15810 25832
rect 16316 25820 16344 25928
rect 16684 25928 18552 25956
rect 16390 25848 16396 25900
rect 16448 25888 16454 25900
rect 16684 25897 16712 25928
rect 18524 25900 18552 25928
rect 18598 25916 18604 25968
rect 18656 25956 18662 25968
rect 18754 25959 18812 25965
rect 18754 25956 18766 25959
rect 18656 25928 18766 25956
rect 18656 25916 18662 25928
rect 18754 25925 18766 25928
rect 18800 25925 18812 25959
rect 19306 25956 19334 25996
rect 21269 25993 21281 26027
rect 21315 26024 21327 26027
rect 22186 26024 22192 26036
rect 21315 25996 22192 26024
rect 21315 25993 21327 25996
rect 21269 25987 21327 25993
rect 22186 25984 22192 25996
rect 22244 25984 22250 26036
rect 27338 26024 27344 26036
rect 22572 25996 27344 26024
rect 19306 25928 21772 25956
rect 18754 25919 18812 25925
rect 16669 25891 16727 25897
rect 16669 25888 16681 25891
rect 16448 25860 16681 25888
rect 16448 25848 16454 25860
rect 16669 25857 16681 25860
rect 16715 25857 16727 25891
rect 16925 25891 16983 25897
rect 16925 25888 16937 25891
rect 16669 25851 16727 25857
rect 16776 25860 16937 25888
rect 16776 25820 16804 25860
rect 16925 25857 16937 25860
rect 16971 25857 16983 25891
rect 16925 25851 16983 25857
rect 17678 25848 17684 25900
rect 17736 25888 17742 25900
rect 18322 25888 18328 25900
rect 17736 25860 18328 25888
rect 17736 25848 17742 25860
rect 18322 25848 18328 25860
rect 18380 25848 18386 25900
rect 18506 25888 18512 25900
rect 18467 25860 18512 25888
rect 18506 25848 18512 25860
rect 18564 25848 18570 25900
rect 19150 25848 19156 25900
rect 19208 25888 19214 25900
rect 19208 25860 20714 25888
rect 19208 25848 19214 25860
rect 15804 25792 15849 25820
rect 16316 25792 16804 25820
rect 20686 25820 20714 25860
rect 20806 25848 20812 25900
rect 20864 25888 20870 25900
rect 20864 25860 20909 25888
rect 20864 25848 20870 25860
rect 21634 25820 21640 25832
rect 20686 25792 21640 25820
rect 15804 25780 15810 25792
rect 21634 25780 21640 25792
rect 21692 25780 21698 25832
rect 16022 25752 16028 25764
rect 15983 25724 16028 25752
rect 16022 25712 16028 25724
rect 16080 25752 16086 25764
rect 16080 25724 16574 25752
rect 16080 25712 16086 25724
rect 13780 25656 14504 25684
rect 13780 25644 13786 25656
rect 14550 25644 14556 25696
rect 14608 25684 14614 25696
rect 14921 25687 14979 25693
rect 14921 25684 14933 25687
rect 14608 25656 14933 25684
rect 14608 25644 14614 25656
rect 14921 25653 14933 25656
rect 14967 25684 14979 25687
rect 15654 25684 15660 25696
rect 14967 25656 15660 25684
rect 14967 25653 14979 25656
rect 14921 25647 14979 25653
rect 15654 25644 15660 25656
rect 15712 25644 15718 25696
rect 16546 25684 16574 25724
rect 20990 25712 20996 25764
rect 21048 25752 21054 25764
rect 21085 25755 21143 25761
rect 21085 25752 21097 25755
rect 21048 25724 21097 25752
rect 21048 25712 21054 25724
rect 21085 25721 21097 25724
rect 21131 25721 21143 25755
rect 21744 25752 21772 25928
rect 21818 25916 21824 25968
rect 21876 25956 21882 25968
rect 21876 25928 22324 25956
rect 21876 25916 21882 25928
rect 21913 25891 21971 25897
rect 21913 25857 21925 25891
rect 21959 25888 21971 25891
rect 22002 25888 22008 25900
rect 21959 25860 22008 25888
rect 21959 25857 21971 25860
rect 21913 25851 21971 25857
rect 22002 25848 22008 25860
rect 22060 25848 22066 25900
rect 22094 25848 22100 25900
rect 22152 25888 22158 25900
rect 22296 25897 22324 25928
rect 22281 25891 22339 25897
rect 22152 25860 22197 25888
rect 22152 25848 22158 25860
rect 22281 25857 22293 25891
rect 22327 25857 22339 25891
rect 22281 25851 22339 25857
rect 22370 25848 22376 25900
rect 22428 25888 22434 25900
rect 22465 25891 22523 25897
rect 22465 25888 22477 25891
rect 22428 25860 22477 25888
rect 22428 25848 22434 25860
rect 22465 25857 22477 25860
rect 22511 25857 22523 25891
rect 22465 25851 22523 25857
rect 22186 25780 22192 25832
rect 22244 25820 22250 25832
rect 22244 25792 22289 25820
rect 22244 25780 22250 25792
rect 22572 25752 22600 25996
rect 27338 25984 27344 25996
rect 27396 25984 27402 26036
rect 27614 25984 27620 26036
rect 27672 26024 27678 26036
rect 28169 26027 28227 26033
rect 28169 26024 28181 26027
rect 27672 25996 28181 26024
rect 27672 25984 27678 25996
rect 28169 25993 28181 25996
rect 28215 25993 28227 26027
rect 28169 25987 28227 25993
rect 27062 25916 27068 25968
rect 27120 25956 27126 25968
rect 27801 25959 27859 25965
rect 27801 25956 27813 25959
rect 27120 25928 27813 25956
rect 27120 25916 27126 25928
rect 27801 25925 27813 25928
rect 27847 25925 27859 25959
rect 28001 25959 28059 25965
rect 28001 25956 28013 25959
rect 27801 25919 27859 25925
rect 27908 25928 28013 25956
rect 23385 25891 23443 25897
rect 23385 25857 23397 25891
rect 23431 25857 23443 25891
rect 23385 25851 23443 25857
rect 22646 25780 22652 25832
rect 22704 25820 22710 25832
rect 22830 25820 22836 25832
rect 22704 25792 22836 25820
rect 22704 25780 22710 25792
rect 22830 25780 22836 25792
rect 22888 25820 22894 25832
rect 23293 25823 23351 25829
rect 23293 25820 23305 25823
rect 22888 25792 23305 25820
rect 22888 25780 22894 25792
rect 23293 25789 23305 25792
rect 23339 25789 23351 25823
rect 23400 25820 23428 25851
rect 23566 25848 23572 25900
rect 23624 25888 23630 25900
rect 24213 25891 24271 25897
rect 24213 25888 24225 25891
rect 23624 25860 24225 25888
rect 23624 25848 23630 25860
rect 24213 25857 24225 25860
rect 24259 25857 24271 25891
rect 24213 25851 24271 25857
rect 24397 25891 24455 25897
rect 24397 25857 24409 25891
rect 24443 25888 24455 25891
rect 24486 25888 24492 25900
rect 24443 25860 24492 25888
rect 24443 25857 24455 25860
rect 24397 25851 24455 25857
rect 24486 25848 24492 25860
rect 24544 25848 24550 25900
rect 24670 25848 24676 25900
rect 24728 25888 24734 25900
rect 25297 25891 25355 25897
rect 25297 25888 25309 25891
rect 24728 25860 25309 25888
rect 24728 25848 24734 25860
rect 25297 25857 25309 25860
rect 25343 25857 25355 25891
rect 25297 25851 25355 25857
rect 25774 25848 25780 25900
rect 25832 25888 25838 25900
rect 27157 25891 27215 25897
rect 27157 25888 27169 25891
rect 25832 25860 27169 25888
rect 25832 25848 25838 25860
rect 27157 25857 27169 25860
rect 27203 25888 27215 25891
rect 27908 25888 27936 25928
rect 28001 25925 28013 25928
rect 28047 25925 28059 25959
rect 28001 25919 28059 25925
rect 27203 25860 27936 25888
rect 27203 25857 27215 25860
rect 27157 25851 27215 25857
rect 23658 25820 23664 25832
rect 23400 25792 23664 25820
rect 23293 25783 23351 25789
rect 23658 25780 23664 25792
rect 23716 25820 23722 25832
rect 24026 25820 24032 25832
rect 23716 25792 24032 25820
rect 23716 25780 23722 25792
rect 24026 25780 24032 25792
rect 24084 25780 24090 25832
rect 25038 25820 25044 25832
rect 24999 25792 25044 25820
rect 25038 25780 25044 25792
rect 25096 25780 25102 25832
rect 26050 25780 26056 25832
rect 26108 25820 26114 25832
rect 26973 25823 27031 25829
rect 26973 25820 26985 25823
rect 26108 25792 26985 25820
rect 26108 25780 26114 25792
rect 26973 25789 26985 25792
rect 27019 25789 27031 25823
rect 26973 25783 27031 25789
rect 21744 25724 22600 25752
rect 21085 25715 21143 25721
rect 22922 25712 22928 25764
rect 22980 25752 22986 25764
rect 26418 25752 26424 25764
rect 22980 25724 24716 25752
rect 26379 25724 26424 25752
rect 22980 25712 22986 25724
rect 16850 25684 16856 25696
rect 16546 25656 16856 25684
rect 16850 25644 16856 25656
rect 16908 25644 16914 25696
rect 18046 25684 18052 25696
rect 18007 25656 18052 25684
rect 18046 25644 18052 25656
rect 18104 25644 18110 25696
rect 18230 25644 18236 25696
rect 18288 25684 18294 25696
rect 19889 25687 19947 25693
rect 19889 25684 19901 25687
rect 18288 25656 19901 25684
rect 18288 25644 18294 25656
rect 19889 25653 19901 25656
rect 19935 25653 19947 25687
rect 19889 25647 19947 25653
rect 22462 25644 22468 25696
rect 22520 25684 22526 25696
rect 22649 25687 22707 25693
rect 22649 25684 22661 25687
rect 22520 25656 22661 25684
rect 22520 25644 22526 25656
rect 22649 25653 22661 25656
rect 22695 25653 22707 25687
rect 22649 25647 22707 25653
rect 23474 25644 23480 25696
rect 23532 25684 23538 25696
rect 23753 25687 23811 25693
rect 23753 25684 23765 25687
rect 23532 25656 23765 25684
rect 23532 25644 23538 25656
rect 23753 25653 23765 25656
rect 23799 25684 23811 25687
rect 23842 25684 23848 25696
rect 23799 25656 23848 25684
rect 23799 25653 23811 25656
rect 23753 25647 23811 25653
rect 23842 25644 23848 25656
rect 23900 25644 23906 25696
rect 24578 25684 24584 25696
rect 24539 25656 24584 25684
rect 24578 25644 24584 25656
rect 24636 25644 24642 25696
rect 24688 25684 24716 25724
rect 26418 25712 26424 25724
rect 26476 25712 26482 25764
rect 25222 25684 25228 25696
rect 24688 25656 25228 25684
rect 25222 25644 25228 25656
rect 25280 25644 25286 25696
rect 26988 25684 27016 25783
rect 27985 25687 28043 25693
rect 27985 25684 27997 25687
rect 26988 25656 27997 25684
rect 27985 25653 27997 25656
rect 28031 25653 28043 25687
rect 27985 25647 28043 25653
rect 1104 25594 28888 25616
rect 1104 25542 5582 25594
rect 5634 25542 5646 25594
rect 5698 25542 5710 25594
rect 5762 25542 5774 25594
rect 5826 25542 5838 25594
rect 5890 25542 14846 25594
rect 14898 25542 14910 25594
rect 14962 25542 14974 25594
rect 15026 25542 15038 25594
rect 15090 25542 15102 25594
rect 15154 25542 24110 25594
rect 24162 25542 24174 25594
rect 24226 25542 24238 25594
rect 24290 25542 24302 25594
rect 24354 25542 24366 25594
rect 24418 25542 28888 25594
rect 1104 25520 28888 25542
rect 9493 25483 9551 25489
rect 9493 25449 9505 25483
rect 9539 25480 9551 25483
rect 11054 25480 11060 25492
rect 9539 25452 11060 25480
rect 9539 25449 9551 25452
rect 9493 25443 9551 25449
rect 11054 25440 11060 25452
rect 11112 25440 11118 25492
rect 11330 25440 11336 25492
rect 11388 25480 11394 25492
rect 19886 25480 19892 25492
rect 11388 25452 19892 25480
rect 11388 25440 11394 25452
rect 19886 25440 19892 25452
rect 19944 25440 19950 25492
rect 21082 25440 21088 25492
rect 21140 25480 21146 25492
rect 21361 25483 21419 25489
rect 21361 25480 21373 25483
rect 21140 25452 21373 25480
rect 21140 25440 21146 25452
rect 21361 25449 21373 25452
rect 21407 25449 21419 25483
rect 21361 25443 21419 25449
rect 21634 25440 21640 25492
rect 21692 25480 21698 25492
rect 23293 25483 23351 25489
rect 21692 25452 22600 25480
rect 21692 25440 21698 25452
rect 12710 25372 12716 25424
rect 12768 25412 12774 25424
rect 12805 25415 12863 25421
rect 12805 25412 12817 25415
rect 12768 25384 12817 25412
rect 12768 25372 12774 25384
rect 12805 25381 12817 25384
rect 12851 25412 12863 25415
rect 12986 25412 12992 25424
rect 12851 25384 12992 25412
rect 12851 25381 12863 25384
rect 12805 25375 12863 25381
rect 12986 25372 12992 25384
rect 13044 25372 13050 25424
rect 13998 25372 14004 25424
rect 14056 25412 14062 25424
rect 14056 25384 16252 25412
rect 14056 25372 14062 25384
rect 10873 25347 10931 25353
rect 10873 25313 10885 25347
rect 10919 25344 10931 25347
rect 11422 25344 11428 25356
rect 10919 25316 11284 25344
rect 11383 25316 11428 25344
rect 10919 25313 10931 25316
rect 10873 25307 10931 25313
rect 9677 25279 9735 25285
rect 9677 25245 9689 25279
rect 9723 25245 9735 25279
rect 9677 25239 9735 25245
rect 10321 25279 10379 25285
rect 10321 25245 10333 25279
rect 10367 25276 10379 25279
rect 10594 25276 10600 25288
rect 10367 25248 10600 25276
rect 10367 25245 10379 25248
rect 10321 25239 10379 25245
rect 9692 25208 9720 25239
rect 10594 25236 10600 25248
rect 10652 25236 10658 25288
rect 10778 25276 10784 25288
rect 10739 25248 10784 25276
rect 10778 25236 10784 25248
rect 10836 25236 10842 25288
rect 10965 25279 11023 25285
rect 10965 25245 10977 25279
rect 11011 25276 11023 25279
rect 11146 25276 11152 25288
rect 11011 25248 11152 25276
rect 11011 25245 11023 25248
rect 10965 25239 11023 25245
rect 11146 25236 11152 25248
rect 11204 25236 11210 25288
rect 11256 25276 11284 25316
rect 11422 25304 11428 25316
rect 11480 25304 11486 25356
rect 15010 25344 15016 25356
rect 14568 25316 15016 25344
rect 14274 25276 14280 25288
rect 11256 25248 14280 25276
rect 14274 25236 14280 25248
rect 14332 25236 14338 25288
rect 14369 25279 14427 25285
rect 14369 25245 14381 25279
rect 14415 25276 14427 25279
rect 14458 25276 14464 25288
rect 14415 25248 14464 25276
rect 14415 25245 14427 25248
rect 14369 25239 14427 25245
rect 14458 25236 14464 25248
rect 14516 25236 14522 25288
rect 14568 25285 14596 25316
rect 15010 25304 15016 25316
rect 15068 25304 15074 25356
rect 15394 25353 15400 25356
rect 15390 25344 15400 25353
rect 15355 25316 15400 25344
rect 15390 25307 15400 25316
rect 15394 25304 15400 25307
rect 15452 25304 15458 25356
rect 16114 25344 16120 25356
rect 15534 25316 16120 25344
rect 14553 25279 14611 25285
rect 14553 25245 14565 25279
rect 14599 25245 14611 25279
rect 14553 25239 14611 25245
rect 14642 25236 14648 25288
rect 14700 25276 14706 25288
rect 15105 25279 15163 25285
rect 15105 25276 15117 25279
rect 14700 25248 15117 25276
rect 14700 25236 14706 25248
rect 15105 25245 15117 25248
rect 15151 25245 15163 25279
rect 15105 25239 15163 25245
rect 11054 25208 11060 25220
rect 9692 25180 11060 25208
rect 11054 25168 11060 25180
rect 11112 25168 11118 25220
rect 11514 25168 11520 25220
rect 11572 25208 11578 25220
rect 11670 25211 11728 25217
rect 11670 25208 11682 25211
rect 11572 25180 11682 25208
rect 11572 25168 11578 25180
rect 11670 25177 11682 25180
rect 11716 25177 11728 25211
rect 11670 25171 11728 25177
rect 12526 25168 12532 25220
rect 12584 25208 12590 25220
rect 13170 25208 13176 25220
rect 12584 25180 13176 25208
rect 12584 25168 12590 25180
rect 13170 25168 13176 25180
rect 13228 25168 13234 25220
rect 13354 25208 13360 25220
rect 13315 25180 13360 25208
rect 13354 25168 13360 25180
rect 13412 25168 13418 25220
rect 13541 25211 13599 25217
rect 13541 25177 13553 25211
rect 13587 25208 13599 25211
rect 15120 25208 15148 25239
rect 15194 25236 15200 25288
rect 15252 25276 15258 25288
rect 15534 25285 15562 25316
rect 16114 25304 16120 25316
rect 16172 25304 16178 25356
rect 15289 25279 15347 25285
rect 15289 25276 15301 25279
rect 15252 25248 15301 25276
rect 15252 25236 15258 25248
rect 15289 25245 15301 25248
rect 15335 25245 15347 25279
rect 15289 25239 15347 25245
rect 15519 25279 15577 25285
rect 15519 25245 15531 25279
rect 15565 25245 15577 25279
rect 15519 25239 15577 25245
rect 15657 25279 15715 25285
rect 15657 25245 15669 25279
rect 15703 25276 15715 25279
rect 15930 25276 15936 25288
rect 15703 25248 15936 25276
rect 15703 25245 15715 25248
rect 15657 25239 15715 25245
rect 15930 25236 15936 25248
rect 15988 25236 15994 25288
rect 16224 25276 16252 25384
rect 17954 25372 17960 25424
rect 18012 25412 18018 25424
rect 18693 25415 18751 25421
rect 18693 25412 18705 25415
rect 18012 25384 18705 25412
rect 18012 25372 18018 25384
rect 18693 25381 18705 25384
rect 18739 25381 18751 25415
rect 18693 25375 18751 25381
rect 22278 25372 22284 25424
rect 22336 25412 22342 25424
rect 22572 25412 22600 25452
rect 23293 25449 23305 25483
rect 23339 25480 23351 25483
rect 23382 25480 23388 25492
rect 23339 25452 23388 25480
rect 23339 25449 23351 25452
rect 23293 25443 23351 25449
rect 23382 25440 23388 25452
rect 23440 25440 23446 25492
rect 24670 25480 24676 25492
rect 24631 25452 24676 25480
rect 24670 25440 24676 25452
rect 24728 25440 24734 25492
rect 22336 25384 22508 25412
rect 22572 25384 23704 25412
rect 22336 25372 22342 25384
rect 16390 25344 16396 25356
rect 16351 25316 16396 25344
rect 16390 25304 16396 25316
rect 16448 25304 16454 25356
rect 18138 25304 18144 25356
rect 18196 25344 18202 25356
rect 18196 25316 18460 25344
rect 18196 25304 18202 25316
rect 16649 25279 16707 25285
rect 16649 25276 16661 25279
rect 16224 25248 16661 25276
rect 16649 25245 16661 25248
rect 16695 25245 16707 25279
rect 17034 25276 17040 25288
rect 16649 25239 16707 25245
rect 16868 25248 17040 25276
rect 13587 25180 15056 25208
rect 15120 25180 15969 25208
rect 13587 25177 13599 25180
rect 13541 25171 13599 25177
rect 10137 25143 10195 25149
rect 10137 25109 10149 25143
rect 10183 25140 10195 25143
rect 13998 25140 14004 25152
rect 10183 25112 14004 25140
rect 10183 25109 10195 25112
rect 10137 25103 10195 25109
rect 13998 25100 14004 25112
rect 14056 25100 14062 25152
rect 14093 25143 14151 25149
rect 14093 25109 14105 25143
rect 14139 25140 14151 25143
rect 14918 25140 14924 25152
rect 14139 25112 14924 25140
rect 14139 25109 14151 25112
rect 14093 25103 14151 25109
rect 14918 25100 14924 25112
rect 14976 25100 14982 25152
rect 15028 25140 15056 25180
rect 15562 25140 15568 25152
rect 15028 25112 15568 25140
rect 15562 25100 15568 25112
rect 15620 25100 15626 25152
rect 15838 25140 15844 25152
rect 15799 25112 15844 25140
rect 15838 25100 15844 25112
rect 15896 25100 15902 25152
rect 15941 25140 15969 25180
rect 16206 25168 16212 25220
rect 16264 25208 16270 25220
rect 16868 25208 16896 25248
rect 17034 25236 17040 25248
rect 17092 25236 17098 25288
rect 18432 25285 18460 25316
rect 19150 25304 19156 25356
rect 19208 25344 19214 25356
rect 19981 25347 20039 25353
rect 19981 25344 19993 25347
rect 19208 25316 19993 25344
rect 19208 25304 19214 25316
rect 19981 25313 19993 25316
rect 20027 25313 20039 25347
rect 19981 25307 20039 25313
rect 18417 25279 18475 25285
rect 18417 25245 18429 25279
rect 18463 25245 18475 25279
rect 18417 25239 18475 25245
rect 18512 25279 18570 25285
rect 18512 25245 18524 25279
rect 18558 25276 18570 25279
rect 18598 25276 18604 25288
rect 18558 25248 18604 25276
rect 18558 25245 18570 25248
rect 18512 25239 18570 25245
rect 18598 25236 18604 25248
rect 18656 25236 18662 25288
rect 18690 25236 18696 25288
rect 18748 25276 18754 25288
rect 19245 25279 19303 25285
rect 19245 25276 19257 25279
rect 18748 25248 19257 25276
rect 18748 25236 18754 25248
rect 19245 25245 19257 25248
rect 19291 25245 19303 25279
rect 19996 25276 20024 25307
rect 20622 25276 20628 25288
rect 19996 25248 20628 25276
rect 19245 25239 19303 25245
rect 20622 25236 20628 25248
rect 20680 25236 20686 25288
rect 22094 25236 22100 25288
rect 22152 25276 22158 25288
rect 22370 25285 22376 25288
rect 22189 25279 22247 25285
rect 22189 25276 22201 25279
rect 22152 25248 22201 25276
rect 22152 25236 22158 25248
rect 22189 25245 22201 25248
rect 22235 25245 22247 25279
rect 22189 25239 22247 25245
rect 22354 25279 22376 25285
rect 22354 25245 22366 25279
rect 22354 25239 22376 25245
rect 22370 25236 22376 25239
rect 22428 25236 22434 25288
rect 22480 25285 22508 25384
rect 23676 25353 23704 25384
rect 23661 25347 23719 25353
rect 23661 25313 23673 25347
rect 23707 25313 23719 25347
rect 28166 25344 28172 25356
rect 28127 25316 28172 25344
rect 23661 25307 23719 25313
rect 28166 25304 28172 25316
rect 28224 25304 28230 25356
rect 22465 25279 22523 25285
rect 22465 25245 22477 25279
rect 22511 25245 22523 25279
rect 22465 25239 22523 25245
rect 22554 25236 22560 25288
rect 22612 25276 22618 25288
rect 23474 25276 23480 25288
rect 22612 25248 22657 25276
rect 23435 25248 23480 25276
rect 22612 25236 22618 25248
rect 23474 25236 23480 25248
rect 23532 25236 23538 25288
rect 23569 25279 23627 25285
rect 23569 25245 23581 25279
rect 23615 25245 23627 25279
rect 23753 25279 23811 25285
rect 23753 25276 23765 25279
rect 23569 25239 23627 25245
rect 23676 25248 23765 25276
rect 16264 25180 16896 25208
rect 16264 25168 16270 25180
rect 16942 25168 16948 25220
rect 17000 25208 17006 25220
rect 20226 25211 20284 25217
rect 20226 25208 20238 25211
rect 17000 25180 20238 25208
rect 17000 25168 17006 25180
rect 20226 25177 20238 25180
rect 20272 25177 20284 25211
rect 20226 25171 20284 25177
rect 17218 25140 17224 25152
rect 15941 25112 17224 25140
rect 17218 25100 17224 25112
rect 17276 25100 17282 25152
rect 17770 25140 17776 25152
rect 17683 25112 17776 25140
rect 17770 25100 17776 25112
rect 17828 25140 17834 25152
rect 19242 25140 19248 25152
rect 17828 25112 19248 25140
rect 17828 25100 17834 25112
rect 19242 25100 19248 25112
rect 19300 25100 19306 25152
rect 19429 25143 19487 25149
rect 19429 25109 19441 25143
rect 19475 25140 19487 25143
rect 19886 25140 19892 25152
rect 19475 25112 19892 25140
rect 19475 25109 19487 25112
rect 19429 25103 19487 25109
rect 19886 25100 19892 25112
rect 19944 25100 19950 25152
rect 22005 25143 22063 25149
rect 22005 25109 22017 25143
rect 22051 25140 22063 25143
rect 22646 25140 22652 25152
rect 22051 25112 22652 25140
rect 22051 25109 22063 25112
rect 22005 25103 22063 25109
rect 22646 25100 22652 25112
rect 22704 25100 22710 25152
rect 23474 25100 23480 25152
rect 23532 25140 23538 25152
rect 23584 25140 23612 25239
rect 23676 25220 23704 25248
rect 23753 25245 23765 25248
rect 23799 25245 23811 25279
rect 23753 25239 23811 25245
rect 24949 25279 25007 25285
rect 24949 25245 24961 25279
rect 24995 25245 25007 25279
rect 24949 25239 25007 25245
rect 25041 25279 25099 25285
rect 25041 25245 25053 25279
rect 25087 25245 25099 25279
rect 25041 25239 25099 25245
rect 25133 25279 25191 25285
rect 25133 25245 25145 25279
rect 25179 25276 25191 25279
rect 25222 25276 25228 25288
rect 25179 25248 25228 25276
rect 25179 25245 25191 25248
rect 25133 25239 25191 25245
rect 23658 25168 23664 25220
rect 23716 25168 23722 25220
rect 23532 25112 23612 25140
rect 23532 25100 23538 25112
rect 24854 25100 24860 25152
rect 24912 25140 24918 25152
rect 24964 25140 24992 25239
rect 25056 25208 25084 25239
rect 25222 25236 25228 25248
rect 25280 25236 25286 25288
rect 25314 25236 25320 25288
rect 25372 25276 25378 25288
rect 26326 25276 26332 25288
rect 25372 25248 25417 25276
rect 26287 25248 26332 25276
rect 25372 25236 25378 25248
rect 26326 25236 26332 25248
rect 26384 25236 26390 25288
rect 25498 25208 25504 25220
rect 25056 25180 25504 25208
rect 25498 25168 25504 25180
rect 25556 25168 25562 25220
rect 26510 25208 26516 25220
rect 26471 25180 26516 25208
rect 26510 25168 26516 25180
rect 26568 25168 26574 25220
rect 24912 25112 24992 25140
rect 24912 25100 24918 25112
rect 1104 25050 28888 25072
rect 1104 24998 10214 25050
rect 10266 24998 10278 25050
rect 10330 24998 10342 25050
rect 10394 24998 10406 25050
rect 10458 24998 10470 25050
rect 10522 24998 19478 25050
rect 19530 24998 19542 25050
rect 19594 24998 19606 25050
rect 19658 24998 19670 25050
rect 19722 24998 19734 25050
rect 19786 24998 28888 25050
rect 1104 24976 28888 24998
rect 11606 24896 11612 24948
rect 11664 24936 11670 24948
rect 12066 24936 12072 24948
rect 11664 24908 12072 24936
rect 11664 24896 11670 24908
rect 12066 24896 12072 24908
rect 12124 24896 12130 24948
rect 12986 24896 12992 24948
rect 13044 24936 13050 24948
rect 13081 24939 13139 24945
rect 13081 24936 13093 24939
rect 13044 24908 13093 24936
rect 13044 24896 13050 24908
rect 13081 24905 13093 24908
rect 13127 24905 13139 24939
rect 13722 24936 13728 24948
rect 13683 24908 13728 24936
rect 13081 24899 13139 24905
rect 13722 24896 13728 24908
rect 13780 24896 13786 24948
rect 14182 24896 14188 24948
rect 14240 24936 14246 24948
rect 14550 24936 14556 24948
rect 14240 24908 14556 24936
rect 14240 24896 14246 24908
rect 14550 24896 14556 24908
rect 14608 24896 14614 24948
rect 14734 24896 14740 24948
rect 14792 24936 14798 24948
rect 15010 24936 15016 24948
rect 14792 24908 15016 24936
rect 14792 24896 14798 24908
rect 15010 24896 15016 24908
rect 15068 24896 15074 24948
rect 15746 24936 15752 24948
rect 15120 24908 15752 24936
rect 10594 24828 10600 24880
rect 10652 24868 10658 24880
rect 13998 24868 14004 24880
rect 10652 24840 14004 24868
rect 10652 24828 10658 24840
rect 13998 24828 14004 24840
rect 14056 24828 14062 24880
rect 14369 24871 14427 24877
rect 14369 24837 14381 24871
rect 14415 24868 14427 24871
rect 15120 24868 15148 24908
rect 15746 24896 15752 24908
rect 15804 24896 15810 24948
rect 15930 24896 15936 24948
rect 15988 24936 15994 24948
rect 17037 24939 17095 24945
rect 17037 24936 17049 24939
rect 15988 24908 17049 24936
rect 15988 24896 15994 24908
rect 17037 24905 17049 24908
rect 17083 24905 17095 24939
rect 17037 24899 17095 24905
rect 17126 24896 17132 24948
rect 17184 24936 17190 24948
rect 22094 24936 22100 24948
rect 17184 24908 22100 24936
rect 17184 24896 17190 24908
rect 22094 24896 22100 24908
rect 22152 24896 22158 24948
rect 22278 24896 22284 24948
rect 22336 24936 22342 24948
rect 26329 24939 26387 24945
rect 26329 24936 26341 24939
rect 22336 24908 26341 24936
rect 22336 24896 22342 24908
rect 16022 24868 16028 24880
rect 14415 24840 15148 24868
rect 15212 24840 16028 24868
rect 14415 24837 14427 24840
rect 14369 24831 14427 24837
rect 10318 24800 10324 24812
rect 10279 24772 10324 24800
rect 10318 24760 10324 24772
rect 10376 24760 10382 24812
rect 10781 24803 10839 24809
rect 10781 24769 10793 24803
rect 10827 24769 10839 24803
rect 10781 24763 10839 24769
rect 10965 24803 11023 24809
rect 10965 24769 10977 24803
rect 11011 24800 11023 24803
rect 11011 24772 12020 24800
rect 11011 24769 11023 24772
rect 10965 24763 11023 24769
rect 10796 24732 10824 24763
rect 11422 24732 11428 24744
rect 10796 24704 11428 24732
rect 11422 24692 11428 24704
rect 11480 24692 11486 24744
rect 11882 24732 11888 24744
rect 11843 24704 11888 24732
rect 11882 24692 11888 24704
rect 11940 24692 11946 24744
rect 10137 24667 10195 24673
rect 10137 24633 10149 24667
rect 10183 24664 10195 24667
rect 11330 24664 11336 24676
rect 10183 24636 11336 24664
rect 10183 24633 10195 24636
rect 10137 24627 10195 24633
rect 11330 24624 11336 24636
rect 11388 24624 11394 24676
rect 11992 24664 12020 24772
rect 12066 24760 12072 24812
rect 12124 24800 12130 24812
rect 12897 24803 12955 24809
rect 12897 24800 12909 24803
rect 12124 24772 12909 24800
rect 12124 24760 12130 24772
rect 12897 24769 12909 24772
rect 12943 24769 12955 24803
rect 12897 24763 12955 24769
rect 13633 24803 13691 24809
rect 13633 24769 13645 24803
rect 13679 24769 13691 24803
rect 13633 24763 13691 24769
rect 12710 24732 12716 24744
rect 12671 24704 12716 24732
rect 12710 24692 12716 24704
rect 12768 24692 12774 24744
rect 12802 24692 12808 24744
rect 12860 24732 12866 24744
rect 13639 24732 13667 24763
rect 13906 24760 13912 24812
rect 13964 24800 13970 24812
rect 15212 24809 15240 24840
rect 16022 24828 16028 24840
rect 16080 24828 16086 24880
rect 16114 24828 16120 24880
rect 16172 24868 16178 24880
rect 19429 24871 19487 24877
rect 19429 24868 19441 24871
rect 16172 24840 19441 24868
rect 16172 24828 16178 24840
rect 19429 24837 19441 24840
rect 19475 24837 19487 24871
rect 22557 24871 22615 24877
rect 22557 24868 22569 24871
rect 19429 24831 19487 24837
rect 21008 24840 22569 24868
rect 15013 24803 15071 24809
rect 15013 24800 15025 24803
rect 13964 24772 15025 24800
rect 13964 24760 13970 24772
rect 15013 24769 15025 24772
rect 15059 24769 15071 24803
rect 15013 24763 15071 24769
rect 15197 24803 15255 24809
rect 15197 24769 15209 24803
rect 15243 24769 15255 24803
rect 15197 24763 15255 24769
rect 15289 24803 15347 24809
rect 15289 24769 15301 24803
rect 15335 24769 15347 24803
rect 15289 24763 15347 24769
rect 12860 24704 13667 24732
rect 12860 24692 12866 24704
rect 14274 24692 14280 24744
rect 14332 24732 14338 24744
rect 14826 24732 14832 24744
rect 14332 24704 14832 24732
rect 14332 24692 14338 24704
rect 14826 24692 14832 24704
rect 14884 24732 14890 24744
rect 15304 24732 15332 24763
rect 15378 24760 15384 24812
rect 15436 24800 15442 24812
rect 15565 24803 15623 24809
rect 15565 24800 15577 24803
rect 15436 24772 15577 24800
rect 15436 24760 15442 24772
rect 15565 24769 15577 24772
rect 15611 24800 15623 24803
rect 15930 24800 15936 24812
rect 15611 24772 15936 24800
rect 15611 24769 15623 24772
rect 15565 24763 15623 24769
rect 15930 24760 15936 24772
rect 15988 24760 15994 24812
rect 16850 24800 16856 24812
rect 16811 24772 16856 24800
rect 16850 24760 16856 24772
rect 16908 24760 16914 24812
rect 17129 24803 17187 24809
rect 17129 24769 17141 24803
rect 17175 24769 17187 24803
rect 17129 24763 17187 24769
rect 17144 24732 17172 24763
rect 17402 24760 17408 24812
rect 17460 24800 17466 24812
rect 17589 24803 17647 24809
rect 17589 24800 17601 24803
rect 17460 24772 17601 24800
rect 17460 24760 17466 24772
rect 17589 24769 17601 24772
rect 17635 24769 17647 24803
rect 18230 24800 18236 24812
rect 18191 24772 18236 24800
rect 17589 24763 17647 24769
rect 18230 24760 18236 24772
rect 18288 24760 18294 24812
rect 18414 24800 18420 24812
rect 18375 24772 18420 24800
rect 18414 24760 18420 24772
rect 18472 24800 18478 24812
rect 19245 24803 19303 24809
rect 19245 24800 19257 24803
rect 18472 24772 19257 24800
rect 18472 24760 18478 24772
rect 19245 24769 19257 24772
rect 19291 24769 19303 24803
rect 19245 24763 19303 24769
rect 19334 24760 19340 24812
rect 19392 24800 19398 24812
rect 20441 24803 20499 24809
rect 20441 24800 20453 24803
rect 19392 24772 20453 24800
rect 19392 24760 19398 24772
rect 20441 24769 20453 24772
rect 20487 24769 20499 24803
rect 20622 24800 20628 24812
rect 20583 24772 20628 24800
rect 20441 24763 20499 24769
rect 20622 24760 20628 24772
rect 20680 24760 20686 24812
rect 20806 24760 20812 24812
rect 20864 24760 20870 24812
rect 14884 24704 17172 24732
rect 14884 24692 14890 24704
rect 18046 24692 18052 24744
rect 18104 24732 18110 24744
rect 19061 24735 19119 24741
rect 19061 24732 19073 24735
rect 18104 24704 19073 24732
rect 18104 24692 18110 24704
rect 19061 24701 19073 24704
rect 19107 24701 19119 24735
rect 19061 24695 19119 24701
rect 20257 24735 20315 24741
rect 20257 24701 20269 24735
rect 20303 24732 20315 24735
rect 20824 24732 20852 24760
rect 20303 24704 20852 24732
rect 21008 24732 21036 24840
rect 22557 24837 22569 24840
rect 22603 24837 22615 24871
rect 22557 24831 22615 24837
rect 23661 24871 23719 24877
rect 23661 24837 23673 24871
rect 23707 24868 23719 24871
rect 25222 24868 25228 24880
rect 23707 24840 25228 24868
rect 23707 24837 23719 24840
rect 23661 24831 23719 24837
rect 25222 24828 25228 24840
rect 25280 24828 25286 24880
rect 21085 24803 21143 24809
rect 21085 24769 21097 24803
rect 21131 24800 21143 24803
rect 21358 24800 21364 24812
rect 21131 24772 21364 24800
rect 21131 24769 21143 24772
rect 21085 24763 21143 24769
rect 21358 24760 21364 24772
rect 21416 24760 21422 24812
rect 22370 24800 22376 24812
rect 22331 24772 22376 24800
rect 22370 24760 22376 24772
rect 22428 24760 22434 24812
rect 22646 24760 22652 24812
rect 22704 24800 22710 24812
rect 22704 24772 22749 24800
rect 22704 24760 22710 24772
rect 22830 24760 22836 24812
rect 22888 24800 22894 24812
rect 23845 24803 23903 24809
rect 23845 24800 23857 24803
rect 22888 24772 23857 24800
rect 22888 24760 22894 24772
rect 23845 24769 23857 24772
rect 23891 24769 23903 24803
rect 23845 24763 23903 24769
rect 23934 24760 23940 24812
rect 23992 24800 23998 24812
rect 25133 24803 25191 24809
rect 23992 24772 24992 24800
rect 23992 24760 23998 24772
rect 21177 24735 21235 24741
rect 21008 24704 21128 24732
rect 20303 24701 20315 24704
rect 20257 24695 20315 24701
rect 21100 24676 21128 24704
rect 21177 24701 21189 24735
rect 21223 24732 21235 24735
rect 21634 24732 21640 24744
rect 21223 24704 21640 24732
rect 21223 24701 21235 24704
rect 21177 24695 21235 24701
rect 21634 24692 21640 24704
rect 21692 24692 21698 24744
rect 23658 24692 23664 24744
rect 23716 24732 23722 24744
rect 24118 24732 24124 24744
rect 23716 24704 23796 24732
rect 24079 24704 24124 24732
rect 23716 24692 23722 24704
rect 13262 24664 13268 24676
rect 11992 24636 13268 24664
rect 13262 24624 13268 24636
rect 13320 24624 13326 24676
rect 16758 24664 16764 24676
rect 14384 24636 16764 24664
rect 10781 24599 10839 24605
rect 10781 24565 10793 24599
rect 10827 24596 10839 24599
rect 10870 24596 10876 24608
rect 10827 24568 10876 24596
rect 10827 24565 10839 24568
rect 10781 24559 10839 24565
rect 10870 24556 10876 24568
rect 10928 24556 10934 24608
rect 11790 24556 11796 24608
rect 11848 24596 11854 24608
rect 12253 24599 12311 24605
rect 12253 24596 12265 24599
rect 11848 24568 12265 24596
rect 11848 24556 11854 24568
rect 12253 24565 12265 24568
rect 12299 24565 12311 24599
rect 12253 24559 12311 24565
rect 12434 24556 12440 24608
rect 12492 24596 12498 24608
rect 14384 24596 14412 24636
rect 16758 24624 16764 24636
rect 16816 24624 16822 24676
rect 17681 24667 17739 24673
rect 17681 24633 17693 24667
rect 17727 24664 17739 24667
rect 20806 24664 20812 24676
rect 17727 24636 20812 24664
rect 17727 24633 17739 24636
rect 17681 24627 17739 24633
rect 20806 24624 20812 24636
rect 20864 24624 20870 24676
rect 21082 24624 21088 24676
rect 21140 24624 21146 24676
rect 22186 24664 22192 24676
rect 22147 24636 22192 24664
rect 22186 24624 22192 24636
rect 22244 24624 22250 24676
rect 12492 24568 14412 24596
rect 12492 24556 12498 24568
rect 14458 24556 14464 24608
rect 14516 24596 14522 24608
rect 15473 24599 15531 24605
rect 14516 24568 14561 24596
rect 14516 24556 14522 24568
rect 15473 24565 15485 24599
rect 15519 24596 15531 24599
rect 15654 24596 15660 24608
rect 15519 24568 15660 24596
rect 15519 24565 15531 24568
rect 15473 24559 15531 24565
rect 15654 24556 15660 24568
rect 15712 24556 15718 24608
rect 15746 24556 15752 24608
rect 15804 24596 15810 24608
rect 16114 24596 16120 24608
rect 15804 24568 16120 24596
rect 15804 24556 15810 24568
rect 16114 24556 16120 24568
rect 16172 24556 16178 24608
rect 16482 24556 16488 24608
rect 16540 24596 16546 24608
rect 16669 24599 16727 24605
rect 16669 24596 16681 24599
rect 16540 24568 16681 24596
rect 16540 24556 16546 24568
rect 16669 24565 16681 24568
rect 16715 24565 16727 24599
rect 16669 24559 16727 24565
rect 17034 24556 17040 24608
rect 17092 24596 17098 24608
rect 18601 24599 18659 24605
rect 18601 24596 18613 24599
rect 17092 24568 18613 24596
rect 17092 24556 17098 24568
rect 18601 24565 18613 24568
rect 18647 24565 18659 24599
rect 18601 24559 18659 24565
rect 18690 24556 18696 24608
rect 18748 24596 18754 24608
rect 23198 24596 23204 24608
rect 18748 24568 23204 24596
rect 18748 24556 18754 24568
rect 23198 24556 23204 24568
rect 23256 24556 23262 24608
rect 23768 24596 23796 24704
rect 24118 24692 24124 24704
rect 24176 24692 24182 24744
rect 24964 24732 24992 24772
rect 25133 24769 25145 24803
rect 25179 24800 25191 24803
rect 25323 24800 25351 24908
rect 26329 24905 26341 24908
rect 26375 24905 26387 24939
rect 26329 24899 26387 24905
rect 26050 24828 26056 24880
rect 26108 24868 26114 24880
rect 26108 24840 26556 24868
rect 26108 24828 26114 24840
rect 26142 24800 26148 24812
rect 25179 24772 25351 24800
rect 26103 24772 26148 24800
rect 25179 24769 25191 24772
rect 25133 24763 25191 24769
rect 26142 24760 26148 24772
rect 26200 24760 26206 24812
rect 26421 24803 26479 24809
rect 26421 24769 26433 24803
rect 26467 24769 26479 24803
rect 26421 24763 26479 24769
rect 25041 24735 25099 24741
rect 25041 24732 25053 24735
rect 24964 24704 25053 24732
rect 25041 24701 25053 24704
rect 25087 24701 25099 24735
rect 25498 24732 25504 24744
rect 25459 24704 25504 24732
rect 25041 24695 25099 24701
rect 25056 24664 25084 24695
rect 25498 24692 25504 24704
rect 25556 24692 25562 24744
rect 26436 24664 26464 24763
rect 26528 24732 26556 24840
rect 26896 24840 27292 24868
rect 26602 24760 26608 24812
rect 26660 24800 26666 24812
rect 26896 24800 26924 24840
rect 26660 24772 26924 24800
rect 26660 24760 26666 24772
rect 26970 24760 26976 24812
rect 27028 24800 27034 24812
rect 27157 24803 27215 24809
rect 27157 24800 27169 24803
rect 27028 24772 27169 24800
rect 27028 24760 27034 24772
rect 27157 24769 27169 24772
rect 27203 24769 27215 24803
rect 27264 24800 27292 24840
rect 27985 24803 28043 24809
rect 27985 24800 27997 24803
rect 27264 24772 27997 24800
rect 27157 24763 27215 24769
rect 27985 24769 27997 24772
rect 28031 24800 28043 24803
rect 28534 24800 28540 24812
rect 28031 24772 28540 24800
rect 28031 24769 28043 24772
rect 27985 24763 28043 24769
rect 28534 24760 28540 24772
rect 28592 24760 28598 24812
rect 27065 24735 27123 24741
rect 27065 24732 27077 24735
rect 26528 24704 27077 24732
rect 27065 24701 27077 24704
rect 27111 24701 27123 24735
rect 27065 24695 27123 24701
rect 25056 24636 26464 24664
rect 26510 24624 26516 24676
rect 26568 24664 26574 24676
rect 28077 24667 28135 24673
rect 28077 24664 28089 24667
rect 26568 24636 28089 24664
rect 26568 24624 26574 24636
rect 28077 24633 28089 24636
rect 28123 24633 28135 24667
rect 28077 24627 28135 24633
rect 24029 24599 24087 24605
rect 24029 24596 24041 24599
rect 23768 24568 24041 24596
rect 24029 24565 24041 24568
rect 24075 24565 24087 24599
rect 24029 24559 24087 24565
rect 24670 24556 24676 24608
rect 24728 24596 24734 24608
rect 25590 24596 25596 24608
rect 24728 24568 25596 24596
rect 24728 24556 24734 24568
rect 25590 24556 25596 24568
rect 25648 24556 25654 24608
rect 25961 24599 26019 24605
rect 25961 24565 25973 24599
rect 26007 24596 26019 24599
rect 27154 24596 27160 24608
rect 26007 24568 27160 24596
rect 26007 24565 26019 24568
rect 25961 24559 26019 24565
rect 27154 24556 27160 24568
rect 27212 24556 27218 24608
rect 27246 24556 27252 24608
rect 27304 24596 27310 24608
rect 27525 24599 27583 24605
rect 27525 24596 27537 24599
rect 27304 24568 27537 24596
rect 27304 24556 27310 24568
rect 27525 24565 27537 24568
rect 27571 24565 27583 24599
rect 27525 24559 27583 24565
rect 1104 24506 28888 24528
rect 1104 24454 5582 24506
rect 5634 24454 5646 24506
rect 5698 24454 5710 24506
rect 5762 24454 5774 24506
rect 5826 24454 5838 24506
rect 5890 24454 14846 24506
rect 14898 24454 14910 24506
rect 14962 24454 14974 24506
rect 15026 24454 15038 24506
rect 15090 24454 15102 24506
rect 15154 24454 24110 24506
rect 24162 24454 24174 24506
rect 24226 24454 24238 24506
rect 24290 24454 24302 24506
rect 24354 24454 24366 24506
rect 24418 24454 28888 24506
rect 1104 24432 28888 24454
rect 10318 24352 10324 24404
rect 10376 24392 10382 24404
rect 10962 24392 10968 24404
rect 10376 24364 10968 24392
rect 10376 24352 10382 24364
rect 10962 24352 10968 24364
rect 11020 24352 11026 24404
rect 11238 24352 11244 24404
rect 11296 24392 11302 24404
rect 11790 24392 11796 24404
rect 11296 24364 11796 24392
rect 11296 24352 11302 24364
rect 11790 24352 11796 24364
rect 11848 24352 11854 24404
rect 12158 24392 12164 24404
rect 11992 24364 12164 24392
rect 11425 24327 11483 24333
rect 11425 24293 11437 24327
rect 11471 24324 11483 24327
rect 11992 24324 12020 24364
rect 12158 24352 12164 24364
rect 12216 24352 12222 24404
rect 12618 24392 12624 24404
rect 12579 24364 12624 24392
rect 12618 24352 12624 24364
rect 12676 24352 12682 24404
rect 14734 24392 14740 24404
rect 12912 24364 14740 24392
rect 11471 24296 12020 24324
rect 11471 24293 11483 24296
rect 11425 24287 11483 24293
rect 12066 24284 12072 24336
rect 12124 24324 12130 24336
rect 12124 24296 12169 24324
rect 12124 24284 12130 24296
rect 12912 24256 12940 24364
rect 14734 24352 14740 24364
rect 14792 24352 14798 24404
rect 16390 24392 16396 24404
rect 14844 24364 15969 24392
rect 13722 24284 13728 24336
rect 13780 24324 13786 24336
rect 14844 24324 14872 24364
rect 15838 24324 15844 24336
rect 13780 24296 14872 24324
rect 14936 24296 15844 24324
rect 13780 24284 13786 24296
rect 11532 24228 12940 24256
rect 10229 24191 10287 24197
rect 10229 24157 10241 24191
rect 10275 24188 10287 24191
rect 10594 24188 10600 24200
rect 10275 24160 10600 24188
rect 10275 24157 10287 24160
rect 10229 24151 10287 24157
rect 10594 24148 10600 24160
rect 10652 24148 10658 24200
rect 10686 24148 10692 24200
rect 10744 24188 10750 24200
rect 10870 24188 10876 24200
rect 10744 24160 10789 24188
rect 10831 24160 10876 24188
rect 10744 24148 10750 24160
rect 10870 24148 10876 24160
rect 10928 24148 10934 24200
rect 11333 24191 11391 24197
rect 11333 24157 11345 24191
rect 11379 24188 11391 24191
rect 11422 24188 11428 24200
rect 11379 24160 11428 24188
rect 11379 24157 11391 24160
rect 11333 24151 11391 24157
rect 11422 24148 11428 24160
rect 11480 24148 11486 24200
rect 11532 24197 11560 24228
rect 12986 24216 12992 24268
rect 13044 24256 13050 24268
rect 13357 24264 13415 24265
rect 13188 24259 13415 24264
rect 13188 24256 13369 24259
rect 13044 24236 13369 24256
rect 13044 24228 13216 24236
rect 13044 24216 13050 24228
rect 13357 24225 13369 24236
rect 13403 24225 13415 24259
rect 13357 24219 13415 24225
rect 13538 24216 13544 24268
rect 13596 24256 13602 24268
rect 13596 24228 13641 24256
rect 13596 24216 13602 24228
rect 11517 24191 11575 24197
rect 11517 24157 11529 24191
rect 11563 24157 11575 24191
rect 11974 24188 11980 24200
rect 11935 24160 11980 24188
rect 11517 24151 11575 24157
rect 11974 24148 11980 24160
rect 12032 24148 12038 24200
rect 12161 24191 12219 24197
rect 12161 24157 12173 24191
rect 12207 24188 12219 24191
rect 12805 24191 12863 24197
rect 12207 24160 12756 24188
rect 12207 24157 12219 24160
rect 12161 24151 12219 24157
rect 10781 24123 10839 24129
rect 10781 24089 10793 24123
rect 10827 24120 10839 24123
rect 12434 24120 12440 24132
rect 10827 24092 12440 24120
rect 10827 24089 10839 24092
rect 10781 24083 10839 24089
rect 12434 24080 12440 24092
rect 12492 24080 12498 24132
rect 12728 24120 12756 24160
rect 12805 24157 12817 24191
rect 12851 24188 12863 24191
rect 12894 24188 12900 24200
rect 12851 24160 12900 24188
rect 12851 24157 12863 24160
rect 12805 24151 12863 24157
rect 12894 24148 12900 24160
rect 12952 24148 12958 24200
rect 13265 24191 13323 24197
rect 13265 24157 13277 24191
rect 13311 24188 13323 24191
rect 14461 24191 14519 24197
rect 13311 24160 14412 24188
rect 13311 24157 13323 24160
rect 13265 24151 13323 24157
rect 14384 24120 14412 24160
rect 14461 24157 14473 24191
rect 14507 24188 14519 24191
rect 14936 24188 14964 24296
rect 15838 24284 15844 24296
rect 15896 24284 15902 24336
rect 15105 24259 15163 24265
rect 15105 24225 15117 24259
rect 15151 24256 15163 24259
rect 15488 24256 15700 24264
rect 15151 24236 15909 24256
rect 15151 24228 15516 24236
rect 15672 24228 15909 24236
rect 15151 24225 15163 24228
rect 15105 24219 15163 24225
rect 14507 24160 14964 24188
rect 14507 24157 14519 24160
rect 14461 24151 14519 24157
rect 15010 24148 15016 24200
rect 15068 24188 15074 24200
rect 15286 24188 15292 24200
rect 15068 24160 15292 24188
rect 15068 24148 15074 24160
rect 15286 24148 15292 24160
rect 15344 24148 15350 24200
rect 15450 24148 15456 24200
rect 15508 24190 15514 24200
rect 15565 24191 15623 24197
rect 15565 24190 15577 24191
rect 15508 24162 15577 24190
rect 15508 24160 15516 24162
rect 15508 24148 15514 24160
rect 15565 24157 15577 24162
rect 15611 24157 15623 24191
rect 15565 24151 15623 24157
rect 15881 24120 15909 24228
rect 15941 24188 15969 24364
rect 16040 24364 16396 24392
rect 16040 24265 16068 24364
rect 16390 24352 16396 24364
rect 16448 24352 16454 24404
rect 16758 24352 16764 24404
rect 16816 24392 16822 24404
rect 22278 24392 22284 24404
rect 16816 24364 22284 24392
rect 16816 24352 16822 24364
rect 22278 24352 22284 24364
rect 22336 24352 22342 24404
rect 22554 24392 22560 24404
rect 22515 24364 22560 24392
rect 22554 24352 22560 24364
rect 22612 24352 22618 24404
rect 25222 24352 25228 24404
rect 25280 24352 25286 24404
rect 17218 24284 17224 24336
rect 17276 24324 17282 24336
rect 17405 24327 17463 24333
rect 17405 24324 17417 24327
rect 17276 24296 17417 24324
rect 17276 24284 17282 24296
rect 17405 24293 17417 24296
rect 17451 24293 17463 24327
rect 17405 24287 17463 24293
rect 17494 24284 17500 24336
rect 17552 24324 17558 24336
rect 18690 24324 18696 24336
rect 17552 24296 18696 24324
rect 17552 24284 17558 24296
rect 18690 24284 18696 24296
rect 18748 24284 18754 24336
rect 20254 24284 20260 24336
rect 20312 24324 20318 24336
rect 20625 24327 20683 24333
rect 20625 24324 20637 24327
rect 20312 24296 20637 24324
rect 20312 24284 20318 24296
rect 20625 24293 20637 24296
rect 20671 24293 20683 24327
rect 20625 24287 20683 24293
rect 16025 24259 16083 24265
rect 16025 24225 16037 24259
rect 16071 24225 16083 24259
rect 16025 24219 16083 24225
rect 17926 24228 18552 24256
rect 17926 24188 17954 24228
rect 15941 24160 17954 24188
rect 18138 24148 18144 24200
rect 18196 24188 18202 24200
rect 18524 24197 18552 24228
rect 22278 24216 22284 24268
rect 22336 24256 22342 24268
rect 22830 24256 22836 24268
rect 22336 24228 22836 24256
rect 22336 24216 22342 24228
rect 22830 24216 22836 24228
rect 22888 24256 22894 24268
rect 23109 24259 23167 24265
rect 23109 24256 23121 24259
rect 22888 24228 23121 24256
rect 22888 24216 22894 24228
rect 23109 24225 23121 24228
rect 23155 24225 23167 24259
rect 23109 24219 23167 24225
rect 23382 24216 23388 24268
rect 23440 24256 23446 24268
rect 23569 24259 23627 24265
rect 23569 24256 23581 24259
rect 23440 24228 23581 24256
rect 23440 24216 23446 24228
rect 23569 24225 23581 24228
rect 23615 24225 23627 24259
rect 23569 24219 23627 24225
rect 18325 24191 18383 24197
rect 18325 24188 18337 24191
rect 18196 24160 18337 24188
rect 18196 24148 18202 24160
rect 18325 24157 18337 24160
rect 18371 24157 18383 24191
rect 18325 24151 18383 24157
rect 18414 24191 18472 24197
rect 18414 24157 18426 24191
rect 18460 24157 18472 24191
rect 18414 24151 18472 24157
rect 18509 24191 18567 24197
rect 18509 24157 18521 24191
rect 18555 24157 18567 24191
rect 18509 24151 18567 24157
rect 16022 24120 16028 24132
rect 12728 24092 14320 24120
rect 14384 24092 14964 24120
rect 13541 24055 13599 24061
rect 13541 24021 13553 24055
rect 13587 24052 13599 24055
rect 13722 24052 13728 24064
rect 13587 24024 13728 24052
rect 13587 24021 13599 24024
rect 13541 24015 13599 24021
rect 13722 24012 13728 24024
rect 13780 24012 13786 24064
rect 14292 24052 14320 24092
rect 14366 24052 14372 24064
rect 14292 24024 14372 24052
rect 14366 24012 14372 24024
rect 14424 24012 14430 24064
rect 14550 24052 14556 24064
rect 14511 24024 14556 24052
rect 14550 24012 14556 24024
rect 14608 24012 14614 24064
rect 14936 24052 14964 24092
rect 15405 24092 15655 24120
rect 15881 24092 16028 24120
rect 15405 24052 15433 24092
rect 14936 24024 15433 24052
rect 15470 24012 15476 24064
rect 15528 24052 15534 24064
rect 15627 24052 15655 24092
rect 16022 24080 16028 24092
rect 16080 24080 16086 24132
rect 16114 24080 16120 24132
rect 16172 24120 16178 24132
rect 16270 24123 16328 24129
rect 16270 24120 16282 24123
rect 16172 24092 16282 24120
rect 16172 24080 16178 24092
rect 16270 24089 16282 24092
rect 16316 24089 16328 24123
rect 16270 24083 16328 24089
rect 18049 24123 18107 24129
rect 18049 24089 18061 24123
rect 18095 24120 18107 24123
rect 18230 24120 18236 24132
rect 18095 24092 18236 24120
rect 18095 24089 18107 24092
rect 18049 24083 18107 24089
rect 18230 24080 18236 24092
rect 18288 24080 18294 24132
rect 18432 24120 18460 24151
rect 18690 24148 18696 24200
rect 18748 24188 18754 24200
rect 18966 24188 18972 24200
rect 18748 24160 18972 24188
rect 18748 24148 18754 24160
rect 18966 24148 18972 24160
rect 19024 24148 19030 24200
rect 19150 24148 19156 24200
rect 19208 24188 19214 24200
rect 19245 24191 19303 24197
rect 19245 24188 19257 24191
rect 19208 24160 19257 24188
rect 19208 24148 19214 24160
rect 19245 24157 19257 24160
rect 19291 24188 19303 24191
rect 21177 24191 21235 24197
rect 21177 24188 21189 24191
rect 19291 24160 21189 24188
rect 19291 24157 19303 24160
rect 19245 24151 19303 24157
rect 21177 24157 21189 24160
rect 21223 24157 21235 24191
rect 22646 24188 22652 24200
rect 21177 24151 21235 24157
rect 21376 24160 22652 24188
rect 18598 24120 18604 24132
rect 18432 24092 18604 24120
rect 18598 24080 18604 24092
rect 18656 24080 18662 24132
rect 18782 24080 18788 24132
rect 18840 24120 18846 24132
rect 19490 24123 19548 24129
rect 19490 24120 19502 24123
rect 18840 24092 19502 24120
rect 18840 24080 18846 24092
rect 19490 24089 19502 24092
rect 19536 24089 19548 24123
rect 21376 24120 21404 24160
rect 22646 24148 22652 24160
rect 22704 24148 22710 24200
rect 23014 24148 23020 24200
rect 23072 24188 23078 24200
rect 23201 24191 23259 24197
rect 23201 24188 23213 24191
rect 23072 24160 23213 24188
rect 23072 24148 23078 24160
rect 23201 24157 23213 24160
rect 23247 24157 23259 24191
rect 23201 24151 23259 24157
rect 19490 24083 19548 24089
rect 19628 24092 21404 24120
rect 21444 24123 21502 24129
rect 19628 24052 19656 24092
rect 21444 24089 21456 24123
rect 21490 24120 21502 24123
rect 21818 24120 21824 24132
rect 21490 24092 21824 24120
rect 21490 24089 21502 24092
rect 21444 24083 21502 24089
rect 21818 24080 21824 24092
rect 21876 24080 21882 24132
rect 22462 24080 22468 24132
rect 22520 24120 22526 24132
rect 23290 24120 23296 24132
rect 22520 24092 23296 24120
rect 22520 24080 22526 24092
rect 23290 24080 23296 24092
rect 23348 24080 23354 24132
rect 23584 24120 23612 24219
rect 23842 24216 23848 24268
rect 23900 24256 23906 24268
rect 24573 24259 24631 24265
rect 24573 24256 24585 24259
rect 23900 24228 24585 24256
rect 23900 24216 23906 24228
rect 24573 24225 24585 24228
rect 24619 24225 24631 24259
rect 24573 24219 24631 24225
rect 24673 24259 24731 24265
rect 24673 24225 24685 24259
rect 24719 24225 24731 24259
rect 24673 24219 24731 24225
rect 24857 24259 24915 24265
rect 24857 24225 24869 24259
rect 24903 24256 24915 24259
rect 25240 24256 25268 24352
rect 28166 24256 28172 24268
rect 24903 24228 25268 24256
rect 28127 24228 28172 24256
rect 24903 24225 24915 24228
rect 24857 24219 24915 24225
rect 24688 24120 24716 24219
rect 28166 24216 28172 24228
rect 28224 24216 28230 24268
rect 24765 24191 24823 24197
rect 24765 24157 24777 24191
rect 24811 24188 24823 24191
rect 24946 24188 24952 24200
rect 24811 24160 24952 24188
rect 24811 24157 24823 24160
rect 24765 24151 24823 24157
rect 24946 24148 24952 24160
rect 25004 24188 25010 24200
rect 25593 24191 25651 24197
rect 25593 24188 25605 24191
rect 25004 24160 25605 24188
rect 25004 24148 25010 24160
rect 25593 24157 25605 24160
rect 25639 24157 25651 24191
rect 26326 24188 26332 24200
rect 26287 24160 26332 24188
rect 25593 24151 25651 24157
rect 26326 24148 26332 24160
rect 26384 24148 26390 24200
rect 25409 24123 25467 24129
rect 25409 24120 25421 24123
rect 23584 24092 25421 24120
rect 25409 24089 25421 24092
rect 25455 24089 25467 24123
rect 25409 24083 25467 24089
rect 26513 24123 26571 24129
rect 26513 24089 26525 24123
rect 26559 24120 26571 24123
rect 28074 24120 28080 24132
rect 26559 24092 28080 24120
rect 26559 24089 26571 24092
rect 26513 24083 26571 24089
rect 28074 24080 28080 24092
rect 28132 24080 28138 24132
rect 15528 24024 15573 24052
rect 15627 24024 19656 24052
rect 15528 24012 15534 24024
rect 21634 24012 21640 24064
rect 21692 24052 21698 24064
rect 22278 24052 22284 24064
rect 21692 24024 22284 24052
rect 21692 24012 21698 24024
rect 22278 24012 22284 24024
rect 22336 24012 22342 24064
rect 23658 24012 23664 24064
rect 23716 24052 23722 24064
rect 24397 24055 24455 24061
rect 24397 24052 24409 24055
rect 23716 24024 24409 24052
rect 23716 24012 23722 24024
rect 24397 24021 24409 24024
rect 24443 24052 24455 24055
rect 24486 24052 24492 24064
rect 24443 24024 24492 24052
rect 24443 24021 24455 24024
rect 24397 24015 24455 24021
rect 24486 24012 24492 24024
rect 24544 24012 24550 24064
rect 25774 24052 25780 24064
rect 25735 24024 25780 24052
rect 25774 24012 25780 24024
rect 25832 24012 25838 24064
rect 1104 23962 28888 23984
rect 1104 23910 10214 23962
rect 10266 23910 10278 23962
rect 10330 23910 10342 23962
rect 10394 23910 10406 23962
rect 10458 23910 10470 23962
rect 10522 23910 19478 23962
rect 19530 23910 19542 23962
rect 19594 23910 19606 23962
rect 19658 23910 19670 23962
rect 19722 23910 19734 23962
rect 19786 23910 28888 23962
rect 1104 23888 28888 23910
rect 9677 23851 9735 23857
rect 9677 23817 9689 23851
rect 9723 23848 9735 23851
rect 13630 23848 13636 23860
rect 9723 23820 13636 23848
rect 9723 23817 9735 23820
rect 9677 23811 9735 23817
rect 13630 23808 13636 23820
rect 13688 23808 13694 23860
rect 13823 23851 13881 23857
rect 13823 23817 13835 23851
rect 13869 23848 13881 23851
rect 14090 23848 14096 23860
rect 13869 23820 14096 23848
rect 13869 23817 13881 23820
rect 13823 23811 13881 23817
rect 14090 23808 14096 23820
rect 14148 23808 14154 23860
rect 14182 23808 14188 23860
rect 14240 23848 14246 23860
rect 15749 23851 15807 23857
rect 15749 23848 15761 23851
rect 14240 23820 15761 23848
rect 14240 23808 14246 23820
rect 15749 23817 15761 23820
rect 15795 23817 15807 23851
rect 15749 23811 15807 23817
rect 16022 23808 16028 23860
rect 16080 23848 16086 23860
rect 17678 23848 17684 23860
rect 16080 23820 17684 23848
rect 16080 23808 16086 23820
rect 17678 23808 17684 23820
rect 17736 23808 17742 23860
rect 18509 23851 18567 23857
rect 18509 23817 18521 23851
rect 18555 23848 18567 23851
rect 18555 23820 18736 23848
rect 18555 23817 18567 23820
rect 18509 23811 18567 23817
rect 13170 23780 13176 23792
rect 11808 23752 12940 23780
rect 13131 23752 13176 23780
rect 1486 23672 1492 23724
rect 1544 23712 1550 23724
rect 2038 23712 2044 23724
rect 1544 23684 2044 23712
rect 1544 23672 1550 23684
rect 2038 23672 2044 23684
rect 2096 23672 2102 23724
rect 9490 23712 9496 23724
rect 9451 23684 9496 23712
rect 9490 23672 9496 23684
rect 9548 23672 9554 23724
rect 9677 23715 9735 23721
rect 9677 23681 9689 23715
rect 9723 23681 9735 23715
rect 9677 23675 9735 23681
rect 10137 23715 10195 23721
rect 10137 23681 10149 23715
rect 10183 23712 10195 23715
rect 10226 23712 10232 23724
rect 10183 23684 10232 23712
rect 10183 23681 10195 23684
rect 10137 23675 10195 23681
rect 9692 23644 9720 23675
rect 10226 23672 10232 23684
rect 10284 23672 10290 23724
rect 10318 23672 10324 23724
rect 10376 23712 10382 23724
rect 10778 23712 10784 23724
rect 10376 23684 10421 23712
rect 10739 23684 10784 23712
rect 10376 23672 10382 23684
rect 10778 23672 10784 23684
rect 10836 23672 10842 23724
rect 10965 23715 11023 23721
rect 10965 23681 10977 23715
rect 11011 23712 11023 23715
rect 11330 23712 11336 23724
rect 11011 23684 11336 23712
rect 11011 23681 11023 23684
rect 10965 23675 11023 23681
rect 11330 23672 11336 23684
rect 11388 23672 11394 23724
rect 11808 23721 11836 23752
rect 11793 23715 11851 23721
rect 11793 23681 11805 23715
rect 11839 23681 11851 23715
rect 11793 23675 11851 23681
rect 11977 23715 12035 23721
rect 11977 23681 11989 23715
rect 12023 23681 12035 23715
rect 12434 23712 12440 23724
rect 12395 23684 12440 23712
rect 11977 23675 12035 23681
rect 10336 23644 10364 23672
rect 9692 23616 10364 23644
rect 11992 23644 12020 23675
rect 12434 23672 12440 23684
rect 12492 23672 12498 23724
rect 12621 23715 12679 23721
rect 12621 23681 12633 23715
rect 12667 23712 12679 23715
rect 12710 23712 12716 23724
rect 12667 23684 12716 23712
rect 12667 23681 12679 23684
rect 12621 23675 12679 23681
rect 12710 23672 12716 23684
rect 12768 23672 12774 23724
rect 12529 23647 12587 23653
rect 12529 23644 12541 23647
rect 11992 23616 12541 23644
rect 12529 23613 12541 23616
rect 12575 23613 12587 23647
rect 12912 23644 12940 23752
rect 13170 23740 13176 23752
rect 13228 23740 13234 23792
rect 16758 23780 16764 23792
rect 14016 23752 16764 23780
rect 13078 23712 13084 23724
rect 13039 23684 13084 23712
rect 13078 23672 13084 23684
rect 13136 23672 13142 23724
rect 13262 23712 13268 23724
rect 13223 23684 13268 23712
rect 13262 23672 13268 23684
rect 13320 23672 13326 23724
rect 13722 23712 13728 23724
rect 13683 23684 13728 23712
rect 13722 23672 13728 23684
rect 13780 23672 13786 23724
rect 13906 23712 13912 23724
rect 13867 23684 13912 23712
rect 13906 23672 13912 23684
rect 13964 23672 13970 23724
rect 14016 23721 14044 23752
rect 16758 23740 16764 23752
rect 16816 23740 16822 23792
rect 18598 23780 18604 23792
rect 17880 23752 18604 23780
rect 14001 23715 14059 23721
rect 14001 23681 14013 23715
rect 14047 23681 14059 23715
rect 14550 23712 14556 23724
rect 14511 23684 14556 23712
rect 14001 23675 14059 23681
rect 14550 23672 14556 23684
rect 14608 23672 14614 23724
rect 14734 23672 14740 23724
rect 14792 23712 14798 23724
rect 15194 23712 15200 23724
rect 14792 23684 15200 23712
rect 14792 23672 14798 23684
rect 15194 23672 15200 23684
rect 15252 23672 15258 23724
rect 15378 23712 15384 23724
rect 15339 23684 15384 23712
rect 15378 23672 15384 23684
rect 15436 23672 15442 23724
rect 15838 23672 15844 23724
rect 15896 23712 15902 23724
rect 17494 23712 17500 23724
rect 15896 23684 17500 23712
rect 15896 23672 15902 23684
rect 17494 23672 17500 23684
rect 17552 23672 17558 23724
rect 15010 23644 15016 23656
rect 12912 23616 15016 23644
rect 12529 23607 12587 23613
rect 15010 23604 15016 23616
rect 15068 23604 15074 23656
rect 15289 23647 15347 23653
rect 15289 23644 15301 23647
rect 15120 23616 15301 23644
rect 10781 23579 10839 23585
rect 10781 23545 10793 23579
rect 10827 23576 10839 23579
rect 15120 23576 15148 23616
rect 15289 23613 15301 23616
rect 15335 23613 15347 23647
rect 15289 23607 15347 23613
rect 15654 23604 15660 23656
rect 15712 23644 15718 23656
rect 16669 23647 16727 23653
rect 16669 23644 16681 23647
rect 15712 23616 16681 23644
rect 15712 23604 15718 23616
rect 16669 23613 16681 23616
rect 16715 23644 16727 23647
rect 16850 23644 16856 23656
rect 16715 23616 16856 23644
rect 16715 23613 16727 23616
rect 16669 23607 16727 23613
rect 16850 23604 16856 23616
rect 16908 23604 16914 23656
rect 16942 23604 16948 23656
rect 17000 23644 17006 23656
rect 17880 23644 17908 23752
rect 18598 23740 18604 23752
rect 18656 23740 18662 23792
rect 18708 23780 18736 23820
rect 18782 23808 18788 23860
rect 18840 23848 18846 23860
rect 21634 23848 21640 23860
rect 18840 23820 21640 23848
rect 18840 23808 18846 23820
rect 21634 23808 21640 23820
rect 21692 23808 21698 23860
rect 21818 23848 21824 23860
rect 21779 23820 21824 23848
rect 21818 23808 21824 23820
rect 21876 23808 21882 23860
rect 22094 23808 22100 23860
rect 22152 23808 22158 23860
rect 24302 23848 24308 23860
rect 23400 23820 24308 23848
rect 18969 23783 19027 23789
rect 18969 23780 18981 23783
rect 18708 23752 18981 23780
rect 18969 23749 18981 23752
rect 19015 23749 19027 23783
rect 18969 23743 19027 23749
rect 19058 23740 19064 23792
rect 19116 23780 19122 23792
rect 20901 23783 20959 23789
rect 20901 23780 20913 23783
rect 19116 23752 20913 23780
rect 19116 23740 19122 23752
rect 20901 23749 20913 23752
rect 20947 23749 20959 23783
rect 22112 23780 22140 23808
rect 23400 23780 23428 23820
rect 24302 23808 24308 23820
rect 24360 23808 24366 23860
rect 24489 23851 24547 23857
rect 24489 23817 24501 23851
rect 24535 23848 24547 23851
rect 24578 23848 24584 23860
rect 24535 23820 24584 23848
rect 24535 23817 24547 23820
rect 24489 23811 24547 23817
rect 24578 23808 24584 23820
rect 24636 23808 24642 23860
rect 24670 23808 24676 23860
rect 24728 23848 24734 23860
rect 26421 23851 26479 23857
rect 26421 23848 26433 23851
rect 24728 23820 26433 23848
rect 24728 23808 24734 23820
rect 26421 23817 26433 23820
rect 26467 23848 26479 23851
rect 26602 23848 26608 23860
rect 26467 23820 26608 23848
rect 26467 23817 26479 23820
rect 26421 23811 26479 23817
rect 26602 23808 26608 23820
rect 26660 23848 26666 23860
rect 26970 23848 26976 23860
rect 26660 23820 26976 23848
rect 26660 23808 26666 23820
rect 26970 23808 26976 23820
rect 27028 23808 27034 23860
rect 28074 23848 28080 23860
rect 28035 23820 28080 23848
rect 28074 23808 28080 23820
rect 28132 23808 28138 23860
rect 22112 23752 23428 23780
rect 20901 23743 20959 23749
rect 18138 23712 18144 23724
rect 18099 23684 18144 23712
rect 18138 23672 18144 23684
rect 18196 23672 18202 23724
rect 18414 23672 18420 23724
rect 18472 23712 18478 23724
rect 18616 23712 18644 23740
rect 18874 23712 18880 23724
rect 18472 23684 18555 23712
rect 18616 23684 18880 23712
rect 18472 23672 18478 23684
rect 18046 23644 18052 23656
rect 17000 23616 17908 23644
rect 18007 23616 18052 23644
rect 17000 23604 17006 23616
rect 18046 23604 18052 23616
rect 18104 23604 18110 23656
rect 10827 23548 15148 23576
rect 10827 23545 10839 23548
rect 10781 23539 10839 23545
rect 16758 23536 16764 23588
rect 16816 23576 16822 23588
rect 18322 23576 18328 23588
rect 16816 23548 18328 23576
rect 16816 23536 16822 23548
rect 18322 23536 18328 23548
rect 18380 23536 18386 23588
rect 18527 23576 18555 23684
rect 18874 23672 18880 23684
rect 18932 23712 18938 23724
rect 19153 23715 19211 23721
rect 19153 23712 19165 23715
rect 18932 23684 19165 23712
rect 18932 23672 18938 23684
rect 19153 23681 19165 23684
rect 19199 23681 19211 23715
rect 19153 23675 19211 23681
rect 19240 23684 20208 23712
rect 18598 23604 18604 23656
rect 18656 23644 18662 23656
rect 19240 23644 19268 23684
rect 18656 23616 19268 23644
rect 19337 23647 19395 23653
rect 18656 23604 18662 23616
rect 19337 23613 19349 23647
rect 19383 23644 19395 23647
rect 19886 23644 19892 23656
rect 19383 23616 19892 23644
rect 19383 23613 19395 23616
rect 19337 23607 19395 23613
rect 19886 23604 19892 23616
rect 19944 23604 19950 23656
rect 20070 23644 20076 23656
rect 20031 23616 20076 23644
rect 20070 23604 20076 23616
rect 20128 23604 20134 23656
rect 20180 23644 20208 23684
rect 20254 23672 20260 23724
rect 20312 23712 20318 23724
rect 20312 23684 20357 23712
rect 20312 23672 20318 23684
rect 20438 23672 20444 23724
rect 20496 23712 20502 23724
rect 21082 23712 21088 23724
rect 20496 23684 20541 23712
rect 21043 23684 21088 23712
rect 20496 23672 20502 23684
rect 21082 23672 21088 23684
rect 21140 23672 21146 23724
rect 21726 23672 21732 23724
rect 21784 23712 21790 23724
rect 22002 23712 22008 23724
rect 21784 23684 22008 23712
rect 21784 23672 21790 23684
rect 22002 23672 22008 23684
rect 22060 23712 22066 23724
rect 22097 23715 22155 23721
rect 22097 23712 22109 23715
rect 22060 23684 22109 23712
rect 22060 23672 22066 23684
rect 22097 23681 22109 23684
rect 22143 23681 22155 23715
rect 22097 23675 22155 23681
rect 22189 23715 22247 23721
rect 22189 23681 22201 23715
rect 22235 23681 22247 23715
rect 22189 23675 22247 23681
rect 20456 23644 20484 23672
rect 20180 23616 20484 23644
rect 22204 23644 22232 23675
rect 22278 23672 22284 23724
rect 22336 23712 22342 23724
rect 22465 23715 22523 23721
rect 22336 23684 22381 23712
rect 22336 23672 22342 23684
rect 22465 23681 22477 23715
rect 22511 23712 22523 23715
rect 22554 23712 22560 23724
rect 22511 23684 22560 23712
rect 22511 23681 22523 23684
rect 22465 23675 22523 23681
rect 22554 23672 22560 23684
rect 22612 23672 22618 23724
rect 23400 23721 23428 23752
rect 23569 23783 23627 23789
rect 23569 23749 23581 23783
rect 23615 23780 23627 23783
rect 25774 23780 25780 23792
rect 23615 23752 25780 23780
rect 23615 23749 23627 23752
rect 23569 23743 23627 23749
rect 25774 23740 25780 23752
rect 25832 23740 25838 23792
rect 23385 23715 23443 23721
rect 23385 23681 23397 23715
rect 23431 23681 23443 23715
rect 23385 23675 23443 23681
rect 23474 23672 23480 23724
rect 23532 23712 23538 23724
rect 23661 23715 23719 23721
rect 23661 23712 23673 23715
rect 23532 23684 23673 23712
rect 23532 23672 23538 23684
rect 23661 23681 23673 23684
rect 23707 23681 23719 23715
rect 24302 23712 24308 23724
rect 24263 23684 24308 23712
rect 23661 23675 23719 23681
rect 24302 23672 24308 23684
rect 24360 23672 24366 23724
rect 24581 23715 24639 23721
rect 24581 23681 24593 23715
rect 24627 23712 24639 23715
rect 24854 23712 24860 23724
rect 24627 23684 24860 23712
rect 24627 23681 24639 23684
rect 24581 23675 24639 23681
rect 24854 23672 24860 23684
rect 24912 23672 24918 23724
rect 25038 23712 25044 23724
rect 24999 23684 25044 23712
rect 25038 23672 25044 23684
rect 25096 23672 25102 23724
rect 25308 23715 25366 23721
rect 25308 23681 25320 23715
rect 25354 23712 25366 23715
rect 25590 23712 25596 23724
rect 25354 23684 25596 23712
rect 25354 23681 25366 23684
rect 25308 23675 25366 23681
rect 25590 23672 25596 23684
rect 25648 23672 25654 23724
rect 27154 23712 27160 23724
rect 27115 23684 27160 23712
rect 27154 23672 27160 23684
rect 27212 23672 27218 23724
rect 27982 23712 27988 23724
rect 27943 23684 27988 23712
rect 27982 23672 27988 23684
rect 28040 23672 28046 23724
rect 22646 23644 22652 23656
rect 22204 23616 22652 23644
rect 22646 23604 22652 23616
rect 22704 23604 22710 23656
rect 23198 23604 23204 23656
rect 23256 23644 23262 23656
rect 27246 23644 27252 23656
rect 23256 23616 25084 23644
rect 27207 23616 27252 23644
rect 23256 23604 23262 23616
rect 25056 23588 25084 23616
rect 27246 23604 27252 23616
rect 27304 23604 27310 23656
rect 19245 23579 19303 23585
rect 19245 23576 19257 23579
rect 18527 23548 19257 23576
rect 19245 23545 19257 23548
rect 19291 23545 19303 23579
rect 19245 23539 19303 23545
rect 19429 23579 19487 23585
rect 19429 23545 19441 23579
rect 19475 23576 19487 23579
rect 19475 23548 19625 23576
rect 19475 23545 19487 23548
rect 19429 23539 19487 23545
rect 19597 23520 19625 23548
rect 19702 23536 19708 23588
rect 19760 23576 19766 23588
rect 19760 23548 24707 23576
rect 19760 23536 19766 23548
rect 1946 23508 1952 23520
rect 1907 23480 1952 23508
rect 1946 23468 1952 23480
rect 2004 23468 2010 23520
rect 10229 23511 10287 23517
rect 10229 23477 10241 23511
rect 10275 23508 10287 23511
rect 11698 23508 11704 23520
rect 10275 23480 11704 23508
rect 10275 23477 10287 23480
rect 10229 23471 10287 23477
rect 11698 23468 11704 23480
rect 11756 23468 11762 23520
rect 11793 23511 11851 23517
rect 11793 23477 11805 23511
rect 11839 23508 11851 23511
rect 11974 23508 11980 23520
rect 11839 23480 11980 23508
rect 11839 23477 11851 23480
rect 11793 23471 11851 23477
rect 11974 23468 11980 23480
rect 12032 23508 12038 23520
rect 18782 23508 18788 23520
rect 12032 23480 18788 23508
rect 12032 23468 12038 23480
rect 18782 23468 18788 23480
rect 18840 23468 18846 23520
rect 19597 23480 19616 23520
rect 19610 23468 19616 23480
rect 19668 23468 19674 23520
rect 21269 23511 21327 23517
rect 21269 23477 21281 23511
rect 21315 23508 21327 23511
rect 22278 23508 22284 23520
rect 21315 23480 22284 23508
rect 21315 23477 21327 23480
rect 21269 23471 21327 23477
rect 22278 23468 22284 23480
rect 22336 23468 22342 23520
rect 23201 23511 23259 23517
rect 23201 23477 23213 23511
rect 23247 23508 23259 23511
rect 23382 23508 23388 23520
rect 23247 23480 23388 23508
rect 23247 23477 23259 23480
rect 23201 23471 23259 23477
rect 23382 23468 23388 23480
rect 23440 23468 23446 23520
rect 24121 23511 24179 23517
rect 24121 23477 24133 23511
rect 24167 23508 24179 23511
rect 24578 23508 24584 23520
rect 24167 23480 24584 23508
rect 24167 23477 24179 23480
rect 24121 23471 24179 23477
rect 24578 23468 24584 23480
rect 24636 23468 24642 23520
rect 24679 23508 24707 23548
rect 25038 23536 25044 23588
rect 25096 23536 25102 23588
rect 27433 23511 27491 23517
rect 27433 23508 27445 23511
rect 24679 23480 27445 23508
rect 27433 23477 27445 23480
rect 27479 23477 27491 23511
rect 27433 23471 27491 23477
rect 1104 23418 28888 23440
rect 1104 23366 5582 23418
rect 5634 23366 5646 23418
rect 5698 23366 5710 23418
rect 5762 23366 5774 23418
rect 5826 23366 5838 23418
rect 5890 23366 14846 23418
rect 14898 23366 14910 23418
rect 14962 23366 14974 23418
rect 15026 23366 15038 23418
rect 15090 23366 15102 23418
rect 15154 23366 24110 23418
rect 24162 23366 24174 23418
rect 24226 23366 24238 23418
rect 24290 23366 24302 23418
rect 24354 23366 24366 23418
rect 24418 23366 28888 23418
rect 1104 23344 28888 23366
rect 11330 23304 11336 23316
rect 11291 23276 11336 23304
rect 11330 23264 11336 23276
rect 11388 23264 11394 23316
rect 13354 23264 13360 23316
rect 13412 23304 13418 23316
rect 13449 23307 13507 23313
rect 13449 23304 13461 23307
rect 13412 23276 13461 23304
rect 13412 23264 13418 23276
rect 13449 23273 13461 23276
rect 13495 23304 13507 23307
rect 13630 23304 13636 23316
rect 13495 23276 13636 23304
rect 13495 23273 13507 23276
rect 13449 23267 13507 23273
rect 13630 23264 13636 23276
rect 13688 23264 13694 23316
rect 13740 23276 16692 23304
rect 9490 23196 9496 23248
rect 9548 23236 9554 23248
rect 13740 23236 13768 23276
rect 15470 23236 15476 23248
rect 9548 23208 13768 23236
rect 15431 23208 15476 23236
rect 9548 23196 9554 23208
rect 15470 23196 15476 23208
rect 15528 23196 15534 23248
rect 15838 23236 15844 23248
rect 15627 23208 15844 23236
rect 1397 23171 1455 23177
rect 1397 23137 1409 23171
rect 1443 23168 1455 23171
rect 1946 23168 1952 23180
rect 1443 23140 1952 23168
rect 1443 23137 1455 23140
rect 1397 23131 1455 23137
rect 1946 23128 1952 23140
rect 2004 23128 2010 23180
rect 2774 23128 2780 23180
rect 2832 23168 2838 23180
rect 2832 23140 2877 23168
rect 2832 23128 2838 23140
rect 11698 23128 11704 23180
rect 11756 23168 11762 23180
rect 11756 23140 13578 23168
rect 11756 23128 11762 23140
rect 10689 23103 10747 23109
rect 10689 23069 10701 23103
rect 10735 23069 10747 23103
rect 10689 23063 10747 23069
rect 10873 23103 10931 23109
rect 10873 23069 10885 23103
rect 10919 23100 10931 23103
rect 11054 23100 11060 23112
rect 10919 23072 11060 23100
rect 10919 23069 10931 23072
rect 10873 23063 10931 23069
rect 1581 23035 1639 23041
rect 1581 23001 1593 23035
rect 1627 23032 1639 23035
rect 2498 23032 2504 23044
rect 1627 23004 2504 23032
rect 1627 23001 1639 23004
rect 1581 22995 1639 23001
rect 2498 22992 2504 23004
rect 2556 22992 2562 23044
rect 10704 23032 10732 23063
rect 11054 23060 11060 23072
rect 11112 23060 11118 23112
rect 11330 23100 11336 23112
rect 11291 23072 11336 23100
rect 11330 23060 11336 23072
rect 11388 23060 11394 23112
rect 11514 23100 11520 23112
rect 11475 23072 11520 23100
rect 11514 23060 11520 23072
rect 11572 23060 11578 23112
rect 11974 23100 11980 23112
rect 11935 23072 11980 23100
rect 11974 23060 11980 23072
rect 12032 23060 12038 23112
rect 12158 23100 12164 23112
rect 12119 23072 12164 23100
rect 12158 23060 12164 23072
rect 12216 23060 12222 23112
rect 12434 23060 12440 23112
rect 12492 23100 12498 23112
rect 12621 23103 12679 23109
rect 12621 23100 12633 23103
rect 12492 23072 12633 23100
rect 12492 23060 12498 23072
rect 12621 23069 12633 23072
rect 12667 23100 12679 23103
rect 13262 23100 13268 23112
rect 12667 23072 13268 23100
rect 12667 23069 12679 23072
rect 12621 23063 12679 23069
rect 13262 23060 13268 23072
rect 13320 23060 13326 23112
rect 13357 23103 13415 23109
rect 13357 23069 13369 23103
rect 13403 23100 13415 23103
rect 13446 23100 13452 23112
rect 13403 23072 13452 23100
rect 13403 23069 13415 23072
rect 13357 23063 13415 23069
rect 13446 23060 13452 23072
rect 13504 23060 13510 23112
rect 13550 23100 13578 23140
rect 13814 23128 13820 23180
rect 13872 23168 13878 23180
rect 14093 23171 14151 23177
rect 14093 23168 14105 23171
rect 13872 23140 14105 23168
rect 13872 23128 13878 23140
rect 14093 23137 14105 23140
rect 14139 23137 14151 23171
rect 14093 23131 14151 23137
rect 15378 23128 15384 23180
rect 15436 23168 15442 23180
rect 15627 23168 15655 23208
rect 15838 23196 15844 23208
rect 15896 23196 15902 23248
rect 16114 23196 16120 23248
rect 16172 23236 16178 23248
rect 16664 23236 16692 23276
rect 17494 23264 17500 23316
rect 17552 23304 17558 23316
rect 17552 23276 17954 23304
rect 17552 23264 17558 23276
rect 17773 23239 17831 23245
rect 17773 23236 17785 23239
rect 16172 23208 16217 23236
rect 16664 23208 17785 23236
rect 16172 23196 16178 23208
rect 17773 23205 17785 23208
rect 17819 23205 17831 23239
rect 17926 23236 17954 23276
rect 18138 23264 18144 23316
rect 18196 23304 18202 23316
rect 18233 23307 18291 23313
rect 18233 23304 18245 23307
rect 18196 23276 18245 23304
rect 18196 23264 18202 23276
rect 18233 23273 18245 23276
rect 18279 23273 18291 23307
rect 18233 23267 18291 23273
rect 18782 23264 18788 23316
rect 18840 23304 18846 23316
rect 19058 23304 19064 23316
rect 18840 23276 19064 23304
rect 18840 23264 18846 23276
rect 19058 23264 19064 23276
rect 19116 23264 19122 23316
rect 19426 23264 19432 23316
rect 19484 23304 19490 23316
rect 20622 23304 20628 23316
rect 19484 23276 20628 23304
rect 19484 23264 19490 23276
rect 20622 23264 20628 23276
rect 20680 23264 20686 23316
rect 20714 23264 20720 23316
rect 20772 23304 20778 23316
rect 25682 23304 25688 23316
rect 20772 23276 25688 23304
rect 20772 23264 20778 23276
rect 25682 23264 25688 23276
rect 25740 23264 25746 23316
rect 18414 23236 18420 23248
rect 17926 23208 18420 23236
rect 17773 23199 17831 23205
rect 18414 23196 18420 23208
rect 18472 23196 18478 23248
rect 21913 23239 21971 23245
rect 19536 23208 20024 23236
rect 15436 23140 15655 23168
rect 15436 23128 15442 23140
rect 15746 23128 15752 23180
rect 15804 23168 15810 23180
rect 17034 23168 17040 23180
rect 15804 23140 16252 23168
rect 15804 23128 15810 23140
rect 13550 23072 14596 23100
rect 11348 23032 11376 23060
rect 10704 23004 11376 23032
rect 12069 23035 12127 23041
rect 12069 23001 12081 23035
rect 12115 23032 12127 23035
rect 14360 23035 14418 23041
rect 12115 23004 14320 23032
rect 12115 23001 12127 23004
rect 12069 22995 12127 23001
rect 10781 22967 10839 22973
rect 10781 22933 10793 22967
rect 10827 22964 10839 22967
rect 10962 22964 10968 22976
rect 10827 22936 10968 22964
rect 10827 22933 10839 22936
rect 10781 22927 10839 22933
rect 10962 22924 10968 22936
rect 11020 22924 11026 22976
rect 12713 22967 12771 22973
rect 12713 22933 12725 22967
rect 12759 22964 12771 22967
rect 14182 22964 14188 22976
rect 12759 22936 14188 22964
rect 12759 22933 12771 22936
rect 12713 22927 12771 22933
rect 14182 22924 14188 22936
rect 14240 22924 14246 22976
rect 14292 22964 14320 23004
rect 14360 23001 14372 23035
rect 14406 23032 14418 23035
rect 14458 23032 14464 23044
rect 14406 23004 14464 23032
rect 14406 23001 14418 23004
rect 14360 22995 14418 23001
rect 14458 22992 14464 23004
rect 14516 22992 14522 23044
rect 14568 23032 14596 23072
rect 14642 23060 14648 23112
rect 14700 23100 14706 23112
rect 15838 23100 15844 23112
rect 14700 23072 15844 23100
rect 14700 23060 14706 23072
rect 15838 23060 15844 23072
rect 15896 23060 15902 23112
rect 16224 23044 16252 23140
rect 16408 23140 17040 23168
rect 16408 23109 16436 23140
rect 17034 23128 17040 23140
rect 17092 23128 17098 23180
rect 17310 23168 17316 23180
rect 17271 23140 17316 23168
rect 17310 23128 17316 23140
rect 17368 23168 17374 23180
rect 17368 23140 18736 23168
rect 17368 23128 17374 23140
rect 16393 23103 16451 23109
rect 16393 23069 16405 23103
rect 16439 23069 16451 23103
rect 16393 23063 16451 23069
rect 16485 23103 16543 23109
rect 16485 23069 16497 23103
rect 16531 23069 16543 23103
rect 16485 23063 16543 23069
rect 16577 23103 16635 23109
rect 16577 23069 16589 23103
rect 16623 23069 16635 23103
rect 16577 23063 16635 23069
rect 16773 23103 16831 23109
rect 16773 23069 16785 23103
rect 16819 23100 16831 23103
rect 16942 23100 16948 23112
rect 16819 23072 16948 23100
rect 16819 23069 16831 23072
rect 16773 23063 16831 23069
rect 16114 23032 16120 23044
rect 14568 23004 16120 23032
rect 16114 22992 16120 23004
rect 16172 22992 16178 23044
rect 16206 22992 16212 23044
rect 16264 23032 16270 23044
rect 16500 23032 16528 23063
rect 16264 23004 16528 23032
rect 16592 23032 16620 23063
rect 16942 23060 16948 23072
rect 17000 23060 17006 23112
rect 17126 23060 17132 23112
rect 17184 23100 17190 23112
rect 17405 23103 17463 23109
rect 17405 23100 17417 23103
rect 17184 23072 17417 23100
rect 17184 23060 17190 23072
rect 17405 23069 17417 23072
rect 17451 23069 17463 23103
rect 18414 23100 18420 23112
rect 18375 23072 18420 23100
rect 17405 23063 17463 23069
rect 17034 23032 17040 23044
rect 16592 23004 17040 23032
rect 16264 22992 16270 23004
rect 17034 22992 17040 23004
rect 17092 22992 17098 23044
rect 16022 22964 16028 22976
rect 14292 22936 16028 22964
rect 16022 22924 16028 22936
rect 16080 22924 16086 22976
rect 17420 22964 17448 23063
rect 18414 23060 18420 23072
rect 18472 23060 18478 23112
rect 18708 23109 18736 23140
rect 19150 23128 19156 23180
rect 19208 23168 19214 23180
rect 19536 23168 19564 23208
rect 19794 23168 19800 23180
rect 19208 23140 19564 23168
rect 19711 23140 19800 23168
rect 19208 23128 19214 23140
rect 19711 23134 19739 23140
rect 18693 23103 18751 23109
rect 18693 23069 18705 23103
rect 18739 23069 18751 23103
rect 18693 23063 18751 23069
rect 19058 23060 19064 23112
rect 19116 23100 19122 23112
rect 19426 23100 19432 23112
rect 19116 23072 19432 23100
rect 19116 23060 19122 23072
rect 19426 23060 19432 23072
rect 19484 23060 19490 23112
rect 19521 23103 19579 23109
rect 19521 23069 19533 23103
rect 19567 23094 19579 23103
rect 19628 23106 19739 23134
rect 19794 23128 19800 23140
rect 19852 23128 19858 23180
rect 19996 23177 20024 23208
rect 21913 23205 21925 23239
rect 21959 23236 21971 23239
rect 22186 23236 22192 23248
rect 21959 23208 22192 23236
rect 21959 23205 21971 23208
rect 21913 23199 21971 23205
rect 22186 23196 22192 23208
rect 22244 23196 22250 23248
rect 22462 23196 22468 23248
rect 22520 23236 22526 23248
rect 22922 23236 22928 23248
rect 22520 23208 22928 23236
rect 22520 23196 22526 23208
rect 22922 23196 22928 23208
rect 22980 23196 22986 23248
rect 28442 23236 28448 23248
rect 24688 23208 28448 23236
rect 19981 23171 20039 23177
rect 19981 23137 19993 23171
rect 20027 23137 20039 23171
rect 19981 23131 20039 23137
rect 21008 23140 22416 23168
rect 19628 23094 19656 23106
rect 19567 23069 19656 23094
rect 19521 23066 19656 23069
rect 19521 23063 19579 23066
rect 20622 23060 20628 23112
rect 20680 23100 20686 23112
rect 21008 23100 21036 23140
rect 20680 23072 21036 23100
rect 20680 23060 20686 23072
rect 21358 23060 21364 23112
rect 21416 23100 21422 23112
rect 22094 23100 22100 23112
rect 21416 23072 22100 23100
rect 21416 23060 21422 23072
rect 22094 23060 22100 23072
rect 22152 23060 22158 23112
rect 22278 23100 22284 23112
rect 22239 23072 22284 23100
rect 22278 23060 22284 23072
rect 22336 23060 22342 23112
rect 22388 23109 22416 23140
rect 22738 23128 22744 23180
rect 22796 23168 22802 23180
rect 23658 23168 23664 23180
rect 22796 23140 23664 23168
rect 22796 23128 22802 23140
rect 23658 23128 23664 23140
rect 23716 23128 23722 23180
rect 22373 23103 22431 23109
rect 22373 23069 22385 23103
rect 22419 23069 22431 23103
rect 22373 23063 22431 23069
rect 23290 23060 23296 23112
rect 23348 23100 23354 23112
rect 23477 23103 23535 23109
rect 23477 23100 23489 23103
rect 23348 23072 23489 23100
rect 23348 23060 23354 23072
rect 23477 23069 23489 23072
rect 23523 23069 23535 23103
rect 23477 23063 23535 23069
rect 23566 23060 23572 23112
rect 23624 23100 23630 23112
rect 23750 23100 23756 23112
rect 23624 23072 23669 23100
rect 23711 23072 23756 23100
rect 23624 23060 23630 23072
rect 23750 23060 23756 23072
rect 23808 23060 23814 23112
rect 23842 23060 23848 23112
rect 23900 23100 23906 23112
rect 24118 23100 24124 23112
rect 23900 23072 24124 23100
rect 23900 23060 23906 23072
rect 24118 23060 24124 23072
rect 24176 23060 24182 23112
rect 24394 23100 24400 23112
rect 24355 23072 24400 23100
rect 24394 23060 24400 23072
rect 24452 23060 24458 23112
rect 24489 23103 24547 23109
rect 24489 23069 24501 23103
rect 24535 23100 24547 23103
rect 24688 23100 24716 23208
rect 28442 23196 28448 23208
rect 28500 23196 28506 23248
rect 25038 23128 25044 23180
rect 25096 23168 25102 23180
rect 25593 23171 25651 23177
rect 25593 23168 25605 23171
rect 25096 23140 25605 23168
rect 25096 23128 25102 23140
rect 25593 23137 25605 23140
rect 25639 23168 25651 23171
rect 26050 23168 26056 23180
rect 25639 23140 26056 23168
rect 25639 23137 25651 23140
rect 25593 23131 25651 23137
rect 26050 23128 26056 23140
rect 26108 23128 26114 23180
rect 26329 23171 26387 23177
rect 26329 23137 26341 23171
rect 26375 23168 26387 23171
rect 27154 23168 27160 23180
rect 26375 23140 27160 23168
rect 26375 23137 26387 23140
rect 26329 23131 26387 23137
rect 27154 23128 27160 23140
rect 27212 23128 27218 23180
rect 28169 23171 28227 23177
rect 28169 23137 28181 23171
rect 28215 23168 28227 23171
rect 28718 23168 28724 23180
rect 28215 23140 28724 23168
rect 28215 23137 28227 23140
rect 28169 23131 28227 23137
rect 28718 23128 28724 23140
rect 28776 23128 28782 23180
rect 24535 23072 24716 23100
rect 24535 23069 24547 23072
rect 24489 23063 24547 23069
rect 24762 23060 24768 23112
rect 24820 23100 24826 23112
rect 25501 23103 25559 23109
rect 25501 23100 25513 23103
rect 24820 23072 25513 23100
rect 24820 23060 24826 23072
rect 25501 23069 25513 23072
rect 25547 23069 25559 23103
rect 25501 23063 25559 23069
rect 17862 22992 17868 23044
rect 17920 23032 17926 23044
rect 18322 23032 18328 23044
rect 17920 23004 18328 23032
rect 17920 22992 17926 23004
rect 18322 22992 18328 23004
rect 18380 23032 18386 23044
rect 19245 23035 19303 23041
rect 19245 23032 19257 23035
rect 18380 23004 19257 23032
rect 18380 22992 18386 23004
rect 19245 23001 19257 23004
rect 19291 23001 19303 23035
rect 20070 23032 20076 23044
rect 19245 22995 19303 23001
rect 19352 23004 20076 23032
rect 19352 22973 19380 23004
rect 20070 22992 20076 23004
rect 20128 22992 20134 23044
rect 20248 23035 20306 23041
rect 20248 23001 20260 23035
rect 20294 23032 20306 23035
rect 21818 23032 21824 23044
rect 20294 23004 21824 23032
rect 20294 23001 20306 23004
rect 20248 22995 20306 23001
rect 21818 22992 21824 23004
rect 21876 22992 21882 23044
rect 22922 22992 22928 23044
rect 22980 23032 22986 23044
rect 24670 23032 24676 23044
rect 22980 23004 24532 23032
rect 24631 23004 24676 23032
rect 22980 22992 22986 23004
rect 18601 22967 18659 22973
rect 18601 22964 18613 22967
rect 17420 22936 18613 22964
rect 18601 22933 18613 22936
rect 18647 22933 18659 22967
rect 18601 22927 18659 22933
rect 19343 22967 19401 22973
rect 19343 22933 19355 22967
rect 19389 22933 19401 22967
rect 19343 22927 19401 22933
rect 19429 22967 19487 22973
rect 19429 22933 19441 22967
rect 19475 22964 19487 22967
rect 20898 22964 20904 22976
rect 19475 22936 20904 22964
rect 19475 22933 19487 22936
rect 19429 22927 19487 22933
rect 20898 22924 20904 22936
rect 20956 22964 20962 22976
rect 21361 22967 21419 22973
rect 21361 22964 21373 22967
rect 20956 22936 21373 22964
rect 20956 22924 20962 22936
rect 21361 22933 21373 22936
rect 21407 22933 21419 22967
rect 21361 22927 21419 22933
rect 23293 22967 23351 22973
rect 23293 22933 23305 22967
rect 23339 22964 23351 22967
rect 23934 22964 23940 22976
rect 23339 22936 23940 22964
rect 23339 22933 23351 22936
rect 23293 22927 23351 22933
rect 23934 22924 23940 22936
rect 23992 22924 23998 22976
rect 24118 22924 24124 22976
rect 24176 22964 24182 22976
rect 24397 22967 24455 22973
rect 24397 22964 24409 22967
rect 24176 22936 24409 22964
rect 24176 22924 24182 22936
rect 24397 22933 24409 22936
rect 24443 22933 24455 22967
rect 24504 22964 24532 23004
rect 24670 22992 24676 23004
rect 24728 22992 24734 23044
rect 25222 22992 25228 23044
rect 25280 23032 25286 23044
rect 26513 23035 26571 23041
rect 26513 23032 26525 23035
rect 25280 23004 26525 23032
rect 25280 22992 25286 23004
rect 26513 23001 26525 23004
rect 26559 23001 26571 23035
rect 26513 22995 26571 23001
rect 24854 22964 24860 22976
rect 24504 22936 24860 22964
rect 24397 22927 24455 22933
rect 24854 22924 24860 22936
rect 24912 22964 24918 22976
rect 25133 22967 25191 22973
rect 25133 22964 25145 22967
rect 24912 22936 25145 22964
rect 24912 22924 24918 22936
rect 25133 22933 25145 22936
rect 25179 22933 25191 22967
rect 25133 22927 25191 22933
rect 25777 22967 25835 22973
rect 25777 22933 25789 22967
rect 25823 22964 25835 22967
rect 27062 22964 27068 22976
rect 25823 22936 27068 22964
rect 25823 22933 25835 22936
rect 25777 22927 25835 22933
rect 27062 22924 27068 22936
rect 27120 22924 27126 22976
rect 1104 22874 28888 22896
rect 1104 22822 10214 22874
rect 10266 22822 10278 22874
rect 10330 22822 10342 22874
rect 10394 22822 10406 22874
rect 10458 22822 10470 22874
rect 10522 22822 19478 22874
rect 19530 22822 19542 22874
rect 19594 22822 19606 22874
rect 19658 22822 19670 22874
rect 19722 22822 19734 22874
rect 19786 22822 28888 22874
rect 1104 22800 28888 22822
rect 2498 22760 2504 22772
rect 2459 22732 2504 22760
rect 2498 22720 2504 22732
rect 2556 22720 2562 22772
rect 13449 22763 13507 22769
rect 13449 22729 13461 22763
rect 13495 22760 13507 22763
rect 13538 22760 13544 22772
rect 13495 22732 13544 22760
rect 13495 22729 13507 22732
rect 13449 22723 13507 22729
rect 13538 22720 13544 22732
rect 13596 22760 13602 22772
rect 13596 22732 15240 22760
rect 13596 22720 13602 22732
rect 10873 22695 10931 22701
rect 10873 22661 10885 22695
rect 10919 22692 10931 22695
rect 15212 22692 15240 22732
rect 15286 22720 15292 22772
rect 15344 22760 15350 22772
rect 16117 22763 16175 22769
rect 16117 22760 16129 22763
rect 15344 22732 16129 22760
rect 15344 22720 15350 22732
rect 16117 22729 16129 22732
rect 16163 22760 16175 22763
rect 16942 22760 16948 22772
rect 16163 22732 16948 22760
rect 16163 22729 16175 22732
rect 16117 22723 16175 22729
rect 16942 22720 16948 22732
rect 17000 22720 17006 22772
rect 17865 22763 17923 22769
rect 17865 22729 17877 22763
rect 17911 22760 17923 22763
rect 18046 22760 18052 22772
rect 17911 22732 18052 22760
rect 17911 22729 17923 22732
rect 17865 22723 17923 22729
rect 18046 22720 18052 22732
rect 18104 22720 18110 22772
rect 18138 22720 18144 22772
rect 18196 22760 18202 22772
rect 21634 22760 21640 22772
rect 18196 22732 21640 22760
rect 18196 22720 18202 22732
rect 21634 22720 21640 22732
rect 21692 22720 21698 22772
rect 21818 22760 21824 22772
rect 21779 22732 21824 22760
rect 21818 22720 21824 22732
rect 21876 22720 21882 22772
rect 24486 22760 24492 22772
rect 23308 22732 24492 22760
rect 15470 22692 15476 22704
rect 10919 22664 15056 22692
rect 10919 22661 10931 22664
rect 10873 22655 10931 22661
rect 2409 22627 2467 22633
rect 2409 22593 2421 22627
rect 2455 22624 2467 22627
rect 2590 22624 2596 22636
rect 2455 22596 2596 22624
rect 2455 22593 2467 22596
rect 2409 22587 2467 22593
rect 2590 22584 2596 22596
rect 2648 22624 2654 22636
rect 4982 22624 4988 22636
rect 2648 22596 4988 22624
rect 2648 22584 2654 22596
rect 4982 22584 4988 22596
rect 5040 22584 5046 22636
rect 10778 22624 10784 22636
rect 10739 22596 10784 22624
rect 10778 22584 10784 22596
rect 10836 22584 10842 22636
rect 10962 22624 10968 22636
rect 10923 22596 10968 22624
rect 10962 22584 10968 22596
rect 11020 22584 11026 22636
rect 11054 22584 11060 22636
rect 11112 22624 11118 22636
rect 11974 22624 11980 22636
rect 11112 22596 11980 22624
rect 11112 22584 11118 22596
rect 11974 22584 11980 22596
rect 12032 22584 12038 22636
rect 12618 22624 12624 22636
rect 12579 22596 12624 22624
rect 12618 22584 12624 22596
rect 12676 22584 12682 22636
rect 13170 22584 13176 22636
rect 13228 22624 13234 22636
rect 13265 22627 13323 22633
rect 13265 22624 13277 22627
rect 13228 22596 13277 22624
rect 13228 22584 13234 22596
rect 13265 22593 13277 22596
rect 13311 22593 13323 22627
rect 13265 22587 13323 22593
rect 13541 22627 13599 22633
rect 13541 22593 13553 22627
rect 13587 22593 13599 22627
rect 14090 22624 14096 22636
rect 14051 22596 14096 22624
rect 13541 22587 13599 22593
rect 13556 22556 13584 22587
rect 14090 22584 14096 22596
rect 14148 22624 14154 22636
rect 14826 22624 14832 22636
rect 14148 22596 14832 22624
rect 14148 22584 14154 22596
rect 14826 22584 14832 22596
rect 14884 22584 14890 22636
rect 14921 22627 14979 22633
rect 14921 22593 14933 22627
rect 14967 22593 14979 22627
rect 14921 22587 14979 22593
rect 13906 22556 13912 22568
rect 13556 22528 13912 22556
rect 13906 22516 13912 22528
rect 13964 22556 13970 22568
rect 14277 22559 14335 22565
rect 14277 22556 14289 22559
rect 13964 22528 14289 22556
rect 13964 22516 13970 22528
rect 14277 22525 14289 22528
rect 14323 22525 14335 22559
rect 14277 22519 14335 22525
rect 14458 22516 14464 22568
rect 14516 22556 14522 22568
rect 14737 22559 14795 22565
rect 14737 22556 14749 22559
rect 14516 22528 14749 22556
rect 14516 22516 14522 22528
rect 14737 22525 14749 22528
rect 14783 22525 14795 22559
rect 14737 22519 14795 22525
rect 13265 22491 13323 22497
rect 13265 22457 13277 22491
rect 13311 22488 13323 22491
rect 14936 22488 14964 22587
rect 15028 22556 15056 22664
rect 15212 22664 15476 22692
rect 15212 22633 15240 22664
rect 15470 22652 15476 22664
rect 15528 22652 15534 22704
rect 17126 22692 17132 22704
rect 15856 22664 17132 22692
rect 15197 22627 15255 22633
rect 15197 22593 15209 22627
rect 15243 22593 15255 22627
rect 15746 22624 15752 22636
rect 15707 22596 15752 22624
rect 15197 22587 15255 22593
rect 15746 22584 15752 22596
rect 15804 22584 15810 22636
rect 15856 22556 15884 22664
rect 17126 22652 17132 22664
rect 17184 22652 17190 22704
rect 19150 22692 19156 22704
rect 18616 22664 19156 22692
rect 15933 22627 15991 22633
rect 15933 22593 15945 22627
rect 15979 22593 15991 22627
rect 16666 22624 16672 22636
rect 16627 22596 16672 22624
rect 15933 22587 15991 22593
rect 15028 22528 15884 22556
rect 15948 22556 15976 22587
rect 16666 22584 16672 22596
rect 16724 22584 16730 22636
rect 16758 22584 16764 22636
rect 16816 22624 16822 22636
rect 17497 22627 17555 22633
rect 17497 22624 17509 22627
rect 16816 22596 17509 22624
rect 16816 22584 16822 22596
rect 17497 22593 17509 22596
rect 17543 22624 17555 22627
rect 18506 22624 18512 22636
rect 17543 22596 18512 22624
rect 17543 22593 17555 22596
rect 17497 22587 17555 22593
rect 18506 22584 18512 22596
rect 18564 22584 18570 22636
rect 18616 22633 18644 22664
rect 19150 22652 19156 22664
rect 19208 22652 19214 22704
rect 20070 22652 20076 22704
rect 20128 22692 20134 22704
rect 20128 22664 22048 22692
rect 20128 22652 20134 22664
rect 18601 22627 18659 22633
rect 18601 22593 18613 22627
rect 18647 22593 18659 22627
rect 18601 22587 18659 22593
rect 18868 22627 18926 22633
rect 18868 22593 18880 22627
rect 18914 22624 18926 22627
rect 19334 22624 19340 22636
rect 18914 22596 19340 22624
rect 18914 22593 18926 22596
rect 18868 22587 18926 22593
rect 19334 22584 19340 22596
rect 19392 22584 19398 22636
rect 19426 22584 19432 22636
rect 19484 22624 19490 22636
rect 19484 22596 19656 22624
rect 19484 22584 19490 22596
rect 16022 22556 16028 22568
rect 15948 22528 16028 22556
rect 16022 22516 16028 22528
rect 16080 22516 16086 22568
rect 16114 22516 16120 22568
rect 16172 22556 16178 22568
rect 17034 22556 17040 22568
rect 16172 22528 17040 22556
rect 16172 22516 16178 22528
rect 17034 22516 17040 22528
rect 17092 22516 17098 22568
rect 17589 22559 17647 22565
rect 17589 22525 17601 22559
rect 17635 22556 17647 22559
rect 17770 22556 17776 22568
rect 17635 22528 17776 22556
rect 17635 22525 17647 22528
rect 17589 22519 17647 22525
rect 17770 22516 17776 22528
rect 17828 22516 17834 22568
rect 19628 22556 19656 22596
rect 20254 22584 20260 22636
rect 20312 22624 20318 22636
rect 20625 22627 20683 22633
rect 20625 22624 20637 22627
rect 20312 22596 20637 22624
rect 20312 22584 20318 22596
rect 20625 22593 20637 22596
rect 20671 22593 20683 22627
rect 20625 22587 20683 22593
rect 20717 22627 20775 22633
rect 20717 22593 20729 22627
rect 20763 22593 20775 22627
rect 20990 22624 20996 22636
rect 20951 22596 20996 22624
rect 20717 22587 20775 22593
rect 20732 22556 20760 22587
rect 20990 22584 20996 22596
rect 21048 22584 21054 22636
rect 22020 22633 22048 22664
rect 22646 22652 22652 22704
rect 22704 22692 22710 22704
rect 23308 22692 23336 22732
rect 24486 22720 24492 22732
rect 24544 22720 24550 22772
rect 25130 22692 25136 22704
rect 22704 22664 23336 22692
rect 22704 22652 22710 22664
rect 22005 22627 22063 22633
rect 22005 22593 22017 22627
rect 22051 22593 22063 22627
rect 22005 22587 22063 22593
rect 23014 22584 23020 22636
rect 23072 22624 23078 22636
rect 23198 22624 23204 22636
rect 23072 22596 23204 22624
rect 23072 22584 23078 22596
rect 23198 22584 23204 22596
rect 23256 22584 23262 22636
rect 23308 22633 23336 22664
rect 24136 22664 25136 22692
rect 23293 22627 23351 22633
rect 23293 22593 23305 22627
rect 23339 22593 23351 22627
rect 23293 22587 23351 22593
rect 23382 22584 23388 22636
rect 23440 22624 23446 22636
rect 23569 22627 23627 22633
rect 23440 22596 23485 22624
rect 23440 22584 23446 22596
rect 23569 22593 23581 22627
rect 23615 22624 23627 22627
rect 23658 22624 23664 22636
rect 23615 22596 23664 22624
rect 23615 22593 23627 22596
rect 23569 22587 23627 22593
rect 23658 22584 23664 22596
rect 23716 22584 23722 22636
rect 20898 22556 20904 22568
rect 19628 22528 20760 22556
rect 20859 22528 20904 22556
rect 20898 22516 20904 22528
rect 20956 22556 20962 22568
rect 24136 22565 24164 22664
rect 25130 22652 25136 22664
rect 25188 22652 25194 22704
rect 24213 22627 24271 22633
rect 24213 22593 24225 22627
rect 24259 22624 24271 22627
rect 24762 22624 24768 22636
rect 24259 22596 24768 22624
rect 24259 22594 24287 22596
rect 24259 22593 24271 22594
rect 24213 22587 24271 22593
rect 24762 22584 24768 22596
rect 24820 22584 24826 22636
rect 25297 22627 25355 22633
rect 25297 22624 25309 22627
rect 24872 22596 25309 22624
rect 22281 22559 22339 22565
rect 22281 22556 22293 22559
rect 20956 22528 22293 22556
rect 20956 22516 20962 22528
rect 22281 22525 22293 22528
rect 22327 22525 22339 22559
rect 24121 22559 24179 22565
rect 24121 22556 24133 22559
rect 22281 22519 22339 22525
rect 23584 22528 24133 22556
rect 13311 22460 14964 22488
rect 13311 22457 13323 22460
rect 13265 22451 13323 22457
rect 15010 22448 15016 22500
rect 15068 22488 15074 22500
rect 15562 22488 15568 22500
rect 15068 22460 15568 22488
rect 15068 22448 15074 22460
rect 15562 22448 15568 22460
rect 15620 22448 15626 22500
rect 16224 22460 16896 22488
rect 12066 22420 12072 22432
rect 12027 22392 12072 22420
rect 12066 22380 12072 22392
rect 12124 22380 12130 22432
rect 12713 22423 12771 22429
rect 12713 22389 12725 22423
rect 12759 22420 12771 22423
rect 14642 22420 14648 22432
rect 12759 22392 14648 22420
rect 12759 22389 12771 22392
rect 12713 22383 12771 22389
rect 14642 22380 14648 22392
rect 14700 22380 14706 22432
rect 15105 22423 15163 22429
rect 15105 22389 15117 22423
rect 15151 22420 15163 22423
rect 15378 22420 15384 22432
rect 15151 22392 15384 22420
rect 15151 22389 15163 22392
rect 15105 22383 15163 22389
rect 15378 22380 15384 22392
rect 15436 22420 15442 22432
rect 15654 22420 15660 22432
rect 15436 22392 15660 22420
rect 15436 22380 15442 22392
rect 15654 22380 15660 22392
rect 15712 22380 15718 22432
rect 15838 22380 15844 22432
rect 15896 22420 15902 22432
rect 16224 22420 16252 22460
rect 16758 22420 16764 22432
rect 15896 22392 16252 22420
rect 16719 22392 16764 22420
rect 15896 22380 15902 22392
rect 16758 22380 16764 22392
rect 16816 22380 16822 22432
rect 16868 22420 16896 22460
rect 16942 22448 16948 22500
rect 17000 22488 17006 22500
rect 18414 22488 18420 22500
rect 17000 22460 18420 22488
rect 17000 22448 17006 22460
rect 18414 22448 18420 22460
rect 18472 22448 18478 22500
rect 20162 22488 20168 22500
rect 19536 22460 20168 22488
rect 19536 22420 19564 22460
rect 20162 22448 20168 22460
rect 20220 22488 20226 22500
rect 23584 22488 23612 22528
rect 24121 22525 24133 22528
rect 24167 22525 24179 22559
rect 24121 22519 24179 22525
rect 20220 22460 23612 22488
rect 20220 22448 20226 22460
rect 23658 22448 23664 22500
rect 23716 22488 23722 22500
rect 24581 22491 24639 22497
rect 24581 22488 24593 22491
rect 23716 22460 24593 22488
rect 23716 22448 23722 22460
rect 24581 22457 24593 22460
rect 24627 22457 24639 22491
rect 24581 22451 24639 22457
rect 24670 22448 24676 22500
rect 24728 22488 24734 22500
rect 24872 22488 24900 22596
rect 25297 22593 25309 22596
rect 25343 22593 25355 22627
rect 25297 22587 25355 22593
rect 25682 22584 25688 22636
rect 25740 22624 25746 22636
rect 27157 22627 27215 22633
rect 27157 22624 27169 22627
rect 25740 22596 27169 22624
rect 25740 22584 25746 22596
rect 27157 22593 27169 22596
rect 27203 22593 27215 22627
rect 27157 22587 27215 22593
rect 27706 22584 27712 22636
rect 27764 22624 27770 22636
rect 27985 22627 28043 22633
rect 27985 22624 27997 22627
rect 27764 22596 27997 22624
rect 27764 22584 27770 22596
rect 27985 22593 27997 22596
rect 28031 22624 28043 22627
rect 28350 22624 28356 22636
rect 28031 22596 28356 22624
rect 28031 22593 28043 22596
rect 27985 22587 28043 22593
rect 28350 22584 28356 22596
rect 28408 22584 28414 22636
rect 25038 22556 25044 22568
rect 24999 22528 25044 22556
rect 25038 22516 25044 22528
rect 25096 22516 25102 22568
rect 27062 22556 27068 22568
rect 27023 22528 27068 22556
rect 27062 22516 27068 22528
rect 27120 22516 27126 22568
rect 24728 22460 24900 22488
rect 24728 22448 24734 22460
rect 16868 22392 19564 22420
rect 19610 22380 19616 22432
rect 19668 22420 19674 22432
rect 19981 22423 20039 22429
rect 19981 22420 19993 22423
rect 19668 22392 19993 22420
rect 19668 22380 19674 22392
rect 19981 22389 19993 22392
rect 20027 22389 20039 22423
rect 20438 22420 20444 22432
rect 20399 22392 20444 22420
rect 19981 22383 20039 22389
rect 20438 22380 20444 22392
rect 20496 22380 20502 22432
rect 20806 22380 20812 22432
rect 20864 22420 20870 22432
rect 22189 22423 22247 22429
rect 22189 22420 22201 22423
rect 20864 22392 22201 22420
rect 20864 22380 20870 22392
rect 22189 22389 22201 22392
rect 22235 22389 22247 22423
rect 22189 22383 22247 22389
rect 22925 22423 22983 22429
rect 22925 22389 22937 22423
rect 22971 22420 22983 22423
rect 23014 22420 23020 22432
rect 22971 22392 23020 22420
rect 22971 22389 22983 22392
rect 22925 22383 22983 22389
rect 23014 22380 23020 22392
rect 23072 22380 23078 22432
rect 23290 22380 23296 22432
rect 23348 22420 23354 22432
rect 25682 22420 25688 22432
rect 23348 22392 25688 22420
rect 23348 22380 23354 22392
rect 25682 22380 25688 22392
rect 25740 22380 25746 22432
rect 26421 22423 26479 22429
rect 26421 22389 26433 22423
rect 26467 22420 26479 22423
rect 27246 22420 27252 22432
rect 26467 22392 27252 22420
rect 26467 22389 26479 22392
rect 26421 22383 26479 22389
rect 27246 22380 27252 22392
rect 27304 22380 27310 22432
rect 27430 22420 27436 22432
rect 27391 22392 27436 22420
rect 27430 22380 27436 22392
rect 27488 22380 27494 22432
rect 27522 22380 27528 22432
rect 27580 22420 27586 22432
rect 28077 22423 28135 22429
rect 28077 22420 28089 22423
rect 27580 22392 28089 22420
rect 27580 22380 27586 22392
rect 28077 22389 28089 22392
rect 28123 22389 28135 22423
rect 28077 22383 28135 22389
rect 1104 22330 28888 22352
rect 1104 22278 5582 22330
rect 5634 22278 5646 22330
rect 5698 22278 5710 22330
rect 5762 22278 5774 22330
rect 5826 22278 5838 22330
rect 5890 22278 14846 22330
rect 14898 22278 14910 22330
rect 14962 22278 14974 22330
rect 15026 22278 15038 22330
rect 15090 22278 15102 22330
rect 15154 22278 24110 22330
rect 24162 22278 24174 22330
rect 24226 22278 24238 22330
rect 24290 22278 24302 22330
rect 24354 22278 24366 22330
rect 24418 22278 28888 22330
rect 1104 22256 28888 22278
rect 10778 22176 10784 22228
rect 10836 22216 10842 22228
rect 14734 22216 14740 22228
rect 10836 22188 14740 22216
rect 10836 22176 10842 22188
rect 14734 22176 14740 22188
rect 14792 22176 14798 22228
rect 15381 22219 15439 22225
rect 15381 22185 15393 22219
rect 15427 22216 15439 22219
rect 15654 22216 15660 22228
rect 15427 22188 15660 22216
rect 15427 22185 15439 22188
rect 15381 22179 15439 22185
rect 15654 22176 15660 22188
rect 15712 22176 15718 22228
rect 16298 22216 16304 22228
rect 15948 22188 16304 22216
rect 12066 22108 12072 22160
rect 12124 22148 12130 22160
rect 15948 22148 15976 22188
rect 16298 22176 16304 22188
rect 16356 22176 16362 22228
rect 16758 22176 16764 22228
rect 16816 22216 16822 22228
rect 24026 22216 24032 22228
rect 16816 22188 24032 22216
rect 16816 22176 16822 22188
rect 24026 22176 24032 22188
rect 24084 22176 24090 22228
rect 24486 22176 24492 22228
rect 24544 22216 24550 22228
rect 25685 22219 25743 22225
rect 24544 22188 24808 22216
rect 24544 22176 24550 22188
rect 17494 22148 17500 22160
rect 12124 22120 15976 22148
rect 16040 22120 17500 22148
rect 12124 22108 12130 22120
rect 11977 22083 12035 22089
rect 11977 22049 11989 22083
rect 12023 22080 12035 22083
rect 14366 22080 14372 22092
rect 12023 22052 14372 22080
rect 12023 22049 12035 22052
rect 11977 22043 12035 22049
rect 14366 22040 14372 22052
rect 14424 22040 14430 22092
rect 14533 22083 14591 22089
rect 14533 22049 14545 22083
rect 14579 22080 14591 22083
rect 15838 22080 15844 22092
rect 14579 22052 15844 22080
rect 14579 22049 14591 22052
rect 14533 22043 14591 22049
rect 15838 22040 15844 22052
rect 15896 22040 15902 22092
rect 11238 22012 11244 22024
rect 11199 21984 11244 22012
rect 11238 21972 11244 21984
rect 11296 21972 11302 22024
rect 11609 22015 11667 22021
rect 11609 21981 11621 22015
rect 11655 22012 11667 22015
rect 11882 22012 11888 22024
rect 11655 21984 11888 22012
rect 11655 21981 11667 21984
rect 11609 21975 11667 21981
rect 11882 21972 11888 21984
rect 11940 21972 11946 22024
rect 12069 22015 12127 22021
rect 12069 21981 12081 22015
rect 12115 21981 12127 22015
rect 12069 21975 12127 21981
rect 12621 22015 12679 22021
rect 12621 21981 12633 22015
rect 12667 22012 12679 22015
rect 12667 21984 13308 22012
rect 12667 21981 12679 21984
rect 12621 21975 12679 21981
rect 12084 21876 12112 21975
rect 12802 21944 12808 21956
rect 12763 21916 12808 21944
rect 12802 21904 12808 21916
rect 12860 21904 12866 21956
rect 13280 21944 13308 21984
rect 13354 21972 13360 22024
rect 13412 22012 13418 22024
rect 13412 21984 13457 22012
rect 13412 21972 13418 21984
rect 13998 21972 14004 22024
rect 14056 22012 14062 22024
rect 14645 22015 14703 22021
rect 14645 22012 14657 22015
rect 14056 21984 14657 22012
rect 14056 21972 14062 21984
rect 14645 21981 14657 21984
rect 14691 21981 14703 22015
rect 15010 22012 15016 22024
rect 14936 22002 15016 22012
rect 14752 21999 15016 22002
rect 14645 21975 14703 21981
rect 14737 21993 15016 21999
rect 14737 21959 14749 21993
rect 14783 21984 15016 21993
rect 14783 21974 14964 21984
rect 14783 21959 14795 21974
rect 15010 21972 15016 21984
rect 15068 21972 15074 22024
rect 15746 22012 15752 22024
rect 15120 21984 15752 22012
rect 13446 21944 13452 21956
rect 13280 21916 13452 21944
rect 13446 21904 13452 21916
rect 13504 21904 13510 21956
rect 13541 21947 13599 21953
rect 13541 21913 13553 21947
rect 13587 21944 13599 21947
rect 13630 21944 13636 21956
rect 13587 21916 13636 21944
rect 13587 21913 13599 21916
rect 13541 21907 13599 21913
rect 13630 21904 13636 21916
rect 13688 21904 13694 21956
rect 14458 21944 14464 21956
rect 14419 21916 14464 21944
rect 14458 21904 14464 21916
rect 14516 21904 14522 21956
rect 14737 21953 14795 21959
rect 15120 21944 15148 21984
rect 15746 21972 15752 21984
rect 15804 21972 15810 22024
rect 16040 21953 16068 22120
rect 17494 22108 17500 22120
rect 17552 22108 17558 22160
rect 17862 22108 17868 22160
rect 17920 22148 17926 22160
rect 18049 22151 18107 22157
rect 18049 22148 18061 22151
rect 17920 22120 18061 22148
rect 17920 22108 17926 22120
rect 18049 22117 18061 22120
rect 18095 22117 18107 22151
rect 20990 22148 20996 22160
rect 18049 22111 18107 22117
rect 20916 22120 20996 22148
rect 16097 22083 16155 22089
rect 16097 22049 16109 22083
rect 16143 22080 16155 22083
rect 19242 22080 19248 22092
rect 16143 22052 17540 22080
rect 16143 22049 16155 22052
rect 16097 22043 16155 22049
rect 16301 22015 16359 22021
rect 16301 21981 16313 22015
rect 16347 22012 16359 22015
rect 16574 22012 16580 22024
rect 16347 21984 16580 22012
rect 16347 21981 16359 21984
rect 16301 21975 16359 21981
rect 16574 21972 16580 21984
rect 16632 21972 16638 22024
rect 14844 21916 15148 21944
rect 15197 21947 15255 21953
rect 14844 21876 14872 21916
rect 15197 21913 15209 21947
rect 15243 21913 15255 21947
rect 15197 21907 15255 21913
rect 16025 21947 16083 21953
rect 16025 21913 16037 21947
rect 16071 21913 16083 21947
rect 16025 21907 16083 21913
rect 12084 21848 14872 21876
rect 15010 21836 15016 21888
rect 15068 21876 15074 21888
rect 15212 21876 15240 21907
rect 16482 21904 16488 21956
rect 16540 21944 16546 21956
rect 16761 21947 16819 21953
rect 16761 21944 16773 21947
rect 16540 21916 16773 21944
rect 16540 21904 16546 21916
rect 16761 21913 16773 21916
rect 16807 21913 16819 21947
rect 16942 21944 16948 21956
rect 16903 21916 16948 21944
rect 16761 21907 16819 21913
rect 16942 21904 16948 21916
rect 17000 21904 17006 21956
rect 17126 21904 17132 21956
rect 17184 21944 17190 21956
rect 17512 21944 17540 22052
rect 18064 22052 18368 22080
rect 19203 22052 19248 22080
rect 17678 22012 17684 22024
rect 17639 21984 17684 22012
rect 17678 21972 17684 21984
rect 17736 21972 17742 22024
rect 17865 22015 17923 22021
rect 17865 21981 17877 22015
rect 17911 22012 17923 22015
rect 18064 22012 18092 22052
rect 18340 22024 18368 22052
rect 19242 22040 19248 22052
rect 19300 22040 19306 22092
rect 19610 22080 19616 22092
rect 19571 22052 19616 22080
rect 19610 22040 19616 22052
rect 19668 22040 19674 22092
rect 20070 22080 20076 22092
rect 20031 22052 20076 22080
rect 20070 22040 20076 22052
rect 20128 22040 20134 22092
rect 20438 22080 20444 22092
rect 20399 22052 20444 22080
rect 20438 22040 20444 22052
rect 20496 22040 20502 22092
rect 17911 21984 18092 22012
rect 18141 22015 18199 22021
rect 17911 21981 17923 21984
rect 17865 21975 17923 21981
rect 18141 21981 18153 22015
rect 18187 22012 18199 22015
rect 18230 22012 18236 22024
rect 18187 21984 18236 22012
rect 18187 21981 18199 21984
rect 18141 21975 18199 21981
rect 18230 21972 18236 21984
rect 18288 21972 18294 22024
rect 18322 21972 18328 22024
rect 18380 21972 18386 22024
rect 18598 21972 18604 22024
rect 18656 22012 18662 22024
rect 19429 22015 19487 22021
rect 19429 22012 19441 22015
rect 18656 21984 19441 22012
rect 18656 21972 18662 21984
rect 19429 21981 19441 21984
rect 19475 21981 19487 22015
rect 19429 21975 19487 21981
rect 19886 21972 19892 22024
rect 19944 21972 19950 22024
rect 20162 21972 20168 22024
rect 20220 22012 20226 22024
rect 20916 22021 20944 22120
rect 20990 22108 20996 22120
rect 21048 22108 21054 22160
rect 22830 22108 22836 22160
rect 22888 22148 22894 22160
rect 23290 22148 23296 22160
rect 22888 22120 23296 22148
rect 22888 22108 22894 22120
rect 23290 22108 23296 22120
rect 23348 22108 23354 22160
rect 21358 22040 21364 22092
rect 21416 22080 21422 22092
rect 23845 22083 23903 22089
rect 23845 22080 23857 22083
rect 21416 22052 21872 22080
rect 21416 22040 21422 22052
rect 20533 22015 20591 22021
rect 20533 22012 20545 22015
rect 20220 21984 20545 22012
rect 20220 21972 20226 21984
rect 20533 21981 20545 21984
rect 20579 21981 20591 22015
rect 20533 21975 20591 21981
rect 20901 22015 20959 22021
rect 20901 21981 20913 22015
rect 20947 21981 20959 22015
rect 20901 21975 20959 21981
rect 20990 21972 20996 22024
rect 21048 22012 21054 22024
rect 21726 22012 21732 22024
rect 21048 21984 21093 22012
rect 21687 21984 21732 22012
rect 21048 21972 21054 21984
rect 21726 21972 21732 21984
rect 21784 21972 21790 22024
rect 21844 22012 21872 22052
rect 22940 22052 23857 22080
rect 22940 22012 22968 22052
rect 23845 22049 23857 22052
rect 23891 22049 23903 22083
rect 23845 22043 23903 22049
rect 23658 22012 23664 22024
rect 21844 21984 22968 22012
rect 23619 21984 23664 22012
rect 23658 21972 23664 21984
rect 23716 21972 23722 22024
rect 24670 22012 24676 22024
rect 24631 21984 24676 22012
rect 24670 21972 24676 21984
rect 24728 21972 24734 22024
rect 24780 22021 24808 22188
rect 25685 22185 25697 22219
rect 25731 22216 25743 22219
rect 26050 22216 26056 22228
rect 25731 22188 26056 22216
rect 25731 22185 25743 22188
rect 25685 22179 25743 22185
rect 26050 22176 26056 22188
rect 26108 22176 26114 22228
rect 25590 22040 25596 22092
rect 25648 22080 25654 22092
rect 26513 22083 26571 22089
rect 26513 22080 26525 22083
rect 25648 22052 26525 22080
rect 25648 22040 25654 22052
rect 26513 22049 26525 22052
rect 26559 22049 26571 22083
rect 28166 22080 28172 22092
rect 28127 22052 28172 22080
rect 26513 22043 26571 22049
rect 28166 22040 28172 22052
rect 28224 22040 28230 22092
rect 24765 22015 24823 22021
rect 24765 21981 24777 22015
rect 24811 21981 24823 22015
rect 24765 21975 24823 21981
rect 24857 22015 24915 22021
rect 24857 21981 24869 22015
rect 24903 21981 24915 22015
rect 24857 21975 24915 21981
rect 19904 21944 19932 21972
rect 20070 21944 20076 21956
rect 17184 21916 17229 21944
rect 17512 21916 19334 21944
rect 19904 21916 20076 21944
rect 17184 21904 17190 21916
rect 15068 21848 15240 21876
rect 15068 21836 15074 21848
rect 15378 21836 15384 21888
rect 15436 21885 15442 21888
rect 15436 21879 15455 21885
rect 15443 21845 15455 21879
rect 15562 21876 15568 21888
rect 15523 21848 15568 21876
rect 15436 21839 15455 21845
rect 15436 21836 15442 21839
rect 15562 21836 15568 21848
rect 15620 21836 15626 21888
rect 16114 21836 16120 21888
rect 16172 21876 16178 21888
rect 16209 21879 16267 21885
rect 16209 21876 16221 21879
rect 16172 21848 16221 21876
rect 16172 21836 16178 21848
rect 16209 21845 16221 21848
rect 16255 21845 16267 21879
rect 16209 21839 16267 21845
rect 16298 21836 16304 21888
rect 16356 21876 16362 21888
rect 19150 21876 19156 21888
rect 16356 21848 19156 21876
rect 16356 21836 16362 21848
rect 19150 21836 19156 21848
rect 19208 21836 19214 21888
rect 19306 21876 19334 21916
rect 20070 21904 20076 21916
rect 20128 21904 20134 21956
rect 20257 21947 20315 21953
rect 20257 21913 20269 21947
rect 20303 21944 20315 21947
rect 20346 21944 20352 21956
rect 20303 21916 20352 21944
rect 20303 21913 20315 21916
rect 20257 21907 20315 21913
rect 20346 21904 20352 21916
rect 20404 21904 20410 21956
rect 21974 21947 22032 21953
rect 21974 21944 21986 21947
rect 20456 21916 21986 21944
rect 20456 21876 20484 21916
rect 21974 21913 21986 21916
rect 22020 21913 22032 21947
rect 23566 21944 23572 21956
rect 21974 21907 22032 21913
rect 22572 21916 23572 21944
rect 19306 21848 20484 21876
rect 21358 21836 21364 21888
rect 21416 21876 21422 21888
rect 22572 21876 22600 21916
rect 23566 21904 23572 21916
rect 23624 21904 23630 21956
rect 24578 21904 24584 21956
rect 24636 21944 24642 21956
rect 24872 21944 24900 21975
rect 24946 21972 24952 22024
rect 25004 22012 25010 22024
rect 25041 22015 25099 22021
rect 25041 22012 25053 22015
rect 25004 21984 25053 22012
rect 25004 21972 25010 21984
rect 25041 21981 25053 21984
rect 25087 21981 25099 22015
rect 25041 21975 25099 21981
rect 25406 21972 25412 22024
rect 25464 22012 25470 22024
rect 26329 22015 26387 22021
rect 26329 22012 26341 22015
rect 25464 21984 26341 22012
rect 25464 21972 25470 21984
rect 26329 21981 26341 21984
rect 26375 21981 26387 22015
rect 26329 21975 26387 21981
rect 25498 21944 25504 21956
rect 24636 21916 24900 21944
rect 25459 21916 25504 21944
rect 24636 21904 24642 21916
rect 25498 21904 25504 21916
rect 25556 21904 25562 21956
rect 25717 21947 25775 21953
rect 25717 21913 25729 21947
rect 25763 21944 25775 21947
rect 25763 21916 26464 21944
rect 25763 21913 25775 21916
rect 25717 21907 25775 21913
rect 21416 21848 22600 21876
rect 21416 21836 21422 21848
rect 22646 21836 22652 21888
rect 22704 21876 22710 21888
rect 23109 21879 23167 21885
rect 23109 21876 23121 21879
rect 22704 21848 23121 21876
rect 22704 21836 22710 21848
rect 23109 21845 23121 21848
rect 23155 21845 23167 21879
rect 23109 21839 23167 21845
rect 24397 21879 24455 21885
rect 24397 21845 24409 21879
rect 24443 21876 24455 21879
rect 24670 21876 24676 21888
rect 24443 21848 24676 21876
rect 24443 21845 24455 21848
rect 24397 21839 24455 21845
rect 24670 21836 24676 21848
rect 24728 21836 24734 21888
rect 25869 21879 25927 21885
rect 25869 21845 25881 21879
rect 25915 21876 25927 21879
rect 25958 21876 25964 21888
rect 25915 21848 25964 21876
rect 25915 21845 25927 21848
rect 25869 21839 25927 21845
rect 25958 21836 25964 21848
rect 26016 21836 26022 21888
rect 26436 21876 26464 21916
rect 27706 21876 27712 21888
rect 26436 21848 27712 21876
rect 27706 21836 27712 21848
rect 27764 21836 27770 21888
rect 1104 21786 28888 21808
rect 1104 21734 10214 21786
rect 10266 21734 10278 21786
rect 10330 21734 10342 21786
rect 10394 21734 10406 21786
rect 10458 21734 10470 21786
rect 10522 21734 19478 21786
rect 19530 21734 19542 21786
rect 19594 21734 19606 21786
rect 19658 21734 19670 21786
rect 19722 21734 19734 21786
rect 19786 21734 28888 21786
rect 1104 21712 28888 21734
rect 11882 21632 11888 21684
rect 11940 21672 11946 21684
rect 16022 21672 16028 21684
rect 11940 21644 16028 21672
rect 11940 21632 11946 21644
rect 16022 21632 16028 21644
rect 16080 21632 16086 21684
rect 16945 21675 17003 21681
rect 16945 21641 16957 21675
rect 16991 21672 17003 21675
rect 17310 21672 17316 21684
rect 16991 21644 17316 21672
rect 16991 21641 17003 21644
rect 16945 21635 17003 21641
rect 17310 21632 17316 21644
rect 17368 21632 17374 21684
rect 17494 21632 17500 21684
rect 17552 21672 17558 21684
rect 18509 21675 18567 21681
rect 17552 21644 18460 21672
rect 17552 21632 17558 21644
rect 12342 21604 12348 21616
rect 11992 21576 12348 21604
rect 11790 21536 11796 21548
rect 11751 21508 11796 21536
rect 11790 21496 11796 21508
rect 11848 21496 11854 21548
rect 11992 21545 12020 21576
rect 12342 21564 12348 21576
rect 12400 21564 12406 21616
rect 13357 21607 13415 21613
rect 13357 21604 13369 21607
rect 12452 21576 13369 21604
rect 12452 21545 12480 21576
rect 13357 21573 13369 21576
rect 13403 21604 13415 21607
rect 13722 21604 13728 21616
rect 13403 21576 13728 21604
rect 13403 21573 13415 21576
rect 13357 21567 13415 21573
rect 13722 21564 13728 21576
rect 13780 21564 13786 21616
rect 14093 21607 14151 21613
rect 14093 21573 14105 21607
rect 14139 21604 14151 21607
rect 15102 21604 15108 21616
rect 14139 21576 15108 21604
rect 14139 21573 14151 21576
rect 14093 21567 14151 21573
rect 11977 21539 12035 21545
rect 11977 21505 11989 21539
rect 12023 21505 12035 21539
rect 11977 21499 12035 21505
rect 12437 21539 12495 21545
rect 12437 21505 12449 21539
rect 12483 21505 12495 21539
rect 12437 21499 12495 21505
rect 12621 21539 12679 21545
rect 12621 21505 12633 21539
rect 12667 21505 12679 21539
rect 12621 21499 12679 21505
rect 13173 21539 13231 21545
rect 13173 21505 13185 21539
rect 13219 21536 13231 21539
rect 13630 21536 13636 21548
rect 13219 21508 13636 21536
rect 13219 21505 13231 21508
rect 13173 21499 13231 21505
rect 11885 21471 11943 21477
rect 11885 21437 11897 21471
rect 11931 21468 11943 21471
rect 12250 21468 12256 21480
rect 11931 21440 12256 21468
rect 11931 21437 11943 21440
rect 11885 21431 11943 21437
rect 12250 21428 12256 21440
rect 12308 21428 12314 21480
rect 12636 21468 12664 21499
rect 13630 21496 13636 21508
rect 13688 21496 13694 21548
rect 13906 21496 13912 21548
rect 13964 21536 13970 21548
rect 14936 21545 14964 21576
rect 15102 21564 15108 21576
rect 15160 21564 15166 21616
rect 15378 21564 15384 21616
rect 15436 21604 15442 21616
rect 15657 21607 15715 21613
rect 15657 21604 15669 21607
rect 15436 21576 15669 21604
rect 15436 21564 15442 21576
rect 15657 21573 15669 21576
rect 15703 21573 15715 21607
rect 15657 21567 15715 21573
rect 15841 21607 15899 21613
rect 15841 21573 15853 21607
rect 15887 21604 15899 21607
rect 15930 21604 15936 21616
rect 15887 21576 15936 21604
rect 15887 21573 15899 21576
rect 15841 21567 15899 21573
rect 15930 21564 15936 21576
rect 15988 21564 15994 21616
rect 17328 21576 18184 21604
rect 14829 21539 14887 21545
rect 13964 21508 14009 21536
rect 14829 21526 14841 21539
rect 13964 21496 13970 21508
rect 14752 21505 14841 21526
rect 14875 21505 14887 21539
rect 14752 21499 14887 21505
rect 14921 21539 14979 21545
rect 14921 21505 14933 21539
rect 14967 21505 14979 21539
rect 14921 21499 14979 21505
rect 15013 21539 15071 21545
rect 15013 21505 15025 21539
rect 15059 21536 15071 21539
rect 15197 21539 15255 21545
rect 15059 21508 15148 21536
rect 15059 21505 15071 21508
rect 15013 21499 15071 21505
rect 14752 21498 14872 21499
rect 12894 21468 12900 21480
rect 12636 21440 12900 21468
rect 12894 21428 12900 21440
rect 12952 21428 12958 21480
rect 12529 21403 12587 21409
rect 12529 21369 12541 21403
rect 12575 21400 12587 21403
rect 14642 21400 14648 21412
rect 12575 21372 14648 21400
rect 12575 21369 12587 21372
rect 12529 21363 12587 21369
rect 14642 21360 14648 21372
rect 14700 21360 14706 21412
rect 14752 21344 14780 21498
rect 15120 21468 15148 21508
rect 15197 21505 15209 21539
rect 15243 21536 15255 21539
rect 16114 21536 16120 21548
rect 15243 21508 16120 21536
rect 15243 21505 15255 21508
rect 15197 21499 15255 21505
rect 16114 21496 16120 21508
rect 16172 21496 16178 21548
rect 16482 21496 16488 21548
rect 16540 21536 16546 21548
rect 17121 21542 17179 21545
rect 17328 21542 17356 21576
rect 18156 21548 18184 21576
rect 17121 21539 17356 21542
rect 16540 21508 16896 21536
rect 16540 21496 16546 21508
rect 15470 21468 15476 21480
rect 15120 21440 15476 21468
rect 15470 21428 15476 21440
rect 15528 21428 15534 21480
rect 16868 21468 16896 21508
rect 17121 21505 17133 21539
rect 17167 21514 17356 21539
rect 17405 21539 17463 21545
rect 17167 21505 17179 21514
rect 17121 21499 17179 21505
rect 17405 21505 17417 21539
rect 17451 21536 17463 21539
rect 17678 21536 17684 21548
rect 17451 21508 17684 21536
rect 17451 21505 17463 21508
rect 17405 21499 17463 21505
rect 17678 21496 17684 21508
rect 17736 21496 17742 21548
rect 18138 21536 18144 21548
rect 18099 21508 18144 21536
rect 18138 21496 18144 21508
rect 18196 21496 18202 21548
rect 18432 21536 18460 21644
rect 18509 21641 18521 21675
rect 18555 21641 18567 21675
rect 18509 21635 18567 21641
rect 18524 21604 18552 21635
rect 18874 21632 18880 21684
rect 18932 21672 18938 21684
rect 19061 21675 19119 21681
rect 19061 21672 19073 21675
rect 18932 21644 19073 21672
rect 18932 21632 18938 21644
rect 19061 21641 19073 21644
rect 19107 21641 19119 21675
rect 19061 21635 19119 21641
rect 19150 21632 19156 21684
rect 19208 21672 19214 21684
rect 21358 21672 21364 21684
rect 19208 21644 21364 21672
rect 19208 21632 19214 21644
rect 21358 21632 21364 21644
rect 21416 21632 21422 21684
rect 22002 21632 22008 21684
rect 22060 21672 22066 21684
rect 23658 21672 23664 21684
rect 22060 21644 23664 21672
rect 22060 21632 22066 21644
rect 23658 21632 23664 21644
rect 23716 21632 23722 21684
rect 24026 21632 24032 21684
rect 24084 21672 24090 21684
rect 24762 21672 24768 21684
rect 24084 21644 24768 21672
rect 24084 21632 24090 21644
rect 24762 21632 24768 21644
rect 24820 21632 24826 21684
rect 26970 21672 26976 21684
rect 26931 21644 26976 21672
rect 26970 21632 26976 21644
rect 27028 21632 27034 21684
rect 18969 21607 19027 21613
rect 18969 21604 18981 21607
rect 18524 21576 18981 21604
rect 18969 21573 18981 21576
rect 19015 21573 19027 21607
rect 18969 21567 19027 21573
rect 19352 21576 19625 21604
rect 19352 21539 19380 21576
rect 19306 21536 19380 21539
rect 18432 21511 19380 21536
rect 19597 21536 19625 21576
rect 20254 21564 20260 21616
rect 20312 21604 20318 21616
rect 20349 21607 20407 21613
rect 20349 21604 20361 21607
rect 20312 21576 20361 21604
rect 20312 21564 20318 21576
rect 20349 21573 20361 21576
rect 20395 21573 20407 21607
rect 20349 21567 20407 21573
rect 20438 21564 20444 21616
rect 20496 21604 20502 21616
rect 20549 21607 20607 21613
rect 20549 21604 20561 21607
rect 20496 21576 20561 21604
rect 20496 21564 20502 21576
rect 20549 21573 20561 21576
rect 20595 21573 20607 21607
rect 20549 21567 20607 21573
rect 21266 21564 21272 21616
rect 21324 21604 21330 21616
rect 21726 21604 21732 21616
rect 21324 21576 21732 21604
rect 21324 21564 21330 21576
rect 21726 21564 21732 21576
rect 21784 21604 21790 21616
rect 25038 21604 25044 21616
rect 21784 21576 25044 21604
rect 21784 21564 21790 21576
rect 21821 21539 21879 21545
rect 21821 21536 21833 21539
rect 18432 21508 19334 21511
rect 19597 21508 21833 21536
rect 21821 21505 21833 21508
rect 21867 21505 21879 21539
rect 21821 21499 21879 21505
rect 21910 21496 21916 21548
rect 21968 21536 21974 21548
rect 22005 21539 22063 21545
rect 22005 21536 22017 21539
rect 21968 21508 22017 21536
rect 21968 21496 21974 21508
rect 22005 21505 22017 21508
rect 22051 21505 22063 21539
rect 22005 21499 22063 21505
rect 22189 21539 22247 21545
rect 22189 21505 22201 21539
rect 22235 21505 22247 21539
rect 22189 21499 22247 21505
rect 22281 21539 22339 21545
rect 22281 21505 22293 21539
rect 22327 21536 22339 21539
rect 22370 21536 22376 21548
rect 22327 21508 22376 21536
rect 22327 21505 22339 21508
rect 22281 21499 22339 21505
rect 17221 21471 17279 21477
rect 16868 21452 17080 21468
rect 17221 21452 17233 21471
rect 16868 21440 17233 21452
rect 17052 21437 17233 21440
rect 17267 21437 17279 21471
rect 17052 21431 17279 21437
rect 17052 21424 17264 21431
rect 17310 21428 17316 21480
rect 17368 21468 17374 21480
rect 17368 21440 17413 21468
rect 17368 21428 17374 21440
rect 17954 21428 17960 21480
rect 18012 21468 18018 21480
rect 18049 21471 18107 21477
rect 18049 21468 18061 21471
rect 18012 21440 18061 21468
rect 18012 21428 18018 21440
rect 18049 21437 18061 21440
rect 18095 21437 18107 21471
rect 18049 21431 18107 21437
rect 19337 21471 19395 21477
rect 19337 21437 19349 21471
rect 19383 21468 19395 21471
rect 20070 21468 20076 21480
rect 19383 21440 20076 21468
rect 19383 21437 19395 21440
rect 19337 21431 19395 21437
rect 20070 21428 20076 21440
rect 20128 21468 20134 21480
rect 20714 21468 20720 21480
rect 20128 21440 20720 21468
rect 20128 21428 20134 21440
rect 20714 21428 20720 21440
rect 20772 21428 20778 21480
rect 21082 21428 21088 21480
rect 21140 21468 21146 21480
rect 22204 21468 22232 21499
rect 22370 21496 22376 21508
rect 22428 21496 22434 21548
rect 22664 21536 22692 21576
rect 25038 21564 25044 21576
rect 25096 21564 25102 21616
rect 27338 21564 27344 21616
rect 27396 21604 27402 21616
rect 28077 21607 28135 21613
rect 28077 21604 28089 21607
rect 27396 21576 28089 21604
rect 27396 21564 27402 21576
rect 28077 21573 28089 21576
rect 28123 21573 28135 21607
rect 28077 21567 28135 21573
rect 22741 21539 22799 21545
rect 22741 21536 22753 21539
rect 22664 21508 22753 21536
rect 22741 21505 22753 21508
rect 22787 21505 22799 21539
rect 22741 21499 22799 21505
rect 22830 21496 22836 21548
rect 22888 21496 22894 21548
rect 23014 21545 23020 21548
rect 23008 21536 23020 21545
rect 22975 21508 23020 21536
rect 23008 21499 23020 21508
rect 23014 21496 23020 21499
rect 23072 21496 23078 21548
rect 27157 21539 27215 21545
rect 27157 21536 27169 21539
rect 25976 21508 27169 21536
rect 22646 21468 22652 21480
rect 21140 21440 22652 21468
rect 21140 21428 21146 21440
rect 22646 21428 22652 21440
rect 22704 21428 22710 21480
rect 22848 21468 22876 21496
rect 22756 21440 22876 21468
rect 24581 21471 24639 21477
rect 14918 21360 14924 21412
rect 14976 21400 14982 21412
rect 16758 21400 16764 21412
rect 14976 21372 16764 21400
rect 14976 21360 14982 21372
rect 16758 21360 16764 21372
rect 16816 21360 16822 21412
rect 18506 21360 18512 21412
rect 18564 21400 18570 21412
rect 18564 21372 21487 21400
rect 18564 21360 18570 21372
rect 14550 21332 14556 21344
rect 14511 21304 14556 21332
rect 14550 21292 14556 21304
rect 14608 21292 14614 21344
rect 14734 21292 14740 21344
rect 14792 21292 14798 21344
rect 15194 21292 15200 21344
rect 15252 21332 15258 21344
rect 16025 21335 16083 21341
rect 16025 21332 16037 21335
rect 15252 21304 16037 21332
rect 15252 21292 15258 21304
rect 16025 21301 16037 21304
rect 16071 21301 16083 21335
rect 16025 21295 16083 21301
rect 16298 21292 16304 21344
rect 16356 21332 16362 21344
rect 19245 21335 19303 21341
rect 19245 21332 19257 21335
rect 16356 21304 19257 21332
rect 16356 21292 16362 21304
rect 19245 21301 19257 21304
rect 19291 21301 19303 21335
rect 19245 21295 19303 21301
rect 19334 21292 19340 21344
rect 19392 21332 19398 21344
rect 19392 21304 19437 21332
rect 19392 21292 19398 21304
rect 20346 21292 20352 21344
rect 20404 21332 20410 21344
rect 20533 21335 20591 21341
rect 20533 21332 20545 21335
rect 20404 21304 20545 21332
rect 20404 21292 20410 21304
rect 20533 21301 20545 21304
rect 20579 21332 20591 21335
rect 20622 21332 20628 21344
rect 20579 21304 20628 21332
rect 20579 21301 20591 21304
rect 20533 21295 20591 21301
rect 20622 21292 20628 21304
rect 20680 21292 20686 21344
rect 20717 21335 20775 21341
rect 20717 21301 20729 21335
rect 20763 21332 20775 21335
rect 20806 21332 20812 21344
rect 20763 21304 20812 21332
rect 20763 21301 20775 21304
rect 20717 21295 20775 21301
rect 20806 21292 20812 21304
rect 20864 21332 20870 21344
rect 21358 21332 21364 21344
rect 20864 21304 21364 21332
rect 20864 21292 20870 21304
rect 21358 21292 21364 21304
rect 21416 21292 21422 21344
rect 21459 21332 21487 21372
rect 22186 21360 22192 21412
rect 22244 21400 22250 21412
rect 22370 21400 22376 21412
rect 22244 21372 22376 21400
rect 22244 21360 22250 21372
rect 22370 21360 22376 21372
rect 22428 21400 22434 21412
rect 22756 21400 22784 21440
rect 24581 21437 24593 21471
rect 24627 21437 24639 21471
rect 24762 21468 24768 21480
rect 24723 21440 24768 21468
rect 24581 21431 24639 21437
rect 24596 21400 24624 21431
rect 24762 21428 24768 21440
rect 24820 21428 24826 21480
rect 25222 21428 25228 21480
rect 25280 21468 25286 21480
rect 25976 21468 26004 21508
rect 27157 21505 27169 21508
rect 27203 21505 27215 21539
rect 27890 21536 27896 21548
rect 27851 21508 27896 21536
rect 27157 21499 27215 21505
rect 27890 21496 27896 21508
rect 27948 21496 27954 21548
rect 28169 21539 28227 21545
rect 28169 21505 28181 21539
rect 28215 21505 28227 21539
rect 28169 21499 28227 21505
rect 26142 21468 26148 21480
rect 25280 21440 26004 21468
rect 26103 21440 26148 21468
rect 25280 21428 25286 21440
rect 26142 21428 26148 21440
rect 26200 21428 26206 21480
rect 26234 21428 26240 21480
rect 26292 21468 26298 21480
rect 27246 21468 27252 21480
rect 26292 21440 27252 21468
rect 26292 21428 26298 21440
rect 27246 21428 27252 21440
rect 27304 21468 27310 21480
rect 27433 21471 27491 21477
rect 27433 21468 27445 21471
rect 27304 21440 27445 21468
rect 27304 21428 27310 21440
rect 27433 21437 27445 21440
rect 27479 21437 27491 21471
rect 27433 21431 27491 21437
rect 22428 21372 22784 21400
rect 23673 21372 24624 21400
rect 22428 21360 22434 21372
rect 23673 21332 23701 21372
rect 27062 21360 27068 21412
rect 27120 21400 27126 21412
rect 28184 21400 28212 21499
rect 27120 21372 28212 21400
rect 27120 21360 27126 21372
rect 21459 21304 23701 21332
rect 23750 21292 23756 21344
rect 23808 21332 23814 21344
rect 24121 21335 24179 21341
rect 24121 21332 24133 21335
rect 23808 21304 24133 21332
rect 23808 21292 23814 21304
rect 24121 21301 24133 21304
rect 24167 21301 24179 21335
rect 24121 21295 24179 21301
rect 24854 21292 24860 21344
rect 24912 21332 24918 21344
rect 27246 21332 27252 21344
rect 24912 21304 27252 21332
rect 24912 21292 24918 21304
rect 27246 21292 27252 21304
rect 27304 21332 27310 21344
rect 27341 21335 27399 21341
rect 27341 21332 27353 21335
rect 27304 21304 27353 21332
rect 27304 21292 27310 21304
rect 27341 21301 27353 21304
rect 27387 21301 27399 21335
rect 27341 21295 27399 21301
rect 27614 21292 27620 21344
rect 27672 21332 27678 21344
rect 27893 21335 27951 21341
rect 27893 21332 27905 21335
rect 27672 21304 27905 21332
rect 27672 21292 27678 21304
rect 27893 21301 27905 21304
rect 27939 21301 27951 21335
rect 27893 21295 27951 21301
rect 1104 21242 28888 21264
rect 1104 21190 5582 21242
rect 5634 21190 5646 21242
rect 5698 21190 5710 21242
rect 5762 21190 5774 21242
rect 5826 21190 5838 21242
rect 5890 21190 14846 21242
rect 14898 21190 14910 21242
rect 14962 21190 14974 21242
rect 15026 21190 15038 21242
rect 15090 21190 15102 21242
rect 15154 21190 24110 21242
rect 24162 21190 24174 21242
rect 24226 21190 24238 21242
rect 24290 21190 24302 21242
rect 24354 21190 24366 21242
rect 24418 21190 28888 21242
rect 1104 21168 28888 21190
rect 13170 21088 13176 21140
rect 13228 21128 13234 21140
rect 13357 21131 13415 21137
rect 13357 21128 13369 21131
rect 13228 21100 13369 21128
rect 13228 21088 13234 21100
rect 13357 21097 13369 21100
rect 13403 21097 13415 21131
rect 13906 21128 13912 21140
rect 13357 21091 13415 21097
rect 13464 21100 13912 21128
rect 12066 21060 12072 21072
rect 12027 21032 12072 21060
rect 12066 21020 12072 21032
rect 12124 21020 12130 21072
rect 11790 20952 11796 21004
rect 11848 20992 11854 21004
rect 13464 20992 13492 21100
rect 13906 21088 13912 21100
rect 13964 21128 13970 21140
rect 15470 21128 15476 21140
rect 13964 21100 14872 21128
rect 15431 21100 15476 21128
rect 13964 21088 13970 21100
rect 14090 21060 14096 21072
rect 14051 21032 14096 21060
rect 14090 21020 14096 21032
rect 14148 21020 14154 21072
rect 11848 20964 13492 20992
rect 11848 20952 11854 20964
rect 12084 20933 12112 20964
rect 13630 20952 13636 21004
rect 13688 20952 13694 21004
rect 13998 20952 14004 21004
rect 14056 20992 14062 21004
rect 14550 20992 14556 21004
rect 14056 20964 14556 20992
rect 14056 20952 14062 20964
rect 14550 20952 14556 20964
rect 14608 20952 14614 21004
rect 14844 21001 14872 21100
rect 15470 21088 15476 21100
rect 15528 21088 15534 21140
rect 15654 21128 15660 21140
rect 15580 21100 15660 21128
rect 14829 20995 14887 21001
rect 14829 20961 14841 20995
rect 14875 20961 14887 20995
rect 15194 20992 15200 21004
rect 15155 20964 15200 20992
rect 14829 20955 14887 20961
rect 15194 20952 15200 20964
rect 15252 20952 15258 21004
rect 15289 20995 15347 21001
rect 15289 20961 15301 20995
rect 15335 20992 15347 20995
rect 15580 20992 15608 21100
rect 15654 21088 15660 21100
rect 15712 21088 15718 21140
rect 15838 21088 15844 21140
rect 15896 21128 15902 21140
rect 19886 21128 19892 21140
rect 15896 21100 19892 21128
rect 15896 21088 15902 21100
rect 19886 21088 19892 21100
rect 19944 21088 19950 21140
rect 20162 21128 20168 21140
rect 20123 21100 20168 21128
rect 20162 21088 20168 21100
rect 20220 21088 20226 21140
rect 22002 21128 22008 21140
rect 20640 21100 22008 21128
rect 16114 21020 16120 21072
rect 16172 21060 16178 21072
rect 16172 21032 17908 21060
rect 16172 21020 16178 21032
rect 15335 20964 15608 20992
rect 15335 20961 15347 20964
rect 15289 20955 15347 20961
rect 12069 20927 12127 20933
rect 12069 20893 12081 20927
rect 12115 20893 12127 20927
rect 12069 20887 12127 20893
rect 12253 20927 12311 20933
rect 12253 20893 12265 20927
rect 12299 20924 12311 20927
rect 12713 20927 12771 20933
rect 12299 20896 12434 20924
rect 12299 20893 12311 20896
rect 12253 20887 12311 20893
rect 12406 20868 12434 20896
rect 12713 20893 12725 20927
rect 12759 20893 12771 20927
rect 12713 20887 12771 20893
rect 12897 20927 12955 20933
rect 12897 20893 12909 20927
rect 12943 20924 12955 20927
rect 13078 20924 13084 20936
rect 12943 20896 13084 20924
rect 12943 20893 12955 20896
rect 12897 20887 12955 20893
rect 12406 20828 12440 20868
rect 12434 20816 12440 20828
rect 12492 20816 12498 20868
rect 9858 20748 9864 20800
rect 9916 20788 9922 20800
rect 12618 20788 12624 20800
rect 9916 20760 12624 20788
rect 9916 20748 9922 20760
rect 12618 20748 12624 20760
rect 12676 20748 12682 20800
rect 12728 20788 12756 20887
rect 13078 20884 13084 20896
rect 13136 20884 13142 20936
rect 13262 20884 13268 20936
rect 13320 20924 13326 20936
rect 13357 20927 13415 20933
rect 13357 20924 13369 20927
rect 13320 20896 13369 20924
rect 13320 20884 13326 20896
rect 13357 20893 13369 20896
rect 13403 20893 13415 20927
rect 13357 20887 13415 20893
rect 13535 20927 13593 20933
rect 13535 20893 13547 20927
rect 13581 20921 13593 20927
rect 13648 20921 13676 20952
rect 14369 20927 14427 20933
rect 14369 20924 14381 20927
rect 13581 20893 13676 20921
rect 14016 20896 14381 20924
rect 13535 20887 13593 20893
rect 12805 20859 12863 20865
rect 12805 20825 12817 20859
rect 12851 20856 12863 20859
rect 14016 20856 14044 20896
rect 14369 20893 14381 20896
rect 14415 20924 14427 20927
rect 15304 20924 15332 20955
rect 16022 20952 16028 21004
rect 16080 20992 16086 21004
rect 16206 20992 16212 21004
rect 16080 20964 16212 20992
rect 16080 20952 16086 20964
rect 16206 20952 16212 20964
rect 16264 20992 16270 21004
rect 16264 20964 16620 20992
rect 16264 20952 16270 20964
rect 16592 20933 16620 20964
rect 16868 20933 16896 21032
rect 16942 20952 16948 21004
rect 17000 20992 17006 21004
rect 17310 20992 17316 21004
rect 17000 20964 17316 20992
rect 17000 20952 17006 20964
rect 17310 20952 17316 20964
rect 17368 20952 17374 21004
rect 17770 20992 17776 21004
rect 17731 20964 17776 20992
rect 17770 20952 17776 20964
rect 17828 20952 17834 21004
rect 17880 20992 17908 21032
rect 18046 21020 18052 21072
rect 18104 21060 18110 21072
rect 20640 21060 20668 21100
rect 22002 21088 22008 21100
rect 22060 21088 22066 21140
rect 22646 21088 22652 21140
rect 22704 21128 22710 21140
rect 23474 21128 23480 21140
rect 22704 21100 23480 21128
rect 22704 21088 22710 21100
rect 23474 21088 23480 21100
rect 23532 21088 23538 21140
rect 23658 21088 23664 21140
rect 23716 21128 23722 21140
rect 25501 21131 25559 21137
rect 23716 21100 25268 21128
rect 23716 21088 23722 21100
rect 18104 21032 20668 21060
rect 25240 21060 25268 21100
rect 25501 21097 25513 21131
rect 25547 21128 25559 21131
rect 25682 21128 25688 21140
rect 25547 21100 25688 21128
rect 25547 21097 25559 21100
rect 25501 21091 25559 21097
rect 25682 21088 25688 21100
rect 25740 21088 25746 21140
rect 27430 21060 27436 21072
rect 25240 21032 27436 21060
rect 18104 21020 18110 21032
rect 27430 21020 27436 21032
rect 27488 21020 27494 21072
rect 18690 20992 18696 21004
rect 17880 20964 18696 20992
rect 18690 20952 18696 20964
rect 18748 20952 18754 21004
rect 19242 20952 19248 21004
rect 19300 20992 19306 21004
rect 23474 20992 23480 21004
rect 19300 20964 19932 20992
rect 19300 20952 19306 20964
rect 14415 20896 15332 20924
rect 16485 20927 16543 20933
rect 14415 20893 14427 20896
rect 14369 20887 14427 20893
rect 16485 20893 16497 20927
rect 16531 20893 16543 20927
rect 16485 20887 16543 20893
rect 16577 20927 16635 20933
rect 16577 20893 16589 20927
rect 16623 20893 16635 20927
rect 16669 20927 16727 20933
rect 16669 20914 16681 20927
rect 16715 20914 16727 20927
rect 16853 20927 16911 20933
rect 16577 20887 16635 20893
rect 12851 20828 14044 20856
rect 14093 20859 14151 20865
rect 12851 20825 12863 20828
rect 12805 20819 12863 20825
rect 14093 20825 14105 20859
rect 14139 20825 14151 20859
rect 14093 20819 14151 20825
rect 14277 20859 14335 20865
rect 14277 20825 14289 20859
rect 14323 20856 14335 20859
rect 14642 20856 14648 20868
rect 14323 20828 14648 20856
rect 14323 20825 14335 20828
rect 14277 20819 14335 20825
rect 13906 20788 13912 20800
rect 12728 20760 13912 20788
rect 13906 20748 13912 20760
rect 13964 20748 13970 20800
rect 14108 20788 14136 20819
rect 14642 20816 14648 20828
rect 14700 20816 14706 20868
rect 15286 20856 15292 20868
rect 14752 20828 15292 20856
rect 14550 20788 14556 20800
rect 14108 20760 14556 20788
rect 14550 20748 14556 20760
rect 14608 20788 14614 20800
rect 14752 20788 14780 20828
rect 15286 20816 15292 20828
rect 15344 20816 15350 20868
rect 15378 20816 15384 20868
rect 15436 20856 15442 20868
rect 15654 20856 15660 20868
rect 15436 20828 15660 20856
rect 15436 20816 15442 20828
rect 15654 20816 15660 20828
rect 15712 20816 15718 20868
rect 16298 20856 16304 20868
rect 15941 20828 16304 20856
rect 14608 20760 14780 20788
rect 14608 20748 14614 20760
rect 14826 20748 14832 20800
rect 14884 20788 14890 20800
rect 15941 20788 15969 20828
rect 16298 20816 16304 20828
rect 16356 20816 16362 20868
rect 16206 20788 16212 20800
rect 14884 20760 15969 20788
rect 16167 20760 16212 20788
rect 14884 20748 14890 20760
rect 16206 20748 16212 20760
rect 16264 20748 16270 20800
rect 16500 20788 16528 20887
rect 16666 20862 16672 20914
rect 16724 20862 16730 20914
rect 16853 20893 16865 20927
rect 16899 20893 16911 20927
rect 17678 20924 17684 20936
rect 17591 20896 17684 20924
rect 16853 20887 16911 20893
rect 17678 20884 17684 20896
rect 17736 20924 17742 20936
rect 17862 20924 17868 20936
rect 17736 20896 17868 20924
rect 17736 20884 17742 20896
rect 17862 20884 17868 20896
rect 17920 20884 17926 20936
rect 17954 20884 17960 20936
rect 18012 20924 18018 20936
rect 18509 20927 18567 20933
rect 18012 20896 18057 20924
rect 18012 20884 18018 20896
rect 18509 20893 18521 20927
rect 18555 20924 18567 20927
rect 18966 20924 18972 20936
rect 18555 20896 18972 20924
rect 18555 20893 18567 20896
rect 18509 20887 18567 20893
rect 18966 20884 18972 20896
rect 19024 20884 19030 20936
rect 19521 20927 19579 20933
rect 19521 20893 19533 20927
rect 19567 20893 19579 20927
rect 19521 20887 19579 20893
rect 17696 20856 17724 20884
rect 16776 20828 17724 20856
rect 16776 20788 16804 20828
rect 16500 20760 16804 20788
rect 17126 20748 17132 20800
rect 17184 20788 17190 20800
rect 17313 20791 17371 20797
rect 17313 20788 17325 20791
rect 17184 20760 17325 20788
rect 17184 20748 17190 20760
rect 17313 20757 17325 20760
rect 17359 20757 17371 20791
rect 17313 20751 17371 20757
rect 18506 20748 18512 20800
rect 18564 20788 18570 20800
rect 18601 20791 18659 20797
rect 18601 20788 18613 20791
rect 18564 20760 18613 20788
rect 18564 20748 18570 20760
rect 18601 20757 18613 20760
rect 18647 20757 18659 20791
rect 19536 20788 19564 20887
rect 19610 20884 19616 20936
rect 19668 20924 19674 20936
rect 19904 20933 19932 20964
rect 22741 20965 22799 20971
rect 19889 20927 19947 20933
rect 19668 20896 19713 20924
rect 19668 20884 19674 20896
rect 19889 20893 19901 20927
rect 19935 20893 19947 20927
rect 19889 20887 19947 20893
rect 20027 20927 20085 20933
rect 20027 20893 20039 20927
rect 20073 20924 20085 20927
rect 20254 20924 20260 20936
rect 20073 20896 20260 20924
rect 20073 20893 20085 20896
rect 20027 20887 20085 20893
rect 20254 20884 20260 20896
rect 20312 20884 20318 20936
rect 20625 20927 20683 20933
rect 20625 20893 20637 20927
rect 20671 20924 20683 20927
rect 21266 20924 21272 20936
rect 20671 20896 21272 20924
rect 20671 20893 20683 20896
rect 20625 20887 20683 20893
rect 21266 20884 21272 20896
rect 21324 20884 21330 20936
rect 22370 20884 22376 20936
rect 22428 20924 22434 20936
rect 22465 20927 22523 20933
rect 22465 20924 22477 20927
rect 22428 20896 22477 20924
rect 22428 20884 22434 20896
rect 22465 20893 22477 20896
rect 22511 20893 22523 20927
rect 22465 20887 22523 20893
rect 22554 20884 22560 20936
rect 22612 20924 22618 20936
rect 22741 20931 22753 20965
rect 22787 20931 22799 20965
rect 23400 20964 23480 20992
rect 23400 20933 23428 20964
rect 23474 20952 23480 20964
rect 23532 20952 23538 21004
rect 25222 20992 25228 21004
rect 22741 20925 22799 20931
rect 23385 20927 23443 20933
rect 22612 20896 22657 20924
rect 22612 20884 22618 20896
rect 19797 20859 19855 20865
rect 19797 20825 19809 20859
rect 19843 20856 19855 20859
rect 20346 20856 20352 20868
rect 19843 20828 20352 20856
rect 19843 20825 19855 20828
rect 19797 20819 19855 20825
rect 20346 20816 20352 20828
rect 20404 20816 20410 20868
rect 20898 20865 20904 20868
rect 20892 20819 20904 20865
rect 20956 20856 20962 20868
rect 22756 20856 22784 20925
rect 23385 20893 23397 20927
rect 23431 20893 23443 20927
rect 23566 20924 23572 20936
rect 23527 20896 23572 20924
rect 23385 20887 23443 20893
rect 23566 20884 23572 20896
rect 23624 20884 23630 20936
rect 23658 20922 23664 20974
rect 23716 20922 23722 20974
rect 25183 20964 25228 20992
rect 25222 20952 25228 20964
rect 25280 20952 25286 21004
rect 26513 20995 26571 21001
rect 26513 20961 26525 20995
rect 26559 20992 26571 20995
rect 27522 20992 27528 21004
rect 26559 20964 27528 20992
rect 26559 20961 26571 20964
rect 26513 20955 26571 20961
rect 27522 20952 27528 20964
rect 27580 20952 27586 21004
rect 28166 20992 28172 21004
rect 28127 20964 28172 20992
rect 28166 20952 28172 20964
rect 28224 20952 28230 21004
rect 25130 20924 25136 20936
rect 23658 20903 23670 20922
rect 23704 20903 23716 20922
rect 23658 20897 23716 20903
rect 25091 20896 25136 20924
rect 25130 20884 25136 20896
rect 25188 20924 25194 20936
rect 26234 20924 26240 20936
rect 25188 20896 26240 20924
rect 25188 20884 25194 20896
rect 26234 20884 26240 20896
rect 26292 20884 26298 20936
rect 26329 20927 26387 20933
rect 26329 20893 26341 20927
rect 26375 20893 26387 20927
rect 26329 20887 26387 20893
rect 23201 20859 23259 20865
rect 20956 20828 20992 20856
rect 22756 20828 22876 20856
rect 20898 20816 20904 20819
rect 20956 20816 20962 20828
rect 20070 20788 20076 20800
rect 19536 20760 20076 20788
rect 18601 20751 18659 20757
rect 20070 20748 20076 20760
rect 20128 20748 20134 20800
rect 20254 20748 20260 20800
rect 20312 20788 20318 20800
rect 22005 20791 22063 20797
rect 22005 20788 22017 20791
rect 20312 20760 22017 20788
rect 20312 20748 20318 20760
rect 22005 20757 22017 20760
rect 22051 20757 22063 20791
rect 22738 20788 22744 20800
rect 22699 20760 22744 20788
rect 22005 20751 22063 20757
rect 22738 20748 22744 20760
rect 22796 20748 22802 20800
rect 22848 20788 22876 20828
rect 23201 20825 23213 20859
rect 23247 20856 23259 20859
rect 24578 20856 24584 20868
rect 23247 20828 24584 20856
rect 23247 20825 23259 20828
rect 23201 20819 23259 20825
rect 24578 20816 24584 20828
rect 24636 20816 24642 20868
rect 26344 20856 26372 20887
rect 26786 20856 26792 20868
rect 26344 20828 26792 20856
rect 26786 20816 26792 20828
rect 26844 20816 26850 20868
rect 26050 20788 26056 20800
rect 22848 20760 26056 20788
rect 26050 20748 26056 20760
rect 26108 20748 26114 20800
rect 1104 20698 28888 20720
rect 1104 20646 10214 20698
rect 10266 20646 10278 20698
rect 10330 20646 10342 20698
rect 10394 20646 10406 20698
rect 10458 20646 10470 20698
rect 10522 20646 19478 20698
rect 19530 20646 19542 20698
rect 19594 20646 19606 20698
rect 19658 20646 19670 20698
rect 19722 20646 19734 20698
rect 19786 20646 28888 20698
rect 1104 20624 28888 20646
rect 14090 20544 14096 20596
rect 14148 20584 14154 20596
rect 15378 20584 15384 20596
rect 14148 20556 15384 20584
rect 14148 20544 14154 20556
rect 15378 20544 15384 20556
rect 15436 20544 15442 20596
rect 16666 20544 16672 20596
rect 16724 20584 16730 20596
rect 17313 20587 17371 20593
rect 17313 20584 17325 20587
rect 16724 20556 17325 20584
rect 16724 20544 16730 20556
rect 17313 20553 17325 20556
rect 17359 20553 17371 20587
rect 17313 20547 17371 20553
rect 17862 20544 17868 20596
rect 17920 20584 17926 20596
rect 18230 20584 18236 20596
rect 17920 20556 18236 20584
rect 17920 20544 17926 20556
rect 18230 20544 18236 20556
rect 18288 20584 18294 20596
rect 19705 20587 19763 20593
rect 19705 20584 19717 20587
rect 18288 20556 19717 20584
rect 18288 20544 18294 20556
rect 19705 20553 19717 20556
rect 19751 20553 19763 20587
rect 19705 20547 19763 20553
rect 21177 20587 21235 20593
rect 21177 20553 21189 20587
rect 21223 20584 21235 20587
rect 23293 20587 23351 20593
rect 21223 20556 23244 20584
rect 21223 20553 21235 20556
rect 21177 20547 21235 20553
rect 15194 20516 15200 20528
rect 13372 20488 15200 20516
rect 13372 20457 13400 20488
rect 15194 20476 15200 20488
rect 15252 20476 15258 20528
rect 16022 20516 16028 20528
rect 15580 20488 16028 20516
rect 13357 20451 13415 20457
rect 13357 20417 13369 20451
rect 13403 20417 13415 20451
rect 13357 20411 13415 20417
rect 13624 20451 13682 20457
rect 13624 20417 13636 20451
rect 13670 20448 13682 20451
rect 13998 20448 14004 20460
rect 13670 20420 14004 20448
rect 13670 20417 13682 20420
rect 13624 20411 13682 20417
rect 13998 20408 14004 20420
rect 14056 20408 14062 20460
rect 15580 20457 15608 20488
rect 16022 20476 16028 20488
rect 16080 20476 16086 20528
rect 19426 20516 19432 20528
rect 18340 20488 19432 20516
rect 15473 20451 15531 20457
rect 15473 20417 15485 20451
rect 15519 20417 15531 20451
rect 15473 20411 15531 20417
rect 15565 20451 15623 20457
rect 15565 20417 15577 20451
rect 15611 20417 15623 20451
rect 15565 20411 15623 20417
rect 15657 20451 15715 20457
rect 15657 20417 15669 20451
rect 15703 20448 15715 20451
rect 15746 20448 15752 20460
rect 15703 20420 15752 20448
rect 15703 20417 15715 20420
rect 15657 20411 15715 20417
rect 14642 20340 14648 20392
rect 14700 20380 14706 20392
rect 15488 20380 15516 20411
rect 15746 20408 15752 20420
rect 15804 20408 15810 20460
rect 15841 20451 15899 20457
rect 15841 20417 15853 20451
rect 15887 20448 15899 20451
rect 16114 20448 16120 20460
rect 15887 20420 16120 20448
rect 15887 20417 15899 20420
rect 15841 20411 15899 20417
rect 16114 20408 16120 20420
rect 16172 20408 16178 20460
rect 16298 20408 16304 20460
rect 16356 20448 16362 20460
rect 18340 20457 18368 20488
rect 19426 20476 19432 20488
rect 19484 20476 19490 20528
rect 22830 20476 22836 20528
rect 22888 20516 22894 20528
rect 23017 20519 23075 20525
rect 23017 20516 23029 20519
rect 22888 20488 23029 20516
rect 22888 20476 22894 20488
rect 23017 20485 23029 20488
rect 23063 20485 23075 20519
rect 23216 20516 23244 20556
rect 23293 20553 23305 20587
rect 23339 20584 23351 20587
rect 23658 20584 23664 20596
rect 23339 20556 23664 20584
rect 23339 20553 23351 20556
rect 23293 20547 23351 20553
rect 23658 20544 23664 20556
rect 23716 20544 23722 20596
rect 25590 20584 25596 20596
rect 23768 20556 25596 20584
rect 23768 20516 23796 20556
rect 25590 20544 25596 20556
rect 25648 20544 25654 20596
rect 27617 20587 27675 20593
rect 27617 20553 27629 20587
rect 27663 20584 27675 20587
rect 27706 20584 27712 20596
rect 27663 20556 27712 20584
rect 27663 20553 27675 20556
rect 27617 20547 27675 20553
rect 27706 20544 27712 20556
rect 27764 20544 27770 20596
rect 23216 20488 23796 20516
rect 23017 20479 23075 20485
rect 25130 20476 25136 20528
rect 25188 20516 25194 20528
rect 26418 20516 26424 20528
rect 25188 20488 25636 20516
rect 25188 20476 25194 20488
rect 18325 20451 18383 20457
rect 18325 20448 18337 20451
rect 16356 20420 18337 20448
rect 16356 20408 16362 20420
rect 18325 20417 18337 20420
rect 18371 20417 18383 20451
rect 18325 20411 18383 20417
rect 18592 20451 18650 20457
rect 18592 20417 18604 20451
rect 18638 20448 18650 20451
rect 19334 20448 19340 20460
rect 18638 20420 19340 20448
rect 18638 20417 18650 20420
rect 18592 20411 18650 20417
rect 19334 20408 19340 20420
rect 19392 20408 19398 20460
rect 20349 20451 20407 20457
rect 20349 20448 20361 20451
rect 19444 20420 20361 20448
rect 14700 20352 15516 20380
rect 16669 20383 16727 20389
rect 14700 20340 14706 20352
rect 16669 20349 16681 20383
rect 16715 20380 16727 20383
rect 16850 20380 16856 20392
rect 16715 20352 16856 20380
rect 16715 20349 16727 20352
rect 16669 20343 16727 20349
rect 16850 20340 16856 20352
rect 16908 20340 16914 20392
rect 17034 20380 17040 20392
rect 16995 20352 17040 20380
rect 17034 20340 17040 20352
rect 17092 20340 17098 20392
rect 17126 20340 17132 20392
rect 17184 20380 17190 20392
rect 17184 20352 17229 20380
rect 17184 20340 17190 20352
rect 14734 20312 14740 20324
rect 14695 20284 14740 20312
rect 14734 20272 14740 20284
rect 14792 20272 14798 20324
rect 15120 20284 16436 20312
rect 13170 20204 13176 20256
rect 13228 20244 13234 20256
rect 15120 20244 15148 20284
rect 13228 20216 15148 20244
rect 15197 20247 15255 20253
rect 13228 20204 13234 20216
rect 15197 20213 15209 20247
rect 15243 20244 15255 20247
rect 15286 20244 15292 20256
rect 15243 20216 15292 20244
rect 15243 20213 15255 20216
rect 15197 20207 15255 20213
rect 15286 20204 15292 20216
rect 15344 20204 15350 20256
rect 16408 20244 16436 20284
rect 19444 20244 19472 20420
rect 20349 20417 20361 20420
rect 20395 20417 20407 20451
rect 20349 20411 20407 20417
rect 20530 20408 20536 20460
rect 20588 20448 20594 20460
rect 21082 20448 21088 20460
rect 20588 20420 21088 20448
rect 20588 20408 20594 20420
rect 21082 20408 21088 20420
rect 21140 20408 21146 20460
rect 22005 20451 22063 20457
rect 22005 20448 22017 20451
rect 21928 20420 22017 20448
rect 20622 20380 20628 20392
rect 20583 20352 20628 20380
rect 20622 20340 20628 20352
rect 20680 20380 20686 20392
rect 21821 20383 21879 20389
rect 21821 20380 21833 20383
rect 20680 20352 21833 20380
rect 20680 20340 20686 20352
rect 21821 20349 21833 20352
rect 21867 20349 21879 20383
rect 21821 20343 21879 20349
rect 21928 20312 21956 20420
rect 22005 20417 22017 20420
rect 22051 20417 22063 20451
rect 22738 20448 22744 20460
rect 22699 20420 22744 20448
rect 22005 20411 22063 20417
rect 22738 20408 22744 20420
rect 22796 20408 22802 20460
rect 22922 20448 22928 20460
rect 22883 20420 22928 20448
rect 22922 20408 22928 20420
rect 22980 20408 22986 20460
rect 23109 20451 23167 20457
rect 23109 20417 23121 20451
rect 23155 20417 23167 20451
rect 23109 20411 23167 20417
rect 23124 20380 23152 20411
rect 23934 20408 23940 20460
rect 23992 20448 23998 20460
rect 24489 20451 24547 20457
rect 24489 20448 24501 20451
rect 23992 20420 24501 20448
rect 23992 20408 23998 20420
rect 24489 20417 24501 20420
rect 24535 20417 24547 20451
rect 24489 20411 24547 20417
rect 24581 20451 24639 20457
rect 24581 20417 24593 20451
rect 24627 20417 24639 20451
rect 24581 20411 24639 20417
rect 24857 20451 24915 20457
rect 24857 20417 24869 20451
rect 24903 20448 24915 20451
rect 25314 20448 25320 20460
rect 24903 20420 25176 20448
rect 25275 20420 25320 20448
rect 24903 20417 24915 20420
rect 24857 20411 24915 20417
rect 23290 20380 23296 20392
rect 23124 20352 23296 20380
rect 23290 20340 23296 20352
rect 23348 20340 23354 20392
rect 23842 20340 23848 20392
rect 23900 20380 23906 20392
rect 24596 20380 24624 20411
rect 23900 20352 24624 20380
rect 23900 20340 23906 20352
rect 20548 20284 21956 20312
rect 20162 20244 20168 20256
rect 16408 20216 19472 20244
rect 20123 20216 20168 20244
rect 20162 20204 20168 20216
rect 20220 20204 20226 20256
rect 20438 20204 20444 20256
rect 20496 20244 20502 20256
rect 20548 20253 20576 20284
rect 22002 20272 22008 20324
rect 22060 20312 22066 20324
rect 22189 20315 22247 20321
rect 22189 20312 22201 20315
rect 22060 20284 22201 20312
rect 22060 20272 22066 20284
rect 22189 20281 22201 20284
rect 22235 20281 22247 20315
rect 25148 20312 25176 20420
rect 25314 20408 25320 20420
rect 25372 20408 25378 20460
rect 25608 20457 25636 20488
rect 25884 20488 26424 20516
rect 25884 20457 25912 20488
rect 26418 20476 26424 20488
rect 26476 20476 26482 20528
rect 26602 20476 26608 20528
rect 26660 20516 26666 20528
rect 27341 20519 27399 20525
rect 27341 20516 27353 20519
rect 26660 20488 27353 20516
rect 26660 20476 26666 20488
rect 27341 20485 27353 20488
rect 27387 20485 27399 20519
rect 27341 20479 27399 20485
rect 25501 20451 25559 20457
rect 25501 20417 25513 20451
rect 25547 20417 25559 20451
rect 25501 20411 25559 20417
rect 25593 20451 25651 20457
rect 25593 20417 25605 20451
rect 25639 20417 25651 20451
rect 25593 20411 25651 20417
rect 25869 20451 25927 20457
rect 25869 20417 25881 20451
rect 25915 20417 25927 20451
rect 25869 20411 25927 20417
rect 26053 20451 26111 20457
rect 26053 20417 26065 20451
rect 26099 20448 26111 20451
rect 26973 20451 27031 20457
rect 26973 20448 26985 20451
rect 26099 20420 26985 20448
rect 26099 20417 26111 20420
rect 26053 20411 26111 20417
rect 26973 20417 26985 20420
rect 27019 20417 27031 20451
rect 26973 20411 27031 20417
rect 27066 20451 27124 20457
rect 27066 20417 27078 20451
rect 27112 20417 27124 20451
rect 27249 20451 27307 20457
rect 27249 20448 27261 20451
rect 27066 20411 27124 20417
rect 27172 20420 27261 20448
rect 25222 20340 25228 20392
rect 25280 20380 25286 20392
rect 25516 20380 25544 20411
rect 25280 20352 25544 20380
rect 25280 20340 25286 20352
rect 25682 20340 25688 20392
rect 25740 20380 25746 20392
rect 25740 20352 26280 20380
rect 25740 20340 25746 20352
rect 25774 20312 25780 20324
rect 25148 20284 25780 20312
rect 22189 20275 22247 20281
rect 25774 20272 25780 20284
rect 25832 20272 25838 20324
rect 26252 20312 26280 20352
rect 26418 20340 26424 20392
rect 26476 20380 26482 20392
rect 27081 20380 27109 20411
rect 26476 20352 27109 20380
rect 26476 20340 26482 20352
rect 27172 20312 27200 20420
rect 27249 20417 27261 20420
rect 27295 20417 27307 20451
rect 27438 20451 27496 20457
rect 27438 20448 27450 20451
rect 27249 20411 27307 20417
rect 27356 20420 27450 20448
rect 26252 20284 27200 20312
rect 20533 20247 20591 20253
rect 20533 20244 20545 20247
rect 20496 20216 20545 20244
rect 20496 20204 20502 20216
rect 20533 20213 20545 20216
rect 20579 20213 20591 20247
rect 20533 20207 20591 20213
rect 21542 20204 21548 20256
rect 21600 20244 21606 20256
rect 24026 20244 24032 20256
rect 21600 20216 24032 20244
rect 21600 20204 21606 20216
rect 24026 20204 24032 20216
rect 24084 20204 24090 20256
rect 24305 20247 24363 20253
rect 24305 20213 24317 20247
rect 24351 20244 24363 20247
rect 24486 20244 24492 20256
rect 24351 20216 24492 20244
rect 24351 20213 24363 20216
rect 24305 20207 24363 20213
rect 24486 20204 24492 20216
rect 24544 20204 24550 20256
rect 24765 20247 24823 20253
rect 24765 20213 24777 20247
rect 24811 20244 24823 20247
rect 24946 20244 24952 20256
rect 24811 20216 24952 20244
rect 24811 20213 24823 20216
rect 24765 20207 24823 20213
rect 24946 20204 24952 20216
rect 25004 20204 25010 20256
rect 25866 20204 25872 20256
rect 25924 20244 25930 20256
rect 27356 20244 27384 20420
rect 27438 20417 27450 20420
rect 27484 20417 27496 20451
rect 27438 20411 27496 20417
rect 25924 20216 27384 20244
rect 25924 20204 25930 20216
rect 1104 20154 28888 20176
rect 1104 20102 5582 20154
rect 5634 20102 5646 20154
rect 5698 20102 5710 20154
rect 5762 20102 5774 20154
rect 5826 20102 5838 20154
rect 5890 20102 14846 20154
rect 14898 20102 14910 20154
rect 14962 20102 14974 20154
rect 15026 20102 15038 20154
rect 15090 20102 15102 20154
rect 15154 20102 24110 20154
rect 24162 20102 24174 20154
rect 24226 20102 24238 20154
rect 24290 20102 24302 20154
rect 24354 20102 24366 20154
rect 24418 20102 28888 20154
rect 1104 20080 28888 20102
rect 12894 20000 12900 20052
rect 12952 20040 12958 20052
rect 14553 20043 14611 20049
rect 14553 20040 14565 20043
rect 12952 20012 14565 20040
rect 12952 20000 12958 20012
rect 14553 20009 14565 20012
rect 14599 20040 14611 20043
rect 14734 20040 14740 20052
rect 14599 20012 14740 20040
rect 14599 20009 14611 20012
rect 14553 20003 14611 20009
rect 14734 20000 14740 20012
rect 14792 20000 14798 20052
rect 15470 20040 15476 20052
rect 15431 20012 15476 20040
rect 15470 20000 15476 20012
rect 15528 20000 15534 20052
rect 15657 20043 15715 20049
rect 15657 20009 15669 20043
rect 15703 20040 15715 20043
rect 15746 20040 15752 20052
rect 15703 20012 15752 20040
rect 15703 20009 15715 20012
rect 15657 20003 15715 20009
rect 15746 20000 15752 20012
rect 15804 20000 15810 20052
rect 17034 20040 17040 20052
rect 16316 20012 17040 20040
rect 13449 19975 13507 19981
rect 13449 19941 13461 19975
rect 13495 19972 13507 19975
rect 16316 19972 16344 20012
rect 17034 20000 17040 20012
rect 17092 20000 17098 20052
rect 17678 20040 17684 20052
rect 17639 20012 17684 20040
rect 17678 20000 17684 20012
rect 17736 20000 17742 20052
rect 18138 20000 18144 20052
rect 18196 20040 18202 20052
rect 18601 20043 18659 20049
rect 18601 20040 18613 20043
rect 18196 20012 18613 20040
rect 18196 20000 18202 20012
rect 18601 20009 18613 20012
rect 18647 20009 18659 20043
rect 18601 20003 18659 20009
rect 18690 20000 18696 20052
rect 18748 20040 18754 20052
rect 21634 20040 21640 20052
rect 18748 20012 21640 20040
rect 18748 20000 18754 20012
rect 21634 20000 21640 20012
rect 21692 20040 21698 20052
rect 22830 20040 22836 20052
rect 21692 20012 22836 20040
rect 21692 20000 21698 20012
rect 22830 20000 22836 20012
rect 22888 20000 22894 20052
rect 23109 20043 23167 20049
rect 23109 20009 23121 20043
rect 23155 20040 23167 20043
rect 23566 20040 23572 20052
rect 23155 20012 23572 20040
rect 23155 20009 23167 20012
rect 23109 20003 23167 20009
rect 23566 20000 23572 20012
rect 23624 20000 23630 20052
rect 13495 19944 16344 19972
rect 13495 19941 13507 19944
rect 13449 19935 13507 19941
rect 18322 19932 18328 19984
rect 18380 19932 18386 19984
rect 16022 19904 16028 19916
rect 13372 19876 16028 19904
rect 13372 19845 13400 19876
rect 16022 19864 16028 19876
rect 16080 19864 16086 19916
rect 16298 19904 16304 19916
rect 16259 19876 16304 19904
rect 16298 19864 16304 19876
rect 16356 19864 16362 19916
rect 18340 19904 18368 19932
rect 18417 19907 18475 19913
rect 18417 19904 18429 19907
rect 17328 19876 18429 19904
rect 13357 19839 13415 19845
rect 13357 19805 13369 19839
rect 13403 19805 13415 19839
rect 13538 19836 13544 19848
rect 13499 19808 13544 19836
rect 13357 19799 13415 19805
rect 13538 19796 13544 19808
rect 13596 19796 13602 19848
rect 14182 19796 14188 19848
rect 14240 19836 14246 19848
rect 14369 19839 14427 19845
rect 14369 19836 14381 19839
rect 14240 19808 14381 19836
rect 14240 19796 14246 19808
rect 14369 19805 14381 19808
rect 14415 19805 14427 19839
rect 14642 19836 14648 19848
rect 14555 19808 14648 19836
rect 14369 19799 14427 19805
rect 14642 19796 14648 19808
rect 14700 19796 14706 19848
rect 15102 19836 15108 19848
rect 15063 19808 15108 19836
rect 15102 19796 15108 19808
rect 15160 19796 15166 19848
rect 15470 19836 15476 19848
rect 15431 19808 15476 19836
rect 15470 19796 15476 19808
rect 15528 19796 15534 19848
rect 16206 19796 16212 19848
rect 16264 19836 16270 19848
rect 16557 19839 16615 19845
rect 16557 19836 16569 19839
rect 16264 19808 16569 19836
rect 16264 19796 16270 19808
rect 16557 19805 16569 19808
rect 16603 19805 16615 19839
rect 16557 19799 16615 19805
rect 16942 19796 16948 19848
rect 17000 19836 17006 19848
rect 17328 19836 17356 19876
rect 18417 19873 18429 19876
rect 18463 19873 18475 19907
rect 19426 19904 19432 19916
rect 19387 19876 19432 19904
rect 18417 19867 18475 19873
rect 19426 19864 19432 19876
rect 19484 19864 19490 19916
rect 21266 19904 21272 19916
rect 21227 19876 21272 19904
rect 21266 19864 21272 19876
rect 21324 19864 21330 19916
rect 22848 19904 22876 20000
rect 23658 19972 23664 19984
rect 23584 19944 23664 19972
rect 23584 19913 23612 19944
rect 23658 19932 23664 19944
rect 23716 19932 23722 19984
rect 23569 19907 23627 19913
rect 22848 19876 23428 19904
rect 17000 19808 17356 19836
rect 17000 19796 17006 19808
rect 17954 19796 17960 19848
rect 18012 19836 18018 19848
rect 18325 19839 18383 19845
rect 18325 19836 18337 19839
rect 18012 19808 18337 19836
rect 18012 19796 18018 19808
rect 18325 19805 18337 19808
rect 18371 19836 18383 19839
rect 19242 19836 19248 19848
rect 18371 19808 19248 19836
rect 18371 19805 18383 19808
rect 18325 19799 18383 19805
rect 19242 19796 19248 19808
rect 19300 19836 19306 19848
rect 19518 19836 19524 19848
rect 19300 19808 19524 19836
rect 19300 19796 19306 19808
rect 19518 19796 19524 19808
rect 19576 19796 19582 19848
rect 19696 19839 19754 19845
rect 19696 19805 19708 19839
rect 19742 19836 19754 19839
rect 20162 19836 20168 19848
rect 19742 19808 20168 19836
rect 19742 19805 19754 19808
rect 19696 19799 19754 19805
rect 20162 19796 20168 19808
rect 20220 19796 20226 19848
rect 22002 19836 22008 19848
rect 21008 19808 22008 19836
rect 14660 19768 14688 19796
rect 21008 19780 21036 19808
rect 22002 19796 22008 19808
rect 22060 19796 22066 19848
rect 23290 19836 23296 19848
rect 23251 19808 23296 19836
rect 23290 19796 23296 19808
rect 23348 19796 23354 19848
rect 23400 19845 23428 19876
rect 23569 19873 23581 19907
rect 23615 19873 23627 19907
rect 26510 19904 26516 19916
rect 26471 19876 26516 19904
rect 23569 19867 23627 19873
rect 26510 19864 26516 19876
rect 26568 19864 26574 19916
rect 23385 19839 23443 19845
rect 23385 19805 23397 19839
rect 23431 19805 23443 19839
rect 23385 19799 23443 19805
rect 23661 19839 23719 19845
rect 23661 19805 23673 19839
rect 23707 19836 23719 19839
rect 23750 19836 23756 19848
rect 23707 19808 23756 19836
rect 23707 19805 23719 19808
rect 23661 19799 23719 19805
rect 23750 19796 23756 19808
rect 23808 19796 23814 19848
rect 24670 19845 24676 19848
rect 24397 19839 24455 19845
rect 24397 19805 24409 19839
rect 24443 19805 24455 19839
rect 24664 19836 24676 19845
rect 24631 19808 24676 19836
rect 24397 19799 24455 19805
rect 24664 19799 24676 19808
rect 15378 19768 15384 19780
rect 14660 19740 15384 19768
rect 15378 19728 15384 19740
rect 15436 19728 15442 19780
rect 18874 19728 18880 19780
rect 18932 19768 18938 19780
rect 20990 19768 20996 19780
rect 18932 19740 20996 19768
rect 18932 19728 18938 19740
rect 20990 19728 20996 19740
rect 21048 19728 21054 19780
rect 21542 19777 21548 19780
rect 21536 19731 21548 19777
rect 21600 19768 21606 19780
rect 24412 19768 24440 19799
rect 24670 19796 24676 19799
rect 24728 19796 24734 19848
rect 26329 19839 26387 19845
rect 26329 19805 26341 19839
rect 26375 19805 26387 19839
rect 28166 19836 28172 19848
rect 28127 19808 28172 19836
rect 26329 19799 26387 19805
rect 25038 19768 25044 19780
rect 21600 19740 21636 19768
rect 24412 19740 25044 19768
rect 21542 19728 21548 19731
rect 21600 19728 21606 19740
rect 25038 19728 25044 19740
rect 25096 19728 25102 19780
rect 26344 19768 26372 19799
rect 28166 19796 28172 19808
rect 28224 19796 28230 19848
rect 27430 19768 27436 19780
rect 26344 19740 27436 19768
rect 27430 19728 27436 19740
rect 27488 19728 27494 19780
rect 14185 19703 14243 19709
rect 14185 19669 14197 19703
rect 14231 19700 14243 19703
rect 15562 19700 15568 19712
rect 14231 19672 15568 19700
rect 14231 19669 14243 19672
rect 14185 19663 14243 19669
rect 15562 19660 15568 19672
rect 15620 19660 15626 19712
rect 16114 19660 16120 19712
rect 16172 19700 16178 19712
rect 18690 19700 18696 19712
rect 16172 19672 18696 19700
rect 16172 19660 16178 19672
rect 18690 19660 18696 19672
rect 18748 19660 18754 19712
rect 19886 19660 19892 19712
rect 19944 19700 19950 19712
rect 20622 19700 20628 19712
rect 19944 19672 20628 19700
rect 19944 19660 19950 19672
rect 20622 19660 20628 19672
rect 20680 19700 20686 19712
rect 20809 19703 20867 19709
rect 20809 19700 20821 19703
rect 20680 19672 20821 19700
rect 20680 19660 20686 19672
rect 20809 19669 20821 19672
rect 20855 19669 20867 19703
rect 20809 19663 20867 19669
rect 22554 19660 22560 19712
rect 22612 19700 22618 19712
rect 22649 19703 22707 19709
rect 22649 19700 22661 19703
rect 22612 19672 22661 19700
rect 22612 19660 22618 19672
rect 22649 19669 22661 19672
rect 22695 19669 22707 19703
rect 25774 19700 25780 19712
rect 25735 19672 25780 19700
rect 22649 19663 22707 19669
rect 25774 19660 25780 19672
rect 25832 19660 25838 19712
rect 1104 19610 28888 19632
rect 1104 19558 10214 19610
rect 10266 19558 10278 19610
rect 10330 19558 10342 19610
rect 10394 19558 10406 19610
rect 10458 19558 10470 19610
rect 10522 19558 19478 19610
rect 19530 19558 19542 19610
rect 19594 19558 19606 19610
rect 19658 19558 19670 19610
rect 19722 19558 19734 19610
rect 19786 19558 28888 19610
rect 1104 19536 28888 19558
rect 13354 19456 13360 19508
rect 13412 19496 13418 19508
rect 17773 19499 17831 19505
rect 13412 19468 16804 19496
rect 13412 19456 13418 19468
rect 16776 19440 16804 19468
rect 17773 19465 17785 19499
rect 17819 19496 17831 19499
rect 18782 19496 18788 19508
rect 17819 19468 18788 19496
rect 17819 19465 17831 19468
rect 17773 19459 17831 19465
rect 18782 19456 18788 19468
rect 18840 19456 18846 19508
rect 18877 19499 18935 19505
rect 18877 19465 18889 19499
rect 18923 19465 18935 19499
rect 18877 19459 18935 19465
rect 13078 19388 13084 19440
rect 13136 19428 13142 19440
rect 13136 19400 15516 19428
rect 13136 19388 13142 19400
rect 14461 19363 14519 19369
rect 14461 19329 14473 19363
rect 14507 19360 14519 19363
rect 14734 19360 14740 19372
rect 14507 19332 14740 19360
rect 14507 19329 14519 19332
rect 14461 19323 14519 19329
rect 14734 19320 14740 19332
rect 14792 19320 14798 19372
rect 15488 19369 15516 19400
rect 16758 19388 16764 19440
rect 16816 19428 16822 19440
rect 18414 19428 18420 19440
rect 16816 19400 18420 19428
rect 16816 19388 16822 19400
rect 18414 19388 18420 19400
rect 18472 19388 18478 19440
rect 18509 19431 18567 19437
rect 18509 19397 18521 19431
rect 18555 19428 18567 19431
rect 18555 19400 18828 19428
rect 18555 19397 18567 19400
rect 18509 19391 18567 19397
rect 15381 19363 15439 19369
rect 15381 19329 15393 19363
rect 15427 19329 15439 19363
rect 15381 19323 15439 19329
rect 15473 19363 15531 19369
rect 15473 19329 15485 19363
rect 15519 19360 15531 19363
rect 15930 19360 15936 19372
rect 15519 19332 15936 19360
rect 15519 19329 15531 19332
rect 15473 19323 15531 19329
rect 13538 19252 13544 19304
rect 13596 19292 13602 19304
rect 15102 19292 15108 19304
rect 13596 19264 15108 19292
rect 13596 19252 13602 19264
rect 15102 19252 15108 19264
rect 15160 19252 15166 19304
rect 15289 19295 15347 19301
rect 15289 19261 15301 19295
rect 15335 19261 15347 19295
rect 15289 19255 15347 19261
rect 14642 19184 14648 19236
rect 14700 19224 14706 19236
rect 15304 19224 15332 19255
rect 14700 19196 15332 19224
rect 15396 19224 15424 19323
rect 15930 19320 15936 19332
rect 15988 19320 15994 19372
rect 16853 19363 16911 19369
rect 16853 19329 16865 19363
rect 16899 19360 16911 19363
rect 17034 19360 17040 19372
rect 16899 19332 17040 19360
rect 16899 19329 16911 19332
rect 16853 19323 16911 19329
rect 17034 19320 17040 19332
rect 17092 19320 17098 19372
rect 17681 19363 17739 19369
rect 17681 19329 17693 19363
rect 17727 19360 17739 19363
rect 18046 19360 18052 19372
rect 17727 19332 18052 19360
rect 17727 19329 17739 19332
rect 17681 19323 17739 19329
rect 18046 19320 18052 19332
rect 18104 19320 18110 19372
rect 18322 19360 18328 19372
rect 18283 19332 18328 19360
rect 18322 19320 18328 19332
rect 18380 19320 18386 19372
rect 18601 19363 18659 19369
rect 18601 19329 18613 19363
rect 18647 19329 18659 19363
rect 18601 19323 18659 19329
rect 18693 19363 18751 19369
rect 18693 19329 18705 19363
rect 18739 19329 18751 19363
rect 18693 19323 18751 19329
rect 15562 19252 15568 19304
rect 15620 19292 15626 19304
rect 16942 19292 16948 19304
rect 15620 19264 15665 19292
rect 16903 19264 16948 19292
rect 15620 19252 15626 19264
rect 16942 19252 16948 19264
rect 17000 19252 17006 19304
rect 17052 19292 17080 19320
rect 18616 19292 18644 19323
rect 17052 19264 18644 19292
rect 15654 19224 15660 19236
rect 15396 19196 15660 19224
rect 14700 19184 14706 19196
rect 14550 19156 14556 19168
rect 14511 19128 14556 19156
rect 14550 19116 14556 19128
rect 14608 19116 14614 19168
rect 15304 19156 15332 19196
rect 15654 19184 15660 19196
rect 15712 19184 15718 19236
rect 16850 19184 16856 19236
rect 16908 19224 16914 19236
rect 17862 19224 17868 19236
rect 16908 19196 17868 19224
rect 16908 19184 16914 19196
rect 17862 19184 17868 19196
rect 17920 19184 17926 19236
rect 15562 19156 15568 19168
rect 15304 19128 15568 19156
rect 15562 19116 15568 19128
rect 15620 19116 15626 19168
rect 16022 19116 16028 19168
rect 16080 19156 16086 19168
rect 16482 19156 16488 19168
rect 16080 19128 16488 19156
rect 16080 19116 16086 19128
rect 16482 19116 16488 19128
rect 16540 19156 16546 19168
rect 17129 19159 17187 19165
rect 17129 19156 17141 19159
rect 16540 19128 17141 19156
rect 16540 19116 16546 19128
rect 17129 19125 17141 19128
rect 17175 19125 17187 19159
rect 18616 19156 18644 19264
rect 18708 19224 18736 19323
rect 18800 19292 18828 19400
rect 18892 19360 18920 19459
rect 18966 19456 18972 19508
rect 19024 19496 19030 19508
rect 19024 19468 20024 19496
rect 19024 19456 19030 19468
rect 19242 19388 19248 19440
rect 19300 19428 19306 19440
rect 19996 19428 20024 19468
rect 20806 19456 20812 19508
rect 20864 19496 20870 19508
rect 21085 19499 21143 19505
rect 21085 19496 21097 19499
rect 20864 19468 21097 19496
rect 20864 19456 20870 19468
rect 21085 19465 21097 19468
rect 21131 19465 21143 19499
rect 21085 19459 21143 19465
rect 23474 19456 23480 19508
rect 23532 19496 23538 19508
rect 24121 19499 24179 19505
rect 24121 19496 24133 19499
rect 23532 19468 24133 19496
rect 23532 19456 23538 19468
rect 24121 19465 24133 19468
rect 24167 19465 24179 19499
rect 24121 19459 24179 19465
rect 26050 19456 26056 19508
rect 26108 19496 26114 19508
rect 27433 19499 27491 19505
rect 27433 19496 27445 19499
rect 26108 19468 27445 19496
rect 26108 19456 26114 19468
rect 27433 19465 27445 19468
rect 27479 19465 27491 19499
rect 27433 19459 27491 19465
rect 23290 19428 23296 19440
rect 19300 19400 19932 19428
rect 19996 19400 23296 19428
rect 19300 19388 19306 19400
rect 19337 19363 19395 19369
rect 19337 19360 19349 19363
rect 18892 19332 19349 19360
rect 19337 19329 19349 19332
rect 19383 19329 19395 19363
rect 19337 19323 19395 19329
rect 19521 19363 19579 19369
rect 19521 19329 19533 19363
rect 19567 19329 19579 19363
rect 19521 19323 19579 19329
rect 19705 19363 19763 19369
rect 19705 19329 19717 19363
rect 19751 19360 19763 19363
rect 19794 19360 19800 19372
rect 19751 19332 19800 19360
rect 19751 19329 19763 19332
rect 19705 19323 19763 19329
rect 19426 19292 19432 19304
rect 18800 19264 19432 19292
rect 19426 19252 19432 19264
rect 19484 19252 19490 19304
rect 19536 19236 19564 19323
rect 19794 19320 19800 19332
rect 19852 19320 19858 19372
rect 19904 19369 19932 19400
rect 23290 19388 23296 19400
rect 23348 19388 23354 19440
rect 23842 19428 23848 19440
rect 23803 19400 23848 19428
rect 23842 19388 23848 19400
rect 23900 19388 23906 19440
rect 25774 19388 25780 19440
rect 25832 19428 25838 19440
rect 27985 19431 28043 19437
rect 27985 19428 27997 19431
rect 25832 19400 27997 19428
rect 25832 19388 25838 19400
rect 27985 19397 27997 19400
rect 28031 19397 28043 19431
rect 27985 19391 28043 19397
rect 19889 19363 19947 19369
rect 19889 19329 19901 19363
rect 19935 19329 19947 19363
rect 19889 19323 19947 19329
rect 20254 19320 20260 19372
rect 20312 19360 20318 19372
rect 20809 19363 20867 19369
rect 20809 19360 20821 19363
rect 20312 19332 20821 19360
rect 20312 19320 20318 19332
rect 20809 19329 20821 19332
rect 20855 19329 20867 19363
rect 20809 19323 20867 19329
rect 22186 19320 22192 19372
rect 22244 19360 22250 19372
rect 22557 19363 22615 19369
rect 22557 19360 22569 19363
rect 22244 19332 22569 19360
rect 22244 19320 22250 19332
rect 22557 19329 22569 19332
rect 22603 19329 22615 19363
rect 22557 19323 22615 19329
rect 23382 19320 23388 19372
rect 23440 19360 23446 19372
rect 23566 19360 23572 19372
rect 23440 19332 23572 19360
rect 23440 19320 23446 19332
rect 23566 19320 23572 19332
rect 23624 19320 23630 19372
rect 23658 19320 23664 19372
rect 23716 19360 23722 19372
rect 23753 19363 23811 19369
rect 23753 19360 23765 19363
rect 23716 19332 23765 19360
rect 23716 19320 23722 19332
rect 23753 19329 23765 19332
rect 23799 19329 23811 19363
rect 23934 19360 23940 19372
rect 23895 19332 23940 19360
rect 23753 19323 23811 19329
rect 23934 19320 23940 19332
rect 23992 19320 23998 19372
rect 25038 19360 25044 19372
rect 24999 19332 25044 19360
rect 25038 19320 25044 19332
rect 25096 19320 25102 19372
rect 25308 19363 25366 19369
rect 25308 19329 25320 19363
rect 25354 19360 25366 19363
rect 26878 19360 26884 19372
rect 25354 19332 26884 19360
rect 25354 19329 25366 19332
rect 25308 19323 25366 19329
rect 26878 19320 26884 19332
rect 26936 19320 26942 19372
rect 26973 19363 27031 19369
rect 26973 19329 26985 19363
rect 27019 19360 27031 19363
rect 27338 19360 27344 19372
rect 27019 19332 27344 19360
rect 27019 19329 27031 19332
rect 26973 19323 27031 19329
rect 19613 19295 19671 19301
rect 19613 19261 19625 19295
rect 19659 19261 19671 19295
rect 20070 19292 20076 19304
rect 20031 19264 20076 19292
rect 19613 19255 19671 19261
rect 19518 19224 19524 19236
rect 18708 19196 19524 19224
rect 19518 19184 19524 19196
rect 19576 19184 19582 19236
rect 19628 19156 19656 19255
rect 20070 19252 20076 19264
rect 20128 19252 20134 19304
rect 20901 19295 20959 19301
rect 20901 19261 20913 19295
rect 20947 19292 20959 19295
rect 20990 19292 20996 19304
rect 20947 19264 20996 19292
rect 20947 19261 20959 19264
rect 20901 19255 20959 19261
rect 20990 19252 20996 19264
rect 21048 19252 21054 19304
rect 21085 19295 21143 19301
rect 21085 19261 21097 19295
rect 21131 19292 21143 19295
rect 22094 19292 22100 19304
rect 21131 19264 22100 19292
rect 21131 19261 21143 19264
rect 21085 19255 21143 19261
rect 22094 19252 22100 19264
rect 22152 19252 22158 19304
rect 22281 19295 22339 19301
rect 22281 19261 22293 19295
rect 22327 19292 22339 19295
rect 26988 19292 27016 19323
rect 27338 19320 27344 19332
rect 27396 19320 27402 19372
rect 22327 19264 22600 19292
rect 22327 19261 22339 19264
rect 22281 19255 22339 19261
rect 22572 19236 22600 19264
rect 26436 19264 27016 19292
rect 22554 19184 22560 19236
rect 22612 19184 22618 19236
rect 23842 19184 23848 19236
rect 23900 19224 23906 19236
rect 24302 19224 24308 19236
rect 23900 19196 24308 19224
rect 23900 19184 23906 19196
rect 24302 19184 24308 19196
rect 24360 19184 24366 19236
rect 18616 19128 19656 19156
rect 17129 19119 17187 19125
rect 21726 19116 21732 19168
rect 21784 19156 21790 19168
rect 23860 19156 23888 19184
rect 26436 19168 26464 19264
rect 21784 19128 23888 19156
rect 21784 19116 21790 19128
rect 24854 19116 24860 19168
rect 24912 19156 24918 19168
rect 25314 19156 25320 19168
rect 24912 19128 25320 19156
rect 24912 19116 24918 19128
rect 25314 19116 25320 19128
rect 25372 19116 25378 19168
rect 26418 19156 26424 19168
rect 26379 19128 26424 19156
rect 26418 19116 26424 19128
rect 26476 19116 26482 19168
rect 26602 19116 26608 19168
rect 26660 19156 26666 19168
rect 27065 19159 27123 19165
rect 27065 19156 27077 19159
rect 26660 19128 27077 19156
rect 26660 19116 26666 19128
rect 27065 19125 27077 19128
rect 27111 19125 27123 19159
rect 27065 19119 27123 19125
rect 27246 19116 27252 19168
rect 27304 19156 27310 19168
rect 28077 19159 28135 19165
rect 28077 19156 28089 19159
rect 27304 19128 28089 19156
rect 27304 19116 27310 19128
rect 28077 19125 28089 19128
rect 28123 19125 28135 19159
rect 28077 19119 28135 19125
rect 1104 19066 28888 19088
rect 1104 19014 5582 19066
rect 5634 19014 5646 19066
rect 5698 19014 5710 19066
rect 5762 19014 5774 19066
rect 5826 19014 5838 19066
rect 5890 19014 14846 19066
rect 14898 19014 14910 19066
rect 14962 19014 14974 19066
rect 15026 19014 15038 19066
rect 15090 19014 15102 19066
rect 15154 19014 24110 19066
rect 24162 19014 24174 19066
rect 24226 19014 24238 19066
rect 24290 19014 24302 19066
rect 24354 19014 24366 19066
rect 24418 19014 28888 19066
rect 1104 18992 28888 19014
rect 15194 18912 15200 18964
rect 15252 18952 15258 18964
rect 16298 18952 16304 18964
rect 15252 18924 16304 18952
rect 15252 18912 15258 18924
rect 16298 18912 16304 18924
rect 16356 18952 16362 18964
rect 16393 18955 16451 18961
rect 16393 18952 16405 18955
rect 16356 18924 16405 18952
rect 16356 18912 16362 18924
rect 16393 18921 16405 18924
rect 16439 18921 16451 18955
rect 18874 18952 18880 18964
rect 16393 18915 16451 18921
rect 16960 18924 18880 18952
rect 12710 18844 12716 18896
rect 12768 18884 12774 18896
rect 15562 18884 15568 18896
rect 12768 18856 15240 18884
rect 15523 18856 15568 18884
rect 12768 18844 12774 18856
rect 14182 18776 14188 18828
rect 14240 18816 14246 18828
rect 14734 18816 14740 18828
rect 14240 18788 14740 18816
rect 14240 18776 14246 18788
rect 14734 18776 14740 18788
rect 14792 18816 14798 18828
rect 15105 18819 15163 18825
rect 15105 18816 15117 18819
rect 14792 18788 15117 18816
rect 14792 18776 14798 18788
rect 15105 18785 15117 18788
rect 15151 18785 15163 18819
rect 15212 18816 15240 18856
rect 15562 18844 15568 18856
rect 15620 18844 15626 18896
rect 16114 18816 16120 18828
rect 15212 18788 16120 18816
rect 15105 18779 15163 18785
rect 16114 18776 16120 18788
rect 16172 18776 16178 18828
rect 14366 18748 14372 18760
rect 14327 18720 14372 18748
rect 14366 18708 14372 18720
rect 14424 18708 14430 18760
rect 14461 18751 14519 18757
rect 14461 18717 14473 18751
rect 14507 18748 14519 18751
rect 15197 18751 15255 18757
rect 15197 18748 15209 18751
rect 14507 18720 15209 18748
rect 14507 18717 14519 18720
rect 14461 18711 14519 18717
rect 15197 18717 15209 18720
rect 15243 18748 15255 18751
rect 16960 18748 16988 18924
rect 18874 18912 18880 18924
rect 18932 18912 18938 18964
rect 19426 18912 19432 18964
rect 19484 18952 19490 18964
rect 19613 18955 19671 18961
rect 19613 18952 19625 18955
rect 19484 18924 19625 18952
rect 19484 18912 19490 18924
rect 19613 18921 19625 18924
rect 19659 18921 19671 18955
rect 19613 18915 19671 18921
rect 19886 18912 19892 18964
rect 19944 18952 19950 18964
rect 20257 18955 20315 18961
rect 20257 18952 20269 18955
rect 19944 18924 20269 18952
rect 19944 18912 19950 18924
rect 20257 18921 20269 18924
rect 20303 18921 20315 18955
rect 20257 18915 20315 18921
rect 20714 18912 20720 18964
rect 20772 18952 20778 18964
rect 21174 18952 21180 18964
rect 20772 18924 21180 18952
rect 20772 18912 20778 18924
rect 21174 18912 21180 18924
rect 21232 18912 21238 18964
rect 22094 18912 22100 18964
rect 22152 18952 22158 18964
rect 22462 18952 22468 18964
rect 22152 18924 22468 18952
rect 22152 18912 22158 18924
rect 22462 18912 22468 18924
rect 22520 18952 22526 18964
rect 23382 18952 23388 18964
rect 22520 18924 23388 18952
rect 22520 18912 22526 18924
rect 23382 18912 23388 18924
rect 23440 18912 23446 18964
rect 23566 18912 23572 18964
rect 23624 18952 23630 18964
rect 23753 18955 23811 18961
rect 23753 18952 23765 18955
rect 23624 18924 23765 18952
rect 23624 18912 23630 18924
rect 23753 18921 23765 18924
rect 23799 18921 23811 18955
rect 27706 18952 27712 18964
rect 23753 18915 23811 18921
rect 23860 18924 27712 18952
rect 17954 18884 17960 18896
rect 17915 18856 17960 18884
rect 17954 18844 17960 18856
rect 18012 18844 18018 18896
rect 18046 18844 18052 18896
rect 18104 18884 18110 18896
rect 18104 18856 21956 18884
rect 18104 18844 18110 18856
rect 18138 18816 18144 18828
rect 17236 18788 18144 18816
rect 17126 18748 17132 18760
rect 15243 18720 16988 18748
rect 17087 18720 17132 18748
rect 15243 18717 15255 18720
rect 15197 18711 15255 18717
rect 17126 18708 17132 18720
rect 17184 18708 17190 18760
rect 17236 18757 17264 18788
rect 18138 18776 18144 18788
rect 18196 18776 18202 18828
rect 21174 18816 21180 18828
rect 21135 18788 21180 18816
rect 21174 18776 21180 18788
rect 21232 18776 21238 18828
rect 17221 18751 17279 18757
rect 17221 18717 17233 18751
rect 17267 18717 17279 18751
rect 17221 18711 17279 18717
rect 17405 18751 17463 18757
rect 17405 18717 17417 18751
rect 17451 18717 17463 18751
rect 17405 18711 17463 18717
rect 12802 18640 12808 18692
rect 12860 18680 12866 18692
rect 16301 18683 16359 18689
rect 16301 18680 16313 18683
rect 12860 18652 16313 18680
rect 12860 18640 12866 18652
rect 16301 18649 16313 18652
rect 16347 18649 16359 18683
rect 16301 18643 16359 18649
rect 16666 18640 16672 18692
rect 16724 18680 16730 18692
rect 17420 18680 17448 18711
rect 17494 18708 17500 18760
rect 17552 18748 17558 18760
rect 18233 18751 18291 18757
rect 17552 18720 17597 18748
rect 17552 18708 17558 18720
rect 18233 18717 18245 18751
rect 18279 18748 18291 18751
rect 18414 18748 18420 18760
rect 18279 18720 18420 18748
rect 18279 18717 18291 18720
rect 18233 18711 18291 18717
rect 18414 18708 18420 18720
rect 18472 18708 18478 18760
rect 18874 18708 18880 18760
rect 18932 18748 18938 18760
rect 19429 18751 19487 18757
rect 19429 18748 19441 18751
rect 18932 18720 19441 18748
rect 18932 18708 18938 18720
rect 19429 18717 19441 18720
rect 19475 18717 19487 18751
rect 20622 18748 20628 18760
rect 19429 18711 19487 18717
rect 20088 18720 20628 18748
rect 16724 18652 17448 18680
rect 17957 18683 18015 18689
rect 16724 18640 16730 18652
rect 17957 18649 17969 18683
rect 18003 18680 18015 18683
rect 18046 18680 18052 18692
rect 18003 18652 18052 18680
rect 18003 18649 18015 18652
rect 17957 18643 18015 18649
rect 18046 18640 18052 18652
rect 18104 18640 18110 18692
rect 19245 18683 19303 18689
rect 19245 18649 19257 18683
rect 19291 18649 19303 18683
rect 19245 18643 19303 18649
rect 14366 18572 14372 18624
rect 14424 18612 14430 18624
rect 15378 18612 15384 18624
rect 14424 18584 15384 18612
rect 14424 18572 14430 18584
rect 15378 18572 15384 18584
rect 15436 18572 15442 18624
rect 16945 18615 17003 18621
rect 16945 18581 16957 18615
rect 16991 18612 17003 18615
rect 17310 18612 17316 18624
rect 16991 18584 17316 18612
rect 16991 18581 17003 18584
rect 16945 18575 17003 18581
rect 17310 18572 17316 18584
rect 17368 18572 17374 18624
rect 18141 18615 18199 18621
rect 18141 18581 18153 18615
rect 18187 18612 18199 18615
rect 18230 18612 18236 18624
rect 18187 18584 18236 18612
rect 18187 18581 18199 18584
rect 18141 18575 18199 18581
rect 18230 18572 18236 18584
rect 18288 18572 18294 18624
rect 19260 18612 19288 18643
rect 19518 18640 19524 18692
rect 19576 18680 19582 18692
rect 20088 18689 20116 18720
rect 20622 18708 20628 18720
rect 20680 18748 20686 18760
rect 20901 18751 20959 18757
rect 20901 18748 20913 18751
rect 20680 18720 20913 18748
rect 20680 18708 20686 18720
rect 20901 18717 20913 18720
rect 20947 18717 20959 18751
rect 20901 18711 20959 18717
rect 20990 18708 20996 18760
rect 21048 18748 21054 18760
rect 21726 18748 21732 18760
rect 21048 18720 21093 18748
rect 21687 18720 21732 18748
rect 21048 18708 21054 18720
rect 21726 18708 21732 18720
rect 21784 18708 21790 18760
rect 21928 18757 21956 18856
rect 23198 18844 23204 18896
rect 23256 18884 23262 18896
rect 23860 18884 23888 18924
rect 27706 18912 27712 18924
rect 27764 18912 27770 18964
rect 27246 18884 27252 18896
rect 23256 18856 23888 18884
rect 25056 18856 27252 18884
rect 23256 18844 23262 18856
rect 22094 18776 22100 18828
rect 22152 18816 22158 18828
rect 22557 18819 22615 18825
rect 22557 18816 22569 18819
rect 22152 18788 22569 18816
rect 22152 18776 22158 18788
rect 22557 18785 22569 18788
rect 22603 18785 22615 18819
rect 22557 18779 22615 18785
rect 21913 18751 21971 18757
rect 21913 18717 21925 18751
rect 21959 18717 21971 18751
rect 21913 18711 21971 18717
rect 22005 18751 22063 18757
rect 22005 18717 22017 18751
rect 22051 18748 22063 18751
rect 22186 18748 22192 18760
rect 22051 18720 22192 18748
rect 22051 18717 22063 18720
rect 22005 18711 22063 18717
rect 20073 18683 20131 18689
rect 20073 18680 20085 18683
rect 19576 18652 20085 18680
rect 19576 18640 19582 18652
rect 20073 18649 20085 18652
rect 20119 18649 20131 18683
rect 20073 18643 20131 18649
rect 20162 18640 20168 18692
rect 20220 18680 20226 18692
rect 21177 18683 21235 18689
rect 21177 18680 21189 18683
rect 20220 18652 21189 18680
rect 20220 18640 20226 18652
rect 21177 18649 21189 18652
rect 21223 18649 21235 18683
rect 21928 18680 21956 18711
rect 22186 18708 22192 18720
rect 22244 18708 22250 18760
rect 22465 18751 22523 18757
rect 22465 18717 22477 18751
rect 22511 18748 22523 18751
rect 22830 18748 22836 18760
rect 22511 18720 22836 18748
rect 22511 18717 22523 18720
rect 22465 18711 22523 18717
rect 22830 18708 22836 18720
rect 22888 18708 22894 18760
rect 23661 18751 23719 18757
rect 23661 18717 23673 18751
rect 23707 18748 23719 18751
rect 23750 18748 23756 18760
rect 23707 18720 23756 18748
rect 23707 18717 23719 18720
rect 23661 18711 23719 18717
rect 23750 18708 23756 18720
rect 23808 18708 23814 18760
rect 24857 18751 24915 18757
rect 24857 18717 24869 18751
rect 24903 18748 24915 18751
rect 25056 18748 25084 18856
rect 27246 18844 27252 18856
rect 27304 18844 27310 18896
rect 25323 18816 25452 18824
rect 25498 18816 25504 18828
rect 25240 18796 25504 18816
rect 25240 18788 25351 18796
rect 25424 18788 25504 18796
rect 25240 18757 25268 18788
rect 25498 18776 25504 18788
rect 25556 18776 25562 18828
rect 28166 18816 28172 18828
rect 28127 18788 28172 18816
rect 28166 18776 28172 18788
rect 28224 18776 28230 18828
rect 24903 18720 25084 18748
rect 25225 18751 25283 18757
rect 24903 18717 24915 18720
rect 24857 18711 24915 18717
rect 25225 18717 25237 18751
rect 25271 18717 25283 18751
rect 26326 18748 26332 18760
rect 26287 18720 26332 18748
rect 25225 18711 25283 18717
rect 26326 18708 26332 18720
rect 26384 18708 26390 18760
rect 22278 18680 22284 18692
rect 21928 18652 22284 18680
rect 21177 18643 21235 18649
rect 22278 18640 22284 18652
rect 22336 18640 22342 18692
rect 22741 18683 22799 18689
rect 22741 18649 22753 18683
rect 22787 18680 22799 18683
rect 23290 18680 23296 18692
rect 22787 18652 23296 18680
rect 22787 18649 22799 18652
rect 22741 18643 22799 18649
rect 23290 18640 23296 18652
rect 23348 18640 23354 18692
rect 24946 18640 24952 18692
rect 25004 18680 25010 18692
rect 25041 18683 25099 18689
rect 25041 18680 25053 18683
rect 25004 18652 25053 18680
rect 25004 18640 25010 18652
rect 25041 18649 25053 18652
rect 25087 18649 25099 18683
rect 25041 18643 25099 18649
rect 25130 18640 25136 18692
rect 25188 18680 25194 18692
rect 25188 18652 25233 18680
rect 25188 18640 25194 18652
rect 26234 18640 26240 18692
rect 26292 18680 26298 18692
rect 26513 18683 26571 18689
rect 26513 18680 26525 18683
rect 26292 18652 26525 18680
rect 26292 18640 26298 18652
rect 26513 18649 26525 18652
rect 26559 18649 26571 18683
rect 26513 18643 26571 18649
rect 19886 18612 19892 18624
rect 19260 18584 19892 18612
rect 19886 18572 19892 18584
rect 19944 18572 19950 18624
rect 20254 18572 20260 18624
rect 20312 18621 20318 18624
rect 20312 18615 20331 18621
rect 20319 18581 20331 18615
rect 20438 18612 20444 18624
rect 20399 18584 20444 18612
rect 20312 18575 20331 18581
rect 20312 18572 20318 18575
rect 20438 18572 20444 18584
rect 20496 18572 20502 18624
rect 21818 18612 21824 18624
rect 21876 18621 21882 18624
rect 21785 18584 21824 18612
rect 21818 18572 21824 18584
rect 21876 18575 21885 18621
rect 22462 18612 22468 18624
rect 22423 18584 22468 18612
rect 21876 18572 21882 18575
rect 22462 18572 22468 18584
rect 22520 18572 22526 18624
rect 24302 18572 24308 18624
rect 24360 18612 24366 18624
rect 25409 18615 25467 18621
rect 25409 18612 25421 18615
rect 24360 18584 25421 18612
rect 24360 18572 24366 18584
rect 25409 18581 25421 18584
rect 25455 18581 25467 18615
rect 25409 18575 25467 18581
rect 1104 18522 28888 18544
rect 1104 18470 10214 18522
rect 10266 18470 10278 18522
rect 10330 18470 10342 18522
rect 10394 18470 10406 18522
rect 10458 18470 10470 18522
rect 10522 18470 19478 18522
rect 19530 18470 19542 18522
rect 19594 18470 19606 18522
rect 19658 18470 19670 18522
rect 19722 18470 19734 18522
rect 19786 18470 28888 18522
rect 1104 18448 28888 18470
rect 13725 18411 13783 18417
rect 13725 18377 13737 18411
rect 13771 18408 13783 18411
rect 17494 18408 17500 18420
rect 13771 18380 17500 18408
rect 13771 18377 13783 18380
rect 13725 18371 13783 18377
rect 17494 18368 17500 18380
rect 17552 18368 17558 18420
rect 17862 18408 17868 18420
rect 17604 18380 17868 18408
rect 14182 18340 14188 18352
rect 2746 18312 14188 18340
rect 2317 18275 2375 18281
rect 2317 18241 2329 18275
rect 2363 18272 2375 18275
rect 2746 18272 2774 18312
rect 14182 18300 14188 18312
rect 14240 18300 14246 18352
rect 15194 18340 15200 18352
rect 14292 18312 15200 18340
rect 13630 18272 13636 18284
rect 2363 18244 2774 18272
rect 13591 18244 13636 18272
rect 2363 18241 2375 18244
rect 2317 18235 2375 18241
rect 13630 18232 13636 18244
rect 13688 18232 13694 18284
rect 14292 18281 14320 18312
rect 15194 18300 15200 18312
rect 15252 18300 15258 18352
rect 16761 18343 16819 18349
rect 16761 18309 16773 18343
rect 16807 18340 16819 18343
rect 17604 18340 17632 18380
rect 17862 18368 17868 18380
rect 17920 18368 17926 18420
rect 18046 18368 18052 18420
rect 18104 18368 18110 18420
rect 18322 18368 18328 18420
rect 18380 18408 18386 18420
rect 19153 18411 19211 18417
rect 19153 18408 19165 18411
rect 18380 18380 19165 18408
rect 18380 18368 18386 18380
rect 19153 18377 19165 18380
rect 19199 18377 19211 18411
rect 19153 18371 19211 18377
rect 20622 18368 20628 18420
rect 20680 18408 20686 18420
rect 21177 18411 21235 18417
rect 21177 18408 21189 18411
rect 20680 18380 21189 18408
rect 20680 18368 20686 18380
rect 21177 18377 21189 18380
rect 21223 18377 21235 18411
rect 21177 18371 21235 18377
rect 22830 18368 22836 18420
rect 22888 18408 22894 18420
rect 23109 18411 23167 18417
rect 23109 18408 23121 18411
rect 22888 18380 23121 18408
rect 22888 18368 22894 18380
rect 23109 18377 23121 18380
rect 23155 18377 23167 18411
rect 24486 18408 24492 18420
rect 24447 18380 24492 18408
rect 23109 18371 23167 18377
rect 24486 18368 24492 18380
rect 24544 18368 24550 18420
rect 26878 18368 26884 18420
rect 26936 18408 26942 18420
rect 26973 18411 27031 18417
rect 26973 18408 26985 18411
rect 26936 18380 26985 18408
rect 26936 18368 26942 18380
rect 26973 18377 26985 18380
rect 27019 18377 27031 18411
rect 26973 18371 27031 18377
rect 18064 18340 18092 18368
rect 18785 18343 18843 18349
rect 18785 18340 18797 18343
rect 16807 18312 17632 18340
rect 17696 18312 18797 18340
rect 16807 18309 16819 18312
rect 16761 18303 16819 18309
rect 14277 18275 14335 18281
rect 14277 18241 14289 18275
rect 14323 18241 14335 18275
rect 14277 18235 14335 18241
rect 14544 18275 14602 18281
rect 14544 18241 14556 18275
rect 14590 18272 14602 18275
rect 15286 18272 15292 18284
rect 14590 18244 15292 18272
rect 14590 18241 14602 18244
rect 14544 18235 14602 18241
rect 15286 18232 15292 18244
rect 15344 18232 15350 18284
rect 16669 18275 16727 18281
rect 16669 18241 16681 18275
rect 16715 18272 16727 18275
rect 16850 18272 16856 18284
rect 16715 18244 16856 18272
rect 16715 18241 16727 18244
rect 16669 18235 16727 18241
rect 16850 18232 16856 18244
rect 16908 18232 16914 18284
rect 17310 18272 17316 18284
rect 17271 18244 17316 18272
rect 17310 18232 17316 18244
rect 17368 18232 17374 18284
rect 17494 18272 17500 18284
rect 17455 18244 17500 18272
rect 17494 18232 17500 18244
rect 17552 18232 17558 18284
rect 17696 18281 17724 18312
rect 18785 18309 18797 18312
rect 18831 18340 18843 18343
rect 19242 18340 19248 18352
rect 18831 18312 19248 18340
rect 18831 18309 18843 18312
rect 18785 18303 18843 18309
rect 19242 18300 19248 18312
rect 19300 18300 19306 18352
rect 22738 18340 22744 18352
rect 22699 18312 22744 18340
rect 22738 18300 22744 18312
rect 22796 18300 22802 18352
rect 22941 18343 22999 18349
rect 22941 18340 22953 18343
rect 22848 18312 22953 18340
rect 17681 18275 17739 18281
rect 17681 18241 17693 18275
rect 17727 18241 17739 18275
rect 17862 18272 17868 18284
rect 17823 18244 17868 18272
rect 17681 18235 17739 18241
rect 17862 18232 17868 18244
rect 17920 18232 17926 18284
rect 18049 18275 18107 18281
rect 18049 18241 18061 18275
rect 18095 18272 18107 18275
rect 18509 18275 18567 18281
rect 18509 18272 18521 18275
rect 18095 18244 18521 18272
rect 18095 18241 18107 18244
rect 18049 18235 18107 18241
rect 18509 18241 18521 18244
rect 18555 18241 18567 18275
rect 18509 18235 18567 18241
rect 18602 18275 18660 18281
rect 18602 18241 18614 18275
rect 18648 18241 18660 18275
rect 18874 18272 18880 18284
rect 18835 18244 18880 18272
rect 18602 18235 18660 18241
rect 17589 18207 17647 18213
rect 17589 18173 17601 18207
rect 17635 18204 17647 18207
rect 18138 18204 18144 18216
rect 17635 18176 18144 18204
rect 17635 18173 17647 18176
rect 17589 18167 17647 18173
rect 18138 18164 18144 18176
rect 18196 18164 18202 18216
rect 15378 18096 15384 18148
rect 15436 18136 15442 18148
rect 15657 18139 15715 18145
rect 15657 18136 15669 18139
rect 15436 18108 15669 18136
rect 15436 18096 15442 18108
rect 15657 18105 15669 18108
rect 15703 18105 15715 18139
rect 18616 18136 18644 18235
rect 18874 18232 18880 18244
rect 18932 18232 18938 18284
rect 19015 18275 19073 18281
rect 19015 18241 19027 18275
rect 19061 18272 19073 18275
rect 19061 18244 19288 18272
rect 19061 18241 19073 18244
rect 19015 18235 19073 18241
rect 19260 18204 19288 18244
rect 19334 18232 19340 18284
rect 19392 18272 19398 18284
rect 19797 18275 19855 18281
rect 19797 18272 19809 18275
rect 19392 18244 19809 18272
rect 19392 18232 19398 18244
rect 19797 18241 19809 18244
rect 19843 18241 19855 18275
rect 19797 18235 19855 18241
rect 19886 18232 19892 18284
rect 19944 18232 19950 18284
rect 20070 18281 20076 18284
rect 20064 18235 20076 18281
rect 20128 18272 20134 18284
rect 20128 18244 20164 18272
rect 20070 18232 20076 18235
rect 20128 18232 20134 18244
rect 21818 18232 21824 18284
rect 21876 18272 21882 18284
rect 22005 18275 22063 18281
rect 22005 18272 22017 18275
rect 21876 18244 22017 18272
rect 21876 18232 21882 18244
rect 22005 18241 22017 18244
rect 22051 18241 22063 18275
rect 22005 18235 22063 18241
rect 22186 18232 22192 18284
rect 22244 18272 22250 18284
rect 22848 18272 22876 18312
rect 22941 18309 22953 18312
rect 22987 18309 22999 18343
rect 22941 18303 22999 18309
rect 24121 18343 24179 18349
rect 24121 18309 24133 18343
rect 24167 18340 24179 18343
rect 24854 18340 24860 18352
rect 24167 18312 24860 18340
rect 24167 18309 24179 18312
rect 24121 18303 24179 18309
rect 24854 18300 24860 18312
rect 24912 18300 24918 18352
rect 27798 18340 27804 18352
rect 26160 18312 27804 18340
rect 24302 18272 24308 18284
rect 22244 18244 22876 18272
rect 24263 18244 24308 18272
rect 22244 18232 22250 18244
rect 24302 18232 24308 18244
rect 24360 18232 24366 18284
rect 24578 18272 24584 18284
rect 24539 18244 24584 18272
rect 24578 18232 24584 18244
rect 24636 18232 24642 18284
rect 24762 18232 24768 18284
rect 24820 18272 24826 18284
rect 25038 18272 25044 18284
rect 24820 18244 25044 18272
rect 24820 18232 24826 18244
rect 25038 18232 25044 18244
rect 25096 18232 25102 18284
rect 25308 18275 25366 18281
rect 25308 18241 25320 18275
rect 25354 18272 25366 18275
rect 26050 18272 26056 18284
rect 25354 18244 26056 18272
rect 25354 18241 25366 18244
rect 25308 18235 25366 18241
rect 26050 18232 26056 18244
rect 26108 18232 26114 18284
rect 19904 18204 19932 18232
rect 22278 18204 22284 18216
rect 19260 18176 19932 18204
rect 22239 18176 22284 18204
rect 22278 18164 22284 18176
rect 22336 18164 22342 18216
rect 15657 18099 15715 18105
rect 17880 18108 18644 18136
rect 17880 18080 17908 18108
rect 1854 18068 1860 18080
rect 1815 18040 1860 18068
rect 1854 18028 1860 18040
rect 1912 18028 1918 18080
rect 2406 18068 2412 18080
rect 2367 18040 2412 18068
rect 2406 18028 2412 18040
rect 2464 18028 2470 18080
rect 14550 18028 14556 18080
rect 14608 18068 14614 18080
rect 17862 18068 17868 18080
rect 14608 18040 17868 18068
rect 14608 18028 14614 18040
rect 17862 18028 17868 18040
rect 17920 18028 17926 18080
rect 18322 18028 18328 18080
rect 18380 18068 18386 18080
rect 21450 18068 21456 18080
rect 18380 18040 21456 18068
rect 18380 18028 18386 18040
rect 21450 18028 21456 18040
rect 21508 18028 21514 18080
rect 21818 18068 21824 18080
rect 21779 18040 21824 18068
rect 21818 18028 21824 18040
rect 21876 18028 21882 18080
rect 22186 18068 22192 18080
rect 22147 18040 22192 18068
rect 22186 18028 22192 18040
rect 22244 18028 22250 18080
rect 22278 18028 22284 18080
rect 22336 18068 22342 18080
rect 22925 18071 22983 18077
rect 22925 18068 22937 18071
rect 22336 18040 22937 18068
rect 22336 18028 22342 18040
rect 22925 18037 22937 18040
rect 22971 18037 22983 18071
rect 22925 18031 22983 18037
rect 23382 18028 23388 18080
rect 23440 18068 23446 18080
rect 26160 18068 26188 18312
rect 27798 18300 27804 18312
rect 27856 18300 27862 18352
rect 27157 18275 27215 18281
rect 27157 18241 27169 18275
rect 27203 18272 27215 18275
rect 27614 18272 27620 18284
rect 27203 18244 27620 18272
rect 27203 18241 27215 18244
rect 27157 18235 27215 18241
rect 27614 18232 27620 18244
rect 27672 18232 27678 18284
rect 27893 18275 27951 18281
rect 27893 18241 27905 18275
rect 27939 18241 27951 18275
rect 27893 18235 27951 18241
rect 26418 18164 26424 18216
rect 26476 18204 26482 18216
rect 27433 18207 27491 18213
rect 27433 18204 27445 18207
rect 26476 18176 27445 18204
rect 26476 18164 26482 18176
rect 27433 18173 27445 18176
rect 27479 18173 27491 18207
rect 27908 18204 27936 18235
rect 27433 18167 27491 18173
rect 27540 18176 27936 18204
rect 28169 18207 28227 18213
rect 27540 18136 27568 18176
rect 28169 18173 28181 18207
rect 28215 18204 28227 18207
rect 28258 18204 28264 18216
rect 28215 18176 28264 18204
rect 28215 18173 28227 18176
rect 28169 18167 28227 18173
rect 28258 18164 28264 18176
rect 28316 18164 28322 18216
rect 26988 18108 27568 18136
rect 26988 18080 27016 18108
rect 27614 18096 27620 18148
rect 27672 18136 27678 18148
rect 28077 18139 28135 18145
rect 28077 18136 28089 18139
rect 27672 18108 28089 18136
rect 27672 18096 27678 18108
rect 28077 18105 28089 18108
rect 28123 18105 28135 18139
rect 28077 18099 28135 18105
rect 23440 18040 26188 18068
rect 26421 18071 26479 18077
rect 23440 18028 23446 18040
rect 26421 18037 26433 18071
rect 26467 18068 26479 18071
rect 26970 18068 26976 18080
rect 26467 18040 26976 18068
rect 26467 18037 26479 18040
rect 26421 18031 26479 18037
rect 26970 18028 26976 18040
rect 27028 18028 27034 18080
rect 27062 18028 27068 18080
rect 27120 18068 27126 18080
rect 27338 18068 27344 18080
rect 27120 18040 27344 18068
rect 27120 18028 27126 18040
rect 27338 18028 27344 18040
rect 27396 18028 27402 18080
rect 27982 18068 27988 18080
rect 27943 18040 27988 18068
rect 27982 18028 27988 18040
rect 28040 18028 28046 18080
rect 1104 17978 28888 18000
rect 1104 17926 5582 17978
rect 5634 17926 5646 17978
rect 5698 17926 5710 17978
rect 5762 17926 5774 17978
rect 5826 17926 5838 17978
rect 5890 17926 14846 17978
rect 14898 17926 14910 17978
rect 14962 17926 14974 17978
rect 15026 17926 15038 17978
rect 15090 17926 15102 17978
rect 15154 17926 24110 17978
rect 24162 17926 24174 17978
rect 24226 17926 24238 17978
rect 24290 17926 24302 17978
rect 24354 17926 24366 17978
rect 24418 17926 28888 17978
rect 1104 17904 28888 17926
rect 6270 17824 6276 17876
rect 6328 17864 6334 17876
rect 6328 17836 17080 17864
rect 6328 17824 6334 17836
rect 15381 17799 15439 17805
rect 15381 17765 15393 17799
rect 15427 17796 15439 17799
rect 15654 17796 15660 17808
rect 15427 17768 15660 17796
rect 15427 17765 15439 17768
rect 15381 17759 15439 17765
rect 15654 17756 15660 17768
rect 15712 17756 15718 17808
rect 1397 17731 1455 17737
rect 1397 17697 1409 17731
rect 1443 17728 1455 17731
rect 1854 17728 1860 17740
rect 1443 17700 1860 17728
rect 1443 17697 1455 17700
rect 1397 17691 1455 17697
rect 1854 17688 1860 17700
rect 1912 17688 1918 17740
rect 2774 17688 2780 17740
rect 2832 17728 2838 17740
rect 2832 17700 2877 17728
rect 2832 17688 2838 17700
rect 14734 17688 14740 17740
rect 14792 17728 14798 17740
rect 14921 17731 14979 17737
rect 14921 17728 14933 17731
rect 14792 17700 14933 17728
rect 14792 17688 14798 17700
rect 14921 17697 14933 17700
rect 14967 17697 14979 17731
rect 14921 17691 14979 17697
rect 15194 17688 15200 17740
rect 15252 17728 15258 17740
rect 15838 17728 15844 17740
rect 15252 17700 15844 17728
rect 15252 17688 15258 17700
rect 15838 17688 15844 17700
rect 15896 17688 15902 17740
rect 14550 17620 14556 17672
rect 14608 17660 14614 17672
rect 15013 17663 15071 17669
rect 15013 17660 15025 17663
rect 14608 17632 15025 17660
rect 14608 17620 14614 17632
rect 15013 17629 15025 17632
rect 15059 17629 15071 17663
rect 17052 17660 17080 17836
rect 17126 17824 17132 17876
rect 17184 17864 17190 17876
rect 17221 17867 17279 17873
rect 17221 17864 17233 17867
rect 17184 17836 17233 17864
rect 17184 17824 17190 17836
rect 17221 17833 17233 17836
rect 17267 17833 17279 17867
rect 17221 17827 17279 17833
rect 17236 17728 17264 17827
rect 18230 17824 18236 17876
rect 18288 17864 18294 17876
rect 19429 17867 19487 17873
rect 19429 17864 19441 17867
rect 18288 17836 19441 17864
rect 18288 17824 18294 17836
rect 19429 17833 19441 17836
rect 19475 17833 19487 17867
rect 19429 17827 19487 17833
rect 20441 17867 20499 17873
rect 20441 17833 20453 17867
rect 20487 17864 20499 17867
rect 20714 17864 20720 17876
rect 20487 17836 20720 17864
rect 20487 17833 20499 17836
rect 20441 17827 20499 17833
rect 20714 17824 20720 17836
rect 20772 17864 20778 17876
rect 20990 17864 20996 17876
rect 20772 17836 20996 17864
rect 20772 17824 20778 17836
rect 20990 17824 20996 17836
rect 21048 17824 21054 17876
rect 24762 17864 24768 17876
rect 24412 17836 24768 17864
rect 19334 17756 19340 17808
rect 19392 17796 19398 17808
rect 19613 17799 19671 17805
rect 19613 17796 19625 17799
rect 19392 17768 19625 17796
rect 19392 17756 19398 17768
rect 19613 17765 19625 17768
rect 19659 17765 19671 17799
rect 20254 17796 20260 17808
rect 19613 17759 19671 17765
rect 20180 17768 20260 17796
rect 17681 17731 17739 17737
rect 17681 17728 17693 17731
rect 17236 17700 17693 17728
rect 17681 17697 17693 17700
rect 17727 17697 17739 17731
rect 19628 17728 19656 17759
rect 20180 17728 20208 17768
rect 20254 17756 20260 17768
rect 20312 17756 20318 17808
rect 24412 17740 24440 17836
rect 24762 17824 24768 17836
rect 24820 17824 24826 17876
rect 25314 17824 25320 17876
rect 25372 17864 25378 17876
rect 26326 17864 26332 17876
rect 25372 17836 26332 17864
rect 25372 17824 25378 17836
rect 26326 17824 26332 17836
rect 26384 17824 26390 17876
rect 25777 17799 25835 17805
rect 25777 17765 25789 17799
rect 25823 17765 25835 17799
rect 25777 17759 25835 17765
rect 24302 17728 24308 17740
rect 17681 17691 17739 17697
rect 17788 17700 19564 17728
rect 19628 17700 20208 17728
rect 17788 17660 17816 17700
rect 17052 17632 17816 17660
rect 17957 17663 18015 17669
rect 15013 17623 15071 17629
rect 17957 17629 17969 17663
rect 18003 17660 18015 17663
rect 18230 17660 18236 17672
rect 18003 17632 18236 17660
rect 18003 17629 18015 17632
rect 17957 17623 18015 17629
rect 1581 17595 1639 17601
rect 1581 17561 1593 17595
rect 1627 17592 1639 17595
rect 2406 17592 2412 17604
rect 1627 17564 2412 17592
rect 1627 17561 1639 17564
rect 1581 17555 1639 17561
rect 2406 17552 2412 17564
rect 2464 17552 2470 17604
rect 15654 17552 15660 17604
rect 15712 17592 15718 17604
rect 16086 17595 16144 17601
rect 16086 17592 16098 17595
rect 15712 17564 16098 17592
rect 15712 17552 15718 17564
rect 16086 17561 16098 17564
rect 16132 17561 16144 17595
rect 16086 17555 16144 17561
rect 16482 17552 16488 17604
rect 16540 17592 16546 17604
rect 17494 17592 17500 17604
rect 16540 17564 17500 17592
rect 16540 17552 16546 17564
rect 17494 17552 17500 17564
rect 17552 17592 17558 17604
rect 17972 17592 18000 17623
rect 18230 17620 18236 17632
rect 18288 17620 18294 17672
rect 18414 17620 18420 17672
rect 18472 17660 18478 17672
rect 18472 17632 19472 17660
rect 18472 17620 18478 17632
rect 19242 17592 19248 17604
rect 17552 17564 18000 17592
rect 19203 17564 19248 17592
rect 17552 17552 17558 17564
rect 19242 17552 19248 17564
rect 19300 17552 19306 17604
rect 19444 17533 19472 17632
rect 19536 17592 19564 17700
rect 19886 17620 19892 17672
rect 19944 17660 19950 17672
rect 20073 17663 20131 17669
rect 20073 17660 20085 17663
rect 19944 17632 20085 17660
rect 19944 17620 19950 17632
rect 20073 17629 20085 17632
rect 20119 17629 20131 17663
rect 20180 17660 20208 17700
rect 22066 17700 24308 17728
rect 20243 17663 20301 17669
rect 20243 17660 20255 17663
rect 20180 17632 20255 17660
rect 20073 17623 20131 17629
rect 20243 17629 20255 17632
rect 20289 17629 20301 17663
rect 20990 17660 20996 17672
rect 20951 17632 20996 17660
rect 20243 17623 20301 17629
rect 20990 17620 20996 17632
rect 21048 17620 21054 17672
rect 21260 17663 21318 17669
rect 21260 17629 21272 17663
rect 21306 17660 21318 17663
rect 21818 17660 21824 17672
rect 21306 17632 21824 17660
rect 21306 17629 21318 17632
rect 21260 17623 21318 17629
rect 21818 17620 21824 17632
rect 21876 17620 21882 17672
rect 22066 17592 22094 17700
rect 24302 17688 24308 17700
rect 24360 17688 24366 17740
rect 24394 17688 24400 17740
rect 24452 17728 24458 17740
rect 24452 17700 24545 17728
rect 24452 17688 24458 17700
rect 23566 17660 23572 17672
rect 23527 17632 23572 17660
rect 23566 17620 23572 17632
rect 23624 17620 23630 17672
rect 23750 17660 23756 17672
rect 23711 17632 23756 17660
rect 23750 17620 23756 17632
rect 23808 17620 23814 17672
rect 23845 17663 23903 17669
rect 23845 17629 23857 17663
rect 23891 17660 23903 17663
rect 25682 17660 25688 17672
rect 23891 17632 25688 17660
rect 23891 17629 23903 17632
rect 23845 17623 23903 17629
rect 25682 17620 25688 17632
rect 25740 17660 25746 17672
rect 25792 17660 25820 17759
rect 28166 17728 28172 17740
rect 28127 17700 28172 17728
rect 28166 17688 28172 17700
rect 28224 17688 28230 17740
rect 25740 17632 25820 17660
rect 26329 17663 26387 17669
rect 25740 17620 25746 17632
rect 26329 17629 26341 17663
rect 26375 17629 26387 17663
rect 26329 17623 26387 17629
rect 19536 17564 22094 17592
rect 23385 17595 23443 17601
rect 23385 17561 23397 17595
rect 23431 17592 23443 17595
rect 24642 17595 24700 17601
rect 24642 17592 24654 17595
rect 23431 17564 24654 17592
rect 23431 17561 23443 17564
rect 23385 17555 23443 17561
rect 24642 17561 24654 17564
rect 24688 17561 24700 17595
rect 24642 17555 24700 17561
rect 24762 17552 24768 17604
rect 24820 17592 24826 17604
rect 26344 17592 26372 17623
rect 24820 17564 26372 17592
rect 26513 17595 26571 17601
rect 24820 17552 24826 17564
rect 26513 17561 26525 17595
rect 26559 17592 26571 17595
rect 27062 17592 27068 17604
rect 26559 17564 27068 17592
rect 26559 17561 26571 17564
rect 26513 17555 26571 17561
rect 27062 17552 27068 17564
rect 27120 17552 27126 17604
rect 19444 17527 19503 17533
rect 19444 17496 19457 17527
rect 19445 17493 19457 17496
rect 19491 17493 19503 17527
rect 19445 17487 19503 17493
rect 22278 17484 22284 17536
rect 22336 17524 22342 17536
rect 22373 17527 22431 17533
rect 22373 17524 22385 17527
rect 22336 17496 22385 17524
rect 22336 17484 22342 17496
rect 22373 17493 22385 17496
rect 22419 17493 22431 17527
rect 22373 17487 22431 17493
rect 23750 17484 23756 17536
rect 23808 17524 23814 17536
rect 25590 17524 25596 17536
rect 23808 17496 25596 17524
rect 23808 17484 23814 17496
rect 25590 17484 25596 17496
rect 25648 17484 25654 17536
rect 1104 17434 28888 17456
rect 1104 17382 10214 17434
rect 10266 17382 10278 17434
rect 10330 17382 10342 17434
rect 10394 17382 10406 17434
rect 10458 17382 10470 17434
rect 10522 17382 19478 17434
rect 19530 17382 19542 17434
rect 19594 17382 19606 17434
rect 19658 17382 19670 17434
rect 19722 17382 19734 17434
rect 19786 17382 28888 17434
rect 1104 17360 28888 17382
rect 15654 17320 15660 17332
rect 15615 17292 15660 17320
rect 15654 17280 15660 17292
rect 15712 17280 15718 17332
rect 19242 17280 19248 17332
rect 19300 17320 19306 17332
rect 19337 17323 19395 17329
rect 19337 17320 19349 17323
rect 19300 17292 19349 17320
rect 19300 17280 19306 17292
rect 19337 17289 19349 17292
rect 19383 17289 19395 17323
rect 19337 17283 19395 17289
rect 19886 17280 19892 17332
rect 19944 17320 19950 17332
rect 21177 17323 21235 17329
rect 21177 17320 21189 17323
rect 19944 17292 21189 17320
rect 19944 17280 19950 17292
rect 21177 17289 21189 17292
rect 21223 17289 21235 17323
rect 21177 17283 21235 17289
rect 22738 17280 22744 17332
rect 22796 17320 22802 17332
rect 23201 17323 23259 17329
rect 23201 17320 23213 17323
rect 22796 17292 23213 17320
rect 22796 17280 22802 17292
rect 23201 17289 23213 17292
rect 23247 17289 23259 17323
rect 23201 17283 23259 17289
rect 23290 17280 23296 17332
rect 23348 17320 23354 17332
rect 23348 17292 25820 17320
rect 23348 17280 23354 17292
rect 16022 17212 16028 17264
rect 16080 17252 16086 17264
rect 17678 17252 17684 17264
rect 16080 17224 17684 17252
rect 16080 17212 16086 17224
rect 17678 17212 17684 17224
rect 17736 17212 17742 17264
rect 18414 17252 18420 17264
rect 18064 17224 18420 17252
rect 15841 17187 15899 17193
rect 15841 17153 15853 17187
rect 15887 17153 15899 17187
rect 15841 17147 15899 17153
rect 1397 17119 1455 17125
rect 1397 17085 1409 17119
rect 1443 17085 1455 17119
rect 1578 17116 1584 17128
rect 1539 17088 1584 17116
rect 1397 17079 1455 17085
rect 1412 17048 1440 17079
rect 1578 17076 1584 17088
rect 1636 17076 1642 17128
rect 1854 17116 1860 17128
rect 1815 17088 1860 17116
rect 1854 17076 1860 17088
rect 1912 17076 1918 17128
rect 2498 17048 2504 17060
rect 1412 17020 2504 17048
rect 2498 17008 2504 17020
rect 2556 17008 2562 17060
rect 15856 17048 15884 17147
rect 15930 17144 15936 17196
rect 15988 17184 15994 17196
rect 17957 17187 18015 17193
rect 17957 17184 17969 17187
rect 15988 17156 17969 17184
rect 15988 17144 15994 17156
rect 17957 17153 17969 17156
rect 18003 17153 18015 17187
rect 17957 17147 18015 17153
rect 16117 17119 16175 17125
rect 16117 17085 16129 17119
rect 16163 17116 16175 17119
rect 16482 17116 16488 17128
rect 16163 17088 16488 17116
rect 16163 17085 16175 17088
rect 16117 17079 16175 17085
rect 16482 17076 16488 17088
rect 16540 17076 16546 17128
rect 16666 17116 16672 17128
rect 16627 17088 16672 17116
rect 16666 17076 16672 17088
rect 16724 17076 16730 17128
rect 16945 17119 17003 17125
rect 16945 17085 16957 17119
rect 16991 17116 17003 17119
rect 18064 17116 18092 17224
rect 18414 17212 18420 17224
rect 18472 17212 18478 17264
rect 20990 17252 20996 17264
rect 19812 17224 20996 17252
rect 18230 17193 18236 17196
rect 18224 17184 18236 17193
rect 18191 17156 18236 17184
rect 18224 17147 18236 17156
rect 18230 17144 18236 17147
rect 18288 17144 18294 17196
rect 19812 17193 19840 17224
rect 20990 17212 20996 17224
rect 21048 17252 21054 17264
rect 24486 17252 24492 17264
rect 21048 17224 24492 17252
rect 21048 17212 21054 17224
rect 19797 17187 19855 17193
rect 19797 17153 19809 17187
rect 19843 17153 19855 17187
rect 19797 17147 19855 17153
rect 20064 17187 20122 17193
rect 20064 17153 20076 17187
rect 20110 17184 20122 17187
rect 20438 17184 20444 17196
rect 20110 17156 20444 17184
rect 20110 17153 20122 17156
rect 20064 17147 20122 17153
rect 20438 17144 20444 17156
rect 20496 17144 20502 17196
rect 21836 17193 21864 17224
rect 21821 17187 21879 17193
rect 21821 17153 21833 17187
rect 21867 17153 21879 17187
rect 21821 17147 21879 17153
rect 22088 17187 22146 17193
rect 22088 17153 22100 17187
rect 22134 17184 22146 17187
rect 22462 17184 22468 17196
rect 22134 17156 22468 17184
rect 22134 17153 22146 17156
rect 22088 17147 22146 17153
rect 22462 17144 22468 17156
rect 22520 17144 22526 17196
rect 23676 17193 23704 17224
rect 24486 17212 24492 17224
rect 24544 17212 24550 17264
rect 25498 17252 25504 17264
rect 25459 17224 25504 17252
rect 25498 17212 25504 17224
rect 25556 17212 25562 17264
rect 25590 17212 25596 17264
rect 25648 17252 25654 17264
rect 25701 17255 25759 17261
rect 25701 17252 25713 17255
rect 25648 17224 25713 17252
rect 25648 17212 25654 17224
rect 25701 17221 25713 17224
rect 25747 17221 25759 17255
rect 25792 17252 25820 17292
rect 28077 17255 28135 17261
rect 28077 17252 28089 17255
rect 25792 17224 28089 17252
rect 25701 17215 25759 17221
rect 28077 17221 28089 17224
rect 28123 17221 28135 17255
rect 28077 17215 28135 17221
rect 23661 17187 23719 17193
rect 23661 17153 23673 17187
rect 23707 17153 23719 17187
rect 23661 17147 23719 17153
rect 23750 17144 23756 17196
rect 23808 17184 23814 17196
rect 23917 17187 23975 17193
rect 23917 17184 23929 17187
rect 23808 17156 23929 17184
rect 23808 17144 23814 17156
rect 23917 17153 23929 17156
rect 23963 17153 23975 17187
rect 27157 17187 27215 17193
rect 27157 17184 27169 17187
rect 23917 17147 23975 17153
rect 25884 17156 27169 17184
rect 16991 17088 18092 17116
rect 16991 17085 17003 17088
rect 16945 17079 17003 17085
rect 16850 17048 16856 17060
rect 15856 17020 16856 17048
rect 16850 17008 16856 17020
rect 16908 17008 16914 17060
rect 16960 16992 16988 17079
rect 16025 16983 16083 16989
rect 16025 16949 16037 16983
rect 16071 16980 16083 16983
rect 16942 16980 16948 16992
rect 16071 16952 16948 16980
rect 16071 16949 16083 16952
rect 16025 16943 16083 16949
rect 16942 16940 16948 16952
rect 17000 16940 17006 16992
rect 17770 16940 17776 16992
rect 17828 16980 17834 16992
rect 21634 16980 21640 16992
rect 17828 16952 21640 16980
rect 17828 16940 17834 16952
rect 21634 16940 21640 16952
rect 21692 16940 21698 16992
rect 23382 16940 23388 16992
rect 23440 16980 23446 16992
rect 25041 16983 25099 16989
rect 25041 16980 25053 16983
rect 23440 16952 25053 16980
rect 23440 16940 23446 16952
rect 25041 16949 25053 16952
rect 25087 16949 25099 16983
rect 25682 16980 25688 16992
rect 25643 16952 25688 16980
rect 25041 16943 25099 16949
rect 25682 16940 25688 16952
rect 25740 16940 25746 16992
rect 25884 16989 25912 17156
rect 27157 17153 27169 17156
rect 27203 17184 27215 17187
rect 27801 17187 27859 17193
rect 27801 17184 27813 17187
rect 27203 17156 27813 17184
rect 27203 17153 27215 17156
rect 27157 17147 27215 17153
rect 27801 17153 27813 17156
rect 27847 17184 27859 17187
rect 27982 17184 27988 17196
rect 27847 17156 27988 17184
rect 27847 17153 27859 17156
rect 27801 17147 27859 17153
rect 27982 17144 27988 17156
rect 28040 17144 28046 17196
rect 26970 17116 26976 17128
rect 26931 17088 26976 17116
rect 26970 17076 26976 17088
rect 27028 17076 27034 17128
rect 27522 17076 27528 17128
rect 27580 17116 27586 17128
rect 27893 17119 27951 17125
rect 27893 17116 27905 17119
rect 27580 17088 27905 17116
rect 27580 17076 27586 17088
rect 27893 17085 27905 17088
rect 27939 17085 27951 17119
rect 27893 17079 27951 17085
rect 26142 17008 26148 17060
rect 26200 17048 26206 17060
rect 27801 17051 27859 17057
rect 27801 17048 27813 17051
rect 26200 17020 27813 17048
rect 26200 17008 26206 17020
rect 27801 17017 27813 17020
rect 27847 17017 27859 17051
rect 27801 17011 27859 17017
rect 25869 16983 25927 16989
rect 25869 16949 25881 16983
rect 25915 16949 25927 16983
rect 25869 16943 25927 16949
rect 26694 16940 26700 16992
rect 26752 16980 26758 16992
rect 27338 16980 27344 16992
rect 26752 16952 27344 16980
rect 26752 16940 26758 16952
rect 27338 16940 27344 16952
rect 27396 16940 27402 16992
rect 1104 16890 28888 16912
rect 1104 16838 5582 16890
rect 5634 16838 5646 16890
rect 5698 16838 5710 16890
rect 5762 16838 5774 16890
rect 5826 16838 5838 16890
rect 5890 16838 14846 16890
rect 14898 16838 14910 16890
rect 14962 16838 14974 16890
rect 15026 16838 15038 16890
rect 15090 16838 15102 16890
rect 15154 16838 24110 16890
rect 24162 16838 24174 16890
rect 24226 16838 24238 16890
rect 24290 16838 24302 16890
rect 24354 16838 24366 16890
rect 24418 16838 28888 16890
rect 1104 16816 28888 16838
rect 1578 16736 1584 16788
rect 1636 16776 1642 16788
rect 1765 16779 1823 16785
rect 1765 16776 1777 16779
rect 1636 16748 1777 16776
rect 1636 16736 1642 16748
rect 1765 16745 1777 16748
rect 1811 16745 1823 16779
rect 2498 16776 2504 16788
rect 2459 16748 2504 16776
rect 1765 16739 1823 16745
rect 2498 16736 2504 16748
rect 2556 16736 2562 16788
rect 17310 16736 17316 16788
rect 17368 16776 17374 16788
rect 20438 16776 20444 16788
rect 17368 16748 18552 16776
rect 20399 16748 20444 16776
rect 17368 16736 17374 16748
rect 15838 16600 15844 16652
rect 15896 16640 15902 16652
rect 16669 16643 16727 16649
rect 16669 16640 16681 16643
rect 15896 16612 16681 16640
rect 15896 16600 15902 16612
rect 16669 16609 16681 16612
rect 16715 16609 16727 16643
rect 16669 16603 16727 16609
rect 1670 16582 1676 16594
rect 1631 16554 1676 16582
rect 1670 16542 1676 16554
rect 1728 16542 1734 16594
rect 16022 16572 16028 16584
rect 15983 16544 16028 16572
rect 16022 16532 16028 16544
rect 16080 16532 16086 16584
rect 16117 16575 16175 16581
rect 16117 16541 16129 16575
rect 16163 16572 16175 16575
rect 17218 16572 17224 16584
rect 16163 16544 17224 16572
rect 16163 16541 16175 16544
rect 16117 16535 16175 16541
rect 17218 16532 17224 16544
rect 17276 16532 17282 16584
rect 18524 16581 18552 16748
rect 20438 16736 20444 16748
rect 20496 16736 20502 16788
rect 21453 16779 21511 16785
rect 21453 16745 21465 16779
rect 21499 16776 21511 16779
rect 21542 16776 21548 16788
rect 21499 16748 21548 16776
rect 21499 16745 21511 16748
rect 21453 16739 21511 16745
rect 21542 16736 21548 16748
rect 21600 16736 21606 16788
rect 22094 16736 22100 16788
rect 22152 16776 22158 16788
rect 22152 16748 22197 16776
rect 22152 16736 22158 16748
rect 23290 16736 23296 16788
rect 23348 16736 23354 16788
rect 21174 16708 21180 16720
rect 20548 16680 21180 16708
rect 19334 16600 19340 16652
rect 19392 16640 19398 16652
rect 19797 16643 19855 16649
rect 19797 16640 19809 16643
rect 19392 16612 19809 16640
rect 19392 16600 19398 16612
rect 19797 16609 19809 16612
rect 19843 16609 19855 16643
rect 19797 16603 19855 16609
rect 19981 16643 20039 16649
rect 19981 16609 19993 16643
rect 20027 16640 20039 16643
rect 20548 16640 20576 16680
rect 21174 16668 21180 16680
rect 21232 16708 21238 16720
rect 22002 16708 22008 16720
rect 21232 16680 22008 16708
rect 21232 16668 21238 16680
rect 22002 16668 22008 16680
rect 22060 16668 22066 16720
rect 23308 16708 23336 16736
rect 22112 16680 23336 16708
rect 20714 16640 20720 16652
rect 20027 16612 20576 16640
rect 20640 16612 20720 16640
rect 20027 16609 20039 16612
rect 19981 16603 20039 16609
rect 18509 16575 18567 16581
rect 18509 16541 18521 16575
rect 18555 16541 18567 16575
rect 18509 16535 18567 16541
rect 19705 16575 19763 16581
rect 19705 16541 19717 16575
rect 19751 16572 19763 16575
rect 19886 16572 19892 16584
rect 19751 16544 19892 16572
rect 19751 16541 19763 16544
rect 19705 16535 19763 16541
rect 19886 16532 19892 16544
rect 19944 16532 19950 16584
rect 20640 16581 20668 16612
rect 20714 16600 20720 16612
rect 20772 16600 20778 16652
rect 22112 16640 22140 16680
rect 21928 16612 22140 16640
rect 20441 16575 20499 16581
rect 20441 16541 20453 16575
rect 20487 16541 20499 16575
rect 20441 16535 20499 16541
rect 20625 16575 20683 16581
rect 20625 16541 20637 16575
rect 20671 16541 20683 16575
rect 20625 16535 20683 16541
rect 21453 16575 21511 16581
rect 21453 16541 21465 16575
rect 21499 16541 21511 16575
rect 21634 16572 21640 16584
rect 21595 16544 21640 16572
rect 21453 16535 21511 16541
rect 16936 16507 16994 16513
rect 16936 16473 16948 16507
rect 16982 16504 16994 16507
rect 17126 16504 17132 16516
rect 16982 16476 17132 16504
rect 16982 16473 16994 16476
rect 16936 16467 16994 16473
rect 17126 16464 17132 16476
rect 17184 16464 17190 16516
rect 18138 16464 18144 16516
rect 18196 16504 18202 16516
rect 18601 16507 18659 16513
rect 18601 16504 18613 16507
rect 18196 16476 18613 16504
rect 18196 16464 18202 16476
rect 18601 16473 18613 16476
rect 18647 16473 18659 16507
rect 18601 16467 18659 16473
rect 19981 16507 20039 16513
rect 19981 16473 19993 16507
rect 20027 16504 20039 16507
rect 20456 16504 20484 16535
rect 20027 16476 20484 16504
rect 21468 16504 21496 16535
rect 21634 16532 21640 16544
rect 21692 16572 21698 16584
rect 21928 16572 21956 16612
rect 22186 16600 22192 16652
rect 22244 16640 22250 16652
rect 22244 16612 22416 16640
rect 22244 16600 22250 16612
rect 22204 16572 22232 16600
rect 22388 16581 22416 16612
rect 22830 16600 22836 16652
rect 22888 16640 22894 16652
rect 23290 16640 23296 16652
rect 22888 16612 23296 16640
rect 22888 16600 22894 16612
rect 23290 16600 23296 16612
rect 23348 16640 23354 16652
rect 24486 16640 24492 16652
rect 23348 16612 23612 16640
rect 24447 16612 24492 16640
rect 23348 16600 23354 16612
rect 21692 16544 21956 16572
rect 22020 16544 22232 16572
rect 22373 16575 22431 16581
rect 21692 16532 21698 16544
rect 22020 16504 22048 16544
rect 22373 16541 22385 16575
rect 22419 16541 22431 16575
rect 23382 16572 23388 16584
rect 23343 16544 23388 16572
rect 22373 16535 22431 16541
rect 23382 16532 23388 16544
rect 23440 16532 23446 16584
rect 23584 16581 23612 16612
rect 24486 16600 24492 16612
rect 24544 16600 24550 16652
rect 23569 16575 23627 16581
rect 23569 16541 23581 16575
rect 23615 16541 23627 16575
rect 23569 16535 23627 16541
rect 24756 16575 24814 16581
rect 24756 16541 24768 16575
rect 24802 16572 24814 16575
rect 26142 16572 26148 16584
rect 24802 16544 26148 16572
rect 24802 16541 24814 16544
rect 24756 16535 24814 16541
rect 26142 16532 26148 16544
rect 26200 16532 26206 16584
rect 26326 16572 26332 16584
rect 26287 16544 26332 16572
rect 26326 16532 26332 16544
rect 26384 16532 26390 16584
rect 21468 16476 22048 16504
rect 22097 16507 22155 16513
rect 20027 16473 20039 16476
rect 19981 16467 20039 16473
rect 22097 16473 22109 16507
rect 22143 16504 22155 16507
rect 22738 16504 22744 16516
rect 22143 16476 22744 16504
rect 22143 16473 22155 16476
rect 22097 16467 22155 16473
rect 22738 16464 22744 16476
rect 22796 16464 22802 16516
rect 23753 16507 23811 16513
rect 23753 16473 23765 16507
rect 23799 16504 23811 16507
rect 25590 16504 25596 16516
rect 23799 16476 25596 16504
rect 23799 16473 23811 16476
rect 23753 16467 23811 16473
rect 25590 16464 25596 16476
rect 25648 16464 25654 16516
rect 26513 16507 26571 16513
rect 26513 16473 26525 16507
rect 26559 16504 26571 16507
rect 26878 16504 26884 16516
rect 26559 16476 26884 16504
rect 26559 16473 26571 16476
rect 26513 16467 26571 16473
rect 26878 16464 26884 16476
rect 26936 16464 26942 16516
rect 28166 16504 28172 16516
rect 28127 16476 28172 16504
rect 28166 16464 28172 16476
rect 28224 16464 28230 16516
rect 16666 16396 16672 16448
rect 16724 16436 16730 16448
rect 18049 16439 18107 16445
rect 18049 16436 18061 16439
rect 16724 16408 18061 16436
rect 16724 16396 16730 16408
rect 18049 16405 18061 16408
rect 18095 16405 18107 16439
rect 22278 16436 22284 16448
rect 22239 16408 22284 16436
rect 18049 16399 18107 16405
rect 22278 16396 22284 16408
rect 22336 16396 22342 16448
rect 23014 16396 23020 16448
rect 23072 16436 23078 16448
rect 24854 16436 24860 16448
rect 23072 16408 24860 16436
rect 23072 16396 23078 16408
rect 24854 16396 24860 16408
rect 24912 16396 24918 16448
rect 25130 16396 25136 16448
rect 25188 16436 25194 16448
rect 25498 16436 25504 16448
rect 25188 16408 25504 16436
rect 25188 16396 25194 16408
rect 25498 16396 25504 16408
rect 25556 16436 25562 16448
rect 25869 16439 25927 16445
rect 25869 16436 25881 16439
rect 25556 16408 25881 16436
rect 25556 16396 25562 16408
rect 25869 16405 25881 16408
rect 25915 16405 25927 16439
rect 25869 16399 25927 16405
rect 1104 16346 28888 16368
rect 1104 16294 10214 16346
rect 10266 16294 10278 16346
rect 10330 16294 10342 16346
rect 10394 16294 10406 16346
rect 10458 16294 10470 16346
rect 10522 16294 19478 16346
rect 19530 16294 19542 16346
rect 19594 16294 19606 16346
rect 19658 16294 19670 16346
rect 19722 16294 19734 16346
rect 19786 16294 28888 16346
rect 1104 16272 28888 16294
rect 16482 16192 16488 16244
rect 16540 16232 16546 16244
rect 17037 16235 17095 16241
rect 17037 16232 17049 16235
rect 16540 16204 17049 16232
rect 16540 16192 16546 16204
rect 17037 16201 17049 16204
rect 17083 16201 17095 16235
rect 17037 16195 17095 16201
rect 18141 16235 18199 16241
rect 18141 16201 18153 16235
rect 18187 16232 18199 16235
rect 18230 16232 18236 16244
rect 18187 16204 18236 16232
rect 18187 16201 18199 16204
rect 18141 16195 18199 16201
rect 18230 16192 18236 16204
rect 18288 16192 18294 16244
rect 20070 16192 20076 16244
rect 20128 16232 20134 16244
rect 20165 16235 20223 16241
rect 20165 16232 20177 16235
rect 20128 16204 20177 16232
rect 20128 16192 20134 16204
rect 20165 16201 20177 16204
rect 20211 16201 20223 16235
rect 20898 16232 20904 16244
rect 20859 16204 20904 16232
rect 20165 16195 20223 16201
rect 20898 16192 20904 16204
rect 20956 16192 20962 16244
rect 22189 16235 22247 16241
rect 22189 16201 22201 16235
rect 22235 16232 22247 16235
rect 22922 16232 22928 16244
rect 22235 16204 22928 16232
rect 22235 16201 22247 16204
rect 22189 16195 22247 16201
rect 22922 16192 22928 16204
rect 22980 16192 22986 16244
rect 24670 16192 24676 16244
rect 24728 16232 24734 16244
rect 27525 16235 27583 16241
rect 27525 16232 27537 16235
rect 24728 16204 27537 16232
rect 24728 16192 24734 16204
rect 27525 16201 27537 16204
rect 27571 16201 27583 16235
rect 27525 16195 27583 16201
rect 16758 16124 16764 16176
rect 16816 16164 16822 16176
rect 16853 16167 16911 16173
rect 16853 16164 16865 16167
rect 16816 16136 16865 16164
rect 16816 16124 16822 16136
rect 16853 16133 16865 16136
rect 16899 16133 16911 16167
rect 16853 16127 16911 16133
rect 18417 16167 18475 16173
rect 18417 16133 18429 16167
rect 18463 16164 18475 16167
rect 20530 16164 20536 16176
rect 18463 16136 20536 16164
rect 18463 16133 18475 16136
rect 18417 16127 18475 16133
rect 20530 16124 20536 16136
rect 20588 16124 20594 16176
rect 22554 16164 22560 16176
rect 22020 16136 22560 16164
rect 16942 16056 16948 16108
rect 17000 16096 17006 16108
rect 17129 16099 17187 16105
rect 17129 16096 17141 16099
rect 17000 16068 17141 16096
rect 17000 16056 17006 16068
rect 17129 16065 17141 16068
rect 17175 16065 17187 16099
rect 17129 16059 17187 16065
rect 18141 16099 18199 16105
rect 18141 16065 18153 16099
rect 18187 16096 18199 16099
rect 19334 16096 19340 16108
rect 18187 16068 19340 16096
rect 18187 16065 18199 16068
rect 18141 16059 18199 16065
rect 19334 16056 19340 16068
rect 19392 16056 19398 16108
rect 20073 16099 20131 16105
rect 20073 16065 20085 16099
rect 20119 16096 20131 16099
rect 20162 16096 20168 16108
rect 20119 16068 20168 16096
rect 20119 16065 20131 16068
rect 20073 16059 20131 16065
rect 20162 16056 20168 16068
rect 20220 16056 20226 16108
rect 20257 16099 20315 16105
rect 20257 16065 20269 16099
rect 20303 16096 20315 16099
rect 20346 16096 20352 16108
rect 20303 16068 20352 16096
rect 20303 16065 20315 16068
rect 20257 16059 20315 16065
rect 20346 16056 20352 16068
rect 20404 16056 20410 16108
rect 20806 16096 20812 16108
rect 20767 16068 20812 16096
rect 20806 16056 20812 16068
rect 20864 16056 20870 16108
rect 20993 16099 21051 16105
rect 20993 16065 21005 16099
rect 21039 16096 21051 16099
rect 21358 16096 21364 16108
rect 21039 16068 21364 16096
rect 21039 16065 21051 16068
rect 20993 16059 21051 16065
rect 21358 16056 21364 16068
rect 21416 16056 21422 16108
rect 22020 16105 22048 16136
rect 22554 16124 22560 16136
rect 22612 16124 22618 16176
rect 23198 16124 23204 16176
rect 23256 16164 23262 16176
rect 24765 16167 24823 16173
rect 23256 16136 23796 16164
rect 23256 16124 23262 16136
rect 22005 16099 22063 16105
rect 22005 16065 22017 16099
rect 22051 16065 22063 16099
rect 22005 16059 22063 16065
rect 22189 16099 22247 16105
rect 22189 16065 22201 16099
rect 22235 16096 22247 16099
rect 22370 16096 22376 16108
rect 22235 16068 22376 16096
rect 22235 16065 22247 16068
rect 22189 16059 22247 16065
rect 22370 16056 22376 16068
rect 22428 16056 22434 16108
rect 22649 16099 22707 16105
rect 22649 16065 22661 16099
rect 22695 16096 22707 16099
rect 22738 16096 22744 16108
rect 22695 16068 22744 16096
rect 22695 16065 22707 16068
rect 22649 16059 22707 16065
rect 22738 16056 22744 16068
rect 22796 16056 22802 16108
rect 23293 16099 23351 16105
rect 23293 16065 23305 16099
rect 23339 16096 23351 16099
rect 23382 16096 23388 16108
rect 23339 16068 23388 16096
rect 23339 16065 23351 16068
rect 23293 16059 23351 16065
rect 23382 16056 23388 16068
rect 23440 16056 23446 16108
rect 23658 16096 23664 16108
rect 23492 16068 23664 16096
rect 17954 15988 17960 16040
rect 18012 16028 18018 16040
rect 18233 16031 18291 16037
rect 18233 16028 18245 16031
rect 18012 16000 18245 16028
rect 18012 15988 18018 16000
rect 18233 15997 18245 16000
rect 18279 15997 18291 16031
rect 23492 16028 23520 16068
rect 23658 16056 23664 16068
rect 23716 16056 23722 16108
rect 18233 15991 18291 15997
rect 22756 16000 23520 16028
rect 23569 16031 23627 16037
rect 16850 15960 16856 15972
rect 16811 15932 16856 15960
rect 16850 15920 16856 15932
rect 16908 15920 16914 15972
rect 22756 15969 22784 16000
rect 23569 15997 23581 16031
rect 23615 16028 23627 16031
rect 23768 16028 23796 16136
rect 24765 16133 24777 16167
rect 24811 16164 24823 16167
rect 27338 16164 27344 16176
rect 24811 16136 27344 16164
rect 24811 16133 24823 16136
rect 24765 16127 24823 16133
rect 27338 16124 27344 16136
rect 27396 16124 27402 16176
rect 27433 16099 27491 16105
rect 27433 16096 27445 16099
rect 25976 16068 27445 16096
rect 24578 16028 24584 16040
rect 23615 16000 23796 16028
rect 24539 16000 24584 16028
rect 23615 15997 23627 16000
rect 23569 15991 23627 15997
rect 22741 15963 22799 15969
rect 22741 15929 22753 15963
rect 22787 15929 22799 15963
rect 22741 15923 22799 15929
rect 23290 15920 23296 15972
rect 23348 15960 23354 15972
rect 23385 15963 23443 15969
rect 23385 15960 23397 15963
rect 23348 15932 23397 15960
rect 23348 15920 23354 15932
rect 23385 15929 23397 15932
rect 23431 15929 23443 15963
rect 23584 15960 23612 15991
rect 24578 15988 24584 16000
rect 24636 15988 24642 16040
rect 24854 15988 24860 16040
rect 24912 16028 24918 16040
rect 25976 16028 26004 16068
rect 27433 16065 27445 16068
rect 27479 16096 27491 16099
rect 27982 16096 27988 16108
rect 27479 16068 27988 16096
rect 27479 16065 27491 16068
rect 27433 16059 27491 16065
rect 27982 16056 27988 16068
rect 28040 16056 28046 16108
rect 26142 16028 26148 16040
rect 24912 16000 26004 16028
rect 26103 16000 26148 16028
rect 24912 15988 24918 16000
rect 26142 15988 26148 16000
rect 26200 15988 26206 16040
rect 28258 15960 28264 15972
rect 23584 15932 28264 15960
rect 23385 15923 23443 15929
rect 28258 15920 28264 15932
rect 28316 15920 28322 15972
rect 1394 15852 1400 15904
rect 1452 15892 1458 15904
rect 1581 15895 1639 15901
rect 1581 15892 1593 15895
rect 1452 15864 1593 15892
rect 1452 15852 1458 15864
rect 1581 15861 1593 15864
rect 1627 15861 1639 15895
rect 1581 15855 1639 15861
rect 23474 15852 23480 15904
rect 23532 15892 23538 15904
rect 23532 15864 23577 15892
rect 23532 15852 23538 15864
rect 1104 15802 28888 15824
rect 1104 15750 5582 15802
rect 5634 15750 5646 15802
rect 5698 15750 5710 15802
rect 5762 15750 5774 15802
rect 5826 15750 5838 15802
rect 5890 15750 14846 15802
rect 14898 15750 14910 15802
rect 14962 15750 14974 15802
rect 15026 15750 15038 15802
rect 15090 15750 15102 15802
rect 15154 15750 24110 15802
rect 24162 15750 24174 15802
rect 24226 15750 24238 15802
rect 24290 15750 24302 15802
rect 24354 15750 24366 15802
rect 24418 15750 28888 15802
rect 1104 15728 28888 15750
rect 17126 15688 17132 15700
rect 17087 15660 17132 15688
rect 17126 15648 17132 15660
rect 17184 15648 17190 15700
rect 22925 15691 22983 15697
rect 22925 15657 22937 15691
rect 22971 15688 22983 15691
rect 23658 15688 23664 15700
rect 22971 15660 23664 15688
rect 22971 15657 22983 15660
rect 22925 15651 22983 15657
rect 23658 15648 23664 15660
rect 23716 15648 23722 15700
rect 25133 15691 25191 15697
rect 25133 15657 25145 15691
rect 25179 15688 25191 15691
rect 27522 15688 27528 15700
rect 25179 15660 27528 15688
rect 25179 15657 25191 15660
rect 25133 15651 25191 15657
rect 27522 15648 27528 15660
rect 27580 15648 27586 15700
rect 22465 15623 22523 15629
rect 22465 15589 22477 15623
rect 22511 15620 22523 15623
rect 23845 15623 23903 15629
rect 22511 15592 23612 15620
rect 22511 15589 22523 15592
rect 22465 15583 22523 15589
rect 1394 15552 1400 15564
rect 1355 15524 1400 15552
rect 1394 15512 1400 15524
rect 1452 15512 1458 15564
rect 2774 15512 2780 15564
rect 2832 15552 2838 15564
rect 23474 15552 23480 15564
rect 2832 15524 2877 15552
rect 22940 15524 23480 15552
rect 2832 15512 2838 15524
rect 16942 15444 16948 15496
rect 17000 15484 17006 15496
rect 17129 15487 17187 15493
rect 17129 15484 17141 15487
rect 17000 15456 17141 15484
rect 17000 15444 17006 15456
rect 17129 15453 17141 15456
rect 17175 15453 17187 15487
rect 17129 15447 17187 15453
rect 17313 15487 17371 15493
rect 17313 15453 17325 15487
rect 17359 15484 17371 15487
rect 17770 15484 17776 15496
rect 17359 15456 17776 15484
rect 17359 15453 17371 15456
rect 17313 15447 17371 15453
rect 17770 15444 17776 15456
rect 17828 15444 17834 15496
rect 22940 15493 22968 15524
rect 23474 15512 23480 15524
rect 23532 15512 23538 15564
rect 23584 15552 23612 15592
rect 23845 15589 23857 15623
rect 23891 15620 23903 15623
rect 24486 15620 24492 15632
rect 23891 15592 24492 15620
rect 23891 15589 23903 15592
rect 23845 15583 23903 15589
rect 24486 15580 24492 15592
rect 24544 15580 24550 15632
rect 26326 15580 26332 15632
rect 26384 15580 26390 15632
rect 26344 15552 26372 15580
rect 23584 15524 26372 15552
rect 22925 15487 22983 15493
rect 22925 15453 22937 15487
rect 22971 15453 22983 15487
rect 22925 15447 22983 15453
rect 23109 15487 23167 15493
rect 23109 15453 23121 15487
rect 23155 15484 23167 15487
rect 24673 15487 24731 15493
rect 24673 15484 24685 15487
rect 23155 15456 24685 15484
rect 23155 15453 23167 15456
rect 23109 15447 23167 15453
rect 24673 15453 24685 15456
rect 24719 15484 24731 15487
rect 25409 15487 25467 15493
rect 25409 15484 25421 15487
rect 24719 15456 25421 15484
rect 24719 15453 24731 15456
rect 24673 15447 24731 15453
rect 25409 15453 25421 15456
rect 25455 15484 25467 15487
rect 25590 15484 25596 15496
rect 25455 15456 25596 15484
rect 25455 15453 25467 15456
rect 25409 15447 25467 15453
rect 25590 15444 25596 15456
rect 25648 15444 25654 15496
rect 26326 15484 26332 15496
rect 26287 15456 26332 15484
rect 26326 15444 26332 15456
rect 26384 15444 26390 15496
rect 1578 15416 1584 15428
rect 1539 15388 1584 15416
rect 1578 15376 1584 15388
rect 1636 15376 1642 15428
rect 13814 15376 13820 15428
rect 13872 15416 13878 15428
rect 23661 15419 23719 15425
rect 23661 15416 23673 15419
rect 13872 15388 23673 15416
rect 13872 15376 13878 15388
rect 23661 15385 23673 15388
rect 23707 15385 23719 15419
rect 23661 15379 23719 15385
rect 23842 15376 23848 15428
rect 23900 15416 23906 15428
rect 24397 15419 24455 15425
rect 24397 15416 24409 15419
rect 23900 15388 24409 15416
rect 23900 15376 23906 15388
rect 24397 15385 24409 15388
rect 24443 15385 24455 15419
rect 25130 15416 25136 15428
rect 25091 15388 25136 15416
rect 24397 15379 24455 15385
rect 25130 15376 25136 15388
rect 25188 15376 25194 15428
rect 25317 15419 25375 15425
rect 25317 15385 25329 15419
rect 25363 15416 25375 15419
rect 25682 15416 25688 15428
rect 25363 15388 25688 15416
rect 25363 15385 25375 15388
rect 25317 15379 25375 15385
rect 23566 15308 23572 15360
rect 23624 15348 23630 15360
rect 24495 15351 24553 15357
rect 24495 15348 24507 15351
rect 23624 15320 24507 15348
rect 23624 15308 23630 15320
rect 24495 15317 24507 15320
rect 24541 15317 24553 15351
rect 24495 15311 24553 15317
rect 24581 15351 24639 15357
rect 24581 15317 24593 15351
rect 24627 15348 24639 15351
rect 24854 15348 24860 15360
rect 24627 15320 24860 15348
rect 24627 15317 24639 15320
rect 24581 15311 24639 15317
rect 24854 15308 24860 15320
rect 24912 15348 24918 15360
rect 25332 15348 25360 15379
rect 25682 15376 25688 15388
rect 25740 15376 25746 15428
rect 26510 15416 26516 15428
rect 26471 15388 26516 15416
rect 26510 15376 26516 15388
rect 26568 15376 26574 15428
rect 28166 15416 28172 15428
rect 28127 15388 28172 15416
rect 28166 15376 28172 15388
rect 28224 15376 28230 15428
rect 24912 15320 25360 15348
rect 24912 15308 24918 15320
rect 1104 15258 28888 15280
rect 1104 15206 10214 15258
rect 10266 15206 10278 15258
rect 10330 15206 10342 15258
rect 10394 15206 10406 15258
rect 10458 15206 10470 15258
rect 10522 15206 19478 15258
rect 19530 15206 19542 15258
rect 19594 15206 19606 15258
rect 19658 15206 19670 15258
rect 19722 15206 19734 15258
rect 19786 15206 28888 15258
rect 1104 15184 28888 15206
rect 1578 15104 1584 15156
rect 1636 15144 1642 15156
rect 1673 15147 1731 15153
rect 1673 15144 1685 15147
rect 1636 15116 1685 15144
rect 1636 15104 1642 15116
rect 1673 15113 1685 15116
rect 1719 15113 1731 15147
rect 1673 15107 1731 15113
rect 23753 15147 23811 15153
rect 23753 15113 23765 15147
rect 23799 15144 23811 15147
rect 23934 15144 23940 15156
rect 23799 15116 23940 15144
rect 23799 15113 23811 15116
rect 23753 15107 23811 15113
rect 23934 15104 23940 15116
rect 23992 15104 23998 15156
rect 25038 15144 25044 15156
rect 24999 15116 25044 15144
rect 25038 15104 25044 15116
rect 25096 15104 25102 15156
rect 25685 15147 25743 15153
rect 25685 15113 25697 15147
rect 25731 15144 25743 15147
rect 26234 15144 26240 15156
rect 25731 15116 26240 15144
rect 25731 15113 25743 15116
rect 25685 15107 25743 15113
rect 26234 15104 26240 15116
rect 26292 15104 26298 15156
rect 26329 15147 26387 15153
rect 26329 15113 26341 15147
rect 26375 15144 26387 15147
rect 26510 15144 26516 15156
rect 26375 15116 26516 15144
rect 26375 15113 26387 15116
rect 26329 15107 26387 15113
rect 26510 15104 26516 15116
rect 26568 15104 26574 15156
rect 27062 15104 27068 15156
rect 27120 15144 27126 15156
rect 27157 15147 27215 15153
rect 27157 15144 27169 15147
rect 27120 15116 27169 15144
rect 27120 15104 27126 15116
rect 27157 15113 27169 15116
rect 27203 15113 27215 15147
rect 27157 15107 27215 15113
rect 25222 15036 25228 15088
rect 25280 15076 25286 15088
rect 28534 15076 28540 15088
rect 25280 15048 25728 15076
rect 25280 15036 25286 15048
rect 1486 14968 1492 15020
rect 1544 15008 1550 15020
rect 1581 15011 1639 15017
rect 1581 15008 1593 15011
rect 1544 14980 1593 15008
rect 1544 14968 1550 14980
rect 1581 14977 1593 14980
rect 1627 14977 1639 15011
rect 1581 14971 1639 14977
rect 23382 14968 23388 15020
rect 23440 15008 23446 15020
rect 23661 15011 23719 15017
rect 23661 15008 23673 15011
rect 23440 14980 23673 15008
rect 23440 14968 23446 14980
rect 23661 14977 23673 14980
rect 23707 14977 23719 15011
rect 23661 14971 23719 14977
rect 24489 15011 24547 15017
rect 24489 14977 24501 15011
rect 24535 15008 24547 15011
rect 24762 15008 24768 15020
rect 24535 14980 24768 15008
rect 24535 14977 24547 14980
rect 24489 14971 24547 14977
rect 24762 14968 24768 14980
rect 24820 14968 24826 15020
rect 24949 15011 25007 15017
rect 24949 14977 24961 15011
rect 24995 15008 25007 15011
rect 25130 15008 25136 15020
rect 24995 14980 25136 15008
rect 24995 14977 25007 14980
rect 24949 14971 25007 14977
rect 25130 14968 25136 14980
rect 25188 14968 25194 15020
rect 25593 15011 25651 15017
rect 25593 14977 25605 15011
rect 25639 14977 25651 15011
rect 25593 14971 25651 14977
rect 25038 14900 25044 14952
rect 25096 14940 25102 14952
rect 25608 14940 25636 14971
rect 25096 14912 25636 14940
rect 25700 14940 25728 15048
rect 26252 15048 28540 15076
rect 26252 15017 26280 15048
rect 28534 15036 28540 15048
rect 28592 15036 28598 15088
rect 26237 15011 26295 15017
rect 26237 14977 26249 15011
rect 26283 14977 26295 15011
rect 26237 14971 26295 14977
rect 27065 15011 27123 15017
rect 27065 14977 27077 15011
rect 27111 15008 27123 15011
rect 27246 15008 27252 15020
rect 27111 14980 27252 15008
rect 27111 14977 27123 14980
rect 27065 14971 27123 14977
rect 27246 14968 27252 14980
rect 27304 14968 27310 15020
rect 27709 15011 27767 15017
rect 27709 14977 27721 15011
rect 27755 14977 27767 15011
rect 27709 14971 27767 14977
rect 27724 14940 27752 14971
rect 25700 14912 27752 14940
rect 25096 14900 25102 14912
rect 27798 14900 27804 14952
rect 27856 14940 27862 14952
rect 27985 14943 28043 14949
rect 27985 14940 27997 14943
rect 27856 14912 27997 14940
rect 27856 14900 27862 14912
rect 27985 14909 27997 14912
rect 28031 14909 28043 14943
rect 27985 14903 28043 14909
rect 14458 14832 14464 14884
rect 14516 14872 14522 14884
rect 27893 14875 27951 14881
rect 27893 14872 27905 14875
rect 14516 14844 27905 14872
rect 14516 14832 14522 14844
rect 27893 14841 27905 14844
rect 27939 14841 27951 14875
rect 27893 14835 27951 14841
rect 1394 14764 1400 14816
rect 1452 14804 1458 14816
rect 2409 14807 2467 14813
rect 2409 14804 2421 14807
rect 1452 14776 2421 14804
rect 1452 14764 1458 14776
rect 2409 14773 2421 14776
rect 2455 14773 2467 14807
rect 2409 14767 2467 14773
rect 27801 14807 27859 14813
rect 27801 14773 27813 14807
rect 27847 14804 27859 14807
rect 27982 14804 27988 14816
rect 27847 14776 27988 14804
rect 27847 14773 27859 14776
rect 27801 14767 27859 14773
rect 27982 14764 27988 14776
rect 28040 14764 28046 14816
rect 1104 14714 28888 14736
rect 1104 14662 5582 14714
rect 5634 14662 5646 14714
rect 5698 14662 5710 14714
rect 5762 14662 5774 14714
rect 5826 14662 5838 14714
rect 5890 14662 14846 14714
rect 14898 14662 14910 14714
rect 14962 14662 14974 14714
rect 15026 14662 15038 14714
rect 15090 14662 15102 14714
rect 15154 14662 24110 14714
rect 24162 14662 24174 14714
rect 24226 14662 24238 14714
rect 24290 14662 24302 14714
rect 24354 14662 24366 14714
rect 24418 14662 28888 14714
rect 1104 14640 28888 14662
rect 24946 14600 24952 14612
rect 24907 14572 24952 14600
rect 24946 14560 24952 14572
rect 25004 14560 25010 14612
rect 25685 14603 25743 14609
rect 25685 14569 25697 14603
rect 25731 14600 25743 14603
rect 25866 14600 25872 14612
rect 25731 14572 25872 14600
rect 25731 14569 25743 14572
rect 25685 14563 25743 14569
rect 25866 14560 25872 14572
rect 25924 14560 25930 14612
rect 23845 14535 23903 14541
rect 23845 14501 23857 14535
rect 23891 14532 23903 14535
rect 25314 14532 25320 14544
rect 23891 14504 25320 14532
rect 23891 14501 23903 14504
rect 23845 14495 23903 14501
rect 25314 14492 25320 14504
rect 25372 14492 25378 14544
rect 26418 14532 26424 14544
rect 25608 14504 26424 14532
rect 1394 14464 1400 14476
rect 1355 14436 1400 14464
rect 1394 14424 1400 14436
rect 1452 14424 1458 14476
rect 1854 14464 1860 14476
rect 1815 14436 1860 14464
rect 1854 14424 1860 14436
rect 1912 14424 1918 14476
rect 7650 14424 7656 14476
rect 7708 14464 7714 14476
rect 9950 14464 9956 14476
rect 7708 14436 9956 14464
rect 7708 14424 7714 14436
rect 9950 14424 9956 14436
rect 10008 14424 10014 14476
rect 24854 14396 24860 14408
rect 24815 14368 24860 14396
rect 24854 14356 24860 14368
rect 24912 14356 24918 14408
rect 25608 14405 25636 14504
rect 26418 14492 26424 14504
rect 26476 14492 26482 14544
rect 26329 14467 26387 14473
rect 26329 14433 26341 14467
rect 26375 14464 26387 14467
rect 28074 14464 28080 14476
rect 26375 14436 28080 14464
rect 26375 14433 26387 14436
rect 26329 14427 26387 14433
rect 28074 14424 28080 14436
rect 28132 14424 28138 14476
rect 25593 14399 25651 14405
rect 25593 14365 25605 14399
rect 25639 14365 25651 14399
rect 25593 14359 25651 14365
rect 1578 14328 1584 14340
rect 1539 14300 1584 14328
rect 1578 14288 1584 14300
rect 1636 14288 1642 14340
rect 26513 14331 26571 14337
rect 26513 14297 26525 14331
rect 26559 14328 26571 14331
rect 27798 14328 27804 14340
rect 26559 14300 27804 14328
rect 26559 14297 26571 14300
rect 26513 14291 26571 14297
rect 27798 14288 27804 14300
rect 27856 14288 27862 14340
rect 28166 14328 28172 14340
rect 28127 14300 28172 14328
rect 28166 14288 28172 14300
rect 28224 14288 28230 14340
rect 1104 14170 28888 14192
rect 1104 14118 10214 14170
rect 10266 14118 10278 14170
rect 10330 14118 10342 14170
rect 10394 14118 10406 14170
rect 10458 14118 10470 14170
rect 10522 14118 19478 14170
rect 19530 14118 19542 14170
rect 19594 14118 19606 14170
rect 19658 14118 19670 14170
rect 19722 14118 19734 14170
rect 19786 14118 28888 14170
rect 1104 14096 28888 14118
rect 1578 14016 1584 14068
rect 1636 14056 1642 14068
rect 1857 14059 1915 14065
rect 1857 14056 1869 14059
rect 1636 14028 1869 14056
rect 1636 14016 1642 14028
rect 1857 14025 1869 14028
rect 1903 14025 1915 14059
rect 25774 14056 25780 14068
rect 25735 14028 25780 14056
rect 1857 14019 1915 14025
rect 25774 14016 25780 14028
rect 25832 14016 25838 14068
rect 26878 14016 26884 14068
rect 26936 14056 26942 14068
rect 27157 14059 27215 14065
rect 27157 14056 27169 14059
rect 26936 14028 27169 14056
rect 26936 14016 26942 14028
rect 27157 14025 27169 14028
rect 27203 14025 27215 14059
rect 27798 14056 27804 14068
rect 27759 14028 27804 14056
rect 27157 14019 27215 14025
rect 27798 14016 27804 14028
rect 27856 14016 27862 14068
rect 1765 13923 1823 13929
rect 1765 13889 1777 13923
rect 1811 13920 1823 13923
rect 1854 13920 1860 13932
rect 1811 13892 1860 13920
rect 1811 13889 1823 13892
rect 1765 13883 1823 13889
rect 1854 13880 1860 13892
rect 1912 13880 1918 13932
rect 25225 13923 25283 13929
rect 25225 13889 25237 13923
rect 25271 13920 25283 13923
rect 25406 13920 25412 13932
rect 25271 13892 25412 13920
rect 25271 13889 25283 13892
rect 25225 13883 25283 13889
rect 25406 13880 25412 13892
rect 25464 13880 25470 13932
rect 25685 13923 25743 13929
rect 25685 13889 25697 13923
rect 25731 13920 25743 13923
rect 26970 13920 26976 13932
rect 25731 13892 26976 13920
rect 25731 13889 25743 13892
rect 25685 13883 25743 13889
rect 26970 13880 26976 13892
rect 27028 13880 27034 13932
rect 27065 13923 27123 13929
rect 27065 13889 27077 13923
rect 27111 13889 27123 13923
rect 27065 13883 27123 13889
rect 12986 13812 12992 13864
rect 13044 13852 13050 13864
rect 20622 13852 20628 13864
rect 13044 13824 20628 13852
rect 13044 13812 13050 13824
rect 20622 13812 20628 13824
rect 20680 13812 20686 13864
rect 25038 13812 25044 13864
rect 25096 13852 25102 13864
rect 27080 13852 27108 13883
rect 27246 13880 27252 13932
rect 27304 13920 27310 13932
rect 27709 13923 27767 13929
rect 27709 13920 27721 13923
rect 27304 13892 27721 13920
rect 27304 13880 27310 13892
rect 27709 13889 27721 13892
rect 27755 13889 27767 13923
rect 27709 13883 27767 13889
rect 27798 13852 27804 13864
rect 25096 13824 27804 13852
rect 25096 13812 25102 13824
rect 27798 13812 27804 13824
rect 27856 13812 27862 13864
rect 1104 13626 28888 13648
rect 1104 13574 5582 13626
rect 5634 13574 5646 13626
rect 5698 13574 5710 13626
rect 5762 13574 5774 13626
rect 5826 13574 5838 13626
rect 5890 13574 14846 13626
rect 14898 13574 14910 13626
rect 14962 13574 14974 13626
rect 15026 13574 15038 13626
rect 15090 13574 15102 13626
rect 15154 13574 24110 13626
rect 24162 13574 24174 13626
rect 24226 13574 24238 13626
rect 24290 13574 24302 13626
rect 24354 13574 24366 13626
rect 24418 13574 28888 13626
rect 1104 13552 28888 13574
rect 24578 13472 24584 13524
rect 24636 13512 24642 13524
rect 25593 13515 25651 13521
rect 25593 13512 25605 13515
rect 24636 13484 25605 13512
rect 24636 13472 24642 13484
rect 25593 13481 25605 13484
rect 25639 13481 25651 13515
rect 26050 13512 26056 13524
rect 26011 13484 26056 13512
rect 25593 13475 25651 13481
rect 26050 13472 26056 13484
rect 26108 13472 26114 13524
rect 27154 13512 27160 13524
rect 27115 13484 27160 13512
rect 27154 13472 27160 13484
rect 27212 13472 27218 13524
rect 27338 13472 27344 13524
rect 27396 13512 27402 13524
rect 27893 13515 27951 13521
rect 27893 13512 27905 13515
rect 27396 13484 27905 13512
rect 27396 13472 27402 13484
rect 27893 13481 27905 13484
rect 27939 13481 27951 13515
rect 27893 13475 27951 13481
rect 27614 13376 27620 13388
rect 26068 13348 27620 13376
rect 1486 13268 1492 13320
rect 1544 13308 1550 13320
rect 1581 13311 1639 13317
rect 1581 13308 1593 13311
rect 1544 13280 1593 13308
rect 1544 13268 1550 13280
rect 1581 13277 1593 13280
rect 1627 13277 1639 13311
rect 2406 13308 2412 13320
rect 2367 13280 2412 13308
rect 1581 13271 1639 13277
rect 2406 13268 2412 13280
rect 2464 13268 2470 13320
rect 26068 13317 26096 13348
rect 27614 13336 27620 13348
rect 27672 13336 27678 13388
rect 3053 13311 3111 13317
rect 3053 13308 3065 13311
rect 2746 13280 3065 13308
rect 1394 13200 1400 13252
rect 1452 13240 1458 13252
rect 2746 13240 2774 13280
rect 3053 13277 3065 13280
rect 3099 13277 3111 13311
rect 3053 13271 3111 13277
rect 26053 13311 26111 13317
rect 26053 13277 26065 13311
rect 26099 13277 26111 13311
rect 26053 13271 26111 13277
rect 26237 13311 26295 13317
rect 26237 13277 26249 13311
rect 26283 13308 26295 13311
rect 26694 13308 26700 13320
rect 26283 13280 26700 13308
rect 26283 13277 26295 13280
rect 26237 13271 26295 13277
rect 26694 13268 26700 13280
rect 26752 13268 26758 13320
rect 27341 13311 27399 13317
rect 27341 13277 27353 13311
rect 27387 13277 27399 13311
rect 27798 13308 27804 13320
rect 27759 13280 27804 13308
rect 27341 13271 27399 13277
rect 1452 13212 2774 13240
rect 1452 13200 1458 13212
rect 25958 13200 25964 13252
rect 26016 13240 26022 13252
rect 27356 13240 27384 13271
rect 27798 13268 27804 13280
rect 27856 13268 27862 13320
rect 26016 13212 27384 13240
rect 26016 13200 26022 13212
rect 1578 13132 1584 13184
rect 1636 13172 1642 13184
rect 1673 13175 1731 13181
rect 1673 13172 1685 13175
rect 1636 13144 1685 13172
rect 1636 13132 1642 13144
rect 1673 13141 1685 13144
rect 1719 13141 1731 13175
rect 1673 13135 1731 13141
rect 1104 13082 28888 13104
rect 1104 13030 10214 13082
rect 10266 13030 10278 13082
rect 10330 13030 10342 13082
rect 10394 13030 10406 13082
rect 10458 13030 10470 13082
rect 10522 13030 19478 13082
rect 19530 13030 19542 13082
rect 19594 13030 19606 13082
rect 19658 13030 19670 13082
rect 19722 13030 19734 13082
rect 19786 13030 28888 13082
rect 1104 13008 28888 13030
rect 1578 12900 1584 12912
rect 1539 12872 1584 12900
rect 1578 12860 1584 12872
rect 1636 12860 1642 12912
rect 1394 12832 1400 12844
rect 1355 12804 1400 12832
rect 1394 12792 1400 12804
rect 1452 12792 1458 12844
rect 26326 12792 26332 12844
rect 26384 12832 26390 12844
rect 26421 12835 26479 12841
rect 26421 12832 26433 12835
rect 26384 12804 26433 12832
rect 26384 12792 26390 12804
rect 26421 12801 26433 12804
rect 26467 12801 26479 12835
rect 27430 12832 27436 12844
rect 27391 12804 27436 12832
rect 26421 12795 26479 12801
rect 27430 12792 27436 12804
rect 27488 12792 27494 12844
rect 2774 12724 2780 12776
rect 2832 12764 2838 12776
rect 2832 12736 2877 12764
rect 2832 12724 2838 12736
rect 26786 12724 26792 12776
rect 26844 12764 26850 12776
rect 28077 12767 28135 12773
rect 28077 12764 28089 12767
rect 26844 12736 28089 12764
rect 26844 12724 26850 12736
rect 28077 12733 28089 12736
rect 28123 12733 28135 12767
rect 28077 12727 28135 12733
rect 1104 12538 28888 12560
rect 1104 12486 5582 12538
rect 5634 12486 5646 12538
rect 5698 12486 5710 12538
rect 5762 12486 5774 12538
rect 5826 12486 5838 12538
rect 5890 12486 14846 12538
rect 14898 12486 14910 12538
rect 14962 12486 14974 12538
rect 15026 12486 15038 12538
rect 15090 12486 15102 12538
rect 15154 12486 24110 12538
rect 24162 12486 24174 12538
rect 24226 12486 24238 12538
rect 24290 12486 24302 12538
rect 24354 12486 24366 12538
rect 24418 12486 28888 12538
rect 1104 12464 28888 12486
rect 28074 12424 28080 12436
rect 28035 12396 28080 12424
rect 28074 12384 28080 12396
rect 28132 12384 28138 12436
rect 1397 12291 1455 12297
rect 1397 12257 1409 12291
rect 1443 12288 1455 12291
rect 2406 12288 2412 12300
rect 1443 12260 2412 12288
rect 1443 12257 1455 12260
rect 1397 12251 1455 12257
rect 2406 12248 2412 12260
rect 2464 12248 2470 12300
rect 2774 12248 2780 12300
rect 2832 12288 2838 12300
rect 2832 12260 2877 12288
rect 2832 12248 2838 12260
rect 26326 12180 26332 12232
rect 26384 12220 26390 12232
rect 27433 12223 27491 12229
rect 27433 12220 27445 12223
rect 26384 12192 27445 12220
rect 26384 12180 26390 12192
rect 27433 12189 27445 12192
rect 27479 12189 27491 12223
rect 27433 12183 27491 12189
rect 1581 12155 1639 12161
rect 1581 12121 1593 12155
rect 1627 12152 1639 12155
rect 2498 12152 2504 12164
rect 1627 12124 2504 12152
rect 1627 12121 1639 12124
rect 1581 12115 1639 12121
rect 2498 12112 2504 12124
rect 2556 12112 2562 12164
rect 1104 11994 28888 12016
rect 1104 11942 10214 11994
rect 10266 11942 10278 11994
rect 10330 11942 10342 11994
rect 10394 11942 10406 11994
rect 10458 11942 10470 11994
rect 10522 11942 19478 11994
rect 19530 11942 19542 11994
rect 19594 11942 19606 11994
rect 19658 11942 19670 11994
rect 19722 11942 19734 11994
rect 19786 11942 28888 11994
rect 1104 11920 28888 11942
rect 2498 11880 2504 11892
rect 2459 11852 2504 11880
rect 2498 11840 2504 11852
rect 2556 11840 2562 11892
rect 1765 11747 1823 11753
rect 1765 11713 1777 11747
rect 1811 11713 1823 11747
rect 1765 11707 1823 11713
rect 2409 11747 2467 11753
rect 2409 11713 2421 11747
rect 2455 11744 2467 11747
rect 3694 11744 3700 11756
rect 2455 11716 3700 11744
rect 2455 11713 2467 11716
rect 2409 11707 2467 11713
rect 1780 11676 1808 11707
rect 3694 11704 3700 11716
rect 3752 11744 3758 11756
rect 7282 11744 7288 11756
rect 3752 11716 7288 11744
rect 3752 11704 3758 11716
rect 7282 11704 7288 11716
rect 7340 11704 7346 11756
rect 23750 11704 23756 11756
rect 23808 11744 23814 11756
rect 27249 11747 27307 11753
rect 27249 11744 27261 11747
rect 23808 11716 27261 11744
rect 23808 11704 23814 11716
rect 27249 11713 27261 11716
rect 27295 11713 27307 11747
rect 27982 11744 27988 11756
rect 27943 11716 27988 11744
rect 27249 11707 27307 11713
rect 27982 11704 27988 11716
rect 28040 11704 28046 11756
rect 1854 11676 1860 11688
rect 1767 11648 1860 11676
rect 1854 11636 1860 11648
rect 1912 11676 1918 11688
rect 12986 11676 12992 11688
rect 1912 11648 12992 11676
rect 1912 11636 1918 11648
rect 12986 11636 12992 11648
rect 13044 11636 13050 11688
rect 10134 11568 10140 11620
rect 10192 11608 10198 11620
rect 28169 11611 28227 11617
rect 28169 11608 28181 11611
rect 10192 11580 28181 11608
rect 10192 11568 10198 11580
rect 28169 11577 28181 11580
rect 28215 11577 28227 11611
rect 28169 11571 28227 11577
rect 1578 11500 1584 11552
rect 1636 11540 1642 11552
rect 1857 11543 1915 11549
rect 1857 11540 1869 11543
rect 1636 11512 1869 11540
rect 1636 11500 1642 11512
rect 1857 11509 1869 11512
rect 1903 11509 1915 11543
rect 3234 11540 3240 11552
rect 3195 11512 3240 11540
rect 1857 11503 1915 11509
rect 3234 11500 3240 11512
rect 3292 11500 3298 11552
rect 26510 11500 26516 11552
rect 26568 11540 26574 11552
rect 27341 11543 27399 11549
rect 27341 11540 27353 11543
rect 26568 11512 27353 11540
rect 26568 11500 26574 11512
rect 27341 11509 27353 11512
rect 27387 11509 27399 11543
rect 27341 11503 27399 11509
rect 1104 11450 28888 11472
rect 1104 11398 5582 11450
rect 5634 11398 5646 11450
rect 5698 11398 5710 11450
rect 5762 11398 5774 11450
rect 5826 11398 5838 11450
rect 5890 11398 14846 11450
rect 14898 11398 14910 11450
rect 14962 11398 14974 11450
rect 15026 11398 15038 11450
rect 15090 11398 15102 11450
rect 15154 11398 24110 11450
rect 24162 11398 24174 11450
rect 24226 11398 24238 11450
rect 24290 11398 24302 11450
rect 24354 11398 24366 11450
rect 24418 11398 28888 11450
rect 1104 11376 28888 11398
rect 3234 11268 3240 11280
rect 1412 11240 3240 11268
rect 1412 11209 1440 11240
rect 3234 11228 3240 11240
rect 3292 11228 3298 11280
rect 1397 11203 1455 11209
rect 1397 11169 1409 11203
rect 1443 11169 1455 11203
rect 1578 11200 1584 11212
rect 1539 11172 1584 11200
rect 1397 11163 1455 11169
rect 1578 11160 1584 11172
rect 1636 11160 1642 11212
rect 1854 11200 1860 11212
rect 1815 11172 1860 11200
rect 1854 11160 1860 11172
rect 1912 11160 1918 11212
rect 26326 11200 26332 11212
rect 26287 11172 26332 11200
rect 26326 11160 26332 11172
rect 26384 11160 26390 11212
rect 26510 11200 26516 11212
rect 26471 11172 26516 11200
rect 26510 11160 26516 11172
rect 26568 11160 26574 11212
rect 3970 11132 3976 11144
rect 3931 11104 3976 11132
rect 3970 11092 3976 11104
rect 4028 11092 4034 11144
rect 28166 11064 28172 11076
rect 28127 11036 28172 11064
rect 28166 11024 28172 11036
rect 28224 11024 28230 11076
rect 1104 10906 28888 10928
rect 1104 10854 10214 10906
rect 10266 10854 10278 10906
rect 10330 10854 10342 10906
rect 10394 10854 10406 10906
rect 10458 10854 10470 10906
rect 10522 10854 19478 10906
rect 19530 10854 19542 10906
rect 19594 10854 19606 10906
rect 19658 10854 19670 10906
rect 19722 10854 19734 10906
rect 19786 10854 28888 10906
rect 1104 10832 28888 10854
rect 3970 10724 3976 10736
rect 1504 10696 3976 10724
rect 1504 10665 1532 10696
rect 3970 10684 3976 10696
rect 4028 10684 4034 10736
rect 1489 10659 1547 10665
rect 1489 10625 1501 10659
rect 1535 10625 1547 10659
rect 1489 10619 1547 10625
rect 17218 10616 17224 10668
rect 17276 10656 17282 10668
rect 27801 10659 27859 10665
rect 27801 10656 27813 10659
rect 17276 10628 27813 10656
rect 17276 10616 17282 10628
rect 27801 10625 27813 10628
rect 27847 10625 27859 10659
rect 27801 10619 27859 10625
rect 1673 10591 1731 10597
rect 1673 10557 1685 10591
rect 1719 10588 1731 10591
rect 1946 10588 1952 10600
rect 1719 10560 1952 10588
rect 1719 10557 1731 10560
rect 1673 10551 1731 10557
rect 1946 10548 1952 10560
rect 2004 10548 2010 10600
rect 2866 10588 2872 10600
rect 2827 10560 2872 10588
rect 2866 10548 2872 10560
rect 2924 10548 2930 10600
rect 27338 10452 27344 10464
rect 27299 10424 27344 10452
rect 27338 10412 27344 10424
rect 27396 10412 27402 10464
rect 27890 10452 27896 10464
rect 27851 10424 27896 10452
rect 27890 10412 27896 10424
rect 27948 10412 27954 10464
rect 1104 10362 28888 10384
rect 1104 10310 5582 10362
rect 5634 10310 5646 10362
rect 5698 10310 5710 10362
rect 5762 10310 5774 10362
rect 5826 10310 5838 10362
rect 5890 10310 14846 10362
rect 14898 10310 14910 10362
rect 14962 10310 14974 10362
rect 15026 10310 15038 10362
rect 15090 10310 15102 10362
rect 15154 10310 24110 10362
rect 24162 10310 24174 10362
rect 24226 10310 24238 10362
rect 24290 10310 24302 10362
rect 24354 10310 24366 10362
rect 24418 10310 28888 10362
rect 1104 10288 28888 10310
rect 1946 10248 1952 10260
rect 1907 10220 1952 10248
rect 1946 10208 1952 10220
rect 2004 10208 2010 10260
rect 26513 10115 26571 10121
rect 26513 10081 26525 10115
rect 26559 10112 26571 10115
rect 27890 10112 27896 10124
rect 26559 10084 27896 10112
rect 26559 10081 26571 10084
rect 26513 10075 26571 10081
rect 27890 10072 27896 10084
rect 27948 10072 27954 10124
rect 1857 10047 1915 10053
rect 1857 10013 1869 10047
rect 1903 10044 1915 10047
rect 2038 10044 2044 10056
rect 1903 10016 2044 10044
rect 1903 10013 1915 10016
rect 1857 10007 1915 10013
rect 2038 10004 2044 10016
rect 2096 10004 2102 10056
rect 26326 10044 26332 10056
rect 26287 10016 26332 10044
rect 26326 10004 26332 10016
rect 26384 10004 26390 10056
rect 27430 9936 27436 9988
rect 27488 9976 27494 9988
rect 28169 9979 28227 9985
rect 28169 9976 28181 9979
rect 27488 9948 28181 9976
rect 27488 9936 27494 9948
rect 28169 9945 28181 9948
rect 28215 9945 28227 9979
rect 28169 9939 28227 9945
rect 1104 9818 28888 9840
rect 1104 9766 10214 9818
rect 10266 9766 10278 9818
rect 10330 9766 10342 9818
rect 10394 9766 10406 9818
rect 10458 9766 10470 9818
rect 10522 9766 19478 9818
rect 19530 9766 19542 9818
rect 19594 9766 19606 9818
rect 19658 9766 19670 9818
rect 19722 9766 19734 9818
rect 19786 9766 28888 9818
rect 1104 9744 28888 9766
rect 5442 9596 5448 9648
rect 5500 9636 5506 9648
rect 24854 9636 24860 9648
rect 5500 9608 24860 9636
rect 5500 9596 5506 9608
rect 24854 9596 24860 9608
rect 24912 9596 24918 9648
rect 1486 9528 1492 9580
rect 1544 9568 1550 9580
rect 1581 9571 1639 9577
rect 1581 9568 1593 9571
rect 1544 9540 1593 9568
rect 1544 9528 1550 9540
rect 1581 9537 1593 9540
rect 1627 9537 1639 9571
rect 1581 9531 1639 9537
rect 26326 9528 26332 9580
rect 26384 9568 26390 9580
rect 27249 9571 27307 9577
rect 27249 9568 27261 9571
rect 26384 9540 27261 9568
rect 26384 9528 26390 9540
rect 27249 9537 27261 9540
rect 27295 9537 27307 9571
rect 27706 9568 27712 9580
rect 27667 9540 27712 9568
rect 27249 9531 27307 9537
rect 27706 9528 27712 9540
rect 27764 9528 27770 9580
rect 1578 9324 1584 9376
rect 1636 9364 1642 9376
rect 1673 9367 1731 9373
rect 1673 9364 1685 9367
rect 1636 9336 1685 9364
rect 1636 9324 1642 9336
rect 1673 9333 1685 9336
rect 1719 9333 1731 9367
rect 2406 9364 2412 9376
rect 2367 9336 2412 9364
rect 1673 9327 1731 9333
rect 2406 9324 2412 9336
rect 2464 9324 2470 9376
rect 27798 9364 27804 9376
rect 27759 9336 27804 9364
rect 27798 9324 27804 9336
rect 27856 9324 27862 9376
rect 1104 9274 28888 9296
rect 1104 9222 5582 9274
rect 5634 9222 5646 9274
rect 5698 9222 5710 9274
rect 5762 9222 5774 9274
rect 5826 9222 5838 9274
rect 5890 9222 14846 9274
rect 14898 9222 14910 9274
rect 14962 9222 14974 9274
rect 15026 9222 15038 9274
rect 15090 9222 15102 9274
rect 15154 9222 24110 9274
rect 24162 9222 24174 9274
rect 24226 9222 24238 9274
rect 24290 9222 24302 9274
rect 24354 9222 24366 9274
rect 24418 9222 28888 9274
rect 1104 9200 28888 9222
rect 2406 9092 2412 9104
rect 1412 9064 2412 9092
rect 1412 9033 1440 9064
rect 2406 9052 2412 9064
rect 2464 9052 2470 9104
rect 27338 9092 27344 9104
rect 26344 9064 27344 9092
rect 1397 9027 1455 9033
rect 1397 8993 1409 9027
rect 1443 8993 1455 9027
rect 1578 9024 1584 9036
rect 1539 8996 1584 9024
rect 1397 8987 1455 8993
rect 1578 8984 1584 8996
rect 1636 8984 1642 9036
rect 2774 8984 2780 9036
rect 2832 9024 2838 9036
rect 26344 9033 26372 9064
rect 27338 9052 27344 9064
rect 27396 9052 27402 9104
rect 26329 9027 26387 9033
rect 2832 8996 2877 9024
rect 2832 8984 2838 8996
rect 26329 8993 26341 9027
rect 26375 8993 26387 9027
rect 26329 8987 26387 8993
rect 26513 9027 26571 9033
rect 26513 8993 26525 9027
rect 26559 9024 26571 9027
rect 27798 9024 27804 9036
rect 26559 8996 27804 9024
rect 26559 8993 26571 8996
rect 26513 8987 26571 8993
rect 27798 8984 27804 8996
rect 27856 8984 27862 9036
rect 28166 9024 28172 9036
rect 28127 8996 28172 9024
rect 28166 8984 28172 8996
rect 28224 8984 28230 9036
rect 1104 8730 28888 8752
rect 1104 8678 10214 8730
rect 10266 8678 10278 8730
rect 10330 8678 10342 8730
rect 10394 8678 10406 8730
rect 10458 8678 10470 8730
rect 10522 8678 19478 8730
rect 19530 8678 19542 8730
rect 19594 8678 19606 8730
rect 19658 8678 19670 8730
rect 19722 8678 19734 8730
rect 19786 8678 28888 8730
rect 1104 8656 28888 8678
rect 1854 8480 1860 8492
rect 1815 8452 1860 8480
rect 1854 8440 1860 8452
rect 1912 8440 1918 8492
rect 2501 8483 2559 8489
rect 2501 8449 2513 8483
rect 2547 8480 2559 8483
rect 5442 8480 5448 8492
rect 2547 8452 5448 8480
rect 2547 8449 2559 8452
rect 2501 8443 2559 8449
rect 5442 8440 5448 8452
rect 5500 8440 5506 8492
rect 21358 8372 21364 8424
rect 21416 8412 21422 8424
rect 27982 8412 27988 8424
rect 21416 8384 27988 8412
rect 21416 8372 21422 8384
rect 27982 8372 27988 8384
rect 28040 8372 28046 8424
rect 27614 8304 27620 8356
rect 27672 8344 27678 8356
rect 27893 8347 27951 8353
rect 27893 8344 27905 8347
rect 27672 8316 27905 8344
rect 27672 8304 27678 8316
rect 27893 8313 27905 8316
rect 27939 8313 27951 8347
rect 27893 8307 27951 8313
rect 1578 8236 1584 8288
rect 1636 8276 1642 8288
rect 1949 8279 2007 8285
rect 1949 8276 1961 8279
rect 1636 8248 1961 8276
rect 1636 8236 1642 8248
rect 1949 8245 1961 8248
rect 1995 8245 2007 8279
rect 1949 8239 2007 8245
rect 2130 8236 2136 8288
rect 2188 8276 2194 8288
rect 2593 8279 2651 8285
rect 2593 8276 2605 8279
rect 2188 8248 2605 8276
rect 2188 8236 2194 8248
rect 2593 8245 2605 8248
rect 2639 8245 2651 8279
rect 3326 8276 3332 8288
rect 3287 8248 3332 8276
rect 2593 8239 2651 8245
rect 3326 8236 3332 8248
rect 3384 8236 3390 8288
rect 27246 8276 27252 8288
rect 27207 8248 27252 8276
rect 27246 8236 27252 8248
rect 27304 8236 27310 8288
rect 1104 8186 28888 8208
rect 1104 8134 5582 8186
rect 5634 8134 5646 8186
rect 5698 8134 5710 8186
rect 5762 8134 5774 8186
rect 5826 8134 5838 8186
rect 5890 8134 14846 8186
rect 14898 8134 14910 8186
rect 14962 8134 14974 8186
rect 15026 8134 15038 8186
rect 15090 8134 15102 8186
rect 15154 8134 24110 8186
rect 24162 8134 24174 8186
rect 24226 8134 24238 8186
rect 24290 8134 24302 8186
rect 24354 8134 24366 8186
rect 24418 8134 28888 8186
rect 1104 8112 28888 8134
rect 3326 8004 3332 8016
rect 1412 7976 3332 8004
rect 1412 7945 1440 7976
rect 3326 7964 3332 7976
rect 3384 7964 3390 8016
rect 1397 7939 1455 7945
rect 1397 7905 1409 7939
rect 1443 7905 1455 7939
rect 1578 7936 1584 7948
rect 1539 7908 1584 7936
rect 1397 7899 1455 7905
rect 1578 7896 1584 7908
rect 1636 7896 1642 7948
rect 2774 7896 2780 7948
rect 2832 7936 2838 7948
rect 26329 7939 26387 7945
rect 2832 7908 2877 7936
rect 2832 7896 2838 7908
rect 26329 7905 26341 7939
rect 26375 7936 26387 7939
rect 27246 7936 27252 7948
rect 26375 7908 27252 7936
rect 26375 7905 26387 7908
rect 26329 7899 26387 7905
rect 27246 7896 27252 7908
rect 27304 7896 27310 7948
rect 3973 7871 4031 7877
rect 3973 7868 3985 7871
rect 3160 7840 3985 7868
rect 1946 7760 1952 7812
rect 2004 7800 2010 7812
rect 3160 7800 3188 7840
rect 3973 7837 3985 7840
rect 4019 7837 4031 7871
rect 3973 7831 4031 7837
rect 2004 7772 3188 7800
rect 26513 7803 26571 7809
rect 2004 7760 2010 7772
rect 26513 7769 26525 7803
rect 26559 7800 26571 7803
rect 27798 7800 27804 7812
rect 26559 7772 27804 7800
rect 26559 7769 26571 7772
rect 26513 7763 26571 7769
rect 27798 7760 27804 7772
rect 27856 7760 27862 7812
rect 28166 7800 28172 7812
rect 28127 7772 28172 7800
rect 28166 7760 28172 7772
rect 28224 7760 28230 7812
rect 1104 7642 28888 7664
rect 1104 7590 10214 7642
rect 10266 7590 10278 7642
rect 10330 7590 10342 7642
rect 10394 7590 10406 7642
rect 10458 7590 10470 7642
rect 10522 7590 19478 7642
rect 19530 7590 19542 7642
rect 19594 7590 19606 7642
rect 19658 7590 19670 7642
rect 19722 7590 19734 7642
rect 19786 7590 28888 7642
rect 1104 7568 28888 7590
rect 27798 7528 27804 7540
rect 27759 7500 27804 7528
rect 27798 7488 27804 7500
rect 27856 7488 27862 7540
rect 2130 7460 2136 7472
rect 2091 7432 2136 7460
rect 2130 7420 2136 7432
rect 2188 7420 2194 7472
rect 1946 7392 1952 7404
rect 1907 7364 1952 7392
rect 1946 7352 1952 7364
rect 2004 7352 2010 7404
rect 27706 7392 27712 7404
rect 27667 7364 27712 7392
rect 27706 7352 27712 7364
rect 27764 7352 27770 7404
rect 2958 7324 2964 7336
rect 2919 7296 2964 7324
rect 2958 7284 2964 7296
rect 3016 7284 3022 7336
rect 4430 7188 4436 7200
rect 4391 7160 4436 7188
rect 4430 7148 4436 7160
rect 4488 7148 4494 7200
rect 27246 7188 27252 7200
rect 27207 7160 27252 7188
rect 27246 7148 27252 7160
rect 27304 7148 27310 7200
rect 1104 7098 28888 7120
rect 1104 7046 5582 7098
rect 5634 7046 5646 7098
rect 5698 7046 5710 7098
rect 5762 7046 5774 7098
rect 5826 7046 5838 7098
rect 5890 7046 14846 7098
rect 14898 7046 14910 7098
rect 14962 7046 14974 7098
rect 15026 7046 15038 7098
rect 15090 7046 15102 7098
rect 15154 7046 24110 7098
rect 24162 7046 24174 7098
rect 24226 7046 24238 7098
rect 24290 7046 24302 7098
rect 24354 7046 24366 7098
rect 24418 7046 28888 7098
rect 1104 7024 28888 7046
rect 1397 6851 1455 6857
rect 1397 6817 1409 6851
rect 1443 6848 1455 6851
rect 1443 6820 2820 6848
rect 1443 6817 1455 6820
rect 1397 6811 1455 6817
rect 1581 6715 1639 6721
rect 1581 6681 1593 6715
rect 1627 6712 1639 6715
rect 2590 6712 2596 6724
rect 1627 6684 2596 6712
rect 1627 6681 1639 6684
rect 1581 6675 1639 6681
rect 2590 6672 2596 6684
rect 2648 6672 2654 6724
rect 2792 6712 2820 6820
rect 2866 6808 2872 6860
rect 2924 6848 2930 6860
rect 26329 6851 26387 6857
rect 2924 6820 2969 6848
rect 3804 6820 12434 6848
rect 2924 6808 2930 6820
rect 3804 6789 3832 6820
rect 3789 6783 3847 6789
rect 3789 6749 3801 6783
rect 3835 6749 3847 6783
rect 3789 6743 3847 6749
rect 4617 6783 4675 6789
rect 4617 6749 4629 6783
rect 4663 6749 4675 6783
rect 12406 6780 12434 6820
rect 26329 6817 26341 6851
rect 26375 6848 26387 6851
rect 27246 6848 27252 6860
rect 26375 6820 27252 6848
rect 26375 6817 26387 6820
rect 26329 6811 26387 6817
rect 27246 6808 27252 6820
rect 27304 6808 27310 6860
rect 28166 6848 28172 6860
rect 28127 6820 28172 6848
rect 28166 6808 28172 6820
rect 28224 6808 28230 6860
rect 13998 6780 14004 6792
rect 12406 6752 14004 6780
rect 4617 6743 4675 6749
rect 4632 6712 4660 6743
rect 13998 6740 14004 6752
rect 14056 6740 14062 6792
rect 2792 6684 4660 6712
rect 26513 6715 26571 6721
rect 26513 6681 26525 6715
rect 26559 6712 26571 6715
rect 27890 6712 27896 6724
rect 26559 6684 27896 6712
rect 26559 6681 26571 6684
rect 26513 6675 26571 6681
rect 27890 6672 27896 6684
rect 27948 6672 27954 6724
rect 3602 6604 3608 6656
rect 3660 6644 3666 6656
rect 3881 6647 3939 6653
rect 3881 6644 3893 6647
rect 3660 6616 3893 6644
rect 3660 6604 3666 6616
rect 3881 6613 3893 6616
rect 3927 6613 3939 6647
rect 3881 6607 3939 6613
rect 1104 6554 28888 6576
rect 1104 6502 10214 6554
rect 10266 6502 10278 6554
rect 10330 6502 10342 6554
rect 10394 6502 10406 6554
rect 10458 6502 10470 6554
rect 10522 6502 19478 6554
rect 19530 6502 19542 6554
rect 19594 6502 19606 6554
rect 19658 6502 19670 6554
rect 19722 6502 19734 6554
rect 19786 6502 28888 6554
rect 1104 6480 28888 6502
rect 1762 6400 1768 6452
rect 1820 6440 1826 6452
rect 1949 6443 2007 6449
rect 1949 6440 1961 6443
rect 1820 6412 1961 6440
rect 1820 6400 1826 6412
rect 1949 6409 1961 6412
rect 1995 6409 2007 6443
rect 2590 6440 2596 6452
rect 2551 6412 2596 6440
rect 1949 6403 2007 6409
rect 2590 6400 2596 6412
rect 2648 6400 2654 6452
rect 4706 6400 4712 6452
rect 4764 6400 4770 6452
rect 27890 6440 27896 6452
rect 27851 6412 27896 6440
rect 27890 6400 27896 6412
rect 27948 6400 27954 6452
rect 3602 6372 3608 6384
rect 3563 6344 3608 6372
rect 3602 6332 3608 6344
rect 3660 6332 3666 6384
rect 4154 6332 4160 6384
rect 4212 6372 4218 6384
rect 4724 6372 4752 6400
rect 4212 6344 27844 6372
rect 4212 6332 4218 6344
rect 1949 6307 2007 6313
rect 1949 6273 1961 6307
rect 1995 6304 2007 6307
rect 2501 6307 2559 6313
rect 2501 6304 2513 6307
rect 1995 6276 2513 6304
rect 1995 6273 2007 6276
rect 1949 6267 2007 6273
rect 2501 6273 2513 6276
rect 2547 6304 2559 6307
rect 2590 6304 2596 6316
rect 2547 6276 2596 6304
rect 2547 6273 2559 6276
rect 2501 6267 2559 6273
rect 2590 6264 2596 6276
rect 2648 6264 2654 6316
rect 27816 6313 27844 6344
rect 27157 6307 27215 6313
rect 27157 6273 27169 6307
rect 27203 6304 27215 6307
rect 27801 6307 27859 6313
rect 27203 6276 27752 6304
rect 27203 6273 27215 6276
rect 27157 6267 27215 6273
rect 3421 6239 3479 6245
rect 3421 6205 3433 6239
rect 3467 6236 3479 6239
rect 4430 6236 4436 6248
rect 3467 6208 4436 6236
rect 3467 6205 3479 6208
rect 3421 6199 3479 6205
rect 4430 6196 4436 6208
rect 4488 6196 4494 6248
rect 4522 6196 4528 6248
rect 4580 6236 4586 6248
rect 24578 6236 24584 6248
rect 4580 6208 4625 6236
rect 24539 6208 24584 6236
rect 4580 6196 4586 6208
rect 24578 6196 24584 6208
rect 24636 6196 24642 6248
rect 24765 6239 24823 6245
rect 24765 6205 24777 6239
rect 24811 6236 24823 6239
rect 24946 6236 24952 6248
rect 24811 6208 24952 6236
rect 24811 6205 24823 6208
rect 24765 6199 24823 6205
rect 24946 6196 24952 6208
rect 25004 6196 25010 6248
rect 26050 6236 26056 6248
rect 26011 6208 26056 6236
rect 26050 6196 26056 6208
rect 26108 6196 26114 6248
rect 2682 6128 2688 6180
rect 2740 6168 2746 6180
rect 8662 6168 8668 6180
rect 2740 6140 8668 6168
rect 2740 6128 2746 6140
rect 8662 6128 8668 6140
rect 8720 6128 8726 6180
rect 27724 6168 27752 6276
rect 27801 6273 27813 6307
rect 27847 6273 27859 6307
rect 27801 6267 27859 6273
rect 27798 6168 27804 6180
rect 27724 6140 27804 6168
rect 27798 6128 27804 6140
rect 27856 6128 27862 6180
rect 26510 6060 26516 6112
rect 26568 6100 26574 6112
rect 27249 6103 27307 6109
rect 27249 6100 27261 6103
rect 26568 6072 27261 6100
rect 26568 6060 26574 6072
rect 27249 6069 27261 6072
rect 27295 6069 27307 6103
rect 27249 6063 27307 6069
rect 1104 6010 28888 6032
rect 1104 5958 5582 6010
rect 5634 5958 5646 6010
rect 5698 5958 5710 6010
rect 5762 5958 5774 6010
rect 5826 5958 5838 6010
rect 5890 5958 14846 6010
rect 14898 5958 14910 6010
rect 14962 5958 14974 6010
rect 15026 5958 15038 6010
rect 15090 5958 15102 6010
rect 15154 5958 24110 6010
rect 24162 5958 24174 6010
rect 24226 5958 24238 6010
rect 24290 5958 24302 6010
rect 24354 5958 24366 6010
rect 24418 5958 28888 6010
rect 1104 5936 28888 5958
rect 24578 5856 24584 5908
rect 24636 5896 24642 5908
rect 25225 5899 25283 5905
rect 25225 5896 25237 5899
rect 24636 5868 25237 5896
rect 24636 5856 24642 5868
rect 25225 5865 25237 5868
rect 25271 5865 25283 5899
rect 25225 5859 25283 5865
rect 5905 5831 5963 5837
rect 5905 5828 5917 5831
rect 1412 5800 5917 5828
rect 1412 5769 1440 5800
rect 5905 5797 5917 5800
rect 5951 5797 5963 5831
rect 27614 5828 27620 5840
rect 5905 5791 5963 5797
rect 26344 5800 27620 5828
rect 1397 5763 1455 5769
rect 1397 5729 1409 5763
rect 1443 5729 1455 5763
rect 1854 5760 1860 5772
rect 1815 5732 1860 5760
rect 1397 5723 1455 5729
rect 1854 5720 1860 5732
rect 1912 5720 1918 5772
rect 5350 5720 5356 5772
rect 5408 5760 5414 5772
rect 26344 5769 26372 5800
rect 27614 5788 27620 5800
rect 27672 5788 27678 5840
rect 7193 5763 7251 5769
rect 7193 5760 7205 5763
rect 5408 5732 7205 5760
rect 5408 5720 5414 5732
rect 7193 5729 7205 5732
rect 7239 5729 7251 5763
rect 7193 5723 7251 5729
rect 26329 5763 26387 5769
rect 26329 5729 26341 5763
rect 26375 5729 26387 5763
rect 26510 5760 26516 5772
rect 26471 5732 26516 5760
rect 26329 5723 26387 5729
rect 26510 5720 26516 5732
rect 26568 5720 26574 5772
rect 28166 5760 28172 5772
rect 28127 5732 28172 5760
rect 28166 5720 28172 5732
rect 28224 5720 28230 5772
rect 3789 5695 3847 5701
rect 3789 5661 3801 5695
rect 3835 5692 3847 5695
rect 4154 5692 4160 5704
rect 3835 5664 4160 5692
rect 3835 5661 3847 5664
rect 3789 5655 3847 5661
rect 4154 5652 4160 5664
rect 4212 5652 4218 5704
rect 4614 5692 4620 5704
rect 4575 5664 4620 5692
rect 4614 5652 4620 5664
rect 4672 5652 4678 5704
rect 5261 5695 5319 5701
rect 5261 5661 5273 5695
rect 5307 5692 5319 5695
rect 6362 5692 6368 5704
rect 5307 5664 6368 5692
rect 5307 5661 5319 5664
rect 5261 5655 5319 5661
rect 6362 5652 6368 5664
rect 6420 5652 6426 5704
rect 6546 5692 6552 5704
rect 6507 5664 6552 5692
rect 6546 5652 6552 5664
rect 6604 5652 6610 5704
rect 24854 5652 24860 5704
rect 24912 5692 24918 5704
rect 25869 5695 25927 5701
rect 25869 5692 25881 5695
rect 24912 5664 25881 5692
rect 24912 5652 24918 5664
rect 25869 5661 25881 5664
rect 25915 5661 25927 5695
rect 25869 5655 25927 5661
rect 1578 5624 1584 5636
rect 1539 5596 1584 5624
rect 1578 5584 1584 5596
rect 1636 5584 1642 5636
rect 3878 5556 3884 5568
rect 3839 5528 3884 5556
rect 3878 5516 3884 5528
rect 3936 5516 3942 5568
rect 1104 5466 28888 5488
rect 1104 5414 10214 5466
rect 10266 5414 10278 5466
rect 10330 5414 10342 5466
rect 10394 5414 10406 5466
rect 10458 5414 10470 5466
rect 10522 5414 19478 5466
rect 19530 5414 19542 5466
rect 19594 5414 19606 5466
rect 19658 5414 19670 5466
rect 19722 5414 19734 5466
rect 19786 5414 28888 5466
rect 1104 5392 28888 5414
rect 1489 5355 1547 5361
rect 1489 5321 1501 5355
rect 1535 5352 1547 5355
rect 1578 5352 1584 5364
rect 1535 5324 1584 5352
rect 1535 5321 1547 5324
rect 1489 5315 1547 5321
rect 1578 5312 1584 5324
rect 1636 5312 1642 5364
rect 6546 5352 6552 5364
rect 2056 5324 6552 5352
rect 1397 5219 1455 5225
rect 1397 5185 1409 5219
rect 1443 5216 1455 5219
rect 1670 5216 1676 5228
rect 1443 5188 1676 5216
rect 1443 5185 1455 5188
rect 1397 5179 1455 5185
rect 1670 5176 1676 5188
rect 1728 5176 1734 5228
rect 2056 5225 2084 5324
rect 6546 5312 6552 5324
rect 6604 5312 6610 5364
rect 24946 5312 24952 5364
rect 25004 5352 25010 5364
rect 27893 5355 27951 5361
rect 27893 5352 27905 5355
rect 25004 5324 27905 5352
rect 25004 5312 25010 5324
rect 27893 5321 27905 5324
rect 27939 5321 27951 5355
rect 27893 5315 27951 5321
rect 2225 5287 2283 5293
rect 2225 5253 2237 5287
rect 2271 5284 2283 5287
rect 3878 5284 3884 5296
rect 2271 5256 3884 5284
rect 2271 5253 2283 5256
rect 2225 5247 2283 5253
rect 3878 5244 3884 5256
rect 3936 5244 3942 5296
rect 24765 5287 24823 5293
rect 24765 5253 24777 5287
rect 24811 5284 24823 5287
rect 27249 5287 27307 5293
rect 27249 5284 27261 5287
rect 24811 5256 27261 5284
rect 24811 5253 24823 5256
rect 24765 5247 24823 5253
rect 27249 5253 27261 5256
rect 27295 5253 27307 5287
rect 27249 5247 27307 5253
rect 2041 5219 2099 5225
rect 2041 5185 2053 5219
rect 2087 5185 2099 5219
rect 27154 5216 27160 5228
rect 27115 5188 27160 5216
rect 2041 5179 2099 5185
rect 27154 5176 27160 5188
rect 27212 5176 27218 5228
rect 27801 5219 27859 5225
rect 27801 5185 27813 5219
rect 27847 5216 27859 5219
rect 27982 5216 27988 5228
rect 27847 5188 27988 5216
rect 27847 5185 27859 5188
rect 27801 5179 27859 5185
rect 27982 5176 27988 5188
rect 28040 5176 28046 5228
rect 2774 5108 2780 5160
rect 2832 5148 2838 5160
rect 24581 5151 24639 5157
rect 2832 5120 2877 5148
rect 2832 5108 2838 5120
rect 24581 5117 24593 5151
rect 24627 5148 24639 5151
rect 24854 5148 24860 5160
rect 24627 5120 24860 5148
rect 24627 5117 24639 5120
rect 24581 5111 24639 5117
rect 24854 5108 24860 5120
rect 24912 5108 24918 5160
rect 26142 5148 26148 5160
rect 26103 5120 26148 5148
rect 26142 5108 26148 5120
rect 26200 5108 26206 5160
rect 2314 5040 2320 5092
rect 2372 5080 2378 5092
rect 4430 5080 4436 5092
rect 2372 5052 4436 5080
rect 2372 5040 2378 5052
rect 4430 5040 4436 5052
rect 4488 5040 4494 5092
rect 5074 5040 5080 5092
rect 5132 5080 5138 5092
rect 6549 5083 6607 5089
rect 6549 5080 6561 5083
rect 5132 5052 6561 5080
rect 5132 5040 5138 5052
rect 6549 5049 6561 5052
rect 6595 5049 6607 5083
rect 6549 5043 6607 5049
rect 17126 5040 17132 5092
rect 17184 5080 17190 5092
rect 17586 5080 17592 5092
rect 17184 5052 17592 5080
rect 17184 5040 17190 5052
rect 17586 5040 17592 5052
rect 17644 5080 17650 5092
rect 27706 5080 27712 5092
rect 17644 5052 27712 5080
rect 17644 5040 17650 5052
rect 27706 5040 27712 5052
rect 27764 5040 27770 5092
rect 4246 4972 4252 5024
rect 4304 5012 4310 5024
rect 4525 5015 4583 5021
rect 4525 5012 4537 5015
rect 4304 4984 4537 5012
rect 4304 4972 4310 4984
rect 4525 4981 4537 4984
rect 4571 4981 4583 5015
rect 5166 5012 5172 5024
rect 5127 4984 5172 5012
rect 4525 4975 4583 4981
rect 5166 4972 5172 4984
rect 5224 4972 5230 5024
rect 5813 5015 5871 5021
rect 5813 4981 5825 5015
rect 5859 5012 5871 5015
rect 5902 5012 5908 5024
rect 5859 4984 5908 5012
rect 5859 4981 5871 4984
rect 5813 4975 5871 4981
rect 5902 4972 5908 4984
rect 5960 4972 5966 5024
rect 7190 5012 7196 5024
rect 7151 4984 7196 5012
rect 7190 4972 7196 4984
rect 7248 4972 7254 5024
rect 1104 4922 28888 4944
rect 1104 4870 5582 4922
rect 5634 4870 5646 4922
rect 5698 4870 5710 4922
rect 5762 4870 5774 4922
rect 5826 4870 5838 4922
rect 5890 4870 14846 4922
rect 14898 4870 14910 4922
rect 14962 4870 14974 4922
rect 15026 4870 15038 4922
rect 15090 4870 15102 4922
rect 15154 4870 24110 4922
rect 24162 4870 24174 4922
rect 24226 4870 24238 4922
rect 24290 4870 24302 4922
rect 24354 4870 24366 4922
rect 24418 4870 28888 4922
rect 1104 4848 28888 4870
rect 3789 4675 3847 4681
rect 3789 4641 3801 4675
rect 3835 4672 3847 4675
rect 7190 4672 7196 4684
rect 3835 4644 7196 4672
rect 3835 4641 3847 4644
rect 3789 4635 3847 4641
rect 7190 4632 7196 4644
rect 7248 4632 7254 4684
rect 17126 4672 17132 4684
rect 7392 4644 17132 4672
rect 1765 4607 1823 4613
rect 1765 4573 1777 4607
rect 1811 4604 1823 4607
rect 2406 4604 2412 4616
rect 1811 4576 2412 4604
rect 1811 4573 1823 4576
rect 1765 4567 1823 4573
rect 2406 4564 2412 4576
rect 2464 4564 2470 4616
rect 3050 4604 3056 4616
rect 3011 4576 3056 4604
rect 3050 4564 3056 4576
rect 3108 4564 3114 4616
rect 6270 4604 6276 4616
rect 6231 4576 6276 4604
rect 6270 4564 6276 4576
rect 6328 4564 6334 4616
rect 7282 4604 7288 4616
rect 7195 4576 7288 4604
rect 7282 4564 7288 4576
rect 7340 4604 7346 4616
rect 7392 4604 7420 4644
rect 17126 4632 17132 4644
rect 17184 4632 17190 4684
rect 8110 4604 8116 4616
rect 7340 4576 7420 4604
rect 8071 4576 8116 4604
rect 7340 4564 7346 4576
rect 8110 4564 8116 4576
rect 8168 4564 8174 4616
rect 9030 4564 9036 4616
rect 9088 4604 9094 4616
rect 9217 4607 9275 4613
rect 9217 4604 9229 4607
rect 9088 4576 9229 4604
rect 9088 4564 9094 4576
rect 9217 4573 9229 4576
rect 9263 4573 9275 4607
rect 23842 4604 23848 4616
rect 23803 4576 23848 4604
rect 9217 4567 9275 4573
rect 23842 4564 23848 4576
rect 23900 4564 23906 4616
rect 25869 4607 25927 4613
rect 25869 4573 25881 4607
rect 25915 4604 25927 4607
rect 26329 4607 26387 4613
rect 26329 4604 26341 4607
rect 25915 4576 26341 4604
rect 25915 4573 25927 4576
rect 25869 4567 25927 4573
rect 26329 4573 26341 4576
rect 26375 4573 26387 4607
rect 26329 4567 26387 4573
rect 3145 4539 3203 4545
rect 3145 4505 3157 4539
rect 3191 4536 3203 4539
rect 3973 4539 4031 4545
rect 3973 4536 3985 4539
rect 3191 4508 3985 4536
rect 3191 4505 3203 4508
rect 3145 4499 3203 4505
rect 3973 4505 3985 4508
rect 4019 4505 4031 4539
rect 3973 4499 4031 4505
rect 4338 4496 4344 4548
rect 4396 4536 4402 4548
rect 5629 4539 5687 4545
rect 5629 4536 5641 4539
rect 4396 4508 5641 4536
rect 4396 4496 4402 4508
rect 5629 4505 5641 4508
rect 5675 4505 5687 4539
rect 24854 4536 24860 4548
rect 24815 4508 24860 4536
rect 5629 4499 5687 4505
rect 24854 4496 24860 4508
rect 24912 4496 24918 4548
rect 26513 4539 26571 4545
rect 26513 4505 26525 4539
rect 26559 4536 26571 4539
rect 27706 4536 27712 4548
rect 26559 4508 27712 4536
rect 26559 4505 26571 4508
rect 26513 4499 26571 4505
rect 27706 4496 27712 4508
rect 27764 4496 27770 4548
rect 28169 4539 28227 4545
rect 28169 4505 28181 4539
rect 28215 4536 28227 4539
rect 28350 4536 28356 4548
rect 28215 4508 28356 4536
rect 28215 4505 28227 4508
rect 28169 4499 28227 4505
rect 28350 4496 28356 4508
rect 28408 4496 28414 4548
rect 1578 4428 1584 4480
rect 1636 4468 1642 4480
rect 1857 4471 1915 4477
rect 1857 4468 1869 4471
rect 1636 4440 1869 4468
rect 1636 4428 1642 4440
rect 1857 4437 1869 4440
rect 1903 4437 1915 4471
rect 2498 4468 2504 4480
rect 2459 4440 2504 4468
rect 1857 4431 1915 4437
rect 2498 4428 2504 4440
rect 2556 4428 2562 4480
rect 7374 4468 7380 4480
rect 7335 4440 7380 4468
rect 7374 4428 7380 4440
rect 7432 4428 7438 4480
rect 24946 4468 24952 4480
rect 24907 4440 24952 4468
rect 24946 4428 24952 4440
rect 25004 4428 25010 4480
rect 1104 4378 28888 4400
rect 1104 4326 10214 4378
rect 10266 4326 10278 4378
rect 10330 4326 10342 4378
rect 10394 4326 10406 4378
rect 10458 4326 10470 4378
rect 10522 4326 19478 4378
rect 19530 4326 19542 4378
rect 19594 4326 19606 4378
rect 19658 4326 19670 4378
rect 19722 4326 19734 4378
rect 19786 4326 28888 4378
rect 1104 4304 28888 4326
rect 2406 4224 2412 4276
rect 2464 4264 2470 4276
rect 2464 4236 27568 4264
rect 2464 4224 2470 4236
rect 1578 4196 1584 4208
rect 1539 4168 1584 4196
rect 1578 4156 1584 4168
rect 1636 4156 1642 4208
rect 5074 4196 5080 4208
rect 3712 4168 5080 4196
rect 1394 4128 1400 4140
rect 1355 4100 1400 4128
rect 1394 4088 1400 4100
rect 1452 4088 1458 4140
rect 3712 4137 3740 4168
rect 5074 4156 5080 4168
rect 5132 4156 5138 4208
rect 7374 4196 7380 4208
rect 7335 4168 7380 4196
rect 7374 4156 7380 4168
rect 7432 4156 7438 4208
rect 3697 4131 3755 4137
rect 3697 4097 3709 4131
rect 3743 4097 3755 4131
rect 3697 4091 3755 4097
rect 9493 4131 9551 4137
rect 9493 4097 9505 4131
rect 9539 4128 9551 4131
rect 12894 4128 12900 4140
rect 9539 4100 12900 4128
rect 9539 4097 9551 4100
rect 9493 4091 9551 4097
rect 12894 4088 12900 4100
rect 12952 4088 12958 4140
rect 24854 4088 24860 4140
rect 24912 4128 24918 4140
rect 27154 4128 27160 4140
rect 24912 4100 27160 4128
rect 24912 4088 24918 4100
rect 27154 4088 27160 4100
rect 27212 4088 27218 4140
rect 27540 4137 27568 4236
rect 27525 4131 27583 4137
rect 27525 4097 27537 4131
rect 27571 4128 27583 4131
rect 28258 4128 28264 4140
rect 27571 4100 28264 4128
rect 27571 4097 27583 4100
rect 27525 4091 27583 4097
rect 28258 4088 28264 4100
rect 28316 4088 28322 4140
rect 658 4020 664 4072
rect 716 4060 722 4072
rect 1857 4063 1915 4069
rect 1857 4060 1869 4063
rect 716 4044 1348 4060
rect 1504 4044 1869 4060
rect 716 4032 1869 4044
rect 716 4020 722 4032
rect 1320 4016 1532 4032
rect 1857 4029 1869 4032
rect 1903 4029 1915 4063
rect 1857 4023 1915 4029
rect 3881 4063 3939 4069
rect 3881 4029 3893 4063
rect 3927 4029 3939 4063
rect 4154 4060 4160 4072
rect 4115 4032 4160 4060
rect 3881 4023 3939 4029
rect 3896 3992 3924 4023
rect 4154 4020 4160 4032
rect 4212 4020 4218 4072
rect 7193 4063 7251 4069
rect 7193 4029 7205 4063
rect 7239 4060 7251 4063
rect 8110 4060 8116 4072
rect 7239 4032 8116 4060
rect 7239 4029 7251 4032
rect 7193 4023 7251 4029
rect 8110 4020 8116 4032
rect 8168 4020 8174 4072
rect 8205 4063 8263 4069
rect 8205 4029 8217 4063
rect 8251 4029 8263 4063
rect 8205 4023 8263 4029
rect 3896 3964 7696 3992
rect 1394 3884 1400 3936
rect 1452 3924 1458 3936
rect 5166 3924 5172 3936
rect 1452 3896 5172 3924
rect 1452 3884 1458 3896
rect 5166 3884 5172 3896
rect 5224 3884 5230 3936
rect 6733 3927 6791 3933
rect 6733 3893 6745 3927
rect 6779 3924 6791 3927
rect 6914 3924 6920 3936
rect 6779 3896 6920 3924
rect 6779 3893 6791 3896
rect 6733 3887 6791 3893
rect 6914 3884 6920 3896
rect 6972 3884 6978 3936
rect 7668 3924 7696 3964
rect 7742 3952 7748 4004
rect 7800 3992 7806 4004
rect 8220 3992 8248 4023
rect 12526 4020 12532 4072
rect 12584 4060 12590 4072
rect 12989 4063 13047 4069
rect 12989 4060 13001 4063
rect 12584 4032 13001 4060
rect 12584 4020 12590 4032
rect 12989 4029 13001 4032
rect 13035 4029 13047 4063
rect 13170 4060 13176 4072
rect 13131 4032 13176 4060
rect 12989 4023 13047 4029
rect 13170 4020 13176 4032
rect 13228 4020 13234 4072
rect 13538 4060 13544 4072
rect 13499 4032 13544 4060
rect 13538 4020 13544 4032
rect 13596 4020 13602 4072
rect 17497 4063 17555 4069
rect 17497 4029 17509 4063
rect 17543 4029 17555 4063
rect 17678 4060 17684 4072
rect 17639 4032 17684 4060
rect 17497 4023 17555 4029
rect 17402 3992 17408 4004
rect 7800 3964 8248 3992
rect 8312 3964 17408 3992
rect 7800 3952 7806 3964
rect 8312 3924 8340 3964
rect 17402 3952 17408 3964
rect 17460 3952 17466 4004
rect 17512 3992 17540 4023
rect 17678 4020 17684 4032
rect 17736 4020 17742 4072
rect 18046 4060 18052 4072
rect 18007 4032 18052 4060
rect 18046 4020 18052 4032
rect 18104 4020 18110 4072
rect 23474 4060 23480 4072
rect 23435 4032 23480 4060
rect 23474 4020 23480 4032
rect 23532 4020 23538 4072
rect 23661 4063 23719 4069
rect 23661 4029 23673 4063
rect 23707 4029 23719 4063
rect 23661 4023 23719 4029
rect 25317 4063 25375 4069
rect 25317 4029 25329 4063
rect 25363 4060 25375 4063
rect 25363 4032 26234 4060
rect 25363 4029 25375 4032
rect 25317 4023 25375 4029
rect 17954 3992 17960 4004
rect 17512 3964 17960 3992
rect 17954 3952 17960 3964
rect 18012 3952 18018 4004
rect 23106 3952 23112 4004
rect 23164 3992 23170 4004
rect 23676 3992 23704 4023
rect 23164 3964 23704 3992
rect 26206 3992 26234 4032
rect 28994 3992 29000 4004
rect 26206 3964 29000 3992
rect 23164 3952 23170 3964
rect 28994 3952 29000 3964
rect 29052 3952 29058 4004
rect 7668 3896 8340 3924
rect 9306 3884 9312 3936
rect 9364 3924 9370 3936
rect 9585 3927 9643 3933
rect 9585 3924 9597 3927
rect 9364 3896 9597 3924
rect 9364 3884 9370 3896
rect 9585 3893 9597 3896
rect 9631 3893 9643 3927
rect 10318 3924 10324 3936
rect 10279 3896 10324 3924
rect 9585 3887 9643 3893
rect 10318 3884 10324 3896
rect 10376 3884 10382 3936
rect 15654 3884 15660 3936
rect 15712 3924 15718 3936
rect 15841 3927 15899 3933
rect 15841 3924 15853 3927
rect 15712 3896 15853 3924
rect 15712 3884 15718 3896
rect 15841 3893 15853 3896
rect 15887 3893 15899 3927
rect 15841 3887 15899 3893
rect 22186 3884 22192 3936
rect 22244 3924 22250 3936
rect 23017 3927 23075 3933
rect 23017 3924 23029 3927
rect 22244 3896 23029 3924
rect 22244 3884 22250 3896
rect 23017 3893 23029 3896
rect 23063 3893 23075 3927
rect 23017 3887 23075 3893
rect 25130 3884 25136 3936
rect 25188 3924 25194 3936
rect 25961 3927 26019 3933
rect 25961 3924 25973 3927
rect 25188 3896 25973 3924
rect 25188 3884 25194 3896
rect 25961 3893 25973 3896
rect 26007 3893 26019 3927
rect 25961 3887 26019 3893
rect 1104 3834 28888 3856
rect 1104 3782 5582 3834
rect 5634 3782 5646 3834
rect 5698 3782 5710 3834
rect 5762 3782 5774 3834
rect 5826 3782 5838 3834
rect 5890 3782 14846 3834
rect 14898 3782 14910 3834
rect 14962 3782 14974 3834
rect 15026 3782 15038 3834
rect 15090 3782 15102 3834
rect 15154 3782 24110 3834
rect 24162 3782 24174 3834
rect 24226 3782 24238 3834
rect 24290 3782 24302 3834
rect 24354 3782 24366 3834
rect 24418 3782 28888 3834
rect 1104 3760 28888 3782
rect 5902 3720 5908 3732
rect 2746 3692 5908 3720
rect 2746 3652 2774 3692
rect 5902 3680 5908 3692
rect 5960 3680 5966 3732
rect 12342 3720 12348 3732
rect 6012 3692 12348 3720
rect 1412 3624 2774 3652
rect 1412 3593 1440 3624
rect 3326 3612 3332 3664
rect 3384 3652 3390 3664
rect 4338 3652 4344 3664
rect 3384 3624 4344 3652
rect 3384 3612 3390 3624
rect 4338 3612 4344 3624
rect 4396 3612 4402 3664
rect 6012 3652 6040 3692
rect 12342 3680 12348 3692
rect 12400 3680 12406 3732
rect 12526 3720 12532 3732
rect 12487 3692 12532 3720
rect 12526 3680 12532 3692
rect 12584 3680 12590 3732
rect 13081 3723 13139 3729
rect 13081 3689 13093 3723
rect 13127 3720 13139 3723
rect 13170 3720 13176 3732
rect 13127 3692 13176 3720
rect 13127 3689 13139 3692
rect 13081 3683 13139 3689
rect 13170 3680 13176 3692
rect 13228 3680 13234 3732
rect 17402 3680 17408 3732
rect 17460 3720 17466 3732
rect 19245 3723 19303 3729
rect 19245 3720 19257 3723
rect 17460 3692 19257 3720
rect 17460 3680 17466 3692
rect 19245 3689 19257 3692
rect 19291 3689 19303 3723
rect 23106 3720 23112 3732
rect 23067 3692 23112 3720
rect 19245 3683 19303 3689
rect 23106 3680 23112 3692
rect 23164 3680 23170 3732
rect 23474 3680 23480 3732
rect 23532 3720 23538 3732
rect 23845 3723 23903 3729
rect 23845 3720 23857 3723
rect 23532 3692 23857 3720
rect 23532 3680 23538 3692
rect 23845 3689 23857 3692
rect 23891 3689 23903 3723
rect 23845 3683 23903 3689
rect 10318 3652 10324 3664
rect 4632 3624 6040 3652
rect 9140 3624 10324 3652
rect 1397 3587 1455 3593
rect 1397 3553 1409 3587
rect 1443 3553 1455 3587
rect 1397 3547 1455 3553
rect 1581 3587 1639 3593
rect 1581 3553 1593 3587
rect 1627 3584 1639 3587
rect 3881 3587 3939 3593
rect 3881 3584 3893 3587
rect 1627 3556 3893 3584
rect 1627 3553 1639 3556
rect 1581 3547 1639 3553
rect 3881 3553 3893 3556
rect 3927 3553 3939 3587
rect 3881 3547 3939 3553
rect 3050 3476 3056 3528
rect 3108 3516 3114 3528
rect 3789 3519 3847 3525
rect 3789 3516 3801 3519
rect 3108 3488 3801 3516
rect 3108 3476 3114 3488
rect 3789 3485 3801 3488
rect 3835 3516 3847 3519
rect 4632 3516 4660 3624
rect 5350 3584 5356 3596
rect 5311 3556 5356 3584
rect 5350 3544 5356 3556
rect 5408 3544 5414 3596
rect 5902 3584 5908 3596
rect 5863 3556 5908 3584
rect 5902 3544 5908 3556
rect 5960 3544 5966 3596
rect 9140 3593 9168 3624
rect 10318 3612 10324 3624
rect 10376 3612 10382 3664
rect 12894 3612 12900 3664
rect 12952 3652 12958 3664
rect 16666 3652 16672 3664
rect 12952 3624 16672 3652
rect 12952 3612 12958 3624
rect 16666 3612 16672 3624
rect 16724 3612 16730 3664
rect 19978 3612 19984 3664
rect 20036 3652 20042 3664
rect 24854 3652 24860 3664
rect 20036 3624 24860 3652
rect 20036 3612 20042 3624
rect 24854 3612 24860 3624
rect 24912 3612 24918 3664
rect 9125 3587 9183 3593
rect 9125 3553 9137 3587
rect 9171 3553 9183 3587
rect 9306 3584 9312 3596
rect 9267 3556 9312 3584
rect 9125 3547 9183 3553
rect 9306 3544 9312 3556
rect 9364 3544 9370 3596
rect 9674 3584 9680 3596
rect 9635 3556 9680 3584
rect 9674 3544 9680 3556
rect 9732 3544 9738 3596
rect 15654 3584 15660 3596
rect 15615 3556 15660 3584
rect 15654 3544 15660 3556
rect 15712 3544 15718 3596
rect 16114 3584 16120 3596
rect 16075 3556 16120 3584
rect 16114 3544 16120 3556
rect 16172 3544 16178 3596
rect 20714 3584 20720 3596
rect 19444 3556 20720 3584
rect 3835 3488 4660 3516
rect 4709 3519 4767 3525
rect 3835 3485 3847 3488
rect 3789 3479 3847 3485
rect 4709 3485 4721 3519
rect 4755 3485 4767 3519
rect 7650 3516 7656 3528
rect 7611 3488 7656 3516
rect 4709 3479 4767 3485
rect 3234 3448 3240 3460
rect 3195 3420 3240 3448
rect 3234 3408 3240 3420
rect 3292 3408 3298 3460
rect 3878 3408 3884 3460
rect 3936 3448 3942 3460
rect 4522 3448 4528 3460
rect 3936 3420 4528 3448
rect 3936 3408 3942 3420
rect 4522 3408 4528 3420
rect 4580 3408 4586 3460
rect 2222 3340 2228 3392
rect 2280 3380 2286 3392
rect 4724 3380 4752 3479
rect 7650 3476 7656 3488
rect 7708 3476 7714 3528
rect 11698 3476 11704 3528
rect 11756 3516 11762 3528
rect 11885 3519 11943 3525
rect 11885 3516 11897 3519
rect 11756 3488 11897 3516
rect 11756 3476 11762 3488
rect 11885 3485 11897 3488
rect 11931 3485 11943 3519
rect 12986 3516 12992 3528
rect 12947 3488 12992 3516
rect 11885 3479 11943 3485
rect 12986 3476 12992 3488
rect 13044 3476 13050 3528
rect 14182 3476 14188 3528
rect 14240 3516 14246 3528
rect 14461 3519 14519 3525
rect 14461 3516 14473 3519
rect 14240 3488 14473 3516
rect 14240 3476 14246 3488
rect 14461 3485 14473 3488
rect 14507 3485 14519 3519
rect 14461 3479 14519 3485
rect 18693 3519 18751 3525
rect 18693 3485 18705 3519
rect 18739 3516 18751 3519
rect 18874 3516 18880 3528
rect 18739 3488 18880 3516
rect 18739 3485 18751 3488
rect 18693 3479 18751 3485
rect 18874 3476 18880 3488
rect 18932 3476 18938 3528
rect 19444 3525 19472 3556
rect 20714 3544 20720 3556
rect 20772 3584 20778 3596
rect 25130 3584 25136 3596
rect 20772 3556 22140 3584
rect 25091 3556 25136 3584
rect 20772 3544 20778 3556
rect 19429 3519 19487 3525
rect 19429 3485 19441 3519
rect 19475 3485 19487 3519
rect 19978 3516 19984 3528
rect 19939 3488 19984 3516
rect 19429 3479 19487 3485
rect 5534 3448 5540 3460
rect 5495 3420 5540 3448
rect 5534 3408 5540 3420
rect 5592 3408 5598 3460
rect 7668 3448 7696 3476
rect 15654 3448 15660 3460
rect 7668 3420 15660 3448
rect 15654 3408 15660 3420
rect 15712 3408 15718 3460
rect 15838 3448 15844 3460
rect 15799 3420 15844 3448
rect 15838 3408 15844 3420
rect 15896 3408 15902 3460
rect 18230 3408 18236 3460
rect 18288 3448 18294 3460
rect 19444 3448 19472 3479
rect 19978 3476 19984 3488
rect 20036 3476 20042 3528
rect 20162 3476 20168 3528
rect 20220 3516 20226 3528
rect 20809 3519 20867 3525
rect 20809 3516 20821 3519
rect 20220 3488 20821 3516
rect 20220 3476 20226 3488
rect 20809 3485 20821 3488
rect 20855 3485 20867 3519
rect 20809 3479 20867 3485
rect 21637 3519 21695 3525
rect 21637 3485 21649 3519
rect 21683 3516 21695 3519
rect 21910 3516 21916 3528
rect 21683 3488 21916 3516
rect 21683 3485 21695 3488
rect 21637 3479 21695 3485
rect 21910 3476 21916 3488
rect 21968 3476 21974 3528
rect 22112 3525 22140 3556
rect 25130 3544 25136 3556
rect 25188 3544 25194 3596
rect 26142 3584 26148 3596
rect 26103 3556 26148 3584
rect 26142 3544 26148 3556
rect 26200 3544 26206 3596
rect 22097 3519 22155 3525
rect 22097 3485 22109 3519
rect 22143 3485 22155 3519
rect 23014 3516 23020 3528
rect 22975 3488 23020 3516
rect 22097 3479 22155 3485
rect 23014 3476 23020 3488
rect 23072 3476 23078 3528
rect 24489 3519 24547 3525
rect 24489 3485 24501 3519
rect 24535 3516 24547 3519
rect 24946 3516 24952 3528
rect 24535 3488 24952 3516
rect 24535 3485 24547 3488
rect 24489 3479 24547 3485
rect 24504 3448 24532 3479
rect 24946 3476 24952 3488
rect 25004 3476 25010 3528
rect 27801 3519 27859 3525
rect 27801 3485 27813 3519
rect 27847 3516 27859 3519
rect 27982 3516 27988 3528
rect 27847 3488 27988 3516
rect 27847 3485 27859 3488
rect 27801 3479 27859 3485
rect 27982 3476 27988 3488
rect 28040 3476 28046 3528
rect 18288 3420 19472 3448
rect 19904 3420 24532 3448
rect 24581 3451 24639 3457
rect 18288 3408 18294 3420
rect 2280 3352 4752 3380
rect 4801 3383 4859 3389
rect 2280 3340 2286 3352
rect 4801 3349 4813 3383
rect 4847 3380 4859 3383
rect 6546 3380 6552 3392
rect 4847 3352 6552 3380
rect 4847 3349 4859 3352
rect 4801 3343 4859 3349
rect 6546 3340 6552 3352
rect 6604 3340 6610 3392
rect 7098 3340 7104 3392
rect 7156 3380 7162 3392
rect 7745 3383 7803 3389
rect 7745 3380 7757 3383
rect 7156 3352 7757 3380
rect 7156 3340 7162 3352
rect 7745 3349 7757 3352
rect 7791 3349 7803 3383
rect 7745 3343 7803 3349
rect 14090 3340 14096 3392
rect 14148 3380 14154 3392
rect 19904 3380 19932 3420
rect 24581 3417 24593 3451
rect 24627 3448 24639 3451
rect 25317 3451 25375 3457
rect 25317 3448 25329 3451
rect 24627 3420 25329 3448
rect 24627 3417 24639 3420
rect 24581 3411 24639 3417
rect 25317 3417 25329 3420
rect 25363 3417 25375 3451
rect 25317 3411 25375 3417
rect 20070 3380 20076 3392
rect 14148 3352 19932 3380
rect 20031 3352 20076 3380
rect 14148 3340 14154 3352
rect 20070 3340 20076 3352
rect 20128 3340 20134 3392
rect 22094 3340 22100 3392
rect 22152 3380 22158 3392
rect 22189 3383 22247 3389
rect 22189 3380 22201 3383
rect 22152 3352 22201 3380
rect 22152 3340 22158 3352
rect 22189 3349 22201 3352
rect 22235 3349 22247 3383
rect 22189 3343 22247 3349
rect 23750 3340 23756 3392
rect 23808 3380 23814 3392
rect 27893 3383 27951 3389
rect 27893 3380 27905 3383
rect 23808 3352 27905 3380
rect 23808 3340 23814 3352
rect 27893 3349 27905 3352
rect 27939 3349 27951 3383
rect 27893 3343 27951 3349
rect 1104 3290 28888 3312
rect 1104 3238 10214 3290
rect 10266 3238 10278 3290
rect 10330 3238 10342 3290
rect 10394 3238 10406 3290
rect 10458 3238 10470 3290
rect 10522 3238 19478 3290
rect 19530 3238 19542 3290
rect 19594 3238 19606 3290
rect 19658 3238 19670 3290
rect 19722 3238 19734 3290
rect 19786 3238 28888 3290
rect 1104 3216 28888 3238
rect 4246 3176 4252 3188
rect 2332 3148 4252 3176
rect 2332 3049 2360 3148
rect 4246 3136 4252 3148
rect 4304 3136 4310 3188
rect 5445 3179 5503 3185
rect 5445 3145 5457 3179
rect 5491 3176 5503 3179
rect 5534 3176 5540 3188
rect 5491 3148 5540 3176
rect 5491 3145 5503 3148
rect 5445 3139 5503 3145
rect 5534 3136 5540 3148
rect 5592 3136 5598 3188
rect 5626 3136 5632 3188
rect 5684 3176 5690 3188
rect 27706 3176 27712 3188
rect 5684 3148 27016 3176
rect 27667 3148 27712 3176
rect 5684 3136 5690 3148
rect 2498 3108 2504 3120
rect 2459 3080 2504 3108
rect 2498 3068 2504 3080
rect 2556 3068 2562 3120
rect 2590 3068 2596 3120
rect 2648 3108 2654 3120
rect 7098 3108 7104 3120
rect 2648 3080 5396 3108
rect 7059 3080 7104 3108
rect 2648 3068 2654 3080
rect 1673 3043 1731 3049
rect 1673 3009 1685 3043
rect 1719 3009 1731 3043
rect 1673 3003 1731 3009
rect 2317 3043 2375 3049
rect 2317 3009 2329 3043
rect 2363 3009 2375 3043
rect 2317 3003 2375 3009
rect 1688 2904 1716 3003
rect 4430 3000 4436 3052
rect 4488 3040 4494 3052
rect 5368 3049 5396 3080
rect 7098 3068 7104 3080
rect 7156 3068 7162 3120
rect 14090 3108 14096 3120
rect 8312 3080 14096 3108
rect 4617 3043 4675 3049
rect 4617 3040 4629 3043
rect 4488 3012 4629 3040
rect 4488 3000 4494 3012
rect 4617 3009 4629 3012
rect 4663 3009 4675 3043
rect 4617 3003 4675 3009
rect 5353 3043 5411 3049
rect 5353 3009 5365 3043
rect 5399 3040 5411 3043
rect 6914 3040 6920 3052
rect 5399 3012 5764 3040
rect 6875 3012 6920 3040
rect 5399 3009 5411 3012
rect 5353 3003 5411 3009
rect 2590 2932 2596 2984
rect 2648 2972 2654 2984
rect 2777 2975 2835 2981
rect 2777 2972 2789 2975
rect 2648 2944 2789 2972
rect 2648 2932 2654 2944
rect 2777 2941 2789 2944
rect 2823 2941 2835 2975
rect 4632 2972 4660 3003
rect 5626 2972 5632 2984
rect 4632 2944 5632 2972
rect 2777 2935 2835 2941
rect 5626 2932 5632 2944
rect 5684 2932 5690 2984
rect 3050 2904 3056 2916
rect 1688 2876 3056 2904
rect 3050 2864 3056 2876
rect 3108 2864 3114 2916
rect 5736 2904 5764 3012
rect 6914 3000 6920 3012
rect 6972 3000 6978 3052
rect 7374 2972 7380 2984
rect 7335 2944 7380 2972
rect 7374 2932 7380 2944
rect 7432 2932 7438 2984
rect 8312 2904 8340 3080
rect 14090 3068 14096 3080
rect 14148 3068 14154 3120
rect 17678 3108 17684 3120
rect 17639 3080 17684 3108
rect 17678 3068 17684 3080
rect 17736 3068 17742 3120
rect 22094 3108 22100 3120
rect 22055 3080 22100 3108
rect 22094 3068 22100 3080
rect 22152 3068 22158 3120
rect 24765 3111 24823 3117
rect 24765 3077 24777 3111
rect 24811 3108 24823 3111
rect 24811 3080 26648 3108
rect 24811 3077 24823 3080
rect 24765 3071 24823 3077
rect 9677 3043 9735 3049
rect 9677 3009 9689 3043
rect 9723 3040 9735 3043
rect 9766 3040 9772 3052
rect 9723 3012 9772 3040
rect 9723 3009 9735 3012
rect 9677 3003 9735 3009
rect 9766 3000 9772 3012
rect 9824 3000 9830 3052
rect 11698 3040 11704 3052
rect 11659 3012 11704 3040
rect 11698 3000 11704 3012
rect 11756 3000 11762 3052
rect 14182 3040 14188 3052
rect 14143 3012 14188 3040
rect 14182 3000 14188 3012
rect 14240 3000 14246 3052
rect 17589 3043 17647 3049
rect 17589 3040 17601 3043
rect 16546 3012 17601 3040
rect 11882 2972 11888 2984
rect 11843 2944 11888 2972
rect 11882 2932 11888 2944
rect 11940 2932 11946 2984
rect 12250 2972 12256 2984
rect 12211 2944 12256 2972
rect 12250 2932 12256 2944
rect 12308 2932 12314 2984
rect 14366 2972 14372 2984
rect 14327 2944 14372 2972
rect 14366 2932 14372 2944
rect 14424 2932 14430 2984
rect 14734 2972 14740 2984
rect 14695 2944 14740 2972
rect 14734 2932 14740 2944
rect 14792 2932 14798 2984
rect 5736 2876 8340 2904
rect 8662 2864 8668 2916
rect 8720 2904 8726 2916
rect 16546 2904 16574 3012
rect 17589 3009 17601 3012
rect 17635 3009 17647 3043
rect 18230 3040 18236 3052
rect 18191 3012 18236 3040
rect 17589 3003 17647 3009
rect 8720 2876 16574 2904
rect 8720 2864 8726 2876
rect 1578 2796 1584 2848
rect 1636 2836 1642 2848
rect 1765 2839 1823 2845
rect 1765 2836 1777 2839
rect 1636 2808 1777 2836
rect 1636 2796 1642 2808
rect 1765 2805 1777 2808
rect 1811 2805 1823 2839
rect 1765 2799 1823 2805
rect 4154 2796 4160 2848
rect 4212 2836 4218 2848
rect 4709 2839 4767 2845
rect 4709 2836 4721 2839
rect 4212 2808 4721 2836
rect 4212 2796 4218 2808
rect 4709 2805 4721 2808
rect 4755 2805 4767 2839
rect 9766 2836 9772 2848
rect 9727 2808 9772 2836
rect 4709 2799 4767 2805
rect 9766 2796 9772 2808
rect 9824 2796 9830 2848
rect 17604 2836 17632 3003
rect 18230 3000 18236 3012
rect 18288 3000 18294 3052
rect 18874 3040 18880 3052
rect 18835 3012 18880 3040
rect 18874 3000 18880 3012
rect 18932 3000 18938 3052
rect 21910 3040 21916 3052
rect 21871 3012 21916 3040
rect 21910 3000 21916 3012
rect 21968 3000 21974 3052
rect 26050 3000 26056 3052
rect 26108 3040 26114 3052
rect 26421 3043 26479 3049
rect 26421 3040 26433 3043
rect 26108 3012 26433 3040
rect 26108 3000 26114 3012
rect 26421 3009 26433 3012
rect 26467 3009 26479 3043
rect 26421 3003 26479 3009
rect 18325 2975 18383 2981
rect 18325 2941 18337 2975
rect 18371 2972 18383 2975
rect 19061 2975 19119 2981
rect 19061 2972 19073 2975
rect 18371 2944 19073 2972
rect 18371 2941 18383 2944
rect 18325 2935 18383 2941
rect 19061 2941 19073 2944
rect 19107 2941 19119 2975
rect 19334 2972 19340 2984
rect 19295 2944 19340 2972
rect 19061 2935 19119 2941
rect 19334 2932 19340 2944
rect 19392 2932 19398 2984
rect 22554 2972 22560 2984
rect 22515 2944 22560 2972
rect 22554 2932 22560 2944
rect 22612 2932 22618 2984
rect 24578 2972 24584 2984
rect 24539 2944 24584 2972
rect 24578 2932 24584 2944
rect 24636 2932 24642 2984
rect 24688 2944 25452 2972
rect 24688 2836 24716 2944
rect 24762 2864 24768 2916
rect 24820 2904 24826 2916
rect 25222 2904 25228 2916
rect 24820 2876 25228 2904
rect 24820 2864 24826 2876
rect 25222 2864 25228 2876
rect 25280 2864 25286 2916
rect 25424 2904 25452 2944
rect 25498 2932 25504 2984
rect 25556 2972 25562 2984
rect 26510 2972 26516 2984
rect 25556 2944 26516 2972
rect 25556 2932 25562 2944
rect 26510 2932 26516 2944
rect 26568 2932 26574 2984
rect 26620 2972 26648 3080
rect 26988 3049 27016 3148
rect 27706 3136 27712 3148
rect 27764 3136 27770 3188
rect 26973 3043 27031 3049
rect 26973 3009 26985 3043
rect 27019 3009 27031 3043
rect 26973 3003 27031 3009
rect 27617 3043 27675 3049
rect 27617 3009 27629 3043
rect 27663 3040 27675 3043
rect 27798 3040 27804 3052
rect 27663 3012 27804 3040
rect 27663 3009 27675 3012
rect 27617 3003 27675 3009
rect 27065 2975 27123 2981
rect 27065 2972 27077 2975
rect 26620 2944 27077 2972
rect 27065 2941 27077 2944
rect 27111 2941 27123 2975
rect 27065 2935 27123 2941
rect 27632 2904 27660 3003
rect 27798 3000 27804 3012
rect 27856 3000 27862 3052
rect 25424 2876 27660 2904
rect 17604 2808 24716 2836
rect 25038 2796 25044 2848
rect 25096 2836 25102 2848
rect 29638 2836 29644 2848
rect 25096 2808 29644 2836
rect 25096 2796 25102 2808
rect 29638 2796 29644 2808
rect 29696 2796 29702 2848
rect 1104 2746 28888 2768
rect 1104 2694 5582 2746
rect 5634 2694 5646 2746
rect 5698 2694 5710 2746
rect 5762 2694 5774 2746
rect 5826 2694 5838 2746
rect 5890 2694 14846 2746
rect 14898 2694 14910 2746
rect 14962 2694 14974 2746
rect 15026 2694 15038 2746
rect 15090 2694 15102 2746
rect 15154 2694 24110 2746
rect 24162 2694 24174 2746
rect 24226 2694 24238 2746
rect 24290 2694 24302 2746
rect 24354 2694 24366 2746
rect 24418 2694 28888 2746
rect 1104 2672 28888 2694
rect 6270 2632 6276 2644
rect 1412 2604 6276 2632
rect 1412 2505 1440 2604
rect 6270 2592 6276 2604
rect 6328 2592 6334 2644
rect 11882 2592 11888 2644
rect 11940 2632 11946 2644
rect 11977 2635 12035 2641
rect 11977 2632 11989 2635
rect 11940 2604 11989 2632
rect 11940 2592 11946 2604
rect 11977 2601 11989 2604
rect 12023 2601 12035 2635
rect 11977 2595 12035 2601
rect 14366 2592 14372 2644
rect 14424 2632 14430 2644
rect 14461 2635 14519 2641
rect 14461 2632 14473 2635
rect 14424 2604 14473 2632
rect 14424 2592 14430 2604
rect 14461 2601 14473 2604
rect 14507 2601 14519 2635
rect 15838 2632 15844 2644
rect 15799 2604 15844 2632
rect 14461 2595 14519 2601
rect 15838 2592 15844 2604
rect 15896 2592 15902 2644
rect 16298 2592 16304 2644
rect 16356 2632 16362 2644
rect 17221 2635 17279 2641
rect 17221 2632 17233 2635
rect 16356 2604 17233 2632
rect 16356 2592 16362 2604
rect 17221 2601 17233 2604
rect 17267 2601 17279 2635
rect 17954 2632 17960 2644
rect 17915 2604 17960 2632
rect 17221 2595 17279 2601
rect 17954 2592 17960 2604
rect 18012 2592 18018 2644
rect 18616 2604 26234 2632
rect 4614 2564 4620 2576
rect 3988 2536 4620 2564
rect 1397 2499 1455 2505
rect 1397 2465 1409 2499
rect 1443 2465 1455 2499
rect 1578 2496 1584 2508
rect 1539 2468 1584 2496
rect 1397 2459 1455 2465
rect 1578 2456 1584 2468
rect 1636 2456 1642 2508
rect 2774 2496 2780 2508
rect 2735 2468 2780 2496
rect 2774 2456 2780 2468
rect 2832 2456 2838 2508
rect 3988 2505 4016 2536
rect 4614 2524 4620 2536
rect 4672 2524 4678 2576
rect 5166 2524 5172 2576
rect 5224 2564 5230 2576
rect 5224 2536 6868 2564
rect 5224 2524 5230 2536
rect 3973 2499 4031 2505
rect 3973 2465 3985 2499
rect 4019 2465 4031 2499
rect 4154 2496 4160 2508
rect 4115 2468 4160 2496
rect 3973 2459 4031 2465
rect 4154 2456 4160 2468
rect 4212 2456 4218 2508
rect 4522 2496 4528 2508
rect 4483 2468 4528 2496
rect 4522 2456 4528 2468
rect 4580 2456 4586 2508
rect 6362 2496 6368 2508
rect 6323 2468 6368 2496
rect 6362 2456 6368 2468
rect 6420 2456 6426 2508
rect 6546 2496 6552 2508
rect 6507 2468 6552 2496
rect 6546 2456 6552 2468
rect 6604 2456 6610 2508
rect 6840 2505 6868 2536
rect 9122 2524 9128 2576
rect 9180 2564 9186 2576
rect 9180 2536 9904 2564
rect 9180 2524 9186 2536
rect 6825 2499 6883 2505
rect 6825 2465 6837 2499
rect 6871 2465 6883 2499
rect 9030 2496 9036 2508
rect 8991 2468 9036 2496
rect 6825 2459 6883 2465
rect 9030 2456 9036 2468
rect 9088 2456 9094 2508
rect 9217 2499 9275 2505
rect 9217 2465 9229 2499
rect 9263 2496 9275 2499
rect 9766 2496 9772 2508
rect 9263 2468 9772 2496
rect 9263 2465 9275 2468
rect 9217 2459 9275 2465
rect 9766 2456 9772 2468
rect 9824 2456 9830 2508
rect 9876 2505 9904 2536
rect 9861 2499 9919 2505
rect 9861 2465 9873 2499
rect 9907 2465 9919 2499
rect 9861 2459 9919 2465
rect 11885 2431 11943 2437
rect 11885 2397 11897 2431
rect 11931 2428 11943 2431
rect 12434 2428 12440 2440
rect 11931 2400 12440 2428
rect 11931 2397 11943 2400
rect 11885 2391 11943 2397
rect 12434 2388 12440 2400
rect 12492 2388 12498 2440
rect 14090 2388 14096 2440
rect 14148 2428 14154 2440
rect 14369 2431 14427 2437
rect 14369 2428 14381 2431
rect 14148 2400 14381 2428
rect 14148 2388 14154 2400
rect 14369 2397 14381 2400
rect 14415 2397 14427 2431
rect 14369 2391 14427 2397
rect 15654 2388 15660 2440
rect 15712 2428 15718 2440
rect 15749 2431 15807 2437
rect 15749 2428 15761 2431
rect 15712 2400 15761 2428
rect 15712 2388 15718 2400
rect 15749 2397 15761 2400
rect 15795 2428 15807 2431
rect 18616 2428 18644 2604
rect 18690 2524 18696 2576
rect 18748 2564 18754 2576
rect 26206 2564 26234 2604
rect 26510 2592 26516 2644
rect 26568 2632 26574 2644
rect 27157 2635 27215 2641
rect 27157 2632 27169 2635
rect 26568 2604 27169 2632
rect 26568 2592 26574 2604
rect 27157 2601 27169 2604
rect 27203 2601 27215 2635
rect 27157 2595 27215 2601
rect 27062 2564 27068 2576
rect 18748 2536 20208 2564
rect 26206 2536 27068 2564
rect 18748 2524 18754 2536
rect 19429 2499 19487 2505
rect 19429 2465 19441 2499
rect 19475 2496 19487 2499
rect 20070 2496 20076 2508
rect 19475 2468 20076 2496
rect 19475 2465 19487 2468
rect 19429 2459 19487 2465
rect 20070 2456 20076 2468
rect 20128 2456 20134 2508
rect 20180 2505 20208 2536
rect 27062 2524 27068 2536
rect 27120 2524 27126 2576
rect 20165 2499 20223 2505
rect 20165 2465 20177 2499
rect 20211 2465 20223 2499
rect 20165 2459 20223 2465
rect 22005 2499 22063 2505
rect 22005 2465 22017 2499
rect 22051 2496 22063 2499
rect 22186 2496 22192 2508
rect 22051 2468 22192 2496
rect 22051 2465 22063 2468
rect 22005 2459 22063 2465
rect 22186 2456 22192 2468
rect 22244 2456 22250 2508
rect 23842 2456 23848 2508
rect 23900 2496 23906 2508
rect 24581 2499 24639 2505
rect 24581 2496 24593 2499
rect 23900 2468 24593 2496
rect 23900 2456 23906 2468
rect 24581 2465 24593 2468
rect 24627 2465 24639 2499
rect 24581 2459 24639 2465
rect 24765 2499 24823 2505
rect 24765 2465 24777 2499
rect 24811 2496 24823 2499
rect 27893 2499 27951 2505
rect 27893 2496 27905 2499
rect 24811 2468 27905 2496
rect 24811 2465 24823 2468
rect 24765 2459 24823 2465
rect 27893 2465 27905 2468
rect 27939 2465 27951 2499
rect 27893 2459 27951 2465
rect 15795 2400 18644 2428
rect 19245 2431 19303 2437
rect 15795 2397 15807 2400
rect 15749 2391 15807 2397
rect 19245 2397 19257 2431
rect 19291 2397 19303 2431
rect 19245 2391 19303 2397
rect 27801 2431 27859 2437
rect 27801 2397 27813 2431
rect 27847 2428 27859 2431
rect 27982 2428 27988 2440
rect 27847 2400 27988 2428
rect 27847 2397 27859 2400
rect 27801 2391 27859 2397
rect 16758 2320 16764 2372
rect 16816 2360 16822 2372
rect 17129 2363 17187 2369
rect 17129 2360 17141 2363
rect 16816 2332 17141 2360
rect 16816 2320 16822 2332
rect 17129 2329 17141 2332
rect 17175 2329 17187 2363
rect 19260 2360 19288 2391
rect 27982 2388 27988 2400
rect 28040 2388 28046 2440
rect 20162 2360 20168 2372
rect 19260 2332 20168 2360
rect 17129 2323 17187 2329
rect 20162 2320 20168 2332
rect 20220 2320 20226 2372
rect 22189 2363 22247 2369
rect 22189 2329 22201 2363
rect 22235 2360 22247 2363
rect 23750 2360 23756 2372
rect 22235 2332 23756 2360
rect 22235 2329 22247 2332
rect 22189 2323 22247 2329
rect 23750 2320 23756 2332
rect 23808 2320 23814 2372
rect 23845 2363 23903 2369
rect 23845 2329 23857 2363
rect 23891 2360 23903 2363
rect 25038 2360 25044 2372
rect 23891 2332 25044 2360
rect 23891 2329 23903 2332
rect 23845 2323 23903 2329
rect 25038 2320 25044 2332
rect 25096 2320 25102 2372
rect 26142 2320 26148 2372
rect 26200 2360 26206 2372
rect 26421 2363 26479 2369
rect 26421 2360 26433 2363
rect 26200 2332 26433 2360
rect 26200 2320 26206 2332
rect 26421 2329 26433 2332
rect 26467 2329 26479 2363
rect 26421 2323 26479 2329
rect 1104 2202 28888 2224
rect 1104 2150 10214 2202
rect 10266 2150 10278 2202
rect 10330 2150 10342 2202
rect 10394 2150 10406 2202
rect 10458 2150 10470 2202
rect 10522 2150 19478 2202
rect 19530 2150 19542 2202
rect 19594 2150 19606 2202
rect 19658 2150 19670 2202
rect 19722 2150 19734 2202
rect 19786 2150 28888 2202
rect 1104 2128 28888 2150
rect 3050 1776 3056 1828
rect 3108 1816 3114 1828
rect 7374 1816 7380 1828
rect 3108 1788 7380 1816
rect 3108 1776 3114 1788
rect 7374 1776 7380 1788
rect 7432 1776 7438 1828
<< via1 >>
rect 9036 40808 9088 40860
rect 23572 40808 23624 40860
rect 8852 40740 8904 40792
rect 15936 40740 15988 40792
rect 7564 40672 7616 40724
rect 13912 40672 13964 40724
rect 7656 40604 7708 40656
rect 20352 40604 20404 40656
rect 7472 40536 7524 40588
rect 23940 40536 23992 40588
rect 8944 40468 8996 40520
rect 26884 40468 26936 40520
rect 7380 40400 7432 40452
rect 22284 40400 22336 40452
rect 7196 40332 7248 40384
rect 22008 40332 22060 40384
rect 9312 40264 9364 40316
rect 23664 40264 23716 40316
rect 10324 40196 10376 40248
rect 26332 40196 26384 40248
rect 9864 40128 9916 40180
rect 8392 40060 8444 40112
rect 11060 40060 11112 40112
rect 12624 40128 12676 40180
rect 24768 40128 24820 40180
rect 13084 40060 13136 40112
rect 16580 40060 16632 40112
rect 7932 39992 7984 40044
rect 16948 39992 17000 40044
rect 18052 40060 18104 40112
rect 18880 40060 18932 40112
rect 21272 39992 21324 40044
rect 9680 39924 9732 39976
rect 8484 39856 8536 39908
rect 11888 39856 11940 39908
rect 12440 39856 12492 39908
rect 12716 39924 12768 39976
rect 22192 39924 22244 39976
rect 12992 39856 13044 39908
rect 14004 39856 14056 39908
rect 16580 39856 16632 39908
rect 16672 39856 16724 39908
rect 20812 39856 20864 39908
rect 6644 39788 6696 39840
rect 14280 39788 14332 39840
rect 15568 39788 15620 39840
rect 23480 39788 23532 39840
rect 5582 39686 5634 39738
rect 5646 39686 5698 39738
rect 5710 39686 5762 39738
rect 5774 39686 5826 39738
rect 5838 39686 5890 39738
rect 14846 39686 14898 39738
rect 14910 39686 14962 39738
rect 14974 39686 15026 39738
rect 15038 39686 15090 39738
rect 15102 39686 15154 39738
rect 24110 39686 24162 39738
rect 24174 39686 24226 39738
rect 24238 39686 24290 39738
rect 24302 39686 24354 39738
rect 24366 39686 24418 39738
rect 7104 39627 7156 39636
rect 7104 39593 7113 39627
rect 7113 39593 7147 39627
rect 7147 39593 7156 39627
rect 7104 39584 7156 39593
rect 1768 39423 1820 39432
rect 1768 39389 1777 39423
rect 1777 39389 1811 39423
rect 1811 39389 1820 39423
rect 1768 39380 1820 39389
rect 2412 39423 2464 39432
rect 2412 39389 2421 39423
rect 2421 39389 2455 39423
rect 2455 39389 2464 39423
rect 2412 39380 2464 39389
rect 5448 39516 5500 39568
rect 7012 39516 7064 39568
rect 10876 39584 10928 39636
rect 11060 39584 11112 39636
rect 17500 39584 17552 39636
rect 20168 39516 20220 39568
rect 4160 39448 4212 39500
rect 10140 39448 10192 39500
rect 10324 39491 10376 39500
rect 10324 39457 10333 39491
rect 10333 39457 10367 39491
rect 10367 39457 10376 39491
rect 10324 39448 10376 39457
rect 10692 39448 10744 39500
rect 11796 39491 11848 39500
rect 11796 39457 11805 39491
rect 11805 39457 11839 39491
rect 11839 39457 11848 39491
rect 11796 39448 11848 39457
rect 12256 39448 12308 39500
rect 12532 39448 12584 39500
rect 14096 39448 14148 39500
rect 15476 39491 15528 39500
rect 15476 39457 15485 39491
rect 15485 39457 15519 39491
rect 15519 39457 15528 39491
rect 15476 39448 15528 39457
rect 15660 39448 15712 39500
rect 19984 39491 20036 39500
rect 19984 39457 19993 39491
rect 19993 39457 20027 39491
rect 20027 39457 20036 39491
rect 19984 39448 20036 39457
rect 22008 39491 22060 39500
rect 22008 39457 22017 39491
rect 22017 39457 22051 39491
rect 22051 39457 22060 39491
rect 22008 39448 22060 39457
rect 22192 39491 22244 39500
rect 22192 39457 22201 39491
rect 22201 39457 22235 39491
rect 22235 39457 22244 39491
rect 22192 39448 22244 39457
rect 23848 39491 23900 39500
rect 23848 39457 23857 39491
rect 23857 39457 23891 39491
rect 23891 39457 23900 39491
rect 23848 39448 23900 39457
rect 24768 39491 24820 39500
rect 24768 39457 24777 39491
rect 24777 39457 24811 39491
rect 24811 39457 24820 39491
rect 24768 39448 24820 39457
rect 26056 39491 26108 39500
rect 26056 39457 26065 39491
rect 26065 39457 26099 39491
rect 26099 39457 26108 39491
rect 26056 39448 26108 39457
rect 1676 39244 1728 39296
rect 2504 39287 2556 39296
rect 2504 39253 2513 39287
rect 2513 39253 2547 39287
rect 2547 39253 2556 39287
rect 2504 39244 2556 39253
rect 3148 39287 3200 39296
rect 3148 39253 3157 39287
rect 3157 39253 3191 39287
rect 3191 39253 3200 39287
rect 3148 39244 3200 39253
rect 9680 39423 9732 39432
rect 9680 39389 9689 39423
rect 9689 39389 9723 39423
rect 9723 39389 9732 39423
rect 9680 39380 9732 39389
rect 10048 39380 10100 39432
rect 10784 39423 10836 39432
rect 10784 39389 10793 39423
rect 10793 39389 10827 39423
rect 10827 39389 10836 39423
rect 10784 39380 10836 39389
rect 10876 39380 10928 39432
rect 14280 39423 14332 39432
rect 3976 39355 4028 39364
rect 3976 39321 3985 39355
rect 3985 39321 4019 39355
rect 4019 39321 4028 39355
rect 3976 39312 4028 39321
rect 9772 39312 9824 39364
rect 11520 39312 11572 39364
rect 14280 39389 14289 39423
rect 14289 39389 14323 39423
rect 14323 39389 14332 39423
rect 14280 39380 14332 39389
rect 16672 39423 16724 39432
rect 14004 39312 14056 39364
rect 14464 39355 14516 39364
rect 14464 39321 14473 39355
rect 14473 39321 14507 39355
rect 14507 39321 14516 39355
rect 14464 39312 14516 39321
rect 14556 39312 14608 39364
rect 16672 39389 16681 39423
rect 16681 39389 16715 39423
rect 16715 39389 16724 39423
rect 16672 39380 16724 39389
rect 17592 39380 17644 39432
rect 19340 39380 19392 39432
rect 24584 39423 24636 39432
rect 24584 39389 24593 39423
rect 24593 39389 24627 39423
rect 24627 39389 24636 39423
rect 24584 39380 24636 39389
rect 5264 39244 5316 39296
rect 7104 39244 7156 39296
rect 10692 39244 10744 39296
rect 12348 39244 12400 39296
rect 12808 39244 12860 39296
rect 17316 39244 17368 39296
rect 17684 39244 17736 39296
rect 17868 39312 17920 39364
rect 18972 39312 19024 39364
rect 26792 39312 26844 39364
rect 27620 39355 27672 39364
rect 27620 39321 27629 39355
rect 27629 39321 27663 39355
rect 27663 39321 27672 39355
rect 27620 39312 27672 39321
rect 18604 39244 18656 39296
rect 19892 39244 19944 39296
rect 20996 39244 21048 39296
rect 10214 39142 10266 39194
rect 10278 39142 10330 39194
rect 10342 39142 10394 39194
rect 10406 39142 10458 39194
rect 10470 39142 10522 39194
rect 19478 39142 19530 39194
rect 19542 39142 19594 39194
rect 19606 39142 19658 39194
rect 19670 39142 19722 39194
rect 19734 39142 19786 39194
rect 14464 39040 14516 39092
rect 14556 39040 14608 39092
rect 15292 39040 15344 39092
rect 15476 39040 15528 39092
rect 1676 39015 1728 39024
rect 1676 38981 1685 39015
rect 1685 38981 1719 39015
rect 1719 38981 1728 39015
rect 1676 38972 1728 38981
rect 3148 38972 3200 39024
rect 7380 38947 7432 38956
rect 7380 38913 7389 38947
rect 7389 38913 7423 38947
rect 7423 38913 7432 38947
rect 7380 38904 7432 38913
rect 8668 38947 8720 38956
rect 8668 38913 8677 38947
rect 8677 38913 8711 38947
rect 8711 38913 8720 38947
rect 8668 38904 8720 38913
rect 9312 38947 9364 38956
rect 9312 38913 9321 38947
rect 9321 38913 9355 38947
rect 9355 38913 9364 38947
rect 9312 38904 9364 38913
rect 10876 38972 10928 39024
rect 15660 38972 15712 39024
rect 10232 38904 10284 38956
rect 11888 38904 11940 38956
rect 1492 38879 1544 38888
rect 1492 38845 1501 38879
rect 1501 38845 1535 38879
rect 1535 38845 1544 38879
rect 1492 38836 1544 38845
rect 2872 38879 2924 38888
rect 2872 38845 2881 38879
rect 2881 38845 2915 38879
rect 2915 38845 2924 38879
rect 2872 38836 2924 38845
rect 4620 38836 4672 38888
rect 4712 38879 4764 38888
rect 4712 38845 4721 38879
rect 4721 38845 4755 38879
rect 4755 38845 4764 38879
rect 4712 38836 4764 38845
rect 8576 38836 8628 38888
rect 9220 38836 9272 38888
rect 10324 38836 10376 38888
rect 12716 38904 12768 38956
rect 12992 38947 13044 38956
rect 12992 38913 13001 38947
rect 13001 38913 13035 38947
rect 13035 38913 13044 38947
rect 12992 38904 13044 38913
rect 14648 38904 14700 38956
rect 15568 38947 15620 38956
rect 15568 38913 15577 38947
rect 15577 38913 15611 38947
rect 15611 38913 15620 38947
rect 15568 38904 15620 38913
rect 13176 38879 13228 38888
rect 13176 38845 13185 38879
rect 13185 38845 13219 38879
rect 13219 38845 13228 38879
rect 13176 38836 13228 38845
rect 13544 38879 13596 38888
rect 13544 38845 13553 38879
rect 13553 38845 13587 38879
rect 13587 38845 13596 38879
rect 13544 38836 13596 38845
rect 14096 38836 14148 38888
rect 16764 38972 16816 39024
rect 16948 38972 17000 39024
rect 17684 39015 17736 39024
rect 17684 38981 17690 39015
rect 17690 38981 17724 39015
rect 17724 38981 17736 39015
rect 18420 39040 18472 39092
rect 17684 38972 17736 38981
rect 18328 38972 18380 39024
rect 18880 38972 18932 39024
rect 16488 38904 16540 38956
rect 17500 38947 17552 38956
rect 17500 38913 17509 38947
rect 17509 38913 17543 38947
rect 17543 38913 17552 38947
rect 17500 38904 17552 38913
rect 20076 38972 20128 39024
rect 20352 38972 20404 39024
rect 26976 39015 27028 39024
rect 26976 38981 26985 39015
rect 26985 38981 27019 39015
rect 27019 38981 27028 39015
rect 26976 38972 27028 38981
rect 27160 39015 27212 39024
rect 27160 38981 27185 39015
rect 27185 38981 27212 39015
rect 27160 38972 27212 38981
rect 1676 38768 1728 38820
rect 2412 38768 2464 38820
rect 8024 38811 8076 38820
rect 6552 38743 6604 38752
rect 6552 38709 6561 38743
rect 6561 38709 6595 38743
rect 6595 38709 6604 38743
rect 6552 38700 6604 38709
rect 8024 38777 8033 38811
rect 8033 38777 8067 38811
rect 8067 38777 8076 38811
rect 8024 38768 8076 38777
rect 11336 38768 11388 38820
rect 13268 38768 13320 38820
rect 13360 38768 13412 38820
rect 16212 38768 16264 38820
rect 19064 38836 19116 38888
rect 19800 38836 19852 38888
rect 9128 38700 9180 38752
rect 9220 38700 9272 38752
rect 10324 38700 10376 38752
rect 10508 38743 10560 38752
rect 10508 38709 10517 38743
rect 10517 38709 10551 38743
rect 10551 38709 10560 38743
rect 10508 38700 10560 38709
rect 11244 38700 11296 38752
rect 12532 38700 12584 38752
rect 13084 38700 13136 38752
rect 15476 38700 15528 38752
rect 15752 38700 15804 38752
rect 16304 38700 16356 38752
rect 17592 38700 17644 38752
rect 18328 38768 18380 38820
rect 20260 38904 20312 38956
rect 20720 38904 20772 38956
rect 22284 38947 22336 38956
rect 22284 38913 22293 38947
rect 22293 38913 22327 38947
rect 22327 38913 22336 38947
rect 22284 38904 22336 38913
rect 23664 38904 23716 38956
rect 27988 38947 28040 38956
rect 27988 38913 27997 38947
rect 27997 38913 28031 38947
rect 28031 38913 28040 38947
rect 27988 38904 28040 38913
rect 23204 38879 23256 38888
rect 23204 38845 23213 38879
rect 23213 38845 23247 38879
rect 23247 38845 23256 38879
rect 23204 38836 23256 38845
rect 25964 38836 26016 38888
rect 26148 38879 26200 38888
rect 26148 38845 26157 38879
rect 26157 38845 26191 38879
rect 26191 38845 26200 38879
rect 26148 38836 26200 38845
rect 18420 38700 18472 38752
rect 19892 38700 19944 38752
rect 20628 38700 20680 38752
rect 27436 38768 27488 38820
rect 27344 38743 27396 38752
rect 27344 38709 27353 38743
rect 27353 38709 27387 38743
rect 27387 38709 27396 38743
rect 27344 38700 27396 38709
rect 27528 38700 27580 38752
rect 5582 38598 5634 38650
rect 5646 38598 5698 38650
rect 5710 38598 5762 38650
rect 5774 38598 5826 38650
rect 5838 38598 5890 38650
rect 14846 38598 14898 38650
rect 14910 38598 14962 38650
rect 14974 38598 15026 38650
rect 15038 38598 15090 38650
rect 15102 38598 15154 38650
rect 24110 38598 24162 38650
rect 24174 38598 24226 38650
rect 24238 38598 24290 38650
rect 24302 38598 24354 38650
rect 24366 38598 24418 38650
rect 20 38496 72 38548
rect 1400 38496 1452 38548
rect 3240 38496 3292 38548
rect 4712 38496 4764 38548
rect 8392 38539 8444 38548
rect 8392 38505 8401 38539
rect 8401 38505 8435 38539
rect 8435 38505 8444 38539
rect 8392 38496 8444 38505
rect 9404 38496 9456 38548
rect 6552 38428 6604 38480
rect 7748 38471 7800 38480
rect 7748 38437 7757 38471
rect 7757 38437 7791 38471
rect 7791 38437 7800 38471
rect 7748 38428 7800 38437
rect 12164 38496 12216 38548
rect 12992 38496 13044 38548
rect 13176 38496 13228 38548
rect 18420 38496 18472 38548
rect 2504 38360 2556 38412
rect 2780 38403 2832 38412
rect 2780 38369 2789 38403
rect 2789 38369 2823 38403
rect 2823 38369 2832 38403
rect 2780 38360 2832 38369
rect 5172 38403 5224 38412
rect 5172 38369 5181 38403
rect 5181 38369 5215 38403
rect 5215 38369 5224 38403
rect 5172 38360 5224 38369
rect 5356 38360 5408 38412
rect 8576 38360 8628 38412
rect 4252 38292 4304 38344
rect 9404 38360 9456 38412
rect 9772 38403 9824 38412
rect 9772 38369 9781 38403
rect 9781 38369 9815 38403
rect 9815 38369 9824 38403
rect 9772 38360 9824 38369
rect 10140 38360 10192 38412
rect 10508 38403 10560 38412
rect 10508 38369 10517 38403
rect 10517 38369 10551 38403
rect 10551 38369 10560 38403
rect 10508 38360 10560 38369
rect 10968 38360 11020 38412
rect 14740 38428 14792 38480
rect 23664 38496 23716 38548
rect 26976 38496 27028 38548
rect 1952 38224 2004 38276
rect 2872 38224 2924 38276
rect 9496 38292 9548 38344
rect 10048 38292 10100 38344
rect 11796 38292 11848 38344
rect 12164 38292 12216 38344
rect 12624 38360 12676 38412
rect 15384 38360 15436 38412
rect 15568 38403 15620 38412
rect 15568 38369 15577 38403
rect 15577 38369 15611 38403
rect 15611 38369 15620 38403
rect 15568 38360 15620 38369
rect 15752 38403 15804 38412
rect 15752 38369 15761 38403
rect 15761 38369 15795 38403
rect 15795 38369 15804 38403
rect 15752 38360 15804 38369
rect 16120 38403 16172 38412
rect 16120 38369 16129 38403
rect 16129 38369 16163 38403
rect 16163 38369 16172 38403
rect 16120 38360 16172 38369
rect 16488 38360 16540 38412
rect 17868 38403 17920 38412
rect 12808 38292 12860 38344
rect 13176 38335 13228 38344
rect 13176 38301 13185 38335
rect 13185 38301 13219 38335
rect 13219 38301 13228 38335
rect 13176 38292 13228 38301
rect 13268 38292 13320 38344
rect 14832 38292 14884 38344
rect 15476 38292 15528 38344
rect 17868 38369 17877 38403
rect 17877 38369 17911 38403
rect 17911 38369 17920 38403
rect 17868 38360 17920 38369
rect 18696 38360 18748 38412
rect 20168 38403 20220 38412
rect 20168 38369 20177 38403
rect 20177 38369 20211 38403
rect 20211 38369 20220 38403
rect 20168 38360 20220 38369
rect 20536 38360 20588 38412
rect 21548 38292 21600 38344
rect 22928 38360 22980 38412
rect 23848 38360 23900 38412
rect 23664 38335 23716 38344
rect 5172 38224 5224 38276
rect 6368 38224 6420 38276
rect 8484 38224 8536 38276
rect 9128 38224 9180 38276
rect 10048 38156 10100 38208
rect 11796 38156 11848 38208
rect 11980 38156 12032 38208
rect 13176 38156 13228 38208
rect 14740 38224 14792 38276
rect 22008 38224 22060 38276
rect 22284 38224 22336 38276
rect 18236 38156 18288 38208
rect 18328 38156 18380 38208
rect 20904 38156 20956 38208
rect 23664 38301 23673 38335
rect 23673 38301 23707 38335
rect 23707 38301 23716 38335
rect 23664 38292 23716 38301
rect 23756 38224 23808 38276
rect 24860 38335 24912 38344
rect 24860 38301 24869 38335
rect 24869 38301 24903 38335
rect 24903 38301 24912 38335
rect 25044 38335 25096 38344
rect 24860 38292 24912 38301
rect 25044 38301 25053 38335
rect 25053 38301 25087 38335
rect 25087 38301 25096 38335
rect 25044 38292 25096 38301
rect 25596 38292 25648 38344
rect 26332 38403 26384 38412
rect 26332 38369 26341 38403
rect 26341 38369 26375 38403
rect 26375 38369 26384 38403
rect 26332 38360 26384 38369
rect 27712 38403 27764 38412
rect 27712 38369 27721 38403
rect 27721 38369 27755 38403
rect 27755 38369 27764 38403
rect 27712 38360 27764 38369
rect 25872 38335 25924 38344
rect 25872 38301 25881 38335
rect 25881 38301 25915 38335
rect 25915 38301 25924 38335
rect 25872 38292 25924 38301
rect 24952 38224 25004 38276
rect 22928 38156 22980 38208
rect 23848 38199 23900 38208
rect 23848 38165 23857 38199
rect 23857 38165 23891 38199
rect 23891 38165 23900 38199
rect 23848 38156 23900 38165
rect 24676 38156 24728 38208
rect 24768 38156 24820 38208
rect 25780 38224 25832 38276
rect 10214 38054 10266 38106
rect 10278 38054 10330 38106
rect 10342 38054 10394 38106
rect 10406 38054 10458 38106
rect 10470 38054 10522 38106
rect 19478 38054 19530 38106
rect 19542 38054 19594 38106
rect 19606 38054 19658 38106
rect 19670 38054 19722 38106
rect 19734 38054 19786 38106
rect 3792 37884 3844 37936
rect 6368 37859 6420 37868
rect 6368 37825 6377 37859
rect 6377 37825 6411 37859
rect 6411 37825 6420 37859
rect 6368 37816 6420 37825
rect 18328 37952 18380 38004
rect 19892 37995 19944 38004
rect 19892 37961 19901 37995
rect 19901 37961 19935 37995
rect 19935 37961 19944 37995
rect 19892 37952 19944 37961
rect 23388 37952 23440 38004
rect 25044 37952 25096 38004
rect 25136 37952 25188 38004
rect 2780 37791 2832 37800
rect 2780 37757 2789 37791
rect 2789 37757 2823 37791
rect 2823 37757 2832 37791
rect 3884 37791 3936 37800
rect 2780 37748 2832 37757
rect 3884 37757 3893 37791
rect 3893 37757 3927 37791
rect 3927 37757 3936 37791
rect 3884 37748 3936 37757
rect 4528 37791 4580 37800
rect 4528 37757 4537 37791
rect 4537 37757 4571 37791
rect 4571 37757 4580 37791
rect 4528 37748 4580 37757
rect 6920 37748 6972 37800
rect 9772 37816 9824 37868
rect 10416 37816 10468 37868
rect 10508 37816 10560 37868
rect 11060 37816 11112 37868
rect 11244 37816 11296 37868
rect 11428 37816 11480 37868
rect 11520 37816 11572 37868
rect 11888 37884 11940 37936
rect 12624 37884 12676 37936
rect 12808 37884 12860 37936
rect 14372 37816 14424 37868
rect 9128 37791 9180 37800
rect 9128 37757 9137 37791
rect 9137 37757 9171 37791
rect 9171 37757 9180 37791
rect 9128 37748 9180 37757
rect 9312 37748 9364 37800
rect 10048 37748 10100 37800
rect 10140 37748 10192 37800
rect 11612 37748 11664 37800
rect 11980 37748 12032 37800
rect 12164 37748 12216 37800
rect 12900 37791 12952 37800
rect 12900 37757 12909 37791
rect 12909 37757 12943 37791
rect 12943 37757 12952 37791
rect 12900 37748 12952 37757
rect 12992 37748 13044 37800
rect 13452 37748 13504 37800
rect 14648 37791 14700 37800
rect 14648 37757 14657 37791
rect 14657 37757 14691 37791
rect 14691 37757 14700 37791
rect 14648 37748 14700 37757
rect 15752 37791 15804 37800
rect 15752 37757 15761 37791
rect 15761 37757 15795 37791
rect 15795 37757 15804 37791
rect 15752 37748 15804 37757
rect 16212 37816 16264 37868
rect 27068 37884 27120 37936
rect 27988 37927 28040 37936
rect 27988 37893 27997 37927
rect 27997 37893 28031 37927
rect 28031 37893 28040 37927
rect 27988 37884 28040 37893
rect 17316 37816 17368 37868
rect 19064 37816 19116 37868
rect 16488 37748 16540 37800
rect 4436 37680 4488 37732
rect 8300 37680 8352 37732
rect 8484 37680 8536 37732
rect 16396 37680 16448 37732
rect 8116 37655 8168 37664
rect 8116 37621 8125 37655
rect 8125 37621 8159 37655
rect 8159 37621 8168 37655
rect 8116 37612 8168 37621
rect 8392 37612 8444 37664
rect 15200 37612 15252 37664
rect 18420 37680 18472 37732
rect 18052 37655 18104 37664
rect 18052 37621 18061 37655
rect 18061 37621 18095 37655
rect 18095 37621 18104 37655
rect 18052 37612 18104 37621
rect 19156 37612 19208 37664
rect 20352 37816 20404 37868
rect 20812 37859 20864 37868
rect 20812 37825 20821 37859
rect 20821 37825 20855 37859
rect 20855 37825 20864 37859
rect 20812 37816 20864 37825
rect 21824 37859 21876 37868
rect 21824 37825 21833 37859
rect 21833 37825 21867 37859
rect 21867 37825 21876 37859
rect 21824 37816 21876 37825
rect 24584 37859 24636 37868
rect 24584 37825 24593 37859
rect 24593 37825 24627 37859
rect 24627 37825 24636 37859
rect 24584 37816 24636 37825
rect 26792 37816 26844 37868
rect 19984 37748 20036 37800
rect 21640 37748 21692 37800
rect 22008 37791 22060 37800
rect 22008 37757 22017 37791
rect 22017 37757 22051 37791
rect 22051 37757 22060 37791
rect 22008 37748 22060 37757
rect 19616 37680 19668 37732
rect 21732 37680 21784 37732
rect 21916 37680 21968 37732
rect 23848 37748 23900 37800
rect 25044 37748 25096 37800
rect 25596 37748 25648 37800
rect 26424 37680 26476 37732
rect 20444 37612 20496 37664
rect 20812 37612 20864 37664
rect 22928 37612 22980 37664
rect 25688 37612 25740 37664
rect 28080 37655 28132 37664
rect 28080 37621 28089 37655
rect 28089 37621 28123 37655
rect 28123 37621 28132 37655
rect 28080 37612 28132 37621
rect 5582 37510 5634 37562
rect 5646 37510 5698 37562
rect 5710 37510 5762 37562
rect 5774 37510 5826 37562
rect 5838 37510 5890 37562
rect 14846 37510 14898 37562
rect 14910 37510 14962 37562
rect 14974 37510 15026 37562
rect 15038 37510 15090 37562
rect 15102 37510 15154 37562
rect 24110 37510 24162 37562
rect 24174 37510 24226 37562
rect 24238 37510 24290 37562
rect 24302 37510 24354 37562
rect 24366 37510 24418 37562
rect 3884 37408 3936 37460
rect 7196 37408 7248 37460
rect 7840 37408 7892 37460
rect 8116 37408 8168 37460
rect 17316 37408 17368 37460
rect 17868 37408 17920 37460
rect 18328 37408 18380 37460
rect 25412 37408 25464 37460
rect 25596 37408 25648 37460
rect 1860 37315 1912 37324
rect 1860 37281 1869 37315
rect 1869 37281 1903 37315
rect 1903 37281 1912 37315
rect 1860 37272 1912 37281
rect 5448 37315 5500 37324
rect 5448 37281 5457 37315
rect 5457 37281 5491 37315
rect 5491 37281 5500 37315
rect 5448 37272 5500 37281
rect 9588 37340 9640 37392
rect 9772 37383 9824 37392
rect 9772 37349 9781 37383
rect 9781 37349 9815 37383
rect 9815 37349 9824 37383
rect 9772 37340 9824 37349
rect 11428 37340 11480 37392
rect 11520 37340 11572 37392
rect 12716 37340 12768 37392
rect 11980 37315 12032 37324
rect 4344 37204 4396 37256
rect 8116 37204 8168 37256
rect 9128 37247 9180 37256
rect 9128 37213 9137 37247
rect 9137 37213 9171 37247
rect 9171 37213 9180 37247
rect 9128 37204 9180 37213
rect 9680 37204 9732 37256
rect 9772 37204 9824 37256
rect 10416 37247 10468 37256
rect 10416 37213 10425 37247
rect 10425 37213 10459 37247
rect 10459 37213 10468 37247
rect 10416 37204 10468 37213
rect 11980 37281 11989 37315
rect 11989 37281 12023 37315
rect 12023 37281 12032 37315
rect 11980 37272 12032 37281
rect 12532 37272 12584 37324
rect 12992 37272 13044 37324
rect 14188 37272 14240 37324
rect 16396 37315 16448 37324
rect 16396 37281 16405 37315
rect 16405 37281 16439 37315
rect 16439 37281 16448 37315
rect 16396 37272 16448 37281
rect 1584 37179 1636 37188
rect 1584 37145 1593 37179
rect 1593 37145 1627 37179
rect 1627 37145 1636 37179
rect 1584 37136 1636 37145
rect 4252 37136 4304 37188
rect 4712 37136 4764 37188
rect 10692 37136 10744 37188
rect 10876 37179 10928 37188
rect 10876 37145 10885 37179
rect 10885 37145 10919 37179
rect 10919 37145 10928 37179
rect 10876 37136 10928 37145
rect 11060 37136 11112 37188
rect 12256 37136 12308 37188
rect 13636 37204 13688 37256
rect 14096 37204 14148 37256
rect 13728 37136 13780 37188
rect 3884 37068 3936 37120
rect 13084 37068 13136 37120
rect 13268 37068 13320 37120
rect 16948 37204 17000 37256
rect 21364 37340 21416 37392
rect 18052 37272 18104 37324
rect 18144 37204 18196 37256
rect 18328 37204 18380 37256
rect 18696 37204 18748 37256
rect 20352 37247 20404 37256
rect 19616 37179 19668 37188
rect 15752 37068 15804 37120
rect 16028 37068 16080 37120
rect 19616 37145 19625 37179
rect 19625 37145 19659 37179
rect 19659 37145 19668 37179
rect 19616 37136 19668 37145
rect 20352 37213 20361 37247
rect 20361 37213 20395 37247
rect 20395 37213 20404 37247
rect 20352 37204 20404 37213
rect 21456 37247 21508 37256
rect 20904 37179 20956 37188
rect 20904 37145 20913 37179
rect 20913 37145 20947 37179
rect 20947 37145 20956 37179
rect 20904 37136 20956 37145
rect 21456 37213 21465 37247
rect 21465 37213 21499 37247
rect 21499 37213 21508 37247
rect 21456 37204 21508 37213
rect 23480 37272 23532 37324
rect 23848 37272 23900 37324
rect 26516 37315 26568 37324
rect 26516 37281 26525 37315
rect 26525 37281 26559 37315
rect 26559 37281 26568 37315
rect 26516 37272 26568 37281
rect 22008 37136 22060 37188
rect 17960 37068 18012 37120
rect 19156 37068 19208 37120
rect 24492 37204 24544 37256
rect 24676 37247 24728 37256
rect 24676 37213 24710 37247
rect 24710 37213 24728 37247
rect 24676 37204 24728 37213
rect 26240 37204 26292 37256
rect 28172 37247 28224 37256
rect 28172 37213 28181 37247
rect 28181 37213 28215 37247
rect 28215 37213 28224 37247
rect 28172 37204 28224 37213
rect 22560 37136 22612 37188
rect 22836 37136 22888 37188
rect 23112 37068 23164 37120
rect 23664 37068 23716 37120
rect 28080 37068 28132 37120
rect 10214 36966 10266 37018
rect 10278 36966 10330 37018
rect 10342 36966 10394 37018
rect 10406 36966 10458 37018
rect 10470 36966 10522 37018
rect 19478 36966 19530 37018
rect 19542 36966 19594 37018
rect 19606 36966 19658 37018
rect 19670 36966 19722 37018
rect 19734 36966 19786 37018
rect 1584 36907 1636 36916
rect 1584 36873 1593 36907
rect 1593 36873 1627 36907
rect 1627 36873 1636 36907
rect 1584 36864 1636 36873
rect 2596 36864 2648 36916
rect 1584 36728 1636 36780
rect 4988 36839 5040 36848
rect 4988 36805 4997 36839
rect 4997 36805 5031 36839
rect 5031 36805 5040 36839
rect 4988 36796 5040 36805
rect 5356 36796 5408 36848
rect 2044 36592 2096 36644
rect 4344 36728 4396 36780
rect 5172 36728 5224 36780
rect 7288 36728 7340 36780
rect 3700 36703 3752 36712
rect 3700 36669 3709 36703
rect 3709 36669 3743 36703
rect 3743 36669 3752 36703
rect 3700 36660 3752 36669
rect 9680 36864 9732 36916
rect 12440 36864 12492 36916
rect 12532 36864 12584 36916
rect 8852 36796 8904 36848
rect 8208 36728 8260 36780
rect 8484 36771 8536 36780
rect 8484 36737 8493 36771
rect 8493 36737 8527 36771
rect 8527 36737 8536 36771
rect 8484 36728 8536 36737
rect 8944 36771 8996 36780
rect 8944 36737 8953 36771
rect 8953 36737 8987 36771
rect 8987 36737 8996 36771
rect 8944 36728 8996 36737
rect 7932 36660 7984 36712
rect 9220 36728 9272 36780
rect 11060 36796 11112 36848
rect 12164 36796 12216 36848
rect 12624 36796 12676 36848
rect 13268 36796 13320 36848
rect 14648 36864 14700 36916
rect 15016 36907 15068 36916
rect 15016 36873 15025 36907
rect 15025 36873 15059 36907
rect 15059 36873 15068 36907
rect 15016 36864 15068 36873
rect 15476 36864 15528 36916
rect 18144 36864 18196 36916
rect 20168 36864 20220 36916
rect 21456 36864 21508 36916
rect 22376 36864 22428 36916
rect 22560 36907 22612 36916
rect 22560 36873 22569 36907
rect 22569 36873 22603 36907
rect 22603 36873 22612 36907
rect 22560 36864 22612 36873
rect 22652 36864 22704 36916
rect 24124 36864 24176 36916
rect 26424 36864 26476 36916
rect 26976 36864 27028 36916
rect 9772 36771 9824 36780
rect 9772 36737 9781 36771
rect 9781 36737 9815 36771
rect 9815 36737 9824 36771
rect 9772 36728 9824 36737
rect 10048 36728 10100 36780
rect 10416 36728 10468 36780
rect 10784 36771 10836 36780
rect 9404 36660 9456 36712
rect 10784 36737 10793 36771
rect 10793 36737 10827 36771
rect 10827 36737 10836 36771
rect 10784 36728 10836 36737
rect 10968 36728 11020 36780
rect 11428 36728 11480 36780
rect 11520 36660 11572 36712
rect 8116 36524 8168 36576
rect 10324 36524 10376 36576
rect 11612 36592 11664 36644
rect 13544 36728 13596 36780
rect 13636 36703 13688 36712
rect 11796 36524 11848 36576
rect 13636 36669 13645 36703
rect 13645 36669 13679 36703
rect 13679 36669 13688 36703
rect 13636 36660 13688 36669
rect 15016 36728 15068 36780
rect 15568 36728 15620 36780
rect 15752 36771 15804 36780
rect 15752 36737 15761 36771
rect 15761 36737 15795 36771
rect 15795 36737 15804 36771
rect 15752 36728 15804 36737
rect 15844 36771 15896 36780
rect 15844 36737 15853 36771
rect 15853 36737 15887 36771
rect 15887 36737 15896 36771
rect 15844 36728 15896 36737
rect 16028 36660 16080 36712
rect 16212 36660 16264 36712
rect 18052 36728 18104 36780
rect 19064 36728 19116 36780
rect 20904 36728 20956 36780
rect 21456 36728 21508 36780
rect 21916 36771 21968 36780
rect 21916 36737 21925 36771
rect 21925 36737 21959 36771
rect 21959 36737 21968 36771
rect 21916 36728 21968 36737
rect 23296 36796 23348 36848
rect 24952 36796 25004 36848
rect 17040 36703 17092 36712
rect 17040 36669 17049 36703
rect 17049 36669 17083 36703
rect 17083 36669 17092 36703
rect 17040 36660 17092 36669
rect 13084 36592 13136 36644
rect 16396 36592 16448 36644
rect 19156 36660 19208 36712
rect 20812 36660 20864 36712
rect 23020 36771 23072 36780
rect 23020 36737 23029 36771
rect 23029 36737 23063 36771
rect 23063 36737 23072 36771
rect 23020 36728 23072 36737
rect 23112 36660 23164 36712
rect 23480 36728 23532 36780
rect 24124 36771 24176 36780
rect 24124 36737 24133 36771
rect 24133 36737 24167 36771
rect 24167 36737 24176 36771
rect 24124 36728 24176 36737
rect 24584 36771 24636 36780
rect 24584 36737 24593 36771
rect 24593 36737 24627 36771
rect 24627 36737 24636 36771
rect 24584 36728 24636 36737
rect 28356 36796 28408 36848
rect 27160 36771 27212 36780
rect 27160 36737 27169 36771
rect 27169 36737 27203 36771
rect 27203 36737 27212 36771
rect 27436 36771 27488 36780
rect 27160 36728 27212 36737
rect 27436 36737 27445 36771
rect 27445 36737 27479 36771
rect 27479 36737 27488 36771
rect 27436 36728 27488 36737
rect 23388 36660 23440 36712
rect 23664 36660 23716 36712
rect 18512 36592 18564 36644
rect 19248 36592 19300 36644
rect 13452 36524 13504 36576
rect 21548 36592 21600 36644
rect 21824 36592 21876 36644
rect 26884 36660 26936 36712
rect 27068 36660 27120 36712
rect 28356 36660 28408 36712
rect 27620 36592 27672 36644
rect 20812 36524 20864 36576
rect 24768 36524 24820 36576
rect 27896 36524 27948 36576
rect 5582 36422 5634 36474
rect 5646 36422 5698 36474
rect 5710 36422 5762 36474
rect 5774 36422 5826 36474
rect 5838 36422 5890 36474
rect 14846 36422 14898 36474
rect 14910 36422 14962 36474
rect 14974 36422 15026 36474
rect 15038 36422 15090 36474
rect 15102 36422 15154 36474
rect 24110 36422 24162 36474
rect 24174 36422 24226 36474
rect 24238 36422 24290 36474
rect 24302 36422 24354 36474
rect 24366 36422 24418 36474
rect 1492 36320 1544 36372
rect 3976 36320 4028 36372
rect 4620 36363 4672 36372
rect 4620 36329 4629 36363
rect 4629 36329 4663 36363
rect 4663 36329 4672 36363
rect 4620 36320 4672 36329
rect 5264 36363 5316 36372
rect 5264 36329 5273 36363
rect 5273 36329 5307 36363
rect 5307 36329 5316 36363
rect 5264 36320 5316 36329
rect 6920 36320 6972 36372
rect 7104 36363 7156 36372
rect 7104 36329 7113 36363
rect 7113 36329 7147 36363
rect 7147 36329 7156 36363
rect 7104 36320 7156 36329
rect 6736 36252 6788 36304
rect 9312 36320 9364 36372
rect 9588 36363 9640 36372
rect 9588 36329 9597 36363
rect 9597 36329 9631 36363
rect 9631 36329 9640 36363
rect 9588 36320 9640 36329
rect 7564 36295 7616 36304
rect 7564 36261 7573 36295
rect 7573 36261 7607 36295
rect 7607 36261 7616 36295
rect 7564 36252 7616 36261
rect 8944 36295 8996 36304
rect 1584 36184 1636 36236
rect 6368 36184 6420 36236
rect 8944 36261 8953 36295
rect 8953 36261 8987 36295
rect 8987 36261 8996 36295
rect 8944 36252 8996 36261
rect 9128 36252 9180 36304
rect 10600 36252 10652 36304
rect 13636 36320 13688 36372
rect 13728 36320 13780 36372
rect 14372 36320 14424 36372
rect 14464 36320 14516 36372
rect 15384 36320 15436 36372
rect 15936 36320 15988 36372
rect 12992 36252 13044 36304
rect 14004 36252 14056 36304
rect 15292 36252 15344 36304
rect 15844 36252 15896 36304
rect 17868 36320 17920 36372
rect 18880 36252 18932 36304
rect 19524 36320 19576 36372
rect 21824 36252 21876 36304
rect 22008 36295 22060 36304
rect 22008 36261 22017 36295
rect 22017 36261 22051 36295
rect 22051 36261 22060 36295
rect 22008 36252 22060 36261
rect 23020 36320 23072 36372
rect 23572 36320 23624 36372
rect 24676 36320 24728 36372
rect 24860 36320 24912 36372
rect 27436 36320 27488 36372
rect 25872 36295 25924 36304
rect 10784 36184 10836 36236
rect 11796 36227 11848 36236
rect 11796 36193 11805 36227
rect 11805 36193 11839 36227
rect 11839 36193 11848 36227
rect 11796 36184 11848 36193
rect 14096 36227 14148 36236
rect 14096 36193 14105 36227
rect 14105 36193 14139 36227
rect 14139 36193 14148 36227
rect 14096 36184 14148 36193
rect 15660 36184 15712 36236
rect 16396 36184 16448 36236
rect 2596 36159 2648 36168
rect 2596 36125 2605 36159
rect 2605 36125 2639 36159
rect 2639 36125 2648 36159
rect 2596 36116 2648 36125
rect 3700 36116 3752 36168
rect 7840 36116 7892 36168
rect 8392 36159 8444 36168
rect 8392 36125 8401 36159
rect 8401 36125 8435 36159
rect 8435 36125 8444 36159
rect 8392 36116 8444 36125
rect 9772 36159 9824 36168
rect 9772 36125 9781 36159
rect 9781 36125 9815 36159
rect 9815 36125 9824 36159
rect 9772 36116 9824 36125
rect 10968 36116 11020 36168
rect 11060 36159 11112 36168
rect 11060 36125 11069 36159
rect 11069 36125 11103 36159
rect 11103 36125 11112 36159
rect 11060 36116 11112 36125
rect 9220 36048 9272 36100
rect 11612 36048 11664 36100
rect 12992 36116 13044 36168
rect 14188 36116 14240 36168
rect 16120 36159 16172 36168
rect 16120 36125 16129 36159
rect 16129 36125 16163 36159
rect 16163 36125 16172 36159
rect 16120 36116 16172 36125
rect 16212 36116 16264 36168
rect 18512 36184 18564 36236
rect 19524 36184 19576 36236
rect 19616 36184 19668 36236
rect 9956 35980 10008 36032
rect 10048 35980 10100 36032
rect 10876 35980 10928 36032
rect 10968 35980 11020 36032
rect 12164 35980 12216 36032
rect 12440 35980 12492 36032
rect 13636 36048 13688 36100
rect 13820 35980 13872 36032
rect 13912 35980 13964 36032
rect 17224 36048 17276 36100
rect 20352 36159 20404 36168
rect 18696 36048 18748 36100
rect 19340 36048 19392 36100
rect 20352 36125 20361 36159
rect 20361 36125 20395 36159
rect 20395 36125 20404 36159
rect 20352 36116 20404 36125
rect 19892 36048 19944 36100
rect 19984 36048 20036 36100
rect 21548 36116 21600 36168
rect 21180 36048 21232 36100
rect 21916 36116 21968 36168
rect 22284 36116 22336 36168
rect 22652 36116 22704 36168
rect 22836 36116 22888 36168
rect 22560 36048 22612 36100
rect 23388 36184 23440 36236
rect 23756 36184 23808 36236
rect 25872 36261 25881 36295
rect 25881 36261 25915 36295
rect 25915 36261 25924 36295
rect 25872 36252 25924 36261
rect 25228 36184 25280 36236
rect 28172 36227 28224 36236
rect 28172 36193 28181 36227
rect 28181 36193 28215 36227
rect 28215 36193 28224 36227
rect 28172 36184 28224 36193
rect 23204 36159 23256 36168
rect 23204 36125 23213 36159
rect 23213 36125 23247 36159
rect 23247 36125 23256 36159
rect 23204 36116 23256 36125
rect 25596 36116 25648 36168
rect 26332 36159 26384 36168
rect 26332 36125 26341 36159
rect 26341 36125 26375 36159
rect 26375 36125 26384 36159
rect 26332 36116 26384 36125
rect 14556 35980 14608 36032
rect 16672 35980 16724 36032
rect 17776 35980 17828 36032
rect 18328 35980 18380 36032
rect 20812 35980 20864 36032
rect 22744 35980 22796 36032
rect 23756 35980 23808 36032
rect 25136 35980 25188 36032
rect 25504 36091 25556 36100
rect 25504 36057 25513 36091
rect 25513 36057 25547 36091
rect 25547 36057 25556 36091
rect 25504 36048 25556 36057
rect 27252 35980 27304 36032
rect 10214 35878 10266 35930
rect 10278 35878 10330 35930
rect 10342 35878 10394 35930
rect 10406 35878 10458 35930
rect 10470 35878 10522 35930
rect 19478 35878 19530 35930
rect 19542 35878 19594 35930
rect 19606 35878 19658 35930
rect 19670 35878 19722 35930
rect 19734 35878 19786 35930
rect 3792 35776 3844 35828
rect 8024 35819 8076 35828
rect 8024 35785 8033 35819
rect 8033 35785 8067 35819
rect 8067 35785 8076 35819
rect 8024 35776 8076 35785
rect 9220 35776 9272 35828
rect 11980 35776 12032 35828
rect 12348 35776 12400 35828
rect 7380 35708 7432 35760
rect 4436 35640 4488 35692
rect 6644 35640 6696 35692
rect 7564 35683 7616 35692
rect 7564 35649 7573 35683
rect 7573 35649 7607 35683
rect 7607 35649 7616 35683
rect 7564 35640 7616 35649
rect 1768 35572 1820 35624
rect 2872 35615 2924 35624
rect 2872 35581 2881 35615
rect 2881 35581 2915 35615
rect 2915 35581 2924 35615
rect 2872 35572 2924 35581
rect 4528 35572 4580 35624
rect 8208 35683 8260 35692
rect 8208 35649 8217 35683
rect 8217 35649 8251 35683
rect 8251 35649 8260 35683
rect 8208 35640 8260 35649
rect 9312 35683 9364 35692
rect 5908 35504 5960 35556
rect 8760 35504 8812 35556
rect 9312 35649 9321 35683
rect 9321 35649 9355 35683
rect 9355 35649 9364 35683
rect 9312 35640 9364 35649
rect 9496 35683 9548 35692
rect 9496 35649 9505 35683
rect 9505 35649 9539 35683
rect 9539 35649 9548 35683
rect 9496 35640 9548 35649
rect 9956 35683 10008 35692
rect 9036 35572 9088 35624
rect 9956 35649 9965 35683
rect 9965 35649 9999 35683
rect 9999 35649 10008 35683
rect 9956 35640 10008 35649
rect 9864 35572 9916 35624
rect 10232 35708 10284 35760
rect 11060 35708 11112 35760
rect 12624 35708 12676 35760
rect 12808 35708 12860 35760
rect 12992 35708 13044 35760
rect 13268 35708 13320 35760
rect 11428 35640 11480 35692
rect 12256 35640 12308 35692
rect 12348 35640 12400 35692
rect 13084 35640 13136 35692
rect 13452 35640 13504 35692
rect 13636 35708 13688 35760
rect 13912 35776 13964 35828
rect 15200 35776 15252 35828
rect 16212 35776 16264 35828
rect 16764 35776 16816 35828
rect 18052 35776 18104 35828
rect 18328 35776 18380 35828
rect 10876 35572 10928 35624
rect 11796 35572 11848 35624
rect 12072 35572 12124 35624
rect 12164 35572 12216 35624
rect 14188 35615 14240 35624
rect 13268 35504 13320 35556
rect 13452 35504 13504 35556
rect 3424 35436 3476 35488
rect 10232 35436 10284 35488
rect 10324 35436 10376 35488
rect 11520 35436 11572 35488
rect 12716 35436 12768 35488
rect 12808 35436 12860 35488
rect 14188 35581 14197 35615
rect 14197 35581 14231 35615
rect 14231 35581 14240 35615
rect 14188 35572 14240 35581
rect 14372 35683 14424 35692
rect 14372 35649 14381 35683
rect 14381 35649 14415 35683
rect 14415 35649 14424 35683
rect 15292 35683 15344 35692
rect 14372 35640 14424 35649
rect 15292 35649 15301 35683
rect 15301 35649 15335 35683
rect 15335 35649 15344 35683
rect 15292 35640 15344 35649
rect 15752 35708 15804 35760
rect 15936 35708 15988 35760
rect 17224 35708 17276 35760
rect 18420 35751 18472 35760
rect 18420 35717 18429 35751
rect 18429 35717 18463 35751
rect 18463 35717 18472 35751
rect 18420 35708 18472 35717
rect 18880 35776 18932 35828
rect 18696 35708 18748 35760
rect 15568 35683 15620 35692
rect 15568 35649 15577 35683
rect 15577 35649 15611 35683
rect 15611 35649 15620 35683
rect 16672 35683 16724 35692
rect 15568 35640 15620 35649
rect 16672 35649 16681 35683
rect 16681 35649 16715 35683
rect 16715 35649 16724 35683
rect 16672 35640 16724 35649
rect 17684 35640 17736 35692
rect 18144 35640 18196 35692
rect 20812 35776 20864 35828
rect 19064 35708 19116 35760
rect 19248 35708 19300 35760
rect 19432 35708 19484 35760
rect 19616 35708 19668 35760
rect 19800 35708 19852 35760
rect 20536 35708 20588 35760
rect 22100 35776 22152 35828
rect 23848 35776 23900 35828
rect 21548 35708 21600 35760
rect 25228 35776 25280 35828
rect 19340 35640 19392 35692
rect 20904 35683 20956 35692
rect 20904 35649 20913 35683
rect 20913 35649 20947 35683
rect 20947 35649 20956 35683
rect 20904 35640 20956 35649
rect 13636 35504 13688 35556
rect 15568 35504 15620 35556
rect 17224 35504 17276 35556
rect 19524 35572 19576 35624
rect 13728 35479 13780 35488
rect 13728 35445 13737 35479
rect 13737 35445 13771 35479
rect 13771 35445 13780 35479
rect 13728 35436 13780 35445
rect 14004 35436 14056 35488
rect 14648 35436 14700 35488
rect 15292 35436 15344 35488
rect 15476 35479 15528 35488
rect 15476 35445 15485 35479
rect 15485 35445 15519 35479
rect 15519 35445 15528 35479
rect 15476 35436 15528 35445
rect 16304 35436 16356 35488
rect 17868 35436 17920 35488
rect 19984 35504 20036 35556
rect 20352 35572 20404 35624
rect 19892 35436 19944 35488
rect 20812 35572 20864 35624
rect 21088 35615 21140 35624
rect 21088 35581 21122 35615
rect 21122 35581 21140 35615
rect 21088 35572 21140 35581
rect 21272 35504 21324 35556
rect 21548 35436 21600 35488
rect 21916 35640 21968 35692
rect 22284 35640 22336 35692
rect 22744 35640 22796 35692
rect 23756 35640 23808 35692
rect 24584 35708 24636 35760
rect 24492 35640 24544 35692
rect 26976 35683 27028 35692
rect 26976 35649 26985 35683
rect 26985 35649 27019 35683
rect 27019 35649 27028 35683
rect 26976 35640 27028 35649
rect 27344 35708 27396 35760
rect 27252 35683 27304 35692
rect 27252 35649 27261 35683
rect 27261 35649 27295 35683
rect 27295 35649 27304 35683
rect 27252 35640 27304 35649
rect 22008 35504 22060 35556
rect 22560 35572 22612 35624
rect 23572 35572 23624 35624
rect 27436 35572 27488 35624
rect 22468 35504 22520 35556
rect 23388 35504 23440 35556
rect 24492 35504 24544 35556
rect 24768 35504 24820 35556
rect 26424 35547 26476 35556
rect 26424 35513 26433 35547
rect 26433 35513 26467 35547
rect 26467 35513 26476 35547
rect 26424 35504 26476 35513
rect 22652 35436 22704 35488
rect 22744 35436 22796 35488
rect 23480 35436 23532 35488
rect 23756 35479 23808 35488
rect 23756 35445 23765 35479
rect 23765 35445 23799 35479
rect 23799 35445 23808 35479
rect 23756 35436 23808 35445
rect 23848 35436 23900 35488
rect 25320 35436 25372 35488
rect 27344 35436 27396 35488
rect 5582 35334 5634 35386
rect 5646 35334 5698 35386
rect 5710 35334 5762 35386
rect 5774 35334 5826 35386
rect 5838 35334 5890 35386
rect 14846 35334 14898 35386
rect 14910 35334 14962 35386
rect 14974 35334 15026 35386
rect 15038 35334 15090 35386
rect 15102 35334 15154 35386
rect 24110 35334 24162 35386
rect 24174 35334 24226 35386
rect 24238 35334 24290 35386
rect 24302 35334 24354 35386
rect 24366 35334 24418 35386
rect 1768 35275 1820 35284
rect 1768 35241 1777 35275
rect 1777 35241 1811 35275
rect 1811 35241 1820 35275
rect 1768 35232 1820 35241
rect 3884 35232 3936 35284
rect 4528 35232 4580 35284
rect 6276 35275 6328 35284
rect 6276 35241 6285 35275
rect 6285 35241 6319 35275
rect 6319 35241 6328 35275
rect 6276 35232 6328 35241
rect 9220 35275 9272 35284
rect 9220 35241 9229 35275
rect 9229 35241 9263 35275
rect 9263 35241 9272 35275
rect 9220 35232 9272 35241
rect 9588 35232 9640 35284
rect 10968 35232 11020 35284
rect 11612 35232 11664 35284
rect 5908 35164 5960 35216
rect 8024 35164 8076 35216
rect 10140 35164 10192 35216
rect 10416 35164 10468 35216
rect 11244 35164 11296 35216
rect 11428 35164 11480 35216
rect 13452 35164 13504 35216
rect 7288 35096 7340 35148
rect 2412 35071 2464 35080
rect 2412 35037 2421 35071
rect 2421 35037 2455 35071
rect 2455 35037 2464 35071
rect 2412 35028 2464 35037
rect 3240 35071 3292 35080
rect 3240 35037 3249 35071
rect 3249 35037 3283 35071
rect 3283 35037 3292 35071
rect 3240 35028 3292 35037
rect 4160 35028 4212 35080
rect 6000 35028 6052 35080
rect 6736 35028 6788 35080
rect 7104 35071 7156 35080
rect 7104 35037 7113 35071
rect 7113 35037 7147 35071
rect 7147 35037 7156 35071
rect 7104 35028 7156 35037
rect 8944 35096 8996 35148
rect 8392 35071 8444 35080
rect 8392 35037 8401 35071
rect 8401 35037 8435 35071
rect 8435 35037 8444 35071
rect 8392 35028 8444 35037
rect 9128 35071 9180 35080
rect 9128 35037 9137 35071
rect 9137 35037 9171 35071
rect 9171 35037 9180 35071
rect 9128 35028 9180 35037
rect 9220 35028 9272 35080
rect 9404 35028 9456 35080
rect 12164 35096 12216 35148
rect 12992 35096 13044 35148
rect 15568 35164 15620 35216
rect 16672 35164 16724 35216
rect 17040 35207 17092 35216
rect 17040 35173 17049 35207
rect 17049 35173 17083 35207
rect 17083 35173 17092 35207
rect 17040 35164 17092 35173
rect 17960 35164 18012 35216
rect 18236 35207 18288 35216
rect 18236 35173 18245 35207
rect 18245 35173 18279 35207
rect 18279 35173 18288 35207
rect 18236 35164 18288 35173
rect 18420 35232 18472 35284
rect 18604 35164 18656 35216
rect 19156 35164 19208 35216
rect 19248 35164 19300 35216
rect 19800 35164 19852 35216
rect 15660 35139 15712 35148
rect 10324 35028 10376 35080
rect 2136 34960 2188 35012
rect 3792 34960 3844 35012
rect 7840 34960 7892 35012
rect 10232 34960 10284 35012
rect 11244 35028 11296 35080
rect 11336 35028 11388 35080
rect 12256 35028 12308 35080
rect 12532 35028 12584 35080
rect 12900 35028 12952 35080
rect 13912 35028 13964 35080
rect 14096 35071 14148 35080
rect 14096 35037 14105 35071
rect 14105 35037 14139 35071
rect 14139 35037 14148 35071
rect 14096 35028 14148 35037
rect 14372 35028 14424 35080
rect 14924 35071 14976 35080
rect 14924 35037 14933 35071
rect 14933 35037 14967 35071
rect 14967 35037 14976 35071
rect 14924 35028 14976 35037
rect 15108 35071 15160 35080
rect 15108 35037 15117 35071
rect 15117 35037 15151 35071
rect 15151 35037 15160 35071
rect 15108 35028 15160 35037
rect 15200 35071 15252 35080
rect 15200 35037 15209 35071
rect 15209 35037 15243 35071
rect 15243 35037 15252 35071
rect 15660 35105 15669 35139
rect 15669 35105 15703 35139
rect 15703 35105 15712 35139
rect 15660 35096 15712 35105
rect 17132 35096 17184 35148
rect 15200 35028 15252 35037
rect 17316 35028 17368 35080
rect 18328 35096 18380 35148
rect 22376 35232 22428 35284
rect 22560 35232 22612 35284
rect 22836 35232 22888 35284
rect 25504 35232 25556 35284
rect 25780 35275 25832 35284
rect 25780 35241 25789 35275
rect 25789 35241 25823 35275
rect 25823 35241 25832 35275
rect 25780 35232 25832 35241
rect 26976 35232 27028 35284
rect 27804 35232 27856 35284
rect 18144 35028 18196 35080
rect 11152 34960 11204 35012
rect 11612 34960 11664 35012
rect 11980 34960 12032 35012
rect 14740 34960 14792 35012
rect 1860 34892 1912 34944
rect 7564 34935 7616 34944
rect 7564 34901 7573 34935
rect 7573 34901 7607 34935
rect 7607 34901 7616 34935
rect 7564 34892 7616 34901
rect 8484 34892 8536 34944
rect 9864 34935 9916 34944
rect 9864 34901 9873 34935
rect 9873 34901 9907 34935
rect 9907 34901 9916 34935
rect 9864 34892 9916 34901
rect 10140 34892 10192 34944
rect 10968 34892 11020 34944
rect 12992 34892 13044 34944
rect 13084 34892 13136 34944
rect 13728 34892 13780 34944
rect 13820 34892 13872 34944
rect 16396 34960 16448 35012
rect 18972 35028 19024 35080
rect 21916 35071 21968 35080
rect 21916 35037 21925 35071
rect 21925 35037 21959 35071
rect 21959 35037 21968 35071
rect 22744 35096 22796 35148
rect 24308 35096 24360 35148
rect 24492 35096 24544 35148
rect 25504 35096 25556 35148
rect 21916 35028 21968 35037
rect 14924 34892 14976 34944
rect 17868 34892 17920 34944
rect 19616 34960 19668 35012
rect 20996 34960 21048 35012
rect 22652 35028 22704 35080
rect 22928 35071 22980 35080
rect 22928 35037 22937 35071
rect 22937 35037 22971 35071
rect 22971 35037 22980 35071
rect 22928 35028 22980 35037
rect 24032 35028 24084 35080
rect 22376 34960 22428 35012
rect 25412 35028 25464 35080
rect 27988 35164 28040 35216
rect 26608 35096 26660 35148
rect 28172 35139 28224 35148
rect 28172 35105 28181 35139
rect 28181 35105 28215 35139
rect 28215 35105 28224 35139
rect 28172 35096 28224 35105
rect 20904 34892 20956 34944
rect 21272 34935 21324 34944
rect 21272 34901 21281 34935
rect 21281 34901 21315 34935
rect 21315 34901 21324 34935
rect 21272 34892 21324 34901
rect 22836 34892 22888 34944
rect 23388 34892 23440 34944
rect 24952 34892 25004 34944
rect 10214 34790 10266 34842
rect 10278 34790 10330 34842
rect 10342 34790 10394 34842
rect 10406 34790 10458 34842
rect 10470 34790 10522 34842
rect 19478 34790 19530 34842
rect 19542 34790 19594 34842
rect 19606 34790 19658 34842
rect 19670 34790 19722 34842
rect 19734 34790 19786 34842
rect 3240 34688 3292 34740
rect 3792 34688 3844 34740
rect 9036 34688 9088 34740
rect 9496 34731 9548 34740
rect 9496 34697 9505 34731
rect 9505 34697 9539 34731
rect 9539 34697 9548 34731
rect 9496 34688 9548 34697
rect 11244 34688 11296 34740
rect 11980 34688 12032 34740
rect 17960 34688 18012 34740
rect 20168 34688 20220 34740
rect 1860 34663 1912 34672
rect 1860 34629 1869 34663
rect 1869 34629 1903 34663
rect 1903 34629 1912 34663
rect 1860 34620 1912 34629
rect 8760 34620 8812 34672
rect 8392 34595 8444 34604
rect 8392 34561 8401 34595
rect 8401 34561 8435 34595
rect 8435 34561 8444 34595
rect 8392 34552 8444 34561
rect 2780 34527 2832 34536
rect 2780 34493 2789 34527
rect 2789 34493 2823 34527
rect 2823 34493 2832 34527
rect 2780 34484 2832 34493
rect 7472 34416 7524 34468
rect 11888 34620 11940 34672
rect 13084 34620 13136 34672
rect 9588 34552 9640 34604
rect 10048 34552 10100 34604
rect 11060 34552 11112 34604
rect 1400 34348 1452 34400
rect 7564 34391 7616 34400
rect 7564 34357 7573 34391
rect 7573 34357 7607 34391
rect 7607 34357 7616 34391
rect 7564 34348 7616 34357
rect 9588 34348 9640 34400
rect 10600 34348 10652 34400
rect 10876 34459 10928 34468
rect 10876 34425 10885 34459
rect 10885 34425 10919 34459
rect 10919 34425 10928 34459
rect 10876 34416 10928 34425
rect 11428 34416 11480 34468
rect 13912 34552 13964 34604
rect 15936 34595 15988 34604
rect 13360 34527 13412 34536
rect 13360 34493 13369 34527
rect 13369 34493 13403 34527
rect 13403 34493 13412 34527
rect 13360 34484 13412 34493
rect 14556 34484 14608 34536
rect 12900 34391 12952 34400
rect 12900 34357 12909 34391
rect 12909 34357 12943 34391
rect 12943 34357 12952 34391
rect 12900 34348 12952 34357
rect 12992 34348 13044 34400
rect 15476 34416 15528 34468
rect 14648 34348 14700 34400
rect 15936 34561 15945 34595
rect 15945 34561 15979 34595
rect 15979 34561 15988 34595
rect 15936 34552 15988 34561
rect 16120 34620 16172 34672
rect 18696 34620 18748 34672
rect 20812 34688 20864 34740
rect 22744 34688 22796 34740
rect 23664 34688 23716 34740
rect 24952 34731 25004 34740
rect 24952 34697 24961 34731
rect 24961 34697 24995 34731
rect 24995 34697 25004 34731
rect 24952 34688 25004 34697
rect 25504 34688 25556 34740
rect 26792 34688 26844 34740
rect 16488 34552 16540 34604
rect 16672 34595 16724 34604
rect 16672 34561 16681 34595
rect 16681 34561 16715 34595
rect 16715 34561 16724 34595
rect 16672 34552 16724 34561
rect 17500 34595 17552 34604
rect 16580 34484 16632 34536
rect 16212 34416 16264 34468
rect 17500 34561 17509 34595
rect 17509 34561 17543 34595
rect 17543 34561 17552 34595
rect 17500 34552 17552 34561
rect 17776 34552 17828 34604
rect 18328 34595 18380 34604
rect 18328 34561 18337 34595
rect 18337 34561 18371 34595
rect 18371 34561 18380 34595
rect 18328 34552 18380 34561
rect 19984 34552 20036 34604
rect 22928 34620 22980 34672
rect 17224 34416 17276 34468
rect 20168 34484 20220 34536
rect 20444 34484 20496 34536
rect 18512 34348 18564 34400
rect 20076 34416 20128 34468
rect 20628 34595 20680 34604
rect 20628 34561 20663 34595
rect 20663 34561 20680 34595
rect 20628 34552 20680 34561
rect 20996 34552 21048 34604
rect 21548 34552 21600 34604
rect 21824 34552 21876 34604
rect 22008 34552 22060 34604
rect 22836 34595 22888 34604
rect 22836 34561 22845 34595
rect 22845 34561 22879 34595
rect 22879 34561 22888 34595
rect 22836 34552 22888 34561
rect 23572 34552 23624 34604
rect 20904 34484 20956 34536
rect 20996 34416 21048 34468
rect 21180 34416 21232 34468
rect 23112 34484 23164 34536
rect 24308 34484 24360 34536
rect 24492 34552 24544 34604
rect 24768 34595 24820 34604
rect 24768 34561 24777 34595
rect 24777 34561 24811 34595
rect 24811 34561 24820 34595
rect 24768 34552 24820 34561
rect 25596 34595 25648 34604
rect 25596 34561 25605 34595
rect 25605 34561 25639 34595
rect 25639 34561 25648 34595
rect 25596 34552 25648 34561
rect 24860 34484 24912 34536
rect 25504 34527 25556 34536
rect 25504 34493 25513 34527
rect 25513 34493 25547 34527
rect 25547 34493 25556 34527
rect 25504 34484 25556 34493
rect 28080 34595 28132 34604
rect 28080 34561 28089 34595
rect 28089 34561 28123 34595
rect 28123 34561 28132 34595
rect 28080 34552 28132 34561
rect 28264 34552 28316 34604
rect 19892 34348 19944 34400
rect 20536 34348 20588 34400
rect 20628 34348 20680 34400
rect 22008 34348 22060 34400
rect 22560 34391 22612 34400
rect 22560 34357 22569 34391
rect 22569 34357 22603 34391
rect 22603 34357 22612 34391
rect 22560 34348 22612 34357
rect 23112 34348 23164 34400
rect 24216 34416 24268 34468
rect 26240 34416 26292 34468
rect 27160 34416 27212 34468
rect 27344 34459 27396 34468
rect 27344 34425 27353 34459
rect 27353 34425 27387 34459
rect 27387 34425 27396 34459
rect 27344 34416 27396 34425
rect 24492 34348 24544 34400
rect 24860 34348 24912 34400
rect 25136 34348 25188 34400
rect 28448 34484 28500 34536
rect 5582 34246 5634 34298
rect 5646 34246 5698 34298
rect 5710 34246 5762 34298
rect 5774 34246 5826 34298
rect 5838 34246 5890 34298
rect 14846 34246 14898 34298
rect 14910 34246 14962 34298
rect 14974 34246 15026 34298
rect 15038 34246 15090 34298
rect 15102 34246 15154 34298
rect 24110 34246 24162 34298
rect 24174 34246 24226 34298
rect 24238 34246 24290 34298
rect 24302 34246 24354 34298
rect 24366 34246 24418 34298
rect 7748 34144 7800 34196
rect 1400 34051 1452 34060
rect 1400 34017 1409 34051
rect 1409 34017 1443 34051
rect 1443 34017 1452 34051
rect 1400 34008 1452 34017
rect 2780 34051 2832 34060
rect 2780 34017 2789 34051
rect 2789 34017 2823 34051
rect 2823 34017 2832 34051
rect 8852 34076 8904 34128
rect 9404 34076 9456 34128
rect 2780 34008 2832 34017
rect 9956 34008 10008 34060
rect 7656 33940 7708 33992
rect 7748 33983 7800 33992
rect 7748 33949 7757 33983
rect 7757 33949 7791 33983
rect 7791 33949 7800 33983
rect 7748 33940 7800 33949
rect 8484 33940 8536 33992
rect 9312 33940 9364 33992
rect 9404 33940 9456 33992
rect 2228 33872 2280 33924
rect 9496 33872 9548 33924
rect 10048 33940 10100 33992
rect 10232 34076 10284 34128
rect 10968 34076 11020 34128
rect 12716 34144 12768 34196
rect 10232 33940 10284 33992
rect 10416 33940 10468 33992
rect 10784 34008 10836 34060
rect 11704 34076 11756 34128
rect 11888 34076 11940 34128
rect 12900 34144 12952 34196
rect 14188 34144 14240 34196
rect 14464 34144 14516 34196
rect 15936 34144 15988 34196
rect 16488 34144 16540 34196
rect 16580 34144 16632 34196
rect 17500 34144 17552 34196
rect 18604 34144 18656 34196
rect 19984 34144 20036 34196
rect 20168 34144 20220 34196
rect 20628 34144 20680 34196
rect 21548 34144 21600 34196
rect 21916 34144 21968 34196
rect 23664 34144 23716 34196
rect 12072 34008 12124 34060
rect 12440 34008 12492 34060
rect 13912 34076 13964 34128
rect 14096 34076 14148 34128
rect 17224 34076 17276 34128
rect 18052 34076 18104 34128
rect 21088 34076 21140 34128
rect 22468 34119 22520 34128
rect 22468 34085 22477 34119
rect 22477 34085 22511 34119
rect 22511 34085 22520 34119
rect 22468 34076 22520 34085
rect 23296 34119 23348 34128
rect 12992 34008 13044 34060
rect 11152 33940 11204 33992
rect 11980 33983 12032 33992
rect 9956 33872 10008 33924
rect 11980 33949 11989 33983
rect 11989 33949 12023 33983
rect 12023 33949 12032 33983
rect 11980 33940 12032 33949
rect 12164 33983 12216 33992
rect 12164 33949 12173 33983
rect 12173 33949 12207 33983
rect 12207 33949 12216 33983
rect 12164 33940 12216 33949
rect 12532 33940 12584 33992
rect 12808 33872 12860 33924
rect 7564 33847 7616 33856
rect 7564 33813 7573 33847
rect 7573 33813 7607 33847
rect 7607 33813 7616 33847
rect 7564 33804 7616 33813
rect 13912 33940 13964 33992
rect 14188 33940 14240 33992
rect 14372 33940 14424 33992
rect 14648 33983 14700 33992
rect 14648 33949 14657 33983
rect 14657 33949 14691 33983
rect 14691 33949 14700 33983
rect 14648 33940 14700 33949
rect 14280 33804 14332 33856
rect 14924 33940 14976 33992
rect 14832 33872 14884 33924
rect 18328 34008 18380 34060
rect 19248 34051 19300 34060
rect 19248 34017 19257 34051
rect 19257 34017 19291 34051
rect 19291 34017 19300 34051
rect 19248 34008 19300 34017
rect 15660 33940 15712 33992
rect 16948 33940 17000 33992
rect 15200 33804 15252 33856
rect 17132 33872 17184 33924
rect 20628 33940 20680 33992
rect 21824 34008 21876 34060
rect 23296 34085 23305 34119
rect 23305 34085 23339 34119
rect 23339 34085 23348 34119
rect 23296 34076 23348 34085
rect 23756 34076 23808 34128
rect 23388 34051 23440 34060
rect 23388 34017 23397 34051
rect 23397 34017 23431 34051
rect 23431 34017 23440 34051
rect 23388 34008 23440 34017
rect 23940 34008 23992 34060
rect 24124 34008 24176 34060
rect 26240 34076 26292 34128
rect 25688 34051 25740 34060
rect 25688 34017 25697 34051
rect 25697 34017 25731 34051
rect 25731 34017 25740 34051
rect 25688 34008 25740 34017
rect 26332 34051 26384 34060
rect 26332 34017 26341 34051
rect 26341 34017 26375 34051
rect 26375 34017 26384 34051
rect 26332 34008 26384 34017
rect 28908 34008 28960 34060
rect 22192 33940 22244 33992
rect 22744 33940 22796 33992
rect 25044 33940 25096 33992
rect 18236 33872 18288 33924
rect 18972 33872 19024 33924
rect 19340 33872 19392 33924
rect 18144 33804 18196 33856
rect 18420 33847 18472 33856
rect 18420 33813 18429 33847
rect 18429 33813 18463 33847
rect 18463 33813 18472 33847
rect 18420 33804 18472 33813
rect 18512 33847 18564 33856
rect 18512 33813 18521 33847
rect 18521 33813 18555 33847
rect 18555 33813 18564 33847
rect 18512 33804 18564 33813
rect 18788 33804 18840 33856
rect 20168 33804 20220 33856
rect 20812 33804 20864 33856
rect 24492 33872 24544 33924
rect 26516 33915 26568 33924
rect 22928 33847 22980 33856
rect 22928 33813 22937 33847
rect 22937 33813 22971 33847
rect 22971 33813 22980 33847
rect 22928 33804 22980 33813
rect 23112 33804 23164 33856
rect 26516 33881 26525 33915
rect 26525 33881 26559 33915
rect 26559 33881 26568 33915
rect 26516 33872 26568 33881
rect 25228 33847 25280 33856
rect 25228 33813 25237 33847
rect 25237 33813 25271 33847
rect 25271 33813 25280 33847
rect 25228 33804 25280 33813
rect 10214 33702 10266 33754
rect 10278 33702 10330 33754
rect 10342 33702 10394 33754
rect 10406 33702 10458 33754
rect 10470 33702 10522 33754
rect 19478 33702 19530 33754
rect 19542 33702 19594 33754
rect 19606 33702 19658 33754
rect 19670 33702 19722 33754
rect 19734 33702 19786 33754
rect 2044 33600 2096 33652
rect 2228 33643 2280 33652
rect 2228 33609 2237 33643
rect 2237 33609 2271 33643
rect 2271 33609 2280 33643
rect 2228 33600 2280 33609
rect 9956 33600 10008 33652
rect 11428 33600 11480 33652
rect 11888 33600 11940 33652
rect 12072 33600 12124 33652
rect 15568 33600 15620 33652
rect 18420 33600 18472 33652
rect 20168 33600 20220 33652
rect 21088 33600 21140 33652
rect 25964 33600 26016 33652
rect 1400 33507 1452 33516
rect 1400 33473 1409 33507
rect 1409 33473 1443 33507
rect 1443 33473 1452 33507
rect 1400 33464 1452 33473
rect 1952 33464 2004 33516
rect 7840 33464 7892 33516
rect 8484 33464 8536 33516
rect 9404 33464 9456 33516
rect 9588 33464 9640 33516
rect 10048 33464 10100 33516
rect 12992 33532 13044 33584
rect 18052 33532 18104 33584
rect 18604 33532 18656 33584
rect 10600 33464 10652 33516
rect 10876 33464 10928 33516
rect 11060 33464 11112 33516
rect 11888 33464 11940 33516
rect 12164 33507 12216 33516
rect 12164 33473 12173 33507
rect 12173 33473 12207 33507
rect 12207 33473 12216 33507
rect 12164 33464 12216 33473
rect 12624 33464 12676 33516
rect 13360 33464 13412 33516
rect 10416 33396 10468 33448
rect 10508 33328 10560 33380
rect 10600 33328 10652 33380
rect 12440 33396 12492 33448
rect 12716 33396 12768 33448
rect 12900 33439 12952 33448
rect 12900 33405 12909 33439
rect 12909 33405 12943 33439
rect 12943 33405 12952 33439
rect 12900 33396 12952 33405
rect 12992 33396 13044 33448
rect 14004 33464 14056 33516
rect 15200 33464 15252 33516
rect 15660 33464 15712 33516
rect 19432 33532 19484 33584
rect 19892 33532 19944 33584
rect 23296 33532 23348 33584
rect 14464 33396 14516 33448
rect 10048 33260 10100 33312
rect 13360 33328 13412 33380
rect 14832 33371 14884 33380
rect 14832 33337 14841 33371
rect 14841 33337 14875 33371
rect 14875 33337 14884 33371
rect 14832 33328 14884 33337
rect 15108 33396 15160 33448
rect 19156 33507 19208 33516
rect 19156 33473 19165 33507
rect 19165 33473 19199 33507
rect 19199 33473 19208 33507
rect 19156 33464 19208 33473
rect 19340 33464 19392 33516
rect 19616 33464 19668 33516
rect 22008 33464 22060 33516
rect 22192 33507 22244 33516
rect 22192 33473 22201 33507
rect 22201 33473 22235 33507
rect 22235 33473 22244 33507
rect 22192 33464 22244 33473
rect 22468 33507 22520 33516
rect 22468 33473 22477 33507
rect 22477 33473 22511 33507
rect 22511 33473 22520 33507
rect 23644 33507 23696 33516
rect 22468 33464 22520 33473
rect 23644 33473 23653 33507
rect 23653 33473 23687 33507
rect 23687 33473 23696 33507
rect 23644 33464 23696 33473
rect 24768 33532 24820 33584
rect 27620 33532 27672 33584
rect 23848 33510 23900 33516
rect 23848 33476 23857 33510
rect 23857 33476 23891 33510
rect 23891 33476 23900 33510
rect 23848 33464 23900 33476
rect 15476 33328 15528 33380
rect 16304 33328 16356 33380
rect 18604 33371 18656 33380
rect 18604 33337 18613 33371
rect 18613 33337 18647 33371
rect 18647 33337 18656 33371
rect 18604 33328 18656 33337
rect 11244 33260 11296 33312
rect 14740 33260 14792 33312
rect 15200 33260 15252 33312
rect 22560 33396 22612 33448
rect 22836 33396 22888 33448
rect 26976 33464 27028 33516
rect 19800 33328 19852 33380
rect 24124 33396 24176 33448
rect 24952 33396 25004 33448
rect 25320 33396 25372 33448
rect 26148 33439 26200 33448
rect 26148 33405 26157 33439
rect 26157 33405 26191 33439
rect 26191 33405 26200 33439
rect 26148 33396 26200 33405
rect 27712 33396 27764 33448
rect 19432 33260 19484 33312
rect 21824 33303 21876 33312
rect 21824 33269 21833 33303
rect 21833 33269 21867 33303
rect 21867 33269 21876 33303
rect 21824 33260 21876 33269
rect 22008 33260 22060 33312
rect 22652 33260 22704 33312
rect 23756 33260 23808 33312
rect 27252 33260 27304 33312
rect 27712 33260 27764 33312
rect 28172 33464 28224 33516
rect 5582 33158 5634 33210
rect 5646 33158 5698 33210
rect 5710 33158 5762 33210
rect 5774 33158 5826 33210
rect 5838 33158 5890 33210
rect 14846 33158 14898 33210
rect 14910 33158 14962 33210
rect 14974 33158 15026 33210
rect 15038 33158 15090 33210
rect 15102 33158 15154 33210
rect 24110 33158 24162 33210
rect 24174 33158 24226 33210
rect 24238 33158 24290 33210
rect 24302 33158 24354 33210
rect 24366 33158 24418 33210
rect 3424 33056 3476 33108
rect 10600 33056 10652 33108
rect 10692 33056 10744 33108
rect 11612 33056 11664 33108
rect 12072 33056 12124 33108
rect 9036 32988 9088 33040
rect 9496 32988 9548 33040
rect 10784 32988 10836 33040
rect 11980 32988 12032 33040
rect 13268 33056 13320 33108
rect 13360 33056 13412 33108
rect 13084 32988 13136 33040
rect 18052 33056 18104 33108
rect 18236 33099 18288 33108
rect 18236 33065 18245 33099
rect 18245 33065 18279 33099
rect 18279 33065 18288 33099
rect 18236 33056 18288 33065
rect 1492 32852 1544 32904
rect 7840 32852 7892 32904
rect 8944 32852 8996 32904
rect 10876 32920 10928 32972
rect 12072 32920 12124 32972
rect 14188 32920 14240 32972
rect 8760 32784 8812 32836
rect 9772 32852 9824 32904
rect 9864 32852 9916 32904
rect 10140 32852 10192 32904
rect 10324 32895 10376 32904
rect 10324 32861 10333 32895
rect 10333 32861 10367 32895
rect 10367 32861 10376 32895
rect 10324 32852 10376 32861
rect 10600 32852 10652 32904
rect 11520 32852 11572 32904
rect 9496 32716 9548 32768
rect 11336 32784 11388 32836
rect 11704 32784 11756 32836
rect 12440 32784 12492 32836
rect 12624 32852 12676 32904
rect 12808 32827 12860 32836
rect 12808 32793 12817 32827
rect 12817 32793 12851 32827
rect 12851 32793 12860 32827
rect 12808 32784 12860 32793
rect 13084 32895 13136 32904
rect 13084 32861 13093 32895
rect 13093 32861 13127 32895
rect 13127 32861 13136 32895
rect 14832 32920 14884 32972
rect 13084 32852 13136 32861
rect 15384 32852 15436 32904
rect 15660 32963 15712 32972
rect 15660 32929 15669 32963
rect 15669 32929 15703 32963
rect 15703 32929 15712 32963
rect 15660 32920 15712 32929
rect 21088 32988 21140 33040
rect 22652 33031 22704 33040
rect 22652 32997 22661 33031
rect 22661 32997 22695 33031
rect 22695 32997 22704 33031
rect 22652 32988 22704 32997
rect 19616 32920 19668 32972
rect 23940 33056 23992 33108
rect 17500 32895 17552 32904
rect 17500 32861 17509 32895
rect 17509 32861 17543 32895
rect 17543 32861 17552 32895
rect 17500 32852 17552 32861
rect 18236 32895 18288 32904
rect 18236 32861 18245 32895
rect 18245 32861 18279 32895
rect 18279 32861 18288 32895
rect 18420 32895 18472 32904
rect 18236 32852 18288 32861
rect 18420 32861 18429 32895
rect 18429 32861 18463 32895
rect 18463 32861 18472 32895
rect 18420 32852 18472 32861
rect 18604 32852 18656 32904
rect 19248 32895 19300 32904
rect 19248 32861 19257 32895
rect 19257 32861 19291 32895
rect 19291 32861 19300 32895
rect 19248 32852 19300 32861
rect 19432 32895 19484 32904
rect 19432 32861 19441 32895
rect 19441 32861 19475 32895
rect 19475 32861 19484 32895
rect 19432 32852 19484 32861
rect 19708 32852 19760 32904
rect 19800 32852 19852 32904
rect 20628 32852 20680 32904
rect 21272 32895 21324 32904
rect 21272 32861 21281 32895
rect 21281 32861 21315 32895
rect 21315 32861 21324 32895
rect 21272 32852 21324 32861
rect 21824 32852 21876 32904
rect 21916 32852 21968 32904
rect 24676 32920 24728 32972
rect 23480 32852 23532 32904
rect 27436 33056 27488 33108
rect 25044 32920 25096 32972
rect 25412 32920 25464 32972
rect 25780 32920 25832 32972
rect 28356 32988 28408 33040
rect 26332 32963 26384 32972
rect 26332 32929 26341 32963
rect 26341 32929 26375 32963
rect 26375 32929 26384 32963
rect 26332 32920 26384 32929
rect 28172 32963 28224 32972
rect 28172 32929 28181 32963
rect 28181 32929 28215 32963
rect 28215 32929 28224 32963
rect 28172 32920 28224 32929
rect 25320 32852 25372 32904
rect 25504 32852 25556 32904
rect 13452 32784 13504 32836
rect 13544 32784 13596 32836
rect 14372 32827 14424 32836
rect 12716 32716 12768 32768
rect 13176 32759 13228 32768
rect 13176 32725 13185 32759
rect 13185 32725 13219 32759
rect 13219 32725 13228 32759
rect 13176 32716 13228 32725
rect 14096 32759 14148 32768
rect 14096 32725 14105 32759
rect 14105 32725 14139 32759
rect 14139 32725 14148 32759
rect 14096 32716 14148 32725
rect 14372 32793 14381 32827
rect 14381 32793 14415 32827
rect 14415 32793 14424 32827
rect 14372 32784 14424 32793
rect 14556 32827 14608 32836
rect 14556 32793 14591 32827
rect 14591 32793 14608 32827
rect 14556 32784 14608 32793
rect 14740 32784 14792 32836
rect 16304 32716 16356 32768
rect 17132 32716 17184 32768
rect 18236 32716 18288 32768
rect 18512 32716 18564 32768
rect 18696 32759 18748 32768
rect 18696 32725 18705 32759
rect 18705 32725 18739 32759
rect 18739 32725 18748 32759
rect 18696 32716 18748 32725
rect 19340 32716 19392 32768
rect 19892 32759 19944 32768
rect 19892 32725 19901 32759
rect 19901 32725 19935 32759
rect 19935 32725 19944 32759
rect 19892 32716 19944 32725
rect 20352 32784 20404 32836
rect 21088 32784 21140 32836
rect 24584 32716 24636 32768
rect 24952 32716 25004 32768
rect 10214 32614 10266 32666
rect 10278 32614 10330 32666
rect 10342 32614 10394 32666
rect 10406 32614 10458 32666
rect 10470 32614 10522 32666
rect 19478 32614 19530 32666
rect 19542 32614 19594 32666
rect 19606 32614 19658 32666
rect 19670 32614 19722 32666
rect 19734 32614 19786 32666
rect 9496 32444 9548 32496
rect 8116 32419 8168 32428
rect 8116 32385 8125 32419
rect 8125 32385 8159 32419
rect 8159 32385 8168 32419
rect 8116 32376 8168 32385
rect 8760 32419 8812 32428
rect 1492 32351 1544 32360
rect 1492 32317 1501 32351
rect 1501 32317 1535 32351
rect 1535 32317 1544 32351
rect 1492 32308 1544 32317
rect 1768 32308 1820 32360
rect 2872 32351 2924 32360
rect 2872 32317 2881 32351
rect 2881 32317 2915 32351
rect 2915 32317 2924 32351
rect 2872 32308 2924 32317
rect 8760 32385 8769 32419
rect 8769 32385 8803 32419
rect 8803 32385 8812 32419
rect 8760 32376 8812 32385
rect 9864 32444 9916 32496
rect 10048 32444 10100 32496
rect 10324 32444 10376 32496
rect 12900 32512 12952 32564
rect 13360 32512 13412 32564
rect 8668 32283 8720 32292
rect 8668 32249 8677 32283
rect 8677 32249 8711 32283
rect 8711 32249 8720 32283
rect 8668 32240 8720 32249
rect 9680 32240 9732 32292
rect 10416 32308 10468 32360
rect 10692 32376 10744 32428
rect 10784 32419 10836 32428
rect 10784 32385 10793 32419
rect 10793 32385 10827 32419
rect 10827 32385 10836 32419
rect 12164 32444 12216 32496
rect 12808 32444 12860 32496
rect 10784 32376 10836 32385
rect 11152 32308 11204 32360
rect 10324 32240 10376 32292
rect 13176 32376 13228 32428
rect 13728 32444 13780 32496
rect 14188 32444 14240 32496
rect 14372 32444 14424 32496
rect 13820 32376 13872 32428
rect 11520 32351 11572 32360
rect 11520 32317 11529 32351
rect 11529 32317 11563 32351
rect 11563 32317 11572 32351
rect 11520 32308 11572 32317
rect 13084 32308 13136 32360
rect 17224 32444 17276 32496
rect 17500 32444 17552 32496
rect 18696 32444 18748 32496
rect 20720 32444 20772 32496
rect 21640 32444 21692 32496
rect 16580 32376 16632 32428
rect 16948 32419 17000 32428
rect 16948 32385 16957 32419
rect 16957 32385 16991 32419
rect 16991 32385 17000 32419
rect 16948 32376 17000 32385
rect 17132 32419 17184 32428
rect 17132 32385 17141 32419
rect 17141 32385 17175 32419
rect 17175 32385 17184 32419
rect 17132 32376 17184 32385
rect 18236 32419 18288 32428
rect 18236 32385 18245 32419
rect 18245 32385 18279 32419
rect 18279 32385 18288 32419
rect 18236 32376 18288 32385
rect 19984 32376 20036 32428
rect 20628 32419 20680 32428
rect 20628 32385 20637 32419
rect 20637 32385 20671 32419
rect 20671 32385 20680 32419
rect 20628 32376 20680 32385
rect 21272 32376 21324 32428
rect 21916 32376 21968 32428
rect 22928 32376 22980 32428
rect 23756 32376 23808 32428
rect 24676 32376 24728 32428
rect 25320 32376 25372 32428
rect 27344 32444 27396 32496
rect 27160 32419 27212 32428
rect 27160 32385 27169 32419
rect 27169 32385 27203 32419
rect 27203 32385 27212 32419
rect 27160 32376 27212 32385
rect 27988 32419 28040 32428
rect 27988 32385 27997 32419
rect 27997 32385 28031 32419
rect 28031 32385 28040 32419
rect 27988 32376 28040 32385
rect 12532 32240 12584 32292
rect 19248 32308 19300 32360
rect 25228 32308 25280 32360
rect 25596 32351 25648 32360
rect 25596 32317 25605 32351
rect 25605 32317 25639 32351
rect 25639 32317 25648 32351
rect 25596 32308 25648 32317
rect 27252 32351 27304 32360
rect 27252 32317 27261 32351
rect 27261 32317 27295 32351
rect 27295 32317 27304 32351
rect 27252 32308 27304 32317
rect 13728 32240 13780 32292
rect 14280 32240 14332 32292
rect 9128 32172 9180 32224
rect 9312 32172 9364 32224
rect 11060 32172 11112 32224
rect 12716 32172 12768 32224
rect 12808 32172 12860 32224
rect 13452 32215 13504 32224
rect 13452 32181 13461 32215
rect 13461 32181 13495 32215
rect 13495 32181 13504 32215
rect 13452 32172 13504 32181
rect 13820 32215 13872 32224
rect 13820 32181 13829 32215
rect 13829 32181 13863 32215
rect 13863 32181 13872 32215
rect 13820 32172 13872 32181
rect 14004 32172 14056 32224
rect 16212 32240 16264 32292
rect 15292 32172 15344 32224
rect 15936 32172 15988 32224
rect 17040 32172 17092 32224
rect 19984 32172 20036 32224
rect 23480 32240 23532 32292
rect 24676 32240 24728 32292
rect 24860 32240 24912 32292
rect 25136 32240 25188 32292
rect 24952 32172 25004 32224
rect 25964 32215 26016 32224
rect 25964 32181 25973 32215
rect 25973 32181 26007 32215
rect 26007 32181 26016 32215
rect 25964 32172 26016 32181
rect 26056 32172 26108 32224
rect 27528 32172 27580 32224
rect 5582 32070 5634 32122
rect 5646 32070 5698 32122
rect 5710 32070 5762 32122
rect 5774 32070 5826 32122
rect 5838 32070 5890 32122
rect 14846 32070 14898 32122
rect 14910 32070 14962 32122
rect 14974 32070 15026 32122
rect 15038 32070 15090 32122
rect 15102 32070 15154 32122
rect 24110 32070 24162 32122
rect 24174 32070 24226 32122
rect 24238 32070 24290 32122
rect 24302 32070 24354 32122
rect 24366 32070 24418 32122
rect 1492 31968 1544 32020
rect 10232 31968 10284 32020
rect 10324 31968 10376 32020
rect 10968 31968 11020 32020
rect 11520 31968 11572 32020
rect 13820 31968 13872 32020
rect 1676 31764 1728 31816
rect 6276 31807 6328 31816
rect 6276 31773 6285 31807
rect 6285 31773 6319 31807
rect 6319 31773 6328 31807
rect 6276 31764 6328 31773
rect 9404 31900 9456 31952
rect 11704 31900 11756 31952
rect 12716 31900 12768 31952
rect 13544 31900 13596 31952
rect 9312 31832 9364 31884
rect 7932 31764 7984 31816
rect 9404 31807 9456 31816
rect 9404 31773 9413 31807
rect 9413 31773 9447 31807
rect 9447 31773 9456 31807
rect 9404 31764 9456 31773
rect 9588 31764 9640 31816
rect 10140 31764 10192 31816
rect 10324 31764 10376 31816
rect 2228 31696 2280 31748
rect 6736 31671 6788 31680
rect 6736 31637 6745 31671
rect 6745 31637 6779 31671
rect 6779 31637 6788 31671
rect 6736 31628 6788 31637
rect 9128 31696 9180 31748
rect 9312 31696 9364 31748
rect 9956 31696 10008 31748
rect 10048 31696 10100 31748
rect 10784 31696 10836 31748
rect 11520 31764 11572 31816
rect 11704 31807 11756 31816
rect 11704 31773 11713 31807
rect 11713 31773 11747 31807
rect 11747 31773 11756 31807
rect 11704 31764 11756 31773
rect 13728 31832 13780 31884
rect 12900 31764 12952 31816
rect 14096 31900 14148 31952
rect 15200 31968 15252 32020
rect 18604 31968 18656 32020
rect 19708 31968 19760 32020
rect 20260 31968 20312 32020
rect 20444 31968 20496 32020
rect 23112 31968 23164 32020
rect 23480 32011 23532 32020
rect 23480 31977 23489 32011
rect 23489 31977 23523 32011
rect 23523 31977 23532 32011
rect 23480 31968 23532 31977
rect 25964 31968 26016 32020
rect 14096 31807 14148 31816
rect 14096 31773 14105 31807
rect 14105 31773 14139 31807
rect 14139 31773 14148 31807
rect 14096 31764 14148 31773
rect 15660 31832 15712 31884
rect 17316 31832 17368 31884
rect 19524 31832 19576 31884
rect 19892 31832 19944 31884
rect 14740 31764 14792 31816
rect 8392 31628 8444 31680
rect 9680 31628 9732 31680
rect 11152 31628 11204 31680
rect 14556 31696 14608 31748
rect 14832 31696 14884 31748
rect 16488 31739 16540 31748
rect 16488 31705 16522 31739
rect 16522 31705 16540 31739
rect 17500 31764 17552 31816
rect 19708 31764 19760 31816
rect 20076 31807 20128 31816
rect 20076 31773 20085 31807
rect 20085 31773 20119 31807
rect 20119 31773 20128 31807
rect 20076 31764 20128 31773
rect 20260 31832 20312 31884
rect 26332 31875 26384 31884
rect 20812 31807 20864 31816
rect 20812 31773 20821 31807
rect 20821 31773 20855 31807
rect 20855 31773 20864 31807
rect 20812 31764 20864 31773
rect 22560 31764 22612 31816
rect 23112 31764 23164 31816
rect 23388 31807 23440 31816
rect 23388 31773 23397 31807
rect 23397 31773 23431 31807
rect 23431 31773 23440 31807
rect 23388 31764 23440 31773
rect 16488 31696 16540 31705
rect 17408 31696 17460 31748
rect 18236 31696 18288 31748
rect 12348 31628 12400 31680
rect 13176 31628 13228 31680
rect 13912 31628 13964 31680
rect 16304 31628 16356 31680
rect 16764 31628 16816 31680
rect 17224 31628 17276 31680
rect 18512 31671 18564 31680
rect 18512 31637 18537 31671
rect 18537 31637 18564 31671
rect 18696 31671 18748 31680
rect 18512 31628 18564 31637
rect 18696 31637 18705 31671
rect 18705 31637 18739 31671
rect 18739 31637 18748 31671
rect 18696 31628 18748 31637
rect 19340 31696 19392 31748
rect 19984 31739 20036 31748
rect 19984 31705 19993 31739
rect 19993 31705 20027 31739
rect 20027 31705 20036 31739
rect 19984 31696 20036 31705
rect 20996 31696 21048 31748
rect 21916 31696 21968 31748
rect 20352 31628 20404 31680
rect 20812 31628 20864 31680
rect 22928 31696 22980 31748
rect 23480 31696 23532 31748
rect 26332 31841 26341 31875
rect 26341 31841 26375 31875
rect 26375 31841 26384 31875
rect 26332 31832 26384 31841
rect 28172 31875 28224 31884
rect 28172 31841 28181 31875
rect 28181 31841 28215 31875
rect 28215 31841 28224 31875
rect 28172 31832 28224 31841
rect 24492 31807 24544 31816
rect 24492 31773 24501 31807
rect 24501 31773 24535 31807
rect 24535 31773 24544 31807
rect 24492 31764 24544 31773
rect 24584 31764 24636 31816
rect 23848 31671 23900 31680
rect 23848 31637 23857 31671
rect 23857 31637 23891 31671
rect 23891 31637 23900 31671
rect 23848 31628 23900 31637
rect 24860 31628 24912 31680
rect 25320 31628 25372 31680
rect 10214 31526 10266 31578
rect 10278 31526 10330 31578
rect 10342 31526 10394 31578
rect 10406 31526 10458 31578
rect 10470 31526 10522 31578
rect 19478 31526 19530 31578
rect 19542 31526 19594 31578
rect 19606 31526 19658 31578
rect 19670 31526 19722 31578
rect 19734 31526 19786 31578
rect 9956 31424 10008 31476
rect 10048 31424 10100 31476
rect 14464 31424 14516 31476
rect 1676 31331 1728 31340
rect 1676 31297 1685 31331
rect 1685 31297 1719 31331
rect 1719 31297 1728 31331
rect 1676 31288 1728 31297
rect 9680 31356 9732 31408
rect 2320 31220 2372 31272
rect 2780 31263 2832 31272
rect 2780 31229 2789 31263
rect 2789 31229 2823 31263
rect 2823 31229 2832 31263
rect 8300 31288 8352 31340
rect 8944 31288 8996 31340
rect 9128 31331 9180 31340
rect 9128 31297 9137 31331
rect 9137 31297 9171 31331
rect 9171 31297 9180 31331
rect 9128 31288 9180 31297
rect 10232 31356 10284 31408
rect 12256 31356 12308 31408
rect 12348 31356 12400 31408
rect 2780 31220 2832 31229
rect 8208 31220 8260 31272
rect 8116 31152 8168 31204
rect 9588 31220 9640 31272
rect 10692 31288 10744 31340
rect 10968 31288 11020 31340
rect 11704 31288 11756 31340
rect 12072 31288 12124 31340
rect 13176 31288 13228 31340
rect 13452 31331 13504 31340
rect 13452 31297 13461 31331
rect 13461 31297 13495 31331
rect 13495 31297 13504 31331
rect 13452 31288 13504 31297
rect 13728 31356 13780 31408
rect 15200 31424 15252 31476
rect 14372 31288 14424 31340
rect 14740 31331 14792 31340
rect 14740 31297 14749 31331
rect 14749 31297 14783 31331
rect 14783 31297 14792 31331
rect 14740 31288 14792 31297
rect 10048 31220 10100 31272
rect 10416 31220 10468 31272
rect 12164 31220 12216 31272
rect 12808 31220 12860 31272
rect 10324 31152 10376 31204
rect 10508 31152 10560 31204
rect 13912 31263 13964 31272
rect 13912 31229 13921 31263
rect 13921 31229 13955 31263
rect 13955 31229 13964 31263
rect 13912 31220 13964 31229
rect 14188 31220 14240 31272
rect 14464 31220 14516 31272
rect 15844 31288 15896 31340
rect 16580 31356 16632 31408
rect 20076 31424 20128 31476
rect 22284 31424 22336 31476
rect 16488 31288 16540 31340
rect 22928 31356 22980 31408
rect 17132 31288 17184 31340
rect 23204 31356 23256 31408
rect 23112 31331 23164 31340
rect 23112 31297 23121 31331
rect 23121 31297 23155 31331
rect 23155 31297 23164 31331
rect 23756 31424 23808 31476
rect 23848 31356 23900 31408
rect 24860 31424 24912 31476
rect 25504 31424 25556 31476
rect 26424 31467 26476 31476
rect 26424 31433 26433 31467
rect 26433 31433 26467 31467
rect 26467 31433 26476 31467
rect 26424 31424 26476 31433
rect 27160 31424 27212 31476
rect 27344 31467 27396 31476
rect 27344 31433 27353 31467
rect 27353 31433 27387 31467
rect 27387 31433 27396 31467
rect 27344 31424 27396 31433
rect 28080 31467 28132 31476
rect 28080 31433 28089 31467
rect 28089 31433 28123 31467
rect 28123 31433 28132 31467
rect 28080 31424 28132 31433
rect 23388 31331 23440 31340
rect 23112 31288 23164 31297
rect 23388 31297 23397 31331
rect 23397 31297 23431 31331
rect 23431 31297 23440 31331
rect 23388 31288 23440 31297
rect 24032 31331 24084 31340
rect 24032 31297 24041 31331
rect 24041 31297 24075 31331
rect 24075 31297 24084 31331
rect 24032 31288 24084 31297
rect 24952 31356 25004 31408
rect 24492 31288 24544 31340
rect 16764 31263 16816 31272
rect 16764 31229 16773 31263
rect 16773 31229 16807 31263
rect 16807 31229 16816 31263
rect 16764 31220 16816 31229
rect 17684 31263 17736 31272
rect 17684 31229 17693 31263
rect 17693 31229 17727 31263
rect 17727 31229 17736 31263
rect 17684 31220 17736 31229
rect 19892 31263 19944 31272
rect 19892 31229 19901 31263
rect 19901 31229 19935 31263
rect 19935 31229 19944 31263
rect 19892 31220 19944 31229
rect 24676 31220 24728 31272
rect 25412 31356 25464 31408
rect 25320 31331 25372 31340
rect 25320 31297 25354 31331
rect 25354 31297 25372 31331
rect 25320 31288 25372 31297
rect 25596 31288 25648 31340
rect 26148 31288 26200 31340
rect 27620 31288 27672 31340
rect 28264 31288 28316 31340
rect 8576 31127 8628 31136
rect 8576 31093 8585 31127
rect 8585 31093 8619 31127
rect 8619 31093 8628 31127
rect 8576 31084 8628 31093
rect 8668 31084 8720 31136
rect 10232 31084 10284 31136
rect 10416 31084 10468 31136
rect 11336 31084 11388 31136
rect 11980 31084 12032 31136
rect 12624 31127 12676 31136
rect 12624 31093 12633 31127
rect 12633 31093 12667 31127
rect 12667 31093 12676 31127
rect 12624 31084 12676 31093
rect 16028 31084 16080 31136
rect 16856 31127 16908 31136
rect 16856 31093 16865 31127
rect 16865 31093 16899 31127
rect 16899 31093 16908 31127
rect 16856 31084 16908 31093
rect 16948 31084 17000 31136
rect 19064 31127 19116 31136
rect 19064 31093 19073 31127
rect 19073 31093 19107 31127
rect 19107 31093 19116 31127
rect 19064 31084 19116 31093
rect 21088 31152 21140 31204
rect 21916 31152 21968 31204
rect 20260 31084 20312 31136
rect 20628 31084 20680 31136
rect 21364 31084 21416 31136
rect 22376 31127 22428 31136
rect 22376 31093 22385 31127
rect 22385 31093 22419 31127
rect 22419 31093 22428 31127
rect 22376 31084 22428 31093
rect 22836 31127 22888 31136
rect 22836 31093 22845 31127
rect 22845 31093 22879 31127
rect 22879 31093 22888 31127
rect 22836 31084 22888 31093
rect 23940 31152 23992 31204
rect 23480 31084 23532 31136
rect 25228 31084 25280 31136
rect 25780 31084 25832 31136
rect 5582 30982 5634 31034
rect 5646 30982 5698 31034
rect 5710 30982 5762 31034
rect 5774 30982 5826 31034
rect 5838 30982 5890 31034
rect 14846 30982 14898 31034
rect 14910 30982 14962 31034
rect 14974 30982 15026 31034
rect 15038 30982 15090 31034
rect 15102 30982 15154 31034
rect 24110 30982 24162 31034
rect 24174 30982 24226 31034
rect 24238 30982 24290 31034
rect 24302 30982 24354 31034
rect 24366 30982 24418 31034
rect 2320 30923 2372 30932
rect 2320 30889 2329 30923
rect 2329 30889 2363 30923
rect 2363 30889 2372 30923
rect 2320 30880 2372 30889
rect 7012 30880 7064 30932
rect 11612 30880 11664 30932
rect 11980 30880 12032 30932
rect 12624 30880 12676 30932
rect 12716 30880 12768 30932
rect 15384 30880 15436 30932
rect 17224 30880 17276 30932
rect 19984 30923 20036 30932
rect 19984 30889 19993 30923
rect 19993 30889 20027 30923
rect 20027 30889 20036 30923
rect 19984 30880 20036 30889
rect 20168 30923 20220 30932
rect 20168 30889 20177 30923
rect 20177 30889 20211 30923
rect 20211 30889 20220 30923
rect 20168 30880 20220 30889
rect 20260 30880 20312 30932
rect 9312 30812 9364 30864
rect 8300 30744 8352 30796
rect 12164 30812 12216 30864
rect 12256 30812 12308 30864
rect 16948 30812 17000 30864
rect 17408 30812 17460 30864
rect 22652 30880 22704 30932
rect 23204 30880 23256 30932
rect 25044 30880 25096 30932
rect 2228 30719 2280 30728
rect 2228 30685 2237 30719
rect 2237 30685 2271 30719
rect 2271 30685 2280 30719
rect 2228 30676 2280 30685
rect 8024 30676 8076 30728
rect 8668 30676 8720 30728
rect 9404 30676 9456 30728
rect 10508 30744 10560 30796
rect 10692 30744 10744 30796
rect 11336 30744 11388 30796
rect 12716 30744 12768 30796
rect 14556 30744 14608 30796
rect 10876 30719 10928 30728
rect 10876 30685 10885 30719
rect 10885 30685 10919 30719
rect 10919 30685 10928 30719
rect 10876 30676 10928 30685
rect 12256 30676 12308 30728
rect 12348 30719 12400 30728
rect 12348 30685 12357 30719
rect 12357 30685 12391 30719
rect 12391 30685 12400 30719
rect 12348 30676 12400 30685
rect 12624 30676 12676 30728
rect 13176 30676 13228 30728
rect 9036 30540 9088 30592
rect 9404 30540 9456 30592
rect 12992 30608 13044 30660
rect 13452 30676 13504 30728
rect 13636 30676 13688 30728
rect 14188 30719 14240 30728
rect 14188 30685 14197 30719
rect 14197 30685 14231 30719
rect 14231 30685 14240 30719
rect 14188 30676 14240 30685
rect 14372 30676 14424 30728
rect 14740 30676 14792 30728
rect 15200 30676 15252 30728
rect 15476 30676 15528 30728
rect 15844 30719 15896 30728
rect 15844 30685 15853 30719
rect 15853 30685 15887 30719
rect 15887 30685 15896 30719
rect 15844 30676 15896 30685
rect 17040 30719 17092 30728
rect 17040 30685 17049 30719
rect 17049 30685 17083 30719
rect 17083 30685 17092 30719
rect 17040 30676 17092 30685
rect 17224 30719 17276 30728
rect 17224 30685 17233 30719
rect 17233 30685 17267 30719
rect 17267 30685 17276 30719
rect 17224 30676 17276 30685
rect 17776 30744 17828 30796
rect 18420 30744 18472 30796
rect 17500 30719 17552 30728
rect 17500 30685 17509 30719
rect 17509 30685 17543 30719
rect 17543 30685 17552 30719
rect 17500 30676 17552 30685
rect 19064 30744 19116 30796
rect 19340 30744 19392 30796
rect 12348 30540 12400 30592
rect 12440 30540 12492 30592
rect 12816 30540 12868 30592
rect 15292 30608 15344 30660
rect 16212 30651 16264 30660
rect 16212 30617 16221 30651
rect 16221 30617 16255 30651
rect 16255 30617 16264 30651
rect 16212 30608 16264 30617
rect 19616 30676 19668 30728
rect 20076 30744 20128 30796
rect 23848 30812 23900 30864
rect 28080 30880 28132 30932
rect 25688 30812 25740 30864
rect 20168 30676 20220 30728
rect 21548 30676 21600 30728
rect 22928 30719 22980 30728
rect 22928 30685 22937 30719
rect 22937 30685 22971 30719
rect 22971 30685 22980 30719
rect 22928 30676 22980 30685
rect 23204 30719 23256 30728
rect 18788 30608 18840 30660
rect 18880 30608 18932 30660
rect 19800 30608 19852 30660
rect 20260 30608 20312 30660
rect 22468 30608 22520 30660
rect 23204 30685 23213 30719
rect 23213 30685 23247 30719
rect 23247 30685 23256 30719
rect 23204 30676 23256 30685
rect 23296 30719 23348 30728
rect 23296 30685 23305 30719
rect 23305 30685 23339 30719
rect 23339 30685 23348 30719
rect 23296 30676 23348 30685
rect 23112 30608 23164 30660
rect 24676 30676 24728 30728
rect 24860 30608 24912 30660
rect 16028 30583 16080 30592
rect 16028 30549 16037 30583
rect 16037 30549 16071 30583
rect 16071 30549 16080 30583
rect 16028 30540 16080 30549
rect 16120 30583 16172 30592
rect 16120 30549 16129 30583
rect 16129 30549 16163 30583
rect 16163 30549 16172 30583
rect 16856 30583 16908 30592
rect 16120 30540 16172 30549
rect 16856 30549 16865 30583
rect 16865 30549 16899 30583
rect 16899 30549 16908 30583
rect 16856 30540 16908 30549
rect 16948 30540 17000 30592
rect 18972 30540 19024 30592
rect 23480 30540 23532 30592
rect 25136 30676 25188 30728
rect 27068 30812 27120 30864
rect 27528 30744 27580 30796
rect 28724 30744 28776 30796
rect 26332 30719 26384 30728
rect 26332 30685 26341 30719
rect 26341 30685 26375 30719
rect 26375 30685 26384 30719
rect 26332 30676 26384 30685
rect 25504 30651 25556 30660
rect 25504 30617 25513 30651
rect 25513 30617 25547 30651
rect 25547 30617 25556 30651
rect 25504 30608 25556 30617
rect 27252 30608 27304 30660
rect 26976 30540 27028 30592
rect 10214 30438 10266 30490
rect 10278 30438 10330 30490
rect 10342 30438 10394 30490
rect 10406 30438 10458 30490
rect 10470 30438 10522 30490
rect 19478 30438 19530 30490
rect 19542 30438 19594 30490
rect 19606 30438 19658 30490
rect 19670 30438 19722 30490
rect 19734 30438 19786 30490
rect 9404 30268 9456 30320
rect 9680 30336 9732 30388
rect 10600 30336 10652 30388
rect 6736 30039 6788 30048
rect 6736 30005 6745 30039
rect 6745 30005 6779 30039
rect 6779 30005 6788 30039
rect 6736 29996 6788 30005
rect 8484 30200 8536 30252
rect 8760 30200 8812 30252
rect 9588 30200 9640 30252
rect 10140 30268 10192 30320
rect 10508 30268 10560 30320
rect 12348 30336 12400 30388
rect 12532 30336 12584 30388
rect 15292 30336 15344 30388
rect 15844 30336 15896 30388
rect 16304 30336 16356 30388
rect 18052 30336 18104 30388
rect 18972 30336 19024 30388
rect 11520 30268 11572 30320
rect 11612 30268 11664 30320
rect 12716 30268 12768 30320
rect 12348 30200 12400 30252
rect 14372 30268 14424 30320
rect 13452 30200 13504 30252
rect 14004 30243 14056 30252
rect 14004 30209 14013 30243
rect 14013 30209 14047 30243
rect 14047 30209 14056 30243
rect 14004 30200 14056 30209
rect 11244 30132 11296 30184
rect 12992 30132 13044 30184
rect 15292 30200 15344 30252
rect 15384 30200 15436 30252
rect 15844 30243 15896 30252
rect 15844 30209 15853 30243
rect 15853 30209 15887 30243
rect 15887 30209 15896 30243
rect 15844 30200 15896 30209
rect 16856 30268 16908 30320
rect 18880 30268 18932 30320
rect 19892 30336 19944 30388
rect 20076 30336 20128 30388
rect 20996 30336 21048 30388
rect 22928 30336 22980 30388
rect 25136 30336 25188 30388
rect 17684 30200 17736 30252
rect 19248 30311 19300 30320
rect 19248 30277 19282 30311
rect 19282 30277 19300 30311
rect 19248 30268 19300 30277
rect 19064 30200 19116 30252
rect 20720 30200 20772 30252
rect 16856 30132 16908 30184
rect 17040 30132 17092 30184
rect 8576 29996 8628 30048
rect 8668 30039 8720 30048
rect 8668 30005 8677 30039
rect 8677 30005 8711 30039
rect 8711 30005 8720 30039
rect 8668 29996 8720 30005
rect 9956 29996 10008 30048
rect 10324 30064 10376 30116
rect 11336 30064 11388 30116
rect 12716 30064 12768 30116
rect 13912 30064 13964 30116
rect 12808 29996 12860 30048
rect 13728 29996 13780 30048
rect 16948 30064 17000 30116
rect 18420 29996 18472 30048
rect 20168 30132 20220 30184
rect 20628 30132 20680 30184
rect 20904 30243 20956 30252
rect 20904 30209 20913 30243
rect 20913 30209 20947 30243
rect 20947 30209 20956 30243
rect 23572 30268 23624 30320
rect 24952 30268 25004 30320
rect 25504 30268 25556 30320
rect 20904 30200 20956 30209
rect 22100 30243 22152 30252
rect 22100 30209 22134 30243
rect 22134 30209 22152 30243
rect 22100 30200 22152 30209
rect 22928 30200 22980 30252
rect 25228 30243 25280 30252
rect 25228 30209 25237 30243
rect 25237 30209 25271 30243
rect 25271 30209 25280 30243
rect 25228 30200 25280 30209
rect 25412 30243 25464 30252
rect 25412 30209 25421 30243
rect 25421 30209 25455 30243
rect 25455 30209 25464 30243
rect 26884 30268 26936 30320
rect 25412 30200 25464 30209
rect 25688 30200 25740 30252
rect 26976 30243 27028 30252
rect 26976 30209 26985 30243
rect 26985 30209 27019 30243
rect 27019 30209 27028 30243
rect 26976 30200 27028 30209
rect 27068 30200 27120 30252
rect 27252 30243 27304 30252
rect 27252 30209 27261 30243
rect 27261 30209 27295 30243
rect 27295 30209 27304 30243
rect 27252 30200 27304 30209
rect 21180 30175 21232 30184
rect 21180 30141 21189 30175
rect 21189 30141 21223 30175
rect 21223 30141 21232 30175
rect 21180 30132 21232 30141
rect 23848 30132 23900 30184
rect 19156 29996 19208 30048
rect 20260 29996 20312 30048
rect 21364 30064 21416 30116
rect 23756 30064 23808 30116
rect 25964 30132 26016 30184
rect 26884 30132 26936 30184
rect 25320 29996 25372 30048
rect 27252 29996 27304 30048
rect 5582 29894 5634 29946
rect 5646 29894 5698 29946
rect 5710 29894 5762 29946
rect 5774 29894 5826 29946
rect 5838 29894 5890 29946
rect 14846 29894 14898 29946
rect 14910 29894 14962 29946
rect 14974 29894 15026 29946
rect 15038 29894 15090 29946
rect 15102 29894 15154 29946
rect 24110 29894 24162 29946
rect 24174 29894 24226 29946
rect 24238 29894 24290 29946
rect 24302 29894 24354 29946
rect 24366 29894 24418 29946
rect 9312 29792 9364 29844
rect 9404 29792 9456 29844
rect 10416 29792 10468 29844
rect 10508 29792 10560 29844
rect 12164 29724 12216 29776
rect 13452 29724 13504 29776
rect 6736 29656 6788 29708
rect 1400 29588 1452 29640
rect 3884 29588 3936 29640
rect 7564 29588 7616 29640
rect 8392 29631 8444 29640
rect 8392 29597 8401 29631
rect 8401 29597 8435 29631
rect 8435 29597 8444 29631
rect 8392 29588 8444 29597
rect 9220 29520 9272 29572
rect 10140 29588 10192 29640
rect 9680 29520 9732 29572
rect 10416 29588 10468 29640
rect 10784 29588 10836 29640
rect 11152 29588 11204 29640
rect 11520 29631 11572 29640
rect 11520 29597 11529 29631
rect 11529 29597 11563 29631
rect 11563 29597 11572 29631
rect 11704 29631 11756 29640
rect 11520 29588 11572 29597
rect 11704 29597 11713 29631
rect 11713 29597 11747 29631
rect 11747 29597 11756 29631
rect 11704 29588 11756 29597
rect 11796 29588 11848 29640
rect 12164 29631 12216 29640
rect 12164 29597 12173 29631
rect 12173 29597 12207 29631
rect 12207 29597 12216 29631
rect 12164 29588 12216 29597
rect 13176 29656 13228 29708
rect 14648 29724 14700 29776
rect 15752 29724 15804 29776
rect 16212 29724 16264 29776
rect 14004 29656 14056 29708
rect 17684 29792 17736 29844
rect 17592 29724 17644 29776
rect 18880 29792 18932 29844
rect 19984 29792 20036 29844
rect 20720 29792 20772 29844
rect 20904 29792 20956 29844
rect 21180 29792 21232 29844
rect 22100 29792 22152 29844
rect 24032 29792 24084 29844
rect 18420 29724 18472 29776
rect 21548 29724 21600 29776
rect 22284 29724 22336 29776
rect 25780 29792 25832 29844
rect 25964 29792 26016 29844
rect 25596 29724 25648 29776
rect 28264 29724 28316 29776
rect 17868 29656 17920 29708
rect 21732 29656 21784 29708
rect 21916 29699 21968 29708
rect 21916 29665 21925 29699
rect 21925 29665 21959 29699
rect 21959 29665 21968 29699
rect 21916 29656 21968 29665
rect 22836 29656 22888 29708
rect 13820 29588 13872 29640
rect 14096 29631 14148 29640
rect 14096 29597 14105 29631
rect 14105 29597 14139 29631
rect 14139 29597 14148 29631
rect 14096 29588 14148 29597
rect 9128 29452 9180 29504
rect 9404 29452 9456 29504
rect 10784 29495 10836 29504
rect 10784 29461 10793 29495
rect 10793 29461 10827 29495
rect 10827 29461 10836 29495
rect 10784 29452 10836 29461
rect 12256 29520 12308 29572
rect 12532 29520 12584 29572
rect 12624 29520 12676 29572
rect 15660 29520 15712 29572
rect 17868 29520 17920 29572
rect 19248 29631 19300 29640
rect 19248 29597 19257 29631
rect 19257 29597 19291 29631
rect 19291 29597 19300 29631
rect 19248 29588 19300 29597
rect 19432 29631 19484 29640
rect 19432 29597 19441 29631
rect 19441 29597 19475 29631
rect 19475 29597 19484 29631
rect 20352 29631 20404 29640
rect 19432 29588 19484 29597
rect 20352 29597 20361 29631
rect 20361 29597 20395 29631
rect 20395 29597 20404 29631
rect 20352 29588 20404 29597
rect 22376 29588 22428 29640
rect 24400 29656 24452 29708
rect 25872 29656 25924 29708
rect 23480 29631 23532 29640
rect 23480 29597 23489 29631
rect 23489 29597 23523 29631
rect 23523 29597 23532 29631
rect 23480 29588 23532 29597
rect 23940 29588 23992 29640
rect 25044 29588 25096 29640
rect 26332 29631 26384 29640
rect 26332 29597 26341 29631
rect 26341 29597 26375 29631
rect 26375 29597 26384 29631
rect 26332 29588 26384 29597
rect 17960 29495 18012 29504
rect 17960 29461 17969 29495
rect 17969 29461 18003 29495
rect 18003 29461 18012 29495
rect 17960 29452 18012 29461
rect 18328 29452 18380 29504
rect 18880 29452 18932 29504
rect 19984 29520 20036 29572
rect 23388 29520 23440 29572
rect 10214 29350 10266 29402
rect 10278 29350 10330 29402
rect 10342 29350 10394 29402
rect 10406 29350 10458 29402
rect 10470 29350 10522 29402
rect 19478 29350 19530 29402
rect 19542 29350 19594 29402
rect 19606 29350 19658 29402
rect 19670 29350 19722 29402
rect 19734 29350 19786 29402
rect 9220 29248 9272 29300
rect 10692 29248 10744 29300
rect 10784 29248 10836 29300
rect 13728 29248 13780 29300
rect 13820 29248 13872 29300
rect 18880 29248 18932 29300
rect 19064 29248 19116 29300
rect 21548 29248 21600 29300
rect 21732 29248 21784 29300
rect 24952 29248 25004 29300
rect 26792 29248 26844 29300
rect 1400 29155 1452 29164
rect 1400 29121 1409 29155
rect 1409 29121 1443 29155
rect 1443 29121 1452 29155
rect 1400 29112 1452 29121
rect 10876 29180 10928 29232
rect 1584 29087 1636 29096
rect 1584 29053 1593 29087
rect 1593 29053 1627 29087
rect 1627 29053 1636 29087
rect 1584 29044 1636 29053
rect 2780 29087 2832 29096
rect 2780 29053 2789 29087
rect 2789 29053 2823 29087
rect 2823 29053 2832 29087
rect 10048 29112 10100 29164
rect 10232 29112 10284 29164
rect 10416 29112 10468 29164
rect 10508 29112 10560 29164
rect 11796 29180 11848 29232
rect 11428 29112 11480 29164
rect 12256 29180 12308 29232
rect 12164 29112 12216 29164
rect 14096 29180 14148 29232
rect 14188 29180 14240 29232
rect 15568 29180 15620 29232
rect 15752 29180 15804 29232
rect 2780 29044 2832 29053
rect 7748 29019 7800 29028
rect 7748 28985 7757 29019
rect 7757 28985 7791 29019
rect 7791 28985 7800 29019
rect 7748 28976 7800 28985
rect 11520 29044 11572 29096
rect 11612 29044 11664 29096
rect 13084 29112 13136 29164
rect 15016 29155 15068 29164
rect 15016 29121 15025 29155
rect 15025 29121 15059 29155
rect 15059 29121 15068 29155
rect 16120 29180 16172 29232
rect 17960 29180 18012 29232
rect 18052 29180 18104 29232
rect 22100 29180 22152 29232
rect 23480 29180 23532 29232
rect 15016 29112 15068 29121
rect 16304 29112 16356 29164
rect 16764 29112 16816 29164
rect 18144 29112 18196 29164
rect 22008 29112 22060 29164
rect 22284 29112 22336 29164
rect 11336 28976 11388 29028
rect 12532 28976 12584 29028
rect 13636 28976 13688 29028
rect 9128 28908 9180 28960
rect 9496 28951 9548 28960
rect 9496 28917 9505 28951
rect 9505 28917 9539 28951
rect 9539 28917 9548 28951
rect 9496 28908 9548 28917
rect 10140 28951 10192 28960
rect 10140 28917 10149 28951
rect 10149 28917 10183 28951
rect 10183 28917 10192 28951
rect 10140 28908 10192 28917
rect 11428 28908 11480 28960
rect 13912 28951 13964 28960
rect 13912 28917 13921 28951
rect 13921 28917 13955 28951
rect 13955 28917 13964 28951
rect 15660 28976 15712 29028
rect 13912 28908 13964 28917
rect 15568 28908 15620 28960
rect 16856 29044 16908 29096
rect 17040 29044 17092 29096
rect 18420 29044 18472 29096
rect 17224 28976 17276 29028
rect 18788 29019 18840 29028
rect 18788 28985 18797 29019
rect 18797 28985 18831 29019
rect 18831 28985 18840 29019
rect 18788 28976 18840 28985
rect 16028 28908 16080 28960
rect 16948 28908 17000 28960
rect 17132 28908 17184 28960
rect 18328 28908 18380 28960
rect 19708 29087 19760 29096
rect 19708 29053 19717 29087
rect 19717 29053 19751 29087
rect 19751 29053 19760 29087
rect 19708 29044 19760 29053
rect 21732 29044 21784 29096
rect 21180 28908 21232 28960
rect 21364 28908 21416 28960
rect 21916 28908 21968 28960
rect 22652 29112 22704 29164
rect 22928 29112 22980 29164
rect 23204 29112 23256 29164
rect 23296 29155 23348 29164
rect 23296 29121 23305 29155
rect 23305 29121 23339 29155
rect 23339 29121 23348 29155
rect 23296 29112 23348 29121
rect 23572 29112 23624 29164
rect 24400 29112 24452 29164
rect 24584 29155 24636 29164
rect 24584 29121 24618 29155
rect 24618 29121 24636 29155
rect 24584 29112 24636 29121
rect 22836 29044 22888 29096
rect 23388 29044 23440 29096
rect 26332 29180 26384 29232
rect 26056 29112 26108 29164
rect 26884 29112 26936 29164
rect 27252 29155 27304 29164
rect 27252 29121 27261 29155
rect 27261 29121 27295 29155
rect 27295 29121 27304 29155
rect 27252 29112 27304 29121
rect 22284 28908 22336 28960
rect 22836 28908 22888 28960
rect 22928 28908 22980 28960
rect 23296 28908 23348 28960
rect 25412 28976 25464 29028
rect 25872 28976 25924 29028
rect 26056 28976 26108 29028
rect 28632 28976 28684 29028
rect 27620 28908 27672 28960
rect 5582 28806 5634 28858
rect 5646 28806 5698 28858
rect 5710 28806 5762 28858
rect 5774 28806 5826 28858
rect 5838 28806 5890 28858
rect 14846 28806 14898 28858
rect 14910 28806 14962 28858
rect 14974 28806 15026 28858
rect 15038 28806 15090 28858
rect 15102 28806 15154 28858
rect 24110 28806 24162 28858
rect 24174 28806 24226 28858
rect 24238 28806 24290 28858
rect 24302 28806 24354 28858
rect 24366 28806 24418 28858
rect 1584 28704 1636 28756
rect 1676 28500 1728 28552
rect 8852 28568 8904 28620
rect 8760 28500 8812 28552
rect 10600 28704 10652 28756
rect 10876 28704 10928 28756
rect 11060 28636 11112 28688
rect 10232 28568 10284 28620
rect 10600 28568 10652 28620
rect 11244 28611 11296 28620
rect 11244 28577 11276 28611
rect 11276 28577 11296 28611
rect 11244 28568 11296 28577
rect 12348 28704 12400 28756
rect 12440 28636 12492 28688
rect 17868 28704 17920 28756
rect 18328 28704 18380 28756
rect 19892 28636 19944 28688
rect 22008 28704 22060 28756
rect 21548 28636 21600 28688
rect 21732 28636 21784 28688
rect 23204 28704 23256 28756
rect 27620 28704 27672 28756
rect 13360 28568 13412 28620
rect 13728 28568 13780 28620
rect 14188 28568 14240 28620
rect 10048 28543 10100 28552
rect 8208 28407 8260 28416
rect 8208 28373 8217 28407
rect 8217 28373 8251 28407
rect 8251 28373 8260 28407
rect 8208 28364 8260 28373
rect 9220 28407 9272 28416
rect 9220 28373 9229 28407
rect 9229 28373 9263 28407
rect 9263 28373 9272 28407
rect 9220 28364 9272 28373
rect 10048 28509 10057 28543
rect 10057 28509 10091 28543
rect 10091 28509 10100 28543
rect 10048 28500 10100 28509
rect 10692 28432 10744 28484
rect 11336 28500 11388 28552
rect 12900 28500 12952 28552
rect 13084 28500 13136 28552
rect 13544 28543 13596 28552
rect 13544 28509 13553 28543
rect 13553 28509 13587 28543
rect 13587 28509 13596 28543
rect 13544 28500 13596 28509
rect 14372 28500 14424 28552
rect 14648 28500 14700 28552
rect 14740 28543 14792 28552
rect 14740 28509 14749 28543
rect 14749 28509 14783 28543
rect 14783 28509 14792 28543
rect 14740 28500 14792 28509
rect 17132 28568 17184 28620
rect 17500 28568 17552 28620
rect 16304 28500 16356 28552
rect 17224 28500 17276 28552
rect 18052 28500 18104 28552
rect 18328 28568 18380 28620
rect 19156 28568 19208 28620
rect 19708 28568 19760 28620
rect 11060 28364 11112 28416
rect 11612 28432 11664 28484
rect 11704 28432 11756 28484
rect 17132 28432 17184 28484
rect 20628 28500 20680 28552
rect 20720 28543 20772 28552
rect 20720 28509 20729 28543
rect 20729 28509 20763 28543
rect 20763 28509 20772 28543
rect 21732 28543 21784 28552
rect 20720 28500 20772 28509
rect 21732 28509 21741 28543
rect 21741 28509 21775 28543
rect 21775 28509 21784 28543
rect 21732 28500 21784 28509
rect 23112 28568 23164 28620
rect 28172 28611 28224 28620
rect 19340 28432 19392 28484
rect 19800 28475 19852 28484
rect 19800 28441 19809 28475
rect 19809 28441 19843 28475
rect 19843 28441 19852 28475
rect 19800 28432 19852 28441
rect 20812 28432 20864 28484
rect 12348 28364 12400 28416
rect 12440 28364 12492 28416
rect 13176 28364 13228 28416
rect 16120 28364 16172 28416
rect 16488 28364 16540 28416
rect 18236 28364 18288 28416
rect 19892 28364 19944 28416
rect 22928 28432 22980 28484
rect 23664 28475 23716 28484
rect 23664 28441 23673 28475
rect 23673 28441 23707 28475
rect 23707 28441 23716 28475
rect 23664 28432 23716 28441
rect 23756 28432 23808 28484
rect 24124 28432 24176 28484
rect 28172 28577 28181 28611
rect 28181 28577 28215 28611
rect 28215 28577 28224 28611
rect 28172 28568 28224 28577
rect 24492 28500 24544 28552
rect 24952 28500 25004 28552
rect 25688 28500 25740 28552
rect 26332 28543 26384 28552
rect 26332 28509 26341 28543
rect 26341 28509 26375 28543
rect 26375 28509 26384 28543
rect 26332 28500 26384 28509
rect 26516 28475 26568 28484
rect 26516 28441 26525 28475
rect 26525 28441 26559 28475
rect 26559 28441 26568 28475
rect 26516 28432 26568 28441
rect 22192 28364 22244 28416
rect 25596 28364 25648 28416
rect 25688 28364 25740 28416
rect 10214 28262 10266 28314
rect 10278 28262 10330 28314
rect 10342 28262 10394 28314
rect 10406 28262 10458 28314
rect 10470 28262 10522 28314
rect 19478 28262 19530 28314
rect 19542 28262 19594 28314
rect 19606 28262 19658 28314
rect 19670 28262 19722 28314
rect 19734 28262 19786 28314
rect 8300 28160 8352 28212
rect 12624 28160 12676 28212
rect 12808 28160 12860 28212
rect 13176 28160 13228 28212
rect 13912 28160 13964 28212
rect 14004 28160 14056 28212
rect 9680 28092 9732 28144
rect 11244 28092 11296 28144
rect 11980 28092 12032 28144
rect 9496 28067 9548 28076
rect 9496 28033 9505 28067
rect 9505 28033 9539 28067
rect 9539 28033 9548 28067
rect 9496 28024 9548 28033
rect 9956 28024 10008 28076
rect 8208 27956 8260 28008
rect 11520 28024 11572 28076
rect 11796 27956 11848 28008
rect 12808 28024 12860 28076
rect 13268 28067 13320 28076
rect 13268 28033 13277 28067
rect 13277 28033 13311 28067
rect 13311 28033 13320 28067
rect 13268 28024 13320 28033
rect 13452 28024 13504 28076
rect 12992 27956 13044 28008
rect 13820 27956 13872 28008
rect 11888 27888 11940 27940
rect 12624 27888 12676 27940
rect 14280 28092 14332 28144
rect 14648 28160 14700 28212
rect 15476 28160 15528 28212
rect 15844 28160 15896 28212
rect 16120 28160 16172 28212
rect 26516 28160 26568 28212
rect 28080 28203 28132 28212
rect 28080 28169 28089 28203
rect 28089 28169 28123 28203
rect 28123 28169 28132 28203
rect 28080 28160 28132 28169
rect 15292 28092 15344 28144
rect 18236 28092 18288 28144
rect 21364 28092 21416 28144
rect 22376 28092 22428 28144
rect 25044 28092 25096 28144
rect 27436 28092 27488 28144
rect 17224 28024 17276 28076
rect 17684 28024 17736 28076
rect 19064 28024 19116 28076
rect 21180 28024 21232 28076
rect 21548 28024 21600 28076
rect 23848 28024 23900 28076
rect 14096 27956 14148 28008
rect 17040 27956 17092 28008
rect 18236 27956 18288 28008
rect 18696 27956 18748 28008
rect 20812 27956 20864 28008
rect 12164 27820 12216 27872
rect 14004 27820 14056 27872
rect 15384 27888 15436 27940
rect 16488 27888 16540 27940
rect 18328 27888 18380 27940
rect 18604 27888 18656 27940
rect 20260 27888 20312 27940
rect 20628 27888 20680 27940
rect 21732 27888 21784 27940
rect 23480 27956 23532 28008
rect 24492 28024 24544 28076
rect 25596 28024 25648 28076
rect 27620 28024 27672 28076
rect 25044 27999 25096 28008
rect 23940 27888 23992 27940
rect 24124 27888 24176 27940
rect 25044 27965 25053 27999
rect 25053 27965 25087 27999
rect 25087 27965 25096 27999
rect 25044 27956 25096 27965
rect 26976 27956 27028 28008
rect 20720 27820 20772 27872
rect 21824 27820 21876 27872
rect 22376 27820 22428 27872
rect 23756 27820 23808 27872
rect 26056 27820 26108 27872
rect 27068 27820 27120 27872
rect 5582 27718 5634 27770
rect 5646 27718 5698 27770
rect 5710 27718 5762 27770
rect 5774 27718 5826 27770
rect 5838 27718 5890 27770
rect 14846 27718 14898 27770
rect 14910 27718 14962 27770
rect 14974 27718 15026 27770
rect 15038 27718 15090 27770
rect 15102 27718 15154 27770
rect 24110 27718 24162 27770
rect 24174 27718 24226 27770
rect 24238 27718 24290 27770
rect 24302 27718 24354 27770
rect 24366 27718 24418 27770
rect 9496 27616 9548 27668
rect 10876 27616 10928 27668
rect 12716 27616 12768 27668
rect 13452 27616 13504 27668
rect 15936 27616 15988 27668
rect 15108 27548 15160 27600
rect 16212 27548 16264 27600
rect 9496 27455 9548 27464
rect 9496 27421 9505 27455
rect 9505 27421 9539 27455
rect 9539 27421 9548 27455
rect 9496 27412 9548 27421
rect 10140 27455 10192 27464
rect 10140 27421 10149 27455
rect 10149 27421 10183 27455
rect 10183 27421 10192 27455
rect 10140 27412 10192 27421
rect 10692 27412 10744 27464
rect 10784 27455 10836 27464
rect 10784 27421 10793 27455
rect 10793 27421 10827 27455
rect 10827 27421 10836 27455
rect 11244 27455 11296 27464
rect 10784 27412 10836 27421
rect 11244 27421 11253 27455
rect 11253 27421 11287 27455
rect 11287 27421 11296 27455
rect 11244 27412 11296 27421
rect 9680 27344 9732 27396
rect 6828 27276 6880 27328
rect 9588 27276 9640 27328
rect 11060 27344 11112 27396
rect 11980 27412 12032 27464
rect 12440 27412 12492 27464
rect 15752 27480 15804 27532
rect 17040 27616 17092 27668
rect 17408 27616 17460 27668
rect 21732 27616 21784 27668
rect 22008 27616 22060 27668
rect 23204 27616 23256 27668
rect 23296 27659 23348 27668
rect 23296 27625 23305 27659
rect 23305 27625 23339 27659
rect 23339 27625 23348 27659
rect 23296 27616 23348 27625
rect 23756 27616 23808 27668
rect 17868 27548 17920 27600
rect 18052 27548 18104 27600
rect 13820 27412 13872 27464
rect 14096 27455 14148 27464
rect 14096 27421 14105 27455
rect 14105 27421 14139 27455
rect 14139 27421 14148 27455
rect 18236 27480 18288 27532
rect 18420 27523 18472 27532
rect 18420 27489 18429 27523
rect 18429 27489 18463 27523
rect 18463 27489 18472 27523
rect 18880 27548 18932 27600
rect 23112 27548 23164 27600
rect 25504 27548 25556 27600
rect 25964 27548 26016 27600
rect 18420 27480 18472 27489
rect 21916 27480 21968 27532
rect 14096 27412 14148 27421
rect 11612 27344 11664 27396
rect 12440 27276 12492 27328
rect 12716 27276 12768 27328
rect 12900 27344 12952 27396
rect 14004 27344 14056 27396
rect 18052 27412 18104 27464
rect 18604 27455 18656 27464
rect 18604 27421 18613 27455
rect 18613 27421 18647 27455
rect 18647 27421 18656 27455
rect 24124 27480 24176 27532
rect 22284 27455 22336 27464
rect 18604 27412 18656 27421
rect 15936 27344 15988 27396
rect 16856 27344 16908 27396
rect 22284 27421 22293 27455
rect 22293 27421 22327 27455
rect 22327 27421 22336 27455
rect 22284 27412 22336 27421
rect 22376 27412 22428 27464
rect 23572 27412 23624 27464
rect 25044 27412 25096 27464
rect 26332 27455 26384 27464
rect 26332 27421 26341 27455
rect 26341 27421 26375 27455
rect 26375 27421 26384 27455
rect 26332 27412 26384 27421
rect 19064 27344 19116 27396
rect 19248 27344 19300 27396
rect 19340 27344 19392 27396
rect 20720 27344 20772 27396
rect 20812 27344 20864 27396
rect 21088 27344 21140 27396
rect 22652 27344 22704 27396
rect 23940 27344 23992 27396
rect 25412 27344 25464 27396
rect 28172 27387 28224 27396
rect 28172 27353 28181 27387
rect 28181 27353 28215 27387
rect 28215 27353 28224 27387
rect 28172 27344 28224 27353
rect 14740 27276 14792 27328
rect 15200 27276 15252 27328
rect 17960 27276 18012 27328
rect 18236 27276 18288 27328
rect 22192 27276 22244 27328
rect 22560 27276 22612 27328
rect 24676 27276 24728 27328
rect 24860 27276 24912 27328
rect 10214 27174 10266 27226
rect 10278 27174 10330 27226
rect 10342 27174 10394 27226
rect 10406 27174 10458 27226
rect 10470 27174 10522 27226
rect 19478 27174 19530 27226
rect 19542 27174 19594 27226
rect 19606 27174 19658 27226
rect 19670 27174 19722 27226
rect 19734 27174 19786 27226
rect 9220 27072 9272 27124
rect 11428 27072 11480 27124
rect 12256 27072 12308 27124
rect 13452 27072 13504 27124
rect 18236 27072 18288 27124
rect 10140 27004 10192 27056
rect 11612 27004 11664 27056
rect 10784 26979 10836 26988
rect 9772 26868 9824 26920
rect 9956 26868 10008 26920
rect 9680 26843 9732 26852
rect 9680 26809 9689 26843
rect 9689 26809 9723 26843
rect 9723 26809 9732 26843
rect 9680 26800 9732 26809
rect 10784 26945 10793 26979
rect 10793 26945 10827 26979
rect 10827 26945 10836 26979
rect 10784 26936 10836 26945
rect 11704 26936 11756 26988
rect 12532 26936 12584 26988
rect 11796 26868 11848 26920
rect 12348 26868 12400 26920
rect 14188 27004 14240 27056
rect 16856 27004 16908 27056
rect 17960 27047 18012 27056
rect 17960 27013 17969 27047
rect 17969 27013 18003 27047
rect 18003 27013 18012 27047
rect 17960 27004 18012 27013
rect 18144 27004 18196 27056
rect 12716 26936 12768 26988
rect 12992 26979 13044 26988
rect 12992 26945 13001 26979
rect 13001 26945 13035 26979
rect 13035 26945 13044 26979
rect 12992 26936 13044 26945
rect 13820 26936 13872 26988
rect 14096 26936 14148 26988
rect 14648 26936 14700 26988
rect 14740 26936 14792 26988
rect 15016 26936 15068 26988
rect 15660 26936 15712 26988
rect 15844 26936 15896 26988
rect 16948 26979 17000 26988
rect 16948 26945 16957 26979
rect 16957 26945 16991 26979
rect 16991 26945 17000 26979
rect 16948 26936 17000 26945
rect 12164 26843 12216 26852
rect 12164 26809 12173 26843
rect 12173 26809 12207 26843
rect 12207 26809 12216 26843
rect 12164 26800 12216 26809
rect 12624 26843 12676 26852
rect 12624 26809 12633 26843
rect 12633 26809 12667 26843
rect 12667 26809 12676 26843
rect 12624 26800 12676 26809
rect 13544 26868 13596 26920
rect 13268 26800 13320 26852
rect 14004 26800 14056 26852
rect 15016 26800 15068 26852
rect 15568 26868 15620 26920
rect 16764 26868 16816 26920
rect 17684 26936 17736 26988
rect 17776 26936 17828 26988
rect 18512 27072 18564 27124
rect 19984 27072 20036 27124
rect 18420 27004 18472 27056
rect 22376 27072 22428 27124
rect 24584 27072 24636 27124
rect 27344 27072 27396 27124
rect 27896 27072 27948 27124
rect 22192 27004 22244 27056
rect 27804 27047 27856 27056
rect 27804 27013 27813 27047
rect 27813 27013 27847 27047
rect 27847 27013 27856 27047
rect 27804 27004 27856 27013
rect 17408 26868 17460 26920
rect 18880 26936 18932 26988
rect 21732 26936 21784 26988
rect 21824 26936 21876 26988
rect 22100 26979 22152 26988
rect 22100 26945 22109 26979
rect 22109 26945 22143 26979
rect 22143 26945 22152 26979
rect 22376 26979 22428 26988
rect 22100 26936 22152 26945
rect 22376 26945 22385 26979
rect 22385 26945 22419 26979
rect 22419 26945 22428 26979
rect 22376 26936 22428 26945
rect 22560 26936 22612 26988
rect 23848 26979 23900 26988
rect 23848 26945 23882 26979
rect 23882 26945 23900 26979
rect 23848 26936 23900 26945
rect 24124 26936 24176 26988
rect 25872 26979 25924 26988
rect 25872 26945 25881 26979
rect 25881 26945 25915 26979
rect 25915 26945 25924 26979
rect 25872 26936 25924 26945
rect 27436 26979 27488 26988
rect 27436 26945 27445 26979
rect 27445 26945 27479 26979
rect 27479 26945 27488 26979
rect 27436 26936 27488 26945
rect 9036 26775 9088 26784
rect 9036 26741 9045 26775
rect 9045 26741 9079 26775
rect 9079 26741 9088 26775
rect 9036 26732 9088 26741
rect 10232 26732 10284 26784
rect 11980 26775 12032 26784
rect 11980 26741 11989 26775
rect 11989 26741 12023 26775
rect 12023 26741 12032 26775
rect 11980 26732 12032 26741
rect 12256 26732 12308 26784
rect 12716 26732 12768 26784
rect 13728 26732 13780 26784
rect 14556 26732 14608 26784
rect 17500 26800 17552 26852
rect 18512 26868 18564 26920
rect 20628 26868 20680 26920
rect 23572 26911 23624 26920
rect 23572 26877 23581 26911
rect 23581 26877 23615 26911
rect 23615 26877 23624 26911
rect 23572 26868 23624 26877
rect 24584 26868 24636 26920
rect 15476 26732 15528 26784
rect 16120 26775 16172 26784
rect 16120 26741 16129 26775
rect 16129 26741 16163 26775
rect 16163 26741 16172 26775
rect 16120 26732 16172 26741
rect 19248 26800 19300 26852
rect 22008 26800 22060 26852
rect 24768 26800 24820 26852
rect 18052 26732 18104 26784
rect 18144 26732 18196 26784
rect 20076 26732 20128 26784
rect 20812 26732 20864 26784
rect 21272 26732 21324 26784
rect 21548 26732 21600 26784
rect 21640 26732 21692 26784
rect 22192 26732 22244 26784
rect 23572 26732 23624 26784
rect 25136 26800 25188 26852
rect 25688 26732 25740 26784
rect 5582 26630 5634 26682
rect 5646 26630 5698 26682
rect 5710 26630 5762 26682
rect 5774 26630 5826 26682
rect 5838 26630 5890 26682
rect 14846 26630 14898 26682
rect 14910 26630 14962 26682
rect 14974 26630 15026 26682
rect 15038 26630 15090 26682
rect 15102 26630 15154 26682
rect 24110 26630 24162 26682
rect 24174 26630 24226 26682
rect 24238 26630 24290 26682
rect 24302 26630 24354 26682
rect 24366 26630 24418 26682
rect 13544 26571 13596 26580
rect 9588 26367 9640 26376
rect 9588 26333 9597 26367
rect 9597 26333 9631 26367
rect 9631 26333 9640 26367
rect 9588 26324 9640 26333
rect 9864 26324 9916 26376
rect 12072 26460 12124 26512
rect 13544 26537 13553 26571
rect 13553 26537 13587 26571
rect 13587 26537 13596 26571
rect 13544 26528 13596 26537
rect 18420 26571 18472 26580
rect 15200 26503 15252 26512
rect 12164 26435 12216 26444
rect 12164 26401 12173 26435
rect 12173 26401 12207 26435
rect 12207 26401 12216 26435
rect 12164 26392 12216 26401
rect 13360 26392 13412 26444
rect 13912 26392 13964 26444
rect 11336 26367 11388 26376
rect 11336 26333 11345 26367
rect 11345 26333 11379 26367
rect 11379 26333 11388 26367
rect 11336 26324 11388 26333
rect 11520 26367 11572 26376
rect 11520 26333 11529 26367
rect 11529 26333 11563 26367
rect 11563 26333 11572 26367
rect 11520 26324 11572 26333
rect 11888 26324 11940 26376
rect 11612 26256 11664 26308
rect 11980 26256 12032 26308
rect 12256 26256 12308 26308
rect 12532 26256 12584 26308
rect 12624 26256 12676 26308
rect 13820 26256 13872 26308
rect 14004 26256 14056 26308
rect 14280 26324 14332 26376
rect 15200 26469 15209 26503
rect 15209 26469 15243 26503
rect 15243 26469 15252 26503
rect 15200 26460 15252 26469
rect 17316 26460 17368 26512
rect 17592 26460 17644 26512
rect 17868 26460 17920 26512
rect 18420 26537 18429 26571
rect 18429 26537 18463 26571
rect 18463 26537 18472 26571
rect 18420 26528 18472 26537
rect 18604 26528 18656 26580
rect 19616 26528 19668 26580
rect 20168 26528 20220 26580
rect 22284 26528 22336 26580
rect 23848 26571 23900 26580
rect 14556 26392 14608 26444
rect 14740 26392 14792 26444
rect 14924 26392 14976 26444
rect 15568 26392 15620 26444
rect 15752 26435 15804 26444
rect 15752 26401 15761 26435
rect 15761 26401 15795 26435
rect 15795 26401 15804 26435
rect 15752 26392 15804 26401
rect 18144 26392 18196 26444
rect 18328 26435 18380 26444
rect 18328 26401 18337 26435
rect 18337 26401 18371 26435
rect 18371 26401 18380 26435
rect 18328 26392 18380 26401
rect 17592 26367 17644 26376
rect 17592 26333 17601 26367
rect 17601 26333 17635 26367
rect 17635 26333 17644 26367
rect 17592 26324 17644 26333
rect 18788 26392 18840 26444
rect 18236 26299 18288 26308
rect 10968 26188 11020 26240
rect 12348 26188 12400 26240
rect 13084 26188 13136 26240
rect 13268 26188 13320 26240
rect 15200 26188 15252 26240
rect 15936 26188 15988 26240
rect 18236 26265 18245 26299
rect 18245 26265 18279 26299
rect 18279 26265 18288 26299
rect 18236 26256 18288 26265
rect 18880 26324 18932 26376
rect 21180 26392 21232 26444
rect 20168 26367 20220 26376
rect 20168 26333 20177 26367
rect 20177 26333 20211 26367
rect 20211 26333 20220 26367
rect 20168 26324 20220 26333
rect 20812 26324 20864 26376
rect 22744 26324 22796 26376
rect 23848 26537 23857 26571
rect 23857 26537 23891 26571
rect 23891 26537 23900 26571
rect 23848 26528 23900 26537
rect 24768 26571 24820 26580
rect 24768 26537 24777 26571
rect 24777 26537 24811 26571
rect 24811 26537 24820 26571
rect 24768 26528 24820 26537
rect 24952 26571 25004 26580
rect 24952 26537 24961 26571
rect 24961 26537 24995 26571
rect 24995 26537 25004 26571
rect 25780 26571 25832 26580
rect 24952 26528 25004 26537
rect 25780 26537 25789 26571
rect 25789 26537 25823 26571
rect 25823 26537 25832 26571
rect 25780 26528 25832 26537
rect 23296 26460 23348 26512
rect 23388 26435 23440 26444
rect 23388 26401 23397 26435
rect 23397 26401 23431 26435
rect 23431 26401 23440 26435
rect 23388 26392 23440 26401
rect 23572 26392 23624 26444
rect 28172 26435 28224 26444
rect 28172 26401 28181 26435
rect 28181 26401 28215 26435
rect 28215 26401 28224 26435
rect 28172 26392 28224 26401
rect 23664 26367 23716 26376
rect 23664 26333 23673 26367
rect 23673 26333 23707 26367
rect 23707 26333 23716 26367
rect 23664 26324 23716 26333
rect 25596 26367 25648 26376
rect 19708 26256 19760 26308
rect 20996 26256 21048 26308
rect 24584 26299 24636 26308
rect 24584 26265 24593 26299
rect 24593 26265 24627 26299
rect 24627 26265 24636 26299
rect 24584 26256 24636 26265
rect 25596 26333 25605 26367
rect 25605 26333 25639 26367
rect 25639 26333 25648 26367
rect 25596 26324 25648 26333
rect 25964 26324 26016 26376
rect 26056 26324 26108 26376
rect 24860 26256 24912 26308
rect 18604 26188 18656 26240
rect 18880 26188 18932 26240
rect 19892 26188 19944 26240
rect 21088 26188 21140 26240
rect 22376 26188 22428 26240
rect 25504 26188 25556 26240
rect 10214 26086 10266 26138
rect 10278 26086 10330 26138
rect 10342 26086 10394 26138
rect 10406 26086 10458 26138
rect 10470 26086 10522 26138
rect 19478 26086 19530 26138
rect 19542 26086 19594 26138
rect 19606 26086 19658 26138
rect 19670 26086 19722 26138
rect 19734 26086 19786 26138
rect 10784 25891 10836 25900
rect 10784 25857 10793 25891
rect 10793 25857 10827 25891
rect 10827 25857 10836 25891
rect 10784 25848 10836 25857
rect 11336 25848 11388 25900
rect 11428 25848 11480 25900
rect 13544 25916 13596 25968
rect 12164 25848 12216 25900
rect 13268 25848 13320 25900
rect 11244 25644 11296 25696
rect 12624 25712 12676 25764
rect 13820 25891 13872 25900
rect 13820 25857 13854 25891
rect 13854 25857 13872 25891
rect 13820 25848 13872 25857
rect 14832 25848 14884 25900
rect 13544 25823 13596 25832
rect 13544 25789 13553 25823
rect 13553 25789 13587 25823
rect 13587 25789 13596 25823
rect 13544 25780 13596 25789
rect 16580 25984 16632 26036
rect 15016 25848 15068 25900
rect 15108 25848 15160 25900
rect 16212 25848 16264 25900
rect 13728 25644 13780 25696
rect 15752 25823 15804 25832
rect 15752 25789 15761 25823
rect 15761 25789 15795 25823
rect 15795 25789 15804 25823
rect 16396 25848 16448 25900
rect 18604 25916 18656 25968
rect 22192 25984 22244 26036
rect 27344 26027 27396 26036
rect 17684 25848 17736 25900
rect 18328 25848 18380 25900
rect 18512 25891 18564 25900
rect 18512 25857 18521 25891
rect 18521 25857 18555 25891
rect 18555 25857 18564 25891
rect 18512 25848 18564 25857
rect 19156 25848 19208 25900
rect 20812 25891 20864 25900
rect 20812 25857 20821 25891
rect 20821 25857 20855 25891
rect 20855 25857 20864 25891
rect 20812 25848 20864 25857
rect 15752 25780 15804 25789
rect 21640 25780 21692 25832
rect 16028 25755 16080 25764
rect 16028 25721 16037 25755
rect 16037 25721 16071 25755
rect 16071 25721 16080 25755
rect 16028 25712 16080 25721
rect 14556 25644 14608 25696
rect 15660 25644 15712 25696
rect 20996 25712 21048 25764
rect 21824 25916 21876 25968
rect 22008 25848 22060 25900
rect 22100 25891 22152 25900
rect 22100 25857 22109 25891
rect 22109 25857 22143 25891
rect 22143 25857 22152 25891
rect 22100 25848 22152 25857
rect 22376 25848 22428 25900
rect 22192 25823 22244 25832
rect 22192 25789 22201 25823
rect 22201 25789 22235 25823
rect 22235 25789 22244 25823
rect 22192 25780 22244 25789
rect 27344 25993 27353 26027
rect 27353 25993 27387 26027
rect 27387 25993 27396 26027
rect 27344 25984 27396 25993
rect 27620 25984 27672 26036
rect 27068 25916 27120 25968
rect 22652 25780 22704 25832
rect 22836 25780 22888 25832
rect 23572 25848 23624 25900
rect 24492 25848 24544 25900
rect 24676 25848 24728 25900
rect 25780 25848 25832 25900
rect 23664 25780 23716 25832
rect 24032 25780 24084 25832
rect 25044 25823 25096 25832
rect 25044 25789 25053 25823
rect 25053 25789 25087 25823
rect 25087 25789 25096 25823
rect 25044 25780 25096 25789
rect 26056 25780 26108 25832
rect 22928 25712 22980 25764
rect 26424 25755 26476 25764
rect 16856 25644 16908 25696
rect 18052 25687 18104 25696
rect 18052 25653 18061 25687
rect 18061 25653 18095 25687
rect 18095 25653 18104 25687
rect 18052 25644 18104 25653
rect 18236 25644 18288 25696
rect 22468 25644 22520 25696
rect 23480 25644 23532 25696
rect 23848 25644 23900 25696
rect 24584 25687 24636 25696
rect 24584 25653 24593 25687
rect 24593 25653 24627 25687
rect 24627 25653 24636 25687
rect 24584 25644 24636 25653
rect 26424 25721 26433 25755
rect 26433 25721 26467 25755
rect 26467 25721 26476 25755
rect 26424 25712 26476 25721
rect 25228 25644 25280 25696
rect 5582 25542 5634 25594
rect 5646 25542 5698 25594
rect 5710 25542 5762 25594
rect 5774 25542 5826 25594
rect 5838 25542 5890 25594
rect 14846 25542 14898 25594
rect 14910 25542 14962 25594
rect 14974 25542 15026 25594
rect 15038 25542 15090 25594
rect 15102 25542 15154 25594
rect 24110 25542 24162 25594
rect 24174 25542 24226 25594
rect 24238 25542 24290 25594
rect 24302 25542 24354 25594
rect 24366 25542 24418 25594
rect 11060 25440 11112 25492
rect 11336 25440 11388 25492
rect 19892 25440 19944 25492
rect 21088 25440 21140 25492
rect 21640 25440 21692 25492
rect 12716 25372 12768 25424
rect 12992 25372 13044 25424
rect 14004 25372 14056 25424
rect 11428 25347 11480 25356
rect 10600 25236 10652 25288
rect 10784 25279 10836 25288
rect 10784 25245 10793 25279
rect 10793 25245 10827 25279
rect 10827 25245 10836 25279
rect 10784 25236 10836 25245
rect 11152 25236 11204 25288
rect 11428 25313 11437 25347
rect 11437 25313 11471 25347
rect 11471 25313 11480 25347
rect 11428 25304 11480 25313
rect 14280 25279 14332 25288
rect 14280 25245 14289 25279
rect 14289 25245 14323 25279
rect 14323 25245 14332 25279
rect 14280 25236 14332 25245
rect 14464 25236 14516 25288
rect 15016 25304 15068 25356
rect 15400 25347 15452 25356
rect 15400 25313 15402 25347
rect 15402 25313 15436 25347
rect 15436 25313 15452 25347
rect 15400 25304 15452 25313
rect 14648 25279 14700 25288
rect 14648 25245 14657 25279
rect 14657 25245 14691 25279
rect 14691 25245 14700 25279
rect 14648 25236 14700 25245
rect 11060 25168 11112 25220
rect 11520 25168 11572 25220
rect 12532 25168 12584 25220
rect 13176 25168 13228 25220
rect 13360 25211 13412 25220
rect 13360 25177 13369 25211
rect 13369 25177 13403 25211
rect 13403 25177 13412 25211
rect 13360 25168 13412 25177
rect 15200 25236 15252 25288
rect 16120 25304 16172 25356
rect 15936 25236 15988 25288
rect 17960 25372 18012 25424
rect 22284 25372 22336 25424
rect 23388 25440 23440 25492
rect 24676 25483 24728 25492
rect 24676 25449 24685 25483
rect 24685 25449 24719 25483
rect 24719 25449 24728 25483
rect 24676 25440 24728 25449
rect 16396 25347 16448 25356
rect 16396 25313 16405 25347
rect 16405 25313 16439 25347
rect 16439 25313 16448 25347
rect 16396 25304 16448 25313
rect 18144 25304 18196 25356
rect 14004 25100 14056 25152
rect 14924 25100 14976 25152
rect 15568 25100 15620 25152
rect 15844 25143 15896 25152
rect 15844 25109 15853 25143
rect 15853 25109 15887 25143
rect 15887 25109 15896 25143
rect 15844 25100 15896 25109
rect 16212 25168 16264 25220
rect 17040 25236 17092 25288
rect 19156 25304 19208 25356
rect 18604 25236 18656 25288
rect 18696 25236 18748 25288
rect 20628 25236 20680 25288
rect 22100 25236 22152 25288
rect 22376 25279 22428 25288
rect 22376 25245 22400 25279
rect 22400 25245 22428 25279
rect 22376 25236 22428 25245
rect 28172 25347 28224 25356
rect 28172 25313 28181 25347
rect 28181 25313 28215 25347
rect 28215 25313 28224 25347
rect 28172 25304 28224 25313
rect 22560 25279 22612 25288
rect 22560 25245 22569 25279
rect 22569 25245 22603 25279
rect 22603 25245 22612 25279
rect 23480 25279 23532 25288
rect 22560 25236 22612 25245
rect 23480 25245 23489 25279
rect 23489 25245 23523 25279
rect 23523 25245 23532 25279
rect 23480 25236 23532 25245
rect 16948 25168 17000 25220
rect 17224 25100 17276 25152
rect 17776 25143 17828 25152
rect 17776 25109 17785 25143
rect 17785 25109 17819 25143
rect 17819 25109 17828 25143
rect 17776 25100 17828 25109
rect 19248 25100 19300 25152
rect 19892 25100 19944 25152
rect 22652 25100 22704 25152
rect 23480 25100 23532 25152
rect 23664 25168 23716 25220
rect 24860 25100 24912 25152
rect 25228 25236 25280 25288
rect 25320 25279 25372 25288
rect 25320 25245 25329 25279
rect 25329 25245 25363 25279
rect 25363 25245 25372 25279
rect 26332 25279 26384 25288
rect 25320 25236 25372 25245
rect 26332 25245 26341 25279
rect 26341 25245 26375 25279
rect 26375 25245 26384 25279
rect 26332 25236 26384 25245
rect 25504 25168 25556 25220
rect 26516 25211 26568 25220
rect 26516 25177 26525 25211
rect 26525 25177 26559 25211
rect 26559 25177 26568 25211
rect 26516 25168 26568 25177
rect 10214 24998 10266 25050
rect 10278 24998 10330 25050
rect 10342 24998 10394 25050
rect 10406 24998 10458 25050
rect 10470 24998 10522 25050
rect 19478 24998 19530 25050
rect 19542 24998 19594 25050
rect 19606 24998 19658 25050
rect 19670 24998 19722 25050
rect 19734 24998 19786 25050
rect 11612 24896 11664 24948
rect 12072 24896 12124 24948
rect 12992 24896 13044 24948
rect 13728 24939 13780 24948
rect 13728 24905 13737 24939
rect 13737 24905 13771 24939
rect 13771 24905 13780 24939
rect 13728 24896 13780 24905
rect 14188 24896 14240 24948
rect 14556 24896 14608 24948
rect 14740 24896 14792 24948
rect 15016 24896 15068 24948
rect 10600 24828 10652 24880
rect 14004 24828 14056 24880
rect 15752 24896 15804 24948
rect 15936 24896 15988 24948
rect 17132 24896 17184 24948
rect 22100 24896 22152 24948
rect 22284 24896 22336 24948
rect 10324 24803 10376 24812
rect 10324 24769 10333 24803
rect 10333 24769 10367 24803
rect 10367 24769 10376 24803
rect 10324 24760 10376 24769
rect 11428 24692 11480 24744
rect 11888 24735 11940 24744
rect 11888 24701 11897 24735
rect 11897 24701 11931 24735
rect 11931 24701 11940 24735
rect 11888 24692 11940 24701
rect 11336 24624 11388 24676
rect 12072 24803 12124 24812
rect 12072 24769 12081 24803
rect 12081 24769 12115 24803
rect 12115 24769 12124 24803
rect 12072 24760 12124 24769
rect 12716 24735 12768 24744
rect 12716 24701 12725 24735
rect 12725 24701 12759 24735
rect 12759 24701 12768 24735
rect 12716 24692 12768 24701
rect 12808 24692 12860 24744
rect 13912 24760 13964 24812
rect 16028 24828 16080 24880
rect 16120 24828 16172 24880
rect 14280 24692 14332 24744
rect 14832 24692 14884 24744
rect 15384 24760 15436 24812
rect 15936 24760 15988 24812
rect 16856 24803 16908 24812
rect 16856 24769 16865 24803
rect 16865 24769 16899 24803
rect 16899 24769 16908 24803
rect 16856 24760 16908 24769
rect 17408 24760 17460 24812
rect 18236 24803 18288 24812
rect 18236 24769 18245 24803
rect 18245 24769 18279 24803
rect 18279 24769 18288 24803
rect 18236 24760 18288 24769
rect 18420 24803 18472 24812
rect 18420 24769 18429 24803
rect 18429 24769 18463 24803
rect 18463 24769 18472 24803
rect 18420 24760 18472 24769
rect 19340 24760 19392 24812
rect 20628 24803 20680 24812
rect 20628 24769 20637 24803
rect 20637 24769 20671 24803
rect 20671 24769 20680 24803
rect 20628 24760 20680 24769
rect 20812 24760 20864 24812
rect 18052 24692 18104 24744
rect 25228 24828 25280 24880
rect 21364 24760 21416 24812
rect 22376 24803 22428 24812
rect 22376 24769 22385 24803
rect 22385 24769 22419 24803
rect 22419 24769 22428 24803
rect 22376 24760 22428 24769
rect 22652 24803 22704 24812
rect 22652 24769 22661 24803
rect 22661 24769 22695 24803
rect 22695 24769 22704 24803
rect 22652 24760 22704 24769
rect 22836 24760 22888 24812
rect 23940 24760 23992 24812
rect 21640 24692 21692 24744
rect 23664 24692 23716 24744
rect 24124 24735 24176 24744
rect 13268 24624 13320 24676
rect 10876 24556 10928 24608
rect 11796 24556 11848 24608
rect 12440 24556 12492 24608
rect 16764 24624 16816 24676
rect 20812 24624 20864 24676
rect 21088 24624 21140 24676
rect 22192 24667 22244 24676
rect 22192 24633 22201 24667
rect 22201 24633 22235 24667
rect 22235 24633 22244 24667
rect 22192 24624 22244 24633
rect 14464 24599 14516 24608
rect 14464 24565 14473 24599
rect 14473 24565 14507 24599
rect 14507 24565 14516 24599
rect 14464 24556 14516 24565
rect 15660 24556 15712 24608
rect 15752 24556 15804 24608
rect 16120 24556 16172 24608
rect 16488 24556 16540 24608
rect 17040 24556 17092 24608
rect 18696 24556 18748 24608
rect 23204 24556 23256 24608
rect 24124 24701 24133 24735
rect 24133 24701 24167 24735
rect 24167 24701 24176 24735
rect 24124 24692 24176 24701
rect 26056 24828 26108 24880
rect 26148 24803 26200 24812
rect 26148 24769 26157 24803
rect 26157 24769 26191 24803
rect 26191 24769 26200 24803
rect 26148 24760 26200 24769
rect 25504 24735 25556 24744
rect 25504 24701 25513 24735
rect 25513 24701 25547 24735
rect 25547 24701 25556 24735
rect 25504 24692 25556 24701
rect 26608 24760 26660 24812
rect 26976 24760 27028 24812
rect 28540 24760 28592 24812
rect 26516 24624 26568 24676
rect 24676 24556 24728 24608
rect 25596 24556 25648 24608
rect 27160 24556 27212 24608
rect 27252 24556 27304 24608
rect 5582 24454 5634 24506
rect 5646 24454 5698 24506
rect 5710 24454 5762 24506
rect 5774 24454 5826 24506
rect 5838 24454 5890 24506
rect 14846 24454 14898 24506
rect 14910 24454 14962 24506
rect 14974 24454 15026 24506
rect 15038 24454 15090 24506
rect 15102 24454 15154 24506
rect 24110 24454 24162 24506
rect 24174 24454 24226 24506
rect 24238 24454 24290 24506
rect 24302 24454 24354 24506
rect 24366 24454 24418 24506
rect 10324 24352 10376 24404
rect 10968 24352 11020 24404
rect 11244 24352 11296 24404
rect 11796 24352 11848 24404
rect 12164 24352 12216 24404
rect 12624 24395 12676 24404
rect 12624 24361 12633 24395
rect 12633 24361 12667 24395
rect 12667 24361 12676 24395
rect 12624 24352 12676 24361
rect 12072 24327 12124 24336
rect 12072 24293 12081 24327
rect 12081 24293 12115 24327
rect 12115 24293 12124 24327
rect 12072 24284 12124 24293
rect 14740 24352 14792 24404
rect 13728 24284 13780 24336
rect 10600 24148 10652 24200
rect 10692 24191 10744 24200
rect 10692 24157 10701 24191
rect 10701 24157 10735 24191
rect 10735 24157 10744 24191
rect 10876 24191 10928 24200
rect 10692 24148 10744 24157
rect 10876 24157 10885 24191
rect 10885 24157 10919 24191
rect 10919 24157 10928 24191
rect 10876 24148 10928 24157
rect 11428 24148 11480 24200
rect 12992 24216 13044 24268
rect 13544 24259 13596 24268
rect 13544 24225 13553 24259
rect 13553 24225 13587 24259
rect 13587 24225 13596 24259
rect 13544 24216 13596 24225
rect 11980 24191 12032 24200
rect 11980 24157 11989 24191
rect 11989 24157 12023 24191
rect 12023 24157 12032 24191
rect 11980 24148 12032 24157
rect 12440 24080 12492 24132
rect 12900 24148 12952 24200
rect 15844 24284 15896 24336
rect 15016 24148 15068 24200
rect 15292 24191 15344 24200
rect 15292 24157 15301 24191
rect 15301 24157 15335 24191
rect 15335 24157 15344 24191
rect 15292 24148 15344 24157
rect 15456 24148 15508 24200
rect 16396 24352 16448 24404
rect 16764 24352 16816 24404
rect 22284 24352 22336 24404
rect 22560 24395 22612 24404
rect 22560 24361 22569 24395
rect 22569 24361 22603 24395
rect 22603 24361 22612 24395
rect 22560 24352 22612 24361
rect 25228 24352 25280 24404
rect 17224 24284 17276 24336
rect 17500 24284 17552 24336
rect 18696 24284 18748 24336
rect 20260 24284 20312 24336
rect 18144 24148 18196 24200
rect 22284 24216 22336 24268
rect 22836 24216 22888 24268
rect 23388 24216 23440 24268
rect 13728 24012 13780 24064
rect 14372 24012 14424 24064
rect 14556 24055 14608 24064
rect 14556 24021 14565 24055
rect 14565 24021 14599 24055
rect 14599 24021 14608 24055
rect 14556 24012 14608 24021
rect 15476 24055 15528 24064
rect 15476 24021 15485 24055
rect 15485 24021 15519 24055
rect 15519 24021 15528 24055
rect 16028 24080 16080 24132
rect 16120 24080 16172 24132
rect 18236 24080 18288 24132
rect 18696 24191 18748 24200
rect 18696 24157 18705 24191
rect 18705 24157 18739 24191
rect 18739 24157 18748 24191
rect 18696 24148 18748 24157
rect 18972 24148 19024 24200
rect 19156 24148 19208 24200
rect 18604 24080 18656 24132
rect 18788 24080 18840 24132
rect 22652 24148 22704 24200
rect 23020 24148 23072 24200
rect 21824 24080 21876 24132
rect 22468 24080 22520 24132
rect 23296 24080 23348 24132
rect 23848 24216 23900 24268
rect 28172 24259 28224 24268
rect 28172 24225 28181 24259
rect 28181 24225 28215 24259
rect 28215 24225 28224 24259
rect 28172 24216 28224 24225
rect 24952 24148 25004 24200
rect 26332 24191 26384 24200
rect 26332 24157 26341 24191
rect 26341 24157 26375 24191
rect 26375 24157 26384 24191
rect 26332 24148 26384 24157
rect 28080 24080 28132 24132
rect 15476 24012 15528 24021
rect 21640 24012 21692 24064
rect 22284 24012 22336 24064
rect 23664 24012 23716 24064
rect 24492 24012 24544 24064
rect 25780 24055 25832 24064
rect 25780 24021 25789 24055
rect 25789 24021 25823 24055
rect 25823 24021 25832 24055
rect 25780 24012 25832 24021
rect 10214 23910 10266 23962
rect 10278 23910 10330 23962
rect 10342 23910 10394 23962
rect 10406 23910 10458 23962
rect 10470 23910 10522 23962
rect 19478 23910 19530 23962
rect 19542 23910 19594 23962
rect 19606 23910 19658 23962
rect 19670 23910 19722 23962
rect 19734 23910 19786 23962
rect 13636 23808 13688 23860
rect 14096 23808 14148 23860
rect 14188 23808 14240 23860
rect 16028 23808 16080 23860
rect 17684 23808 17736 23860
rect 13176 23783 13228 23792
rect 1492 23672 1544 23724
rect 2044 23672 2096 23724
rect 9496 23715 9548 23724
rect 9496 23681 9505 23715
rect 9505 23681 9539 23715
rect 9539 23681 9548 23715
rect 9496 23672 9548 23681
rect 10232 23672 10284 23724
rect 10324 23715 10376 23724
rect 10324 23681 10333 23715
rect 10333 23681 10367 23715
rect 10367 23681 10376 23715
rect 10784 23715 10836 23724
rect 10324 23672 10376 23681
rect 10784 23681 10793 23715
rect 10793 23681 10827 23715
rect 10827 23681 10836 23715
rect 10784 23672 10836 23681
rect 11336 23672 11388 23724
rect 12440 23715 12492 23724
rect 12440 23681 12449 23715
rect 12449 23681 12483 23715
rect 12483 23681 12492 23715
rect 12440 23672 12492 23681
rect 12716 23672 12768 23724
rect 13176 23749 13185 23783
rect 13185 23749 13219 23783
rect 13219 23749 13228 23783
rect 13176 23740 13228 23749
rect 13084 23715 13136 23724
rect 13084 23681 13093 23715
rect 13093 23681 13127 23715
rect 13127 23681 13136 23715
rect 13084 23672 13136 23681
rect 13268 23715 13320 23724
rect 13268 23681 13277 23715
rect 13277 23681 13311 23715
rect 13311 23681 13320 23715
rect 13268 23672 13320 23681
rect 13728 23715 13780 23724
rect 13728 23681 13737 23715
rect 13737 23681 13771 23715
rect 13771 23681 13780 23715
rect 13728 23672 13780 23681
rect 13912 23715 13964 23724
rect 13912 23681 13921 23715
rect 13921 23681 13955 23715
rect 13955 23681 13964 23715
rect 13912 23672 13964 23681
rect 16764 23740 16816 23792
rect 14556 23715 14608 23724
rect 14556 23681 14565 23715
rect 14565 23681 14599 23715
rect 14599 23681 14608 23715
rect 14556 23672 14608 23681
rect 14740 23715 14792 23724
rect 14740 23681 14749 23715
rect 14749 23681 14783 23715
rect 14783 23681 14792 23715
rect 14740 23672 14792 23681
rect 15200 23672 15252 23724
rect 15384 23715 15436 23724
rect 15384 23681 15393 23715
rect 15393 23681 15427 23715
rect 15427 23681 15436 23715
rect 15384 23672 15436 23681
rect 15844 23672 15896 23724
rect 17500 23672 17552 23724
rect 15016 23604 15068 23656
rect 15660 23604 15712 23656
rect 16856 23604 16908 23656
rect 16948 23647 17000 23656
rect 16948 23613 16957 23647
rect 16957 23613 16991 23647
rect 16991 23613 17000 23647
rect 18604 23740 18656 23792
rect 18788 23808 18840 23860
rect 21640 23808 21692 23860
rect 21824 23851 21876 23860
rect 21824 23817 21833 23851
rect 21833 23817 21867 23851
rect 21867 23817 21876 23851
rect 21824 23808 21876 23817
rect 22100 23808 22152 23860
rect 19064 23740 19116 23792
rect 24308 23808 24360 23860
rect 24584 23808 24636 23860
rect 24676 23808 24728 23860
rect 26608 23808 26660 23860
rect 26976 23808 27028 23860
rect 28080 23851 28132 23860
rect 28080 23817 28089 23851
rect 28089 23817 28123 23851
rect 28123 23817 28132 23851
rect 28080 23808 28132 23817
rect 18144 23715 18196 23724
rect 18144 23681 18153 23715
rect 18153 23681 18187 23715
rect 18187 23681 18196 23715
rect 18144 23672 18196 23681
rect 18420 23672 18472 23724
rect 18052 23647 18104 23656
rect 16948 23604 17000 23613
rect 18052 23613 18061 23647
rect 18061 23613 18095 23647
rect 18095 23613 18104 23647
rect 18052 23604 18104 23613
rect 16764 23536 16816 23588
rect 18328 23536 18380 23588
rect 18880 23672 18932 23724
rect 18604 23604 18656 23656
rect 19892 23604 19944 23656
rect 20076 23647 20128 23656
rect 20076 23613 20085 23647
rect 20085 23613 20119 23647
rect 20119 23613 20128 23647
rect 20076 23604 20128 23613
rect 20260 23715 20312 23724
rect 20260 23681 20269 23715
rect 20269 23681 20303 23715
rect 20303 23681 20312 23715
rect 20260 23672 20312 23681
rect 20444 23715 20496 23724
rect 20444 23681 20453 23715
rect 20453 23681 20487 23715
rect 20487 23681 20496 23715
rect 21088 23715 21140 23724
rect 20444 23672 20496 23681
rect 21088 23681 21097 23715
rect 21097 23681 21131 23715
rect 21131 23681 21140 23715
rect 21088 23672 21140 23681
rect 21732 23672 21784 23724
rect 22008 23672 22060 23724
rect 22284 23715 22336 23724
rect 22284 23681 22293 23715
rect 22293 23681 22327 23715
rect 22327 23681 22336 23715
rect 22284 23672 22336 23681
rect 22560 23672 22612 23724
rect 25780 23740 25832 23792
rect 23480 23672 23532 23724
rect 24308 23715 24360 23724
rect 24308 23681 24317 23715
rect 24317 23681 24351 23715
rect 24351 23681 24360 23715
rect 24308 23672 24360 23681
rect 24860 23672 24912 23724
rect 25044 23715 25096 23724
rect 25044 23681 25053 23715
rect 25053 23681 25087 23715
rect 25087 23681 25096 23715
rect 25044 23672 25096 23681
rect 25596 23672 25648 23724
rect 27160 23715 27212 23724
rect 27160 23681 27169 23715
rect 27169 23681 27203 23715
rect 27203 23681 27212 23715
rect 27160 23672 27212 23681
rect 27988 23715 28040 23724
rect 27988 23681 27997 23715
rect 27997 23681 28031 23715
rect 28031 23681 28040 23715
rect 27988 23672 28040 23681
rect 22652 23604 22704 23656
rect 23204 23604 23256 23656
rect 27252 23647 27304 23656
rect 27252 23613 27261 23647
rect 27261 23613 27295 23647
rect 27295 23613 27304 23647
rect 27252 23604 27304 23613
rect 19708 23536 19760 23588
rect 1952 23511 2004 23520
rect 1952 23477 1961 23511
rect 1961 23477 1995 23511
rect 1995 23477 2004 23511
rect 1952 23468 2004 23477
rect 11704 23468 11756 23520
rect 11980 23468 12032 23520
rect 18788 23468 18840 23520
rect 19616 23468 19668 23520
rect 22284 23468 22336 23520
rect 23388 23468 23440 23520
rect 24584 23468 24636 23520
rect 25044 23536 25096 23588
rect 5582 23366 5634 23418
rect 5646 23366 5698 23418
rect 5710 23366 5762 23418
rect 5774 23366 5826 23418
rect 5838 23366 5890 23418
rect 14846 23366 14898 23418
rect 14910 23366 14962 23418
rect 14974 23366 15026 23418
rect 15038 23366 15090 23418
rect 15102 23366 15154 23418
rect 24110 23366 24162 23418
rect 24174 23366 24226 23418
rect 24238 23366 24290 23418
rect 24302 23366 24354 23418
rect 24366 23366 24418 23418
rect 11336 23307 11388 23316
rect 11336 23273 11345 23307
rect 11345 23273 11379 23307
rect 11379 23273 11388 23307
rect 11336 23264 11388 23273
rect 13360 23264 13412 23316
rect 13636 23264 13688 23316
rect 9496 23196 9548 23248
rect 15476 23239 15528 23248
rect 15476 23205 15485 23239
rect 15485 23205 15519 23239
rect 15519 23205 15528 23239
rect 15476 23196 15528 23205
rect 1952 23128 2004 23180
rect 2780 23171 2832 23180
rect 2780 23137 2789 23171
rect 2789 23137 2823 23171
rect 2823 23137 2832 23171
rect 2780 23128 2832 23137
rect 11704 23128 11756 23180
rect 2504 22992 2556 23044
rect 11060 23060 11112 23112
rect 11336 23103 11388 23112
rect 11336 23069 11345 23103
rect 11345 23069 11379 23103
rect 11379 23069 11388 23103
rect 11336 23060 11388 23069
rect 11520 23103 11572 23112
rect 11520 23069 11529 23103
rect 11529 23069 11563 23103
rect 11563 23069 11572 23103
rect 11520 23060 11572 23069
rect 11980 23103 12032 23112
rect 11980 23069 11989 23103
rect 11989 23069 12023 23103
rect 12023 23069 12032 23103
rect 11980 23060 12032 23069
rect 12164 23103 12216 23112
rect 12164 23069 12173 23103
rect 12173 23069 12207 23103
rect 12207 23069 12216 23103
rect 12164 23060 12216 23069
rect 12440 23060 12492 23112
rect 13268 23060 13320 23112
rect 13452 23060 13504 23112
rect 13820 23128 13872 23180
rect 15384 23128 15436 23180
rect 15844 23196 15896 23248
rect 16120 23239 16172 23248
rect 16120 23205 16129 23239
rect 16129 23205 16163 23239
rect 16163 23205 16172 23239
rect 17500 23264 17552 23316
rect 16120 23196 16172 23205
rect 18144 23264 18196 23316
rect 18788 23264 18840 23316
rect 19064 23264 19116 23316
rect 19432 23264 19484 23316
rect 20628 23264 20680 23316
rect 20720 23264 20772 23316
rect 25688 23264 25740 23316
rect 18420 23196 18472 23248
rect 15752 23128 15804 23180
rect 10968 22924 11020 22976
rect 14188 22924 14240 22976
rect 14464 22992 14516 23044
rect 14648 23060 14700 23112
rect 15844 23060 15896 23112
rect 17040 23128 17092 23180
rect 17316 23171 17368 23180
rect 17316 23137 17325 23171
rect 17325 23137 17359 23171
rect 17359 23137 17368 23171
rect 17316 23128 17368 23137
rect 16120 22992 16172 23044
rect 16212 22992 16264 23044
rect 16948 23060 17000 23112
rect 17132 23060 17184 23112
rect 18420 23103 18472 23112
rect 17040 22992 17092 23044
rect 16028 22924 16080 22976
rect 18420 23069 18429 23103
rect 18429 23069 18463 23103
rect 18463 23069 18472 23103
rect 18420 23060 18472 23069
rect 19156 23128 19208 23180
rect 19064 23060 19116 23112
rect 19432 23060 19484 23112
rect 19800 23128 19852 23180
rect 22192 23196 22244 23248
rect 22468 23196 22520 23248
rect 22928 23196 22980 23248
rect 20628 23060 20680 23112
rect 21364 23060 21416 23112
rect 22100 23103 22152 23112
rect 22100 23069 22109 23103
rect 22109 23069 22143 23103
rect 22143 23069 22152 23103
rect 22100 23060 22152 23069
rect 22284 23103 22336 23112
rect 22284 23069 22293 23103
rect 22293 23069 22327 23103
rect 22327 23069 22336 23103
rect 22284 23060 22336 23069
rect 22744 23128 22796 23180
rect 23664 23171 23716 23180
rect 23664 23137 23673 23171
rect 23673 23137 23707 23171
rect 23707 23137 23716 23171
rect 23664 23128 23716 23137
rect 23296 23060 23348 23112
rect 23572 23103 23624 23112
rect 23572 23069 23581 23103
rect 23581 23069 23615 23103
rect 23615 23069 23624 23103
rect 23756 23103 23808 23112
rect 23572 23060 23624 23069
rect 23756 23069 23765 23103
rect 23765 23069 23799 23103
rect 23799 23069 23808 23103
rect 23756 23060 23808 23069
rect 23848 23060 23900 23112
rect 24124 23060 24176 23112
rect 24400 23103 24452 23112
rect 24400 23069 24409 23103
rect 24409 23069 24443 23103
rect 24443 23069 24452 23103
rect 24400 23060 24452 23069
rect 28448 23196 28500 23248
rect 25044 23128 25096 23180
rect 26056 23128 26108 23180
rect 27160 23128 27212 23180
rect 28724 23128 28776 23180
rect 24768 23060 24820 23112
rect 17868 22992 17920 23044
rect 18328 22992 18380 23044
rect 20076 22992 20128 23044
rect 21824 22992 21876 23044
rect 22928 22992 22980 23044
rect 24676 23035 24728 23044
rect 20904 22924 20956 22976
rect 23940 22924 23992 22976
rect 24124 22924 24176 22976
rect 24676 23001 24685 23035
rect 24685 23001 24719 23035
rect 24719 23001 24728 23035
rect 24676 22992 24728 23001
rect 25228 22992 25280 23044
rect 24860 22924 24912 22976
rect 27068 22924 27120 22976
rect 10214 22822 10266 22874
rect 10278 22822 10330 22874
rect 10342 22822 10394 22874
rect 10406 22822 10458 22874
rect 10470 22822 10522 22874
rect 19478 22822 19530 22874
rect 19542 22822 19594 22874
rect 19606 22822 19658 22874
rect 19670 22822 19722 22874
rect 19734 22822 19786 22874
rect 2504 22763 2556 22772
rect 2504 22729 2513 22763
rect 2513 22729 2547 22763
rect 2547 22729 2556 22763
rect 2504 22720 2556 22729
rect 13544 22720 13596 22772
rect 15292 22720 15344 22772
rect 16948 22720 17000 22772
rect 18052 22720 18104 22772
rect 18144 22720 18196 22772
rect 21640 22720 21692 22772
rect 21824 22763 21876 22772
rect 21824 22729 21833 22763
rect 21833 22729 21867 22763
rect 21867 22729 21876 22763
rect 21824 22720 21876 22729
rect 2596 22584 2648 22636
rect 4988 22584 5040 22636
rect 10784 22627 10836 22636
rect 10784 22593 10793 22627
rect 10793 22593 10827 22627
rect 10827 22593 10836 22627
rect 10784 22584 10836 22593
rect 10968 22627 11020 22636
rect 10968 22593 10977 22627
rect 10977 22593 11011 22627
rect 11011 22593 11020 22627
rect 10968 22584 11020 22593
rect 11060 22584 11112 22636
rect 11980 22627 12032 22636
rect 11980 22593 11989 22627
rect 11989 22593 12023 22627
rect 12023 22593 12032 22627
rect 11980 22584 12032 22593
rect 12624 22627 12676 22636
rect 12624 22593 12633 22627
rect 12633 22593 12667 22627
rect 12667 22593 12676 22627
rect 12624 22584 12676 22593
rect 13176 22584 13228 22636
rect 14096 22627 14148 22636
rect 14096 22593 14105 22627
rect 14105 22593 14139 22627
rect 14139 22593 14148 22627
rect 14096 22584 14148 22593
rect 14832 22584 14884 22636
rect 13912 22516 13964 22568
rect 14464 22516 14516 22568
rect 15476 22652 15528 22704
rect 15752 22627 15804 22636
rect 15752 22593 15761 22627
rect 15761 22593 15795 22627
rect 15795 22593 15804 22627
rect 15752 22584 15804 22593
rect 17132 22652 17184 22704
rect 16672 22627 16724 22636
rect 16672 22593 16681 22627
rect 16681 22593 16715 22627
rect 16715 22593 16724 22627
rect 16672 22584 16724 22593
rect 16764 22584 16816 22636
rect 18512 22584 18564 22636
rect 19156 22652 19208 22704
rect 20076 22652 20128 22704
rect 19340 22584 19392 22636
rect 19432 22584 19484 22636
rect 16028 22516 16080 22568
rect 16120 22516 16172 22568
rect 17040 22516 17092 22568
rect 17776 22516 17828 22568
rect 20260 22584 20312 22636
rect 20996 22627 21048 22636
rect 20996 22593 21005 22627
rect 21005 22593 21039 22627
rect 21039 22593 21048 22627
rect 20996 22584 21048 22593
rect 22652 22652 22704 22704
rect 24492 22720 24544 22772
rect 23020 22584 23072 22636
rect 23204 22627 23256 22636
rect 23204 22593 23213 22627
rect 23213 22593 23247 22627
rect 23247 22593 23256 22627
rect 23204 22584 23256 22593
rect 23388 22627 23440 22636
rect 23388 22593 23397 22627
rect 23397 22593 23431 22627
rect 23431 22593 23440 22627
rect 23388 22584 23440 22593
rect 23664 22584 23716 22636
rect 20904 22559 20956 22568
rect 20904 22525 20913 22559
rect 20913 22525 20947 22559
rect 20947 22525 20956 22559
rect 25136 22652 25188 22704
rect 24768 22584 24820 22636
rect 20904 22516 20956 22525
rect 15016 22448 15068 22500
rect 15568 22448 15620 22500
rect 12072 22423 12124 22432
rect 12072 22389 12081 22423
rect 12081 22389 12115 22423
rect 12115 22389 12124 22423
rect 12072 22380 12124 22389
rect 14648 22380 14700 22432
rect 15384 22380 15436 22432
rect 15660 22380 15712 22432
rect 15844 22380 15896 22432
rect 16764 22423 16816 22432
rect 16764 22389 16773 22423
rect 16773 22389 16807 22423
rect 16807 22389 16816 22423
rect 16764 22380 16816 22389
rect 16948 22448 17000 22500
rect 18420 22448 18472 22500
rect 20168 22448 20220 22500
rect 23664 22448 23716 22500
rect 24676 22448 24728 22500
rect 25688 22584 25740 22636
rect 27712 22584 27764 22636
rect 28356 22584 28408 22636
rect 25044 22559 25096 22568
rect 25044 22525 25053 22559
rect 25053 22525 25087 22559
rect 25087 22525 25096 22559
rect 25044 22516 25096 22525
rect 27068 22559 27120 22568
rect 27068 22525 27077 22559
rect 27077 22525 27111 22559
rect 27111 22525 27120 22559
rect 27068 22516 27120 22525
rect 19616 22380 19668 22432
rect 20444 22423 20496 22432
rect 20444 22389 20453 22423
rect 20453 22389 20487 22423
rect 20487 22389 20496 22423
rect 20444 22380 20496 22389
rect 20812 22380 20864 22432
rect 23020 22380 23072 22432
rect 23296 22380 23348 22432
rect 25688 22380 25740 22432
rect 27252 22380 27304 22432
rect 27436 22423 27488 22432
rect 27436 22389 27445 22423
rect 27445 22389 27479 22423
rect 27479 22389 27488 22423
rect 27436 22380 27488 22389
rect 27528 22380 27580 22432
rect 5582 22278 5634 22330
rect 5646 22278 5698 22330
rect 5710 22278 5762 22330
rect 5774 22278 5826 22330
rect 5838 22278 5890 22330
rect 14846 22278 14898 22330
rect 14910 22278 14962 22330
rect 14974 22278 15026 22330
rect 15038 22278 15090 22330
rect 15102 22278 15154 22330
rect 24110 22278 24162 22330
rect 24174 22278 24226 22330
rect 24238 22278 24290 22330
rect 24302 22278 24354 22330
rect 24366 22278 24418 22330
rect 10784 22176 10836 22228
rect 14740 22176 14792 22228
rect 15660 22176 15712 22228
rect 12072 22108 12124 22160
rect 16304 22176 16356 22228
rect 16764 22176 16816 22228
rect 24032 22176 24084 22228
rect 24492 22176 24544 22228
rect 14372 22040 14424 22092
rect 15844 22040 15896 22092
rect 11244 22015 11296 22024
rect 11244 21981 11253 22015
rect 11253 21981 11287 22015
rect 11287 21981 11296 22015
rect 11244 21972 11296 21981
rect 11888 22015 11940 22024
rect 11888 21981 11897 22015
rect 11897 21981 11931 22015
rect 11931 21981 11940 22015
rect 11888 21972 11940 21981
rect 12808 21947 12860 21956
rect 12808 21913 12817 21947
rect 12817 21913 12851 21947
rect 12851 21913 12860 21947
rect 12808 21904 12860 21913
rect 13360 22015 13412 22024
rect 13360 21981 13369 22015
rect 13369 21981 13403 22015
rect 13403 21981 13412 22015
rect 13360 21972 13412 21981
rect 14004 21972 14056 22024
rect 15016 21972 15068 22024
rect 13452 21904 13504 21956
rect 13636 21904 13688 21956
rect 14464 21947 14516 21956
rect 14464 21913 14473 21947
rect 14473 21913 14507 21947
rect 14507 21913 14516 21947
rect 14464 21904 14516 21913
rect 15752 21972 15804 22024
rect 17500 22108 17552 22160
rect 17868 22108 17920 22160
rect 19248 22083 19300 22092
rect 16580 21972 16632 22024
rect 15016 21836 15068 21888
rect 16488 21904 16540 21956
rect 16948 21947 17000 21956
rect 16948 21913 16957 21947
rect 16957 21913 16991 21947
rect 16991 21913 17000 21947
rect 16948 21904 17000 21913
rect 17132 21947 17184 21956
rect 17132 21913 17141 21947
rect 17141 21913 17175 21947
rect 17175 21913 17184 21947
rect 17684 22015 17736 22024
rect 17684 21981 17693 22015
rect 17693 21981 17727 22015
rect 17727 21981 17736 22015
rect 17684 21972 17736 21981
rect 19248 22049 19257 22083
rect 19257 22049 19291 22083
rect 19291 22049 19300 22083
rect 19248 22040 19300 22049
rect 19616 22083 19668 22092
rect 19616 22049 19625 22083
rect 19625 22049 19659 22083
rect 19659 22049 19668 22083
rect 19616 22040 19668 22049
rect 20076 22083 20128 22092
rect 20076 22049 20085 22083
rect 20085 22049 20119 22083
rect 20119 22049 20128 22083
rect 20076 22040 20128 22049
rect 20444 22083 20496 22092
rect 20444 22049 20453 22083
rect 20453 22049 20487 22083
rect 20487 22049 20496 22083
rect 20444 22040 20496 22049
rect 18236 21972 18288 22024
rect 18328 21972 18380 22024
rect 18604 21972 18656 22024
rect 19892 21972 19944 22024
rect 20168 21972 20220 22024
rect 20996 22108 21048 22160
rect 22836 22108 22888 22160
rect 23296 22108 23348 22160
rect 21364 22040 21416 22092
rect 20996 22015 21048 22024
rect 20996 21981 21005 22015
rect 21005 21981 21039 22015
rect 21039 21981 21048 22015
rect 21732 22015 21784 22024
rect 20996 21972 21048 21981
rect 21732 21981 21741 22015
rect 21741 21981 21775 22015
rect 21775 21981 21784 22015
rect 21732 21972 21784 21981
rect 23664 22015 23716 22024
rect 23664 21981 23673 22015
rect 23673 21981 23707 22015
rect 23707 21981 23716 22015
rect 23664 21972 23716 21981
rect 24676 22015 24728 22024
rect 24676 21981 24685 22015
rect 24685 21981 24719 22015
rect 24719 21981 24728 22015
rect 24676 21972 24728 21981
rect 26056 22176 26108 22228
rect 25596 22040 25648 22092
rect 28172 22083 28224 22092
rect 28172 22049 28181 22083
rect 28181 22049 28215 22083
rect 28215 22049 28224 22083
rect 28172 22040 28224 22049
rect 17132 21904 17184 21913
rect 15384 21879 15436 21888
rect 15384 21845 15409 21879
rect 15409 21845 15436 21879
rect 15568 21879 15620 21888
rect 15384 21836 15436 21845
rect 15568 21845 15577 21879
rect 15577 21845 15611 21879
rect 15611 21845 15620 21879
rect 15568 21836 15620 21845
rect 16120 21836 16172 21888
rect 16304 21836 16356 21888
rect 19156 21836 19208 21888
rect 20076 21904 20128 21956
rect 20352 21904 20404 21956
rect 21364 21836 21416 21888
rect 23572 21904 23624 21956
rect 24584 21904 24636 21956
rect 24952 21972 25004 22024
rect 25412 21972 25464 22024
rect 25504 21947 25556 21956
rect 25504 21913 25513 21947
rect 25513 21913 25547 21947
rect 25547 21913 25556 21947
rect 25504 21904 25556 21913
rect 22652 21836 22704 21888
rect 24676 21836 24728 21888
rect 25964 21836 26016 21888
rect 27712 21836 27764 21888
rect 10214 21734 10266 21786
rect 10278 21734 10330 21786
rect 10342 21734 10394 21786
rect 10406 21734 10458 21786
rect 10470 21734 10522 21786
rect 19478 21734 19530 21786
rect 19542 21734 19594 21786
rect 19606 21734 19658 21786
rect 19670 21734 19722 21786
rect 19734 21734 19786 21786
rect 11888 21632 11940 21684
rect 16028 21632 16080 21684
rect 17316 21632 17368 21684
rect 17500 21632 17552 21684
rect 11796 21539 11848 21548
rect 11796 21505 11805 21539
rect 11805 21505 11839 21539
rect 11839 21505 11848 21539
rect 11796 21496 11848 21505
rect 12348 21564 12400 21616
rect 13728 21564 13780 21616
rect 12256 21428 12308 21480
rect 13636 21496 13688 21548
rect 13912 21539 13964 21548
rect 13912 21505 13921 21539
rect 13921 21505 13955 21539
rect 13955 21505 13964 21539
rect 15108 21564 15160 21616
rect 15384 21564 15436 21616
rect 15936 21564 15988 21616
rect 13912 21496 13964 21505
rect 12900 21428 12952 21480
rect 14648 21360 14700 21412
rect 16120 21496 16172 21548
rect 16488 21496 16540 21548
rect 15476 21428 15528 21480
rect 17684 21496 17736 21548
rect 18144 21539 18196 21548
rect 18144 21505 18153 21539
rect 18153 21505 18187 21539
rect 18187 21505 18196 21539
rect 18144 21496 18196 21505
rect 18880 21632 18932 21684
rect 19156 21632 19208 21684
rect 21364 21632 21416 21684
rect 22008 21632 22060 21684
rect 23664 21632 23716 21684
rect 24032 21632 24084 21684
rect 24768 21632 24820 21684
rect 26976 21675 27028 21684
rect 26976 21641 26985 21675
rect 26985 21641 27019 21675
rect 27019 21641 27028 21675
rect 26976 21632 27028 21641
rect 20260 21564 20312 21616
rect 20444 21564 20496 21616
rect 21272 21564 21324 21616
rect 21732 21564 21784 21616
rect 21916 21496 21968 21548
rect 17316 21471 17368 21480
rect 17316 21437 17325 21471
rect 17325 21437 17359 21471
rect 17359 21437 17368 21471
rect 17316 21428 17368 21437
rect 17960 21428 18012 21480
rect 20076 21428 20128 21480
rect 20720 21428 20772 21480
rect 21088 21428 21140 21480
rect 22376 21496 22428 21548
rect 25044 21564 25096 21616
rect 27344 21564 27396 21616
rect 22836 21496 22888 21548
rect 23020 21539 23072 21548
rect 23020 21505 23054 21539
rect 23054 21505 23072 21539
rect 23020 21496 23072 21505
rect 22652 21428 22704 21480
rect 14924 21360 14976 21412
rect 16764 21360 16816 21412
rect 18512 21360 18564 21412
rect 14556 21335 14608 21344
rect 14556 21301 14565 21335
rect 14565 21301 14599 21335
rect 14599 21301 14608 21335
rect 14556 21292 14608 21301
rect 14740 21292 14792 21344
rect 15200 21292 15252 21344
rect 16304 21292 16356 21344
rect 19340 21335 19392 21344
rect 19340 21301 19349 21335
rect 19349 21301 19383 21335
rect 19383 21301 19392 21335
rect 19340 21292 19392 21301
rect 20352 21292 20404 21344
rect 20628 21292 20680 21344
rect 20812 21292 20864 21344
rect 21364 21292 21416 21344
rect 22192 21360 22244 21412
rect 22376 21360 22428 21412
rect 24768 21471 24820 21480
rect 24768 21437 24777 21471
rect 24777 21437 24811 21471
rect 24811 21437 24820 21471
rect 24768 21428 24820 21437
rect 25228 21428 25280 21480
rect 27896 21539 27948 21548
rect 27896 21505 27905 21539
rect 27905 21505 27939 21539
rect 27939 21505 27948 21539
rect 27896 21496 27948 21505
rect 26148 21471 26200 21480
rect 26148 21437 26157 21471
rect 26157 21437 26191 21471
rect 26191 21437 26200 21471
rect 26148 21428 26200 21437
rect 26240 21428 26292 21480
rect 27252 21428 27304 21480
rect 27068 21360 27120 21412
rect 23756 21292 23808 21344
rect 24860 21292 24912 21344
rect 27252 21292 27304 21344
rect 27620 21292 27672 21344
rect 5582 21190 5634 21242
rect 5646 21190 5698 21242
rect 5710 21190 5762 21242
rect 5774 21190 5826 21242
rect 5838 21190 5890 21242
rect 14846 21190 14898 21242
rect 14910 21190 14962 21242
rect 14974 21190 15026 21242
rect 15038 21190 15090 21242
rect 15102 21190 15154 21242
rect 24110 21190 24162 21242
rect 24174 21190 24226 21242
rect 24238 21190 24290 21242
rect 24302 21190 24354 21242
rect 24366 21190 24418 21242
rect 13176 21088 13228 21140
rect 12072 21063 12124 21072
rect 12072 21029 12081 21063
rect 12081 21029 12115 21063
rect 12115 21029 12124 21063
rect 12072 21020 12124 21029
rect 11796 20952 11848 21004
rect 13912 21088 13964 21140
rect 15476 21131 15528 21140
rect 14096 21063 14148 21072
rect 14096 21029 14105 21063
rect 14105 21029 14139 21063
rect 14139 21029 14148 21063
rect 14096 21020 14148 21029
rect 13636 20952 13688 21004
rect 14004 20952 14056 21004
rect 14556 20952 14608 21004
rect 15476 21097 15485 21131
rect 15485 21097 15519 21131
rect 15519 21097 15528 21131
rect 15476 21088 15528 21097
rect 15200 20995 15252 21004
rect 15200 20961 15209 20995
rect 15209 20961 15243 20995
rect 15243 20961 15252 20995
rect 15200 20952 15252 20961
rect 15660 21088 15712 21140
rect 15844 21088 15896 21140
rect 19892 21088 19944 21140
rect 20168 21131 20220 21140
rect 20168 21097 20177 21131
rect 20177 21097 20211 21131
rect 20211 21097 20220 21131
rect 20168 21088 20220 21097
rect 16120 21020 16172 21072
rect 12440 20816 12492 20868
rect 9864 20748 9916 20800
rect 12624 20748 12676 20800
rect 13084 20884 13136 20936
rect 13268 20884 13320 20936
rect 16028 20952 16080 21004
rect 16212 20952 16264 21004
rect 16948 20952 17000 21004
rect 17316 20952 17368 21004
rect 17776 20995 17828 21004
rect 17776 20961 17785 20995
rect 17785 20961 17819 20995
rect 17819 20961 17828 20995
rect 17776 20952 17828 20961
rect 18052 21020 18104 21072
rect 22008 21088 22060 21140
rect 22652 21088 22704 21140
rect 23480 21088 23532 21140
rect 23664 21088 23716 21140
rect 25688 21088 25740 21140
rect 27436 21020 27488 21072
rect 18696 20952 18748 21004
rect 19248 20952 19300 21004
rect 13912 20748 13964 20800
rect 14648 20816 14700 20868
rect 14556 20748 14608 20800
rect 15292 20816 15344 20868
rect 15384 20816 15436 20868
rect 15660 20816 15712 20868
rect 14832 20748 14884 20800
rect 16304 20816 16356 20868
rect 16212 20791 16264 20800
rect 16212 20757 16221 20791
rect 16221 20757 16255 20791
rect 16255 20757 16264 20791
rect 16212 20748 16264 20757
rect 16672 20893 16681 20914
rect 16681 20893 16715 20914
rect 16715 20893 16724 20914
rect 16672 20862 16724 20893
rect 17684 20927 17736 20936
rect 17684 20893 17693 20927
rect 17693 20893 17727 20927
rect 17727 20893 17736 20927
rect 17684 20884 17736 20893
rect 17868 20884 17920 20936
rect 17960 20927 18012 20936
rect 17960 20893 17969 20927
rect 17969 20893 18003 20927
rect 18003 20893 18012 20927
rect 17960 20884 18012 20893
rect 18972 20884 19024 20936
rect 17132 20748 17184 20800
rect 18512 20748 18564 20800
rect 19616 20927 19668 20936
rect 19616 20893 19626 20927
rect 19626 20893 19660 20927
rect 19660 20893 19668 20927
rect 19616 20884 19668 20893
rect 20260 20884 20312 20936
rect 21272 20884 21324 20936
rect 22376 20884 22428 20936
rect 22560 20927 22612 20936
rect 22560 20893 22569 20927
rect 22569 20893 22603 20927
rect 22603 20893 22612 20927
rect 23480 20952 23532 21004
rect 25228 20995 25280 21004
rect 22560 20884 22612 20893
rect 20352 20816 20404 20868
rect 20904 20859 20956 20868
rect 20904 20825 20938 20859
rect 20938 20825 20956 20859
rect 23572 20927 23624 20936
rect 23572 20893 23581 20927
rect 23581 20893 23615 20927
rect 23615 20893 23624 20927
rect 23572 20884 23624 20893
rect 23664 20937 23716 20974
rect 23664 20922 23670 20937
rect 23670 20922 23704 20937
rect 23704 20922 23716 20937
rect 25228 20961 25237 20995
rect 25237 20961 25271 20995
rect 25271 20961 25280 20995
rect 25228 20952 25280 20961
rect 27528 20952 27580 21004
rect 28172 20995 28224 21004
rect 28172 20961 28181 20995
rect 28181 20961 28215 20995
rect 28215 20961 28224 20995
rect 28172 20952 28224 20961
rect 25136 20927 25188 20936
rect 25136 20893 25145 20927
rect 25145 20893 25179 20927
rect 25179 20893 25188 20927
rect 25136 20884 25188 20893
rect 26240 20884 26292 20936
rect 20904 20816 20956 20825
rect 20076 20748 20128 20800
rect 20260 20748 20312 20800
rect 22744 20791 22796 20800
rect 22744 20757 22753 20791
rect 22753 20757 22787 20791
rect 22787 20757 22796 20791
rect 22744 20748 22796 20757
rect 24584 20816 24636 20868
rect 26792 20816 26844 20868
rect 26056 20748 26108 20800
rect 10214 20646 10266 20698
rect 10278 20646 10330 20698
rect 10342 20646 10394 20698
rect 10406 20646 10458 20698
rect 10470 20646 10522 20698
rect 19478 20646 19530 20698
rect 19542 20646 19594 20698
rect 19606 20646 19658 20698
rect 19670 20646 19722 20698
rect 19734 20646 19786 20698
rect 14096 20544 14148 20596
rect 15384 20544 15436 20596
rect 16672 20544 16724 20596
rect 17868 20544 17920 20596
rect 18236 20544 18288 20596
rect 15200 20476 15252 20528
rect 14004 20408 14056 20460
rect 16028 20476 16080 20528
rect 14648 20340 14700 20392
rect 15752 20408 15804 20460
rect 16120 20408 16172 20460
rect 16304 20408 16356 20460
rect 19432 20476 19484 20528
rect 22836 20476 22888 20528
rect 23664 20544 23716 20596
rect 25596 20544 25648 20596
rect 27712 20544 27764 20596
rect 25136 20476 25188 20528
rect 19340 20408 19392 20460
rect 16856 20340 16908 20392
rect 17040 20383 17092 20392
rect 17040 20349 17049 20383
rect 17049 20349 17083 20383
rect 17083 20349 17092 20383
rect 17040 20340 17092 20349
rect 17132 20383 17184 20392
rect 17132 20349 17141 20383
rect 17141 20349 17175 20383
rect 17175 20349 17184 20383
rect 17132 20340 17184 20349
rect 14740 20315 14792 20324
rect 14740 20281 14749 20315
rect 14749 20281 14783 20315
rect 14783 20281 14792 20315
rect 14740 20272 14792 20281
rect 13176 20204 13228 20256
rect 15292 20204 15344 20256
rect 20536 20408 20588 20460
rect 21088 20451 21140 20460
rect 21088 20417 21097 20451
rect 21097 20417 21131 20451
rect 21131 20417 21140 20451
rect 21088 20408 21140 20417
rect 20628 20383 20680 20392
rect 20628 20349 20637 20383
rect 20637 20349 20671 20383
rect 20671 20349 20680 20383
rect 20628 20340 20680 20349
rect 22744 20451 22796 20460
rect 22744 20417 22753 20451
rect 22753 20417 22787 20451
rect 22787 20417 22796 20451
rect 22744 20408 22796 20417
rect 22928 20451 22980 20460
rect 22928 20417 22937 20451
rect 22937 20417 22971 20451
rect 22971 20417 22980 20451
rect 22928 20408 22980 20417
rect 23940 20408 23992 20460
rect 25320 20451 25372 20460
rect 23296 20340 23348 20392
rect 23848 20340 23900 20392
rect 20168 20247 20220 20256
rect 20168 20213 20177 20247
rect 20177 20213 20211 20247
rect 20211 20213 20220 20247
rect 20168 20204 20220 20213
rect 20444 20204 20496 20256
rect 22008 20272 22060 20324
rect 25320 20417 25329 20451
rect 25329 20417 25363 20451
rect 25363 20417 25372 20451
rect 25320 20408 25372 20417
rect 26424 20476 26476 20528
rect 26608 20476 26660 20528
rect 25228 20340 25280 20392
rect 25688 20383 25740 20392
rect 25688 20349 25697 20383
rect 25697 20349 25731 20383
rect 25731 20349 25740 20383
rect 25688 20340 25740 20349
rect 25780 20272 25832 20324
rect 26424 20340 26476 20392
rect 21548 20204 21600 20256
rect 24032 20204 24084 20256
rect 24492 20204 24544 20256
rect 24952 20204 25004 20256
rect 25872 20204 25924 20256
rect 5582 20102 5634 20154
rect 5646 20102 5698 20154
rect 5710 20102 5762 20154
rect 5774 20102 5826 20154
rect 5838 20102 5890 20154
rect 14846 20102 14898 20154
rect 14910 20102 14962 20154
rect 14974 20102 15026 20154
rect 15038 20102 15090 20154
rect 15102 20102 15154 20154
rect 24110 20102 24162 20154
rect 24174 20102 24226 20154
rect 24238 20102 24290 20154
rect 24302 20102 24354 20154
rect 24366 20102 24418 20154
rect 12900 20000 12952 20052
rect 14740 20000 14792 20052
rect 15476 20043 15528 20052
rect 15476 20009 15485 20043
rect 15485 20009 15519 20043
rect 15519 20009 15528 20043
rect 15476 20000 15528 20009
rect 15752 20000 15804 20052
rect 17040 20000 17092 20052
rect 17684 20043 17736 20052
rect 17684 20009 17693 20043
rect 17693 20009 17727 20043
rect 17727 20009 17736 20043
rect 17684 20000 17736 20009
rect 18144 20000 18196 20052
rect 18696 20000 18748 20052
rect 21640 20000 21692 20052
rect 22836 20000 22888 20052
rect 23572 20000 23624 20052
rect 18328 19932 18380 19984
rect 16028 19864 16080 19916
rect 16304 19907 16356 19916
rect 16304 19873 16313 19907
rect 16313 19873 16347 19907
rect 16347 19873 16356 19907
rect 16304 19864 16356 19873
rect 13544 19839 13596 19848
rect 13544 19805 13553 19839
rect 13553 19805 13587 19839
rect 13587 19805 13596 19839
rect 13544 19796 13596 19805
rect 14188 19796 14240 19848
rect 14648 19839 14700 19848
rect 14648 19805 14657 19839
rect 14657 19805 14691 19839
rect 14691 19805 14700 19839
rect 14648 19796 14700 19805
rect 15108 19839 15160 19848
rect 15108 19805 15117 19839
rect 15117 19805 15151 19839
rect 15151 19805 15160 19839
rect 15108 19796 15160 19805
rect 15476 19839 15528 19848
rect 15476 19805 15485 19839
rect 15485 19805 15519 19839
rect 15519 19805 15528 19839
rect 15476 19796 15528 19805
rect 16212 19796 16264 19848
rect 16948 19796 17000 19848
rect 19432 19907 19484 19916
rect 19432 19873 19441 19907
rect 19441 19873 19475 19907
rect 19475 19873 19484 19907
rect 19432 19864 19484 19873
rect 21272 19907 21324 19916
rect 21272 19873 21281 19907
rect 21281 19873 21315 19907
rect 21315 19873 21324 19907
rect 21272 19864 21324 19873
rect 23664 19932 23716 19984
rect 17960 19796 18012 19848
rect 19248 19796 19300 19848
rect 19524 19796 19576 19848
rect 20168 19796 20220 19848
rect 22008 19796 22060 19848
rect 23296 19839 23348 19848
rect 23296 19805 23305 19839
rect 23305 19805 23339 19839
rect 23339 19805 23348 19839
rect 23296 19796 23348 19805
rect 26516 19907 26568 19916
rect 26516 19873 26525 19907
rect 26525 19873 26559 19907
rect 26559 19873 26568 19907
rect 26516 19864 26568 19873
rect 23756 19796 23808 19848
rect 24676 19839 24728 19848
rect 24676 19805 24710 19839
rect 24710 19805 24728 19839
rect 15384 19728 15436 19780
rect 18880 19728 18932 19780
rect 20996 19728 21048 19780
rect 21548 19771 21600 19780
rect 21548 19737 21582 19771
rect 21582 19737 21600 19771
rect 24676 19796 24728 19805
rect 28172 19839 28224 19848
rect 21548 19728 21600 19737
rect 25044 19728 25096 19780
rect 28172 19805 28181 19839
rect 28181 19805 28215 19839
rect 28215 19805 28224 19839
rect 28172 19796 28224 19805
rect 27436 19728 27488 19780
rect 15568 19660 15620 19712
rect 16120 19660 16172 19712
rect 18696 19660 18748 19712
rect 19892 19660 19944 19712
rect 20628 19660 20680 19712
rect 22560 19660 22612 19712
rect 25780 19703 25832 19712
rect 25780 19669 25789 19703
rect 25789 19669 25823 19703
rect 25823 19669 25832 19703
rect 25780 19660 25832 19669
rect 10214 19558 10266 19610
rect 10278 19558 10330 19610
rect 10342 19558 10394 19610
rect 10406 19558 10458 19610
rect 10470 19558 10522 19610
rect 19478 19558 19530 19610
rect 19542 19558 19594 19610
rect 19606 19558 19658 19610
rect 19670 19558 19722 19610
rect 19734 19558 19786 19610
rect 13360 19456 13412 19508
rect 18788 19456 18840 19508
rect 13084 19388 13136 19440
rect 14740 19320 14792 19372
rect 16764 19388 16816 19440
rect 18420 19388 18472 19440
rect 13544 19252 13596 19304
rect 15108 19295 15160 19304
rect 15108 19261 15117 19295
rect 15117 19261 15151 19295
rect 15151 19261 15160 19295
rect 15108 19252 15160 19261
rect 14648 19184 14700 19236
rect 15936 19320 15988 19372
rect 17040 19320 17092 19372
rect 18052 19320 18104 19372
rect 18328 19363 18380 19372
rect 18328 19329 18337 19363
rect 18337 19329 18371 19363
rect 18371 19329 18380 19363
rect 18328 19320 18380 19329
rect 15568 19295 15620 19304
rect 15568 19261 15577 19295
rect 15577 19261 15611 19295
rect 15611 19261 15620 19295
rect 16948 19295 17000 19304
rect 15568 19252 15620 19261
rect 16948 19261 16957 19295
rect 16957 19261 16991 19295
rect 16991 19261 17000 19295
rect 16948 19252 17000 19261
rect 14556 19159 14608 19168
rect 14556 19125 14565 19159
rect 14565 19125 14599 19159
rect 14599 19125 14608 19159
rect 14556 19116 14608 19125
rect 15660 19184 15712 19236
rect 16856 19184 16908 19236
rect 17868 19184 17920 19236
rect 15568 19116 15620 19168
rect 16028 19116 16080 19168
rect 16488 19116 16540 19168
rect 18972 19456 19024 19508
rect 19248 19388 19300 19440
rect 20812 19456 20864 19508
rect 23480 19456 23532 19508
rect 26056 19456 26108 19508
rect 19432 19252 19484 19304
rect 19800 19320 19852 19372
rect 23296 19388 23348 19440
rect 23848 19431 23900 19440
rect 23848 19397 23857 19431
rect 23857 19397 23891 19431
rect 23891 19397 23900 19431
rect 23848 19388 23900 19397
rect 25780 19388 25832 19440
rect 20260 19320 20312 19372
rect 22192 19320 22244 19372
rect 23388 19320 23440 19372
rect 23572 19363 23624 19372
rect 23572 19329 23581 19363
rect 23581 19329 23615 19363
rect 23615 19329 23624 19363
rect 23572 19320 23624 19329
rect 23664 19320 23716 19372
rect 23940 19363 23992 19372
rect 23940 19329 23949 19363
rect 23949 19329 23983 19363
rect 23983 19329 23992 19363
rect 23940 19320 23992 19329
rect 25044 19363 25096 19372
rect 25044 19329 25053 19363
rect 25053 19329 25087 19363
rect 25087 19329 25096 19363
rect 25044 19320 25096 19329
rect 26884 19320 26936 19372
rect 20076 19295 20128 19304
rect 19524 19184 19576 19236
rect 20076 19261 20085 19295
rect 20085 19261 20119 19295
rect 20119 19261 20128 19295
rect 20076 19252 20128 19261
rect 20996 19252 21048 19304
rect 22100 19252 22152 19304
rect 27344 19320 27396 19372
rect 22560 19184 22612 19236
rect 23848 19184 23900 19236
rect 24308 19184 24360 19236
rect 21732 19116 21784 19168
rect 24860 19116 24912 19168
rect 25320 19116 25372 19168
rect 26424 19159 26476 19168
rect 26424 19125 26433 19159
rect 26433 19125 26467 19159
rect 26467 19125 26476 19159
rect 26424 19116 26476 19125
rect 26608 19116 26660 19168
rect 27252 19116 27304 19168
rect 5582 19014 5634 19066
rect 5646 19014 5698 19066
rect 5710 19014 5762 19066
rect 5774 19014 5826 19066
rect 5838 19014 5890 19066
rect 14846 19014 14898 19066
rect 14910 19014 14962 19066
rect 14974 19014 15026 19066
rect 15038 19014 15090 19066
rect 15102 19014 15154 19066
rect 24110 19014 24162 19066
rect 24174 19014 24226 19066
rect 24238 19014 24290 19066
rect 24302 19014 24354 19066
rect 24366 19014 24418 19066
rect 15200 18912 15252 18964
rect 16304 18912 16356 18964
rect 12716 18844 12768 18896
rect 15568 18887 15620 18896
rect 14188 18776 14240 18828
rect 14740 18776 14792 18828
rect 15568 18853 15577 18887
rect 15577 18853 15611 18887
rect 15611 18853 15620 18887
rect 15568 18844 15620 18853
rect 16120 18776 16172 18828
rect 14372 18751 14424 18760
rect 14372 18717 14381 18751
rect 14381 18717 14415 18751
rect 14415 18717 14424 18751
rect 14372 18708 14424 18717
rect 18880 18912 18932 18964
rect 19432 18912 19484 18964
rect 19892 18912 19944 18964
rect 20720 18912 20772 18964
rect 21180 18912 21232 18964
rect 22100 18912 22152 18964
rect 22468 18912 22520 18964
rect 23388 18912 23440 18964
rect 23572 18912 23624 18964
rect 17960 18887 18012 18896
rect 17960 18853 17969 18887
rect 17969 18853 18003 18887
rect 18003 18853 18012 18887
rect 17960 18844 18012 18853
rect 18052 18844 18104 18896
rect 17132 18751 17184 18760
rect 17132 18717 17141 18751
rect 17141 18717 17175 18751
rect 17175 18717 17184 18751
rect 17132 18708 17184 18717
rect 18144 18776 18196 18828
rect 21180 18819 21232 18828
rect 21180 18785 21189 18819
rect 21189 18785 21223 18819
rect 21223 18785 21232 18819
rect 21180 18776 21232 18785
rect 12808 18640 12860 18692
rect 16672 18640 16724 18692
rect 17500 18751 17552 18760
rect 17500 18717 17509 18751
rect 17509 18717 17543 18751
rect 17543 18717 17552 18751
rect 17500 18708 17552 18717
rect 18420 18708 18472 18760
rect 18880 18708 18932 18760
rect 18052 18640 18104 18692
rect 14372 18572 14424 18624
rect 15384 18572 15436 18624
rect 17316 18572 17368 18624
rect 18236 18572 18288 18624
rect 19524 18640 19576 18692
rect 20628 18708 20680 18760
rect 20996 18751 21048 18760
rect 20996 18717 21005 18751
rect 21005 18717 21039 18751
rect 21039 18717 21048 18751
rect 21732 18751 21784 18760
rect 20996 18708 21048 18717
rect 21732 18717 21741 18751
rect 21741 18717 21775 18751
rect 21775 18717 21784 18751
rect 21732 18708 21784 18717
rect 23204 18844 23256 18896
rect 27712 18912 27764 18964
rect 22100 18776 22152 18828
rect 20168 18640 20220 18692
rect 22192 18708 22244 18760
rect 22836 18708 22888 18760
rect 23756 18708 23808 18760
rect 27252 18844 27304 18896
rect 25504 18776 25556 18828
rect 28172 18819 28224 18828
rect 28172 18785 28181 18819
rect 28181 18785 28215 18819
rect 28215 18785 28224 18819
rect 28172 18776 28224 18785
rect 26332 18751 26384 18760
rect 26332 18717 26341 18751
rect 26341 18717 26375 18751
rect 26375 18717 26384 18751
rect 26332 18708 26384 18717
rect 22284 18640 22336 18692
rect 23296 18640 23348 18692
rect 24952 18640 25004 18692
rect 25136 18683 25188 18692
rect 25136 18649 25145 18683
rect 25145 18649 25179 18683
rect 25179 18649 25188 18683
rect 25136 18640 25188 18649
rect 26240 18640 26292 18692
rect 19892 18572 19944 18624
rect 20260 18615 20312 18624
rect 20260 18581 20285 18615
rect 20285 18581 20312 18615
rect 20444 18615 20496 18624
rect 20260 18572 20312 18581
rect 20444 18581 20453 18615
rect 20453 18581 20487 18615
rect 20487 18581 20496 18615
rect 20444 18572 20496 18581
rect 21824 18615 21876 18624
rect 21824 18581 21839 18615
rect 21839 18581 21873 18615
rect 21873 18581 21876 18615
rect 21824 18572 21876 18581
rect 22468 18615 22520 18624
rect 22468 18581 22477 18615
rect 22477 18581 22511 18615
rect 22511 18581 22520 18615
rect 22468 18572 22520 18581
rect 24308 18572 24360 18624
rect 10214 18470 10266 18522
rect 10278 18470 10330 18522
rect 10342 18470 10394 18522
rect 10406 18470 10458 18522
rect 10470 18470 10522 18522
rect 19478 18470 19530 18522
rect 19542 18470 19594 18522
rect 19606 18470 19658 18522
rect 19670 18470 19722 18522
rect 19734 18470 19786 18522
rect 17500 18368 17552 18420
rect 14188 18300 14240 18352
rect 13636 18275 13688 18284
rect 13636 18241 13645 18275
rect 13645 18241 13679 18275
rect 13679 18241 13688 18275
rect 13636 18232 13688 18241
rect 15200 18300 15252 18352
rect 17868 18368 17920 18420
rect 18052 18368 18104 18420
rect 18328 18368 18380 18420
rect 20628 18368 20680 18420
rect 22836 18368 22888 18420
rect 24492 18411 24544 18420
rect 24492 18377 24501 18411
rect 24501 18377 24535 18411
rect 24535 18377 24544 18411
rect 24492 18368 24544 18377
rect 26884 18368 26936 18420
rect 15292 18232 15344 18284
rect 16856 18232 16908 18284
rect 17316 18275 17368 18284
rect 17316 18241 17325 18275
rect 17325 18241 17359 18275
rect 17359 18241 17368 18275
rect 17316 18232 17368 18241
rect 17500 18275 17552 18284
rect 17500 18241 17509 18275
rect 17509 18241 17543 18275
rect 17543 18241 17552 18275
rect 17500 18232 17552 18241
rect 19248 18300 19300 18352
rect 22744 18343 22796 18352
rect 22744 18309 22753 18343
rect 22753 18309 22787 18343
rect 22787 18309 22796 18343
rect 22744 18300 22796 18309
rect 17868 18275 17920 18284
rect 17868 18241 17877 18275
rect 17877 18241 17911 18275
rect 17911 18241 17920 18275
rect 17868 18232 17920 18241
rect 18880 18275 18932 18284
rect 18144 18164 18196 18216
rect 15384 18096 15436 18148
rect 18880 18241 18889 18275
rect 18889 18241 18923 18275
rect 18923 18241 18932 18275
rect 18880 18232 18932 18241
rect 19340 18232 19392 18284
rect 19892 18232 19944 18284
rect 20076 18275 20128 18284
rect 20076 18241 20110 18275
rect 20110 18241 20128 18275
rect 20076 18232 20128 18241
rect 21824 18232 21876 18284
rect 22192 18232 22244 18284
rect 24860 18300 24912 18352
rect 24308 18275 24360 18284
rect 24308 18241 24317 18275
rect 24317 18241 24351 18275
rect 24351 18241 24360 18275
rect 24308 18232 24360 18241
rect 24584 18275 24636 18284
rect 24584 18241 24593 18275
rect 24593 18241 24627 18275
rect 24627 18241 24636 18275
rect 24584 18232 24636 18241
rect 24768 18232 24820 18284
rect 25044 18275 25096 18284
rect 25044 18241 25053 18275
rect 25053 18241 25087 18275
rect 25087 18241 25096 18275
rect 25044 18232 25096 18241
rect 26056 18232 26108 18284
rect 22284 18207 22336 18216
rect 22284 18173 22293 18207
rect 22293 18173 22327 18207
rect 22327 18173 22336 18207
rect 22284 18164 22336 18173
rect 1860 18071 1912 18080
rect 1860 18037 1869 18071
rect 1869 18037 1903 18071
rect 1903 18037 1912 18071
rect 1860 18028 1912 18037
rect 2412 18071 2464 18080
rect 2412 18037 2421 18071
rect 2421 18037 2455 18071
rect 2455 18037 2464 18071
rect 2412 18028 2464 18037
rect 14556 18028 14608 18080
rect 17868 18028 17920 18080
rect 18328 18028 18380 18080
rect 21456 18028 21508 18080
rect 21824 18071 21876 18080
rect 21824 18037 21833 18071
rect 21833 18037 21867 18071
rect 21867 18037 21876 18071
rect 21824 18028 21876 18037
rect 22192 18071 22244 18080
rect 22192 18037 22201 18071
rect 22201 18037 22235 18071
rect 22235 18037 22244 18071
rect 22192 18028 22244 18037
rect 22284 18028 22336 18080
rect 23388 18028 23440 18080
rect 27804 18300 27856 18352
rect 27620 18232 27672 18284
rect 26424 18164 26476 18216
rect 28264 18164 28316 18216
rect 27620 18096 27672 18148
rect 26976 18028 27028 18080
rect 27068 18028 27120 18080
rect 27344 18071 27396 18080
rect 27344 18037 27353 18071
rect 27353 18037 27387 18071
rect 27387 18037 27396 18071
rect 27344 18028 27396 18037
rect 27988 18071 28040 18080
rect 27988 18037 27997 18071
rect 27997 18037 28031 18071
rect 28031 18037 28040 18071
rect 27988 18028 28040 18037
rect 5582 17926 5634 17978
rect 5646 17926 5698 17978
rect 5710 17926 5762 17978
rect 5774 17926 5826 17978
rect 5838 17926 5890 17978
rect 14846 17926 14898 17978
rect 14910 17926 14962 17978
rect 14974 17926 15026 17978
rect 15038 17926 15090 17978
rect 15102 17926 15154 17978
rect 24110 17926 24162 17978
rect 24174 17926 24226 17978
rect 24238 17926 24290 17978
rect 24302 17926 24354 17978
rect 24366 17926 24418 17978
rect 6276 17824 6328 17876
rect 15660 17756 15712 17808
rect 1860 17688 1912 17740
rect 2780 17731 2832 17740
rect 2780 17697 2789 17731
rect 2789 17697 2823 17731
rect 2823 17697 2832 17731
rect 2780 17688 2832 17697
rect 14740 17688 14792 17740
rect 15200 17688 15252 17740
rect 15844 17731 15896 17740
rect 15844 17697 15853 17731
rect 15853 17697 15887 17731
rect 15887 17697 15896 17731
rect 15844 17688 15896 17697
rect 14556 17620 14608 17672
rect 17132 17824 17184 17876
rect 18236 17824 18288 17876
rect 20720 17824 20772 17876
rect 20996 17824 21048 17876
rect 19340 17756 19392 17808
rect 20260 17756 20312 17808
rect 24768 17824 24820 17876
rect 25320 17824 25372 17876
rect 26332 17824 26384 17876
rect 2412 17552 2464 17604
rect 15660 17552 15712 17604
rect 16488 17552 16540 17604
rect 17500 17552 17552 17604
rect 18236 17620 18288 17672
rect 18420 17620 18472 17672
rect 19248 17595 19300 17604
rect 19248 17561 19257 17595
rect 19257 17561 19291 17595
rect 19291 17561 19300 17595
rect 19248 17552 19300 17561
rect 19892 17620 19944 17672
rect 20996 17663 21048 17672
rect 20996 17629 21005 17663
rect 21005 17629 21039 17663
rect 21039 17629 21048 17663
rect 20996 17620 21048 17629
rect 21824 17620 21876 17672
rect 24308 17688 24360 17740
rect 24400 17731 24452 17740
rect 24400 17697 24409 17731
rect 24409 17697 24443 17731
rect 24443 17697 24452 17731
rect 24400 17688 24452 17697
rect 23572 17663 23624 17672
rect 23572 17629 23581 17663
rect 23581 17629 23615 17663
rect 23615 17629 23624 17663
rect 23572 17620 23624 17629
rect 23756 17663 23808 17672
rect 23756 17629 23765 17663
rect 23765 17629 23799 17663
rect 23799 17629 23808 17663
rect 23756 17620 23808 17629
rect 25688 17620 25740 17672
rect 28172 17731 28224 17740
rect 28172 17697 28181 17731
rect 28181 17697 28215 17731
rect 28215 17697 28224 17731
rect 28172 17688 28224 17697
rect 24768 17552 24820 17604
rect 27068 17552 27120 17604
rect 22284 17484 22336 17536
rect 23756 17484 23808 17536
rect 25596 17484 25648 17536
rect 10214 17382 10266 17434
rect 10278 17382 10330 17434
rect 10342 17382 10394 17434
rect 10406 17382 10458 17434
rect 10470 17382 10522 17434
rect 19478 17382 19530 17434
rect 19542 17382 19594 17434
rect 19606 17382 19658 17434
rect 19670 17382 19722 17434
rect 19734 17382 19786 17434
rect 15660 17323 15712 17332
rect 15660 17289 15669 17323
rect 15669 17289 15703 17323
rect 15703 17289 15712 17323
rect 15660 17280 15712 17289
rect 19248 17280 19300 17332
rect 19892 17280 19944 17332
rect 22744 17280 22796 17332
rect 23296 17280 23348 17332
rect 16028 17212 16080 17264
rect 17684 17212 17736 17264
rect 1584 17119 1636 17128
rect 1584 17085 1593 17119
rect 1593 17085 1627 17119
rect 1627 17085 1636 17119
rect 1584 17076 1636 17085
rect 1860 17119 1912 17128
rect 1860 17085 1869 17119
rect 1869 17085 1903 17119
rect 1903 17085 1912 17119
rect 1860 17076 1912 17085
rect 2504 17008 2556 17060
rect 15936 17144 15988 17196
rect 16488 17076 16540 17128
rect 16672 17119 16724 17128
rect 16672 17085 16681 17119
rect 16681 17085 16715 17119
rect 16715 17085 16724 17119
rect 16672 17076 16724 17085
rect 18420 17212 18472 17264
rect 18236 17187 18288 17196
rect 18236 17153 18270 17187
rect 18270 17153 18288 17187
rect 18236 17144 18288 17153
rect 20996 17212 21048 17264
rect 20444 17144 20496 17196
rect 22468 17144 22520 17196
rect 24492 17212 24544 17264
rect 25504 17255 25556 17264
rect 25504 17221 25513 17255
rect 25513 17221 25547 17255
rect 25547 17221 25556 17255
rect 25504 17212 25556 17221
rect 25596 17212 25648 17264
rect 23756 17144 23808 17196
rect 16856 17008 16908 17060
rect 16948 16940 17000 16992
rect 17776 16940 17828 16992
rect 21640 16940 21692 16992
rect 23388 16940 23440 16992
rect 25688 16983 25740 16992
rect 25688 16949 25697 16983
rect 25697 16949 25731 16983
rect 25731 16949 25740 16983
rect 25688 16940 25740 16949
rect 27988 17144 28040 17196
rect 26976 17119 27028 17128
rect 26976 17085 26985 17119
rect 26985 17085 27019 17119
rect 27019 17085 27028 17119
rect 26976 17076 27028 17085
rect 27528 17076 27580 17128
rect 26148 17008 26200 17060
rect 26700 16940 26752 16992
rect 27344 16983 27396 16992
rect 27344 16949 27353 16983
rect 27353 16949 27387 16983
rect 27387 16949 27396 16983
rect 27344 16940 27396 16949
rect 5582 16838 5634 16890
rect 5646 16838 5698 16890
rect 5710 16838 5762 16890
rect 5774 16838 5826 16890
rect 5838 16838 5890 16890
rect 14846 16838 14898 16890
rect 14910 16838 14962 16890
rect 14974 16838 15026 16890
rect 15038 16838 15090 16890
rect 15102 16838 15154 16890
rect 24110 16838 24162 16890
rect 24174 16838 24226 16890
rect 24238 16838 24290 16890
rect 24302 16838 24354 16890
rect 24366 16838 24418 16890
rect 1584 16736 1636 16788
rect 2504 16779 2556 16788
rect 2504 16745 2513 16779
rect 2513 16745 2547 16779
rect 2547 16745 2556 16779
rect 2504 16736 2556 16745
rect 17316 16736 17368 16788
rect 20444 16779 20496 16788
rect 15844 16600 15896 16652
rect 1676 16585 1728 16594
rect 1676 16551 1685 16585
rect 1685 16551 1719 16585
rect 1719 16551 1728 16585
rect 1676 16542 1728 16551
rect 16028 16575 16080 16584
rect 16028 16541 16037 16575
rect 16037 16541 16071 16575
rect 16071 16541 16080 16575
rect 16028 16532 16080 16541
rect 17224 16532 17276 16584
rect 20444 16745 20453 16779
rect 20453 16745 20487 16779
rect 20487 16745 20496 16779
rect 20444 16736 20496 16745
rect 21548 16736 21600 16788
rect 22100 16779 22152 16788
rect 22100 16745 22109 16779
rect 22109 16745 22143 16779
rect 22143 16745 22152 16779
rect 22100 16736 22152 16745
rect 23296 16736 23348 16788
rect 19340 16600 19392 16652
rect 21180 16668 21232 16720
rect 22008 16668 22060 16720
rect 19892 16532 19944 16584
rect 20720 16600 20772 16652
rect 21640 16575 21692 16584
rect 17132 16464 17184 16516
rect 18144 16464 18196 16516
rect 21640 16541 21649 16575
rect 21649 16541 21683 16575
rect 21683 16541 21692 16575
rect 22192 16600 22244 16652
rect 22836 16600 22888 16652
rect 23296 16600 23348 16652
rect 24492 16643 24544 16652
rect 21640 16532 21692 16541
rect 23388 16575 23440 16584
rect 23388 16541 23397 16575
rect 23397 16541 23431 16575
rect 23431 16541 23440 16575
rect 23388 16532 23440 16541
rect 24492 16609 24501 16643
rect 24501 16609 24535 16643
rect 24535 16609 24544 16643
rect 24492 16600 24544 16609
rect 26148 16532 26200 16584
rect 26332 16575 26384 16584
rect 26332 16541 26341 16575
rect 26341 16541 26375 16575
rect 26375 16541 26384 16575
rect 26332 16532 26384 16541
rect 22744 16464 22796 16516
rect 25596 16464 25648 16516
rect 26884 16464 26936 16516
rect 28172 16507 28224 16516
rect 28172 16473 28181 16507
rect 28181 16473 28215 16507
rect 28215 16473 28224 16507
rect 28172 16464 28224 16473
rect 16672 16396 16724 16448
rect 22284 16439 22336 16448
rect 22284 16405 22293 16439
rect 22293 16405 22327 16439
rect 22327 16405 22336 16439
rect 22284 16396 22336 16405
rect 23020 16396 23072 16448
rect 24860 16396 24912 16448
rect 25136 16396 25188 16448
rect 25504 16396 25556 16448
rect 10214 16294 10266 16346
rect 10278 16294 10330 16346
rect 10342 16294 10394 16346
rect 10406 16294 10458 16346
rect 10470 16294 10522 16346
rect 19478 16294 19530 16346
rect 19542 16294 19594 16346
rect 19606 16294 19658 16346
rect 19670 16294 19722 16346
rect 19734 16294 19786 16346
rect 16488 16192 16540 16244
rect 18236 16192 18288 16244
rect 20076 16192 20128 16244
rect 20904 16235 20956 16244
rect 20904 16201 20913 16235
rect 20913 16201 20947 16235
rect 20947 16201 20956 16235
rect 20904 16192 20956 16201
rect 22928 16192 22980 16244
rect 24676 16192 24728 16244
rect 16764 16124 16816 16176
rect 20536 16124 20588 16176
rect 16948 16056 17000 16108
rect 19340 16056 19392 16108
rect 20168 16056 20220 16108
rect 20352 16056 20404 16108
rect 20812 16099 20864 16108
rect 20812 16065 20821 16099
rect 20821 16065 20855 16099
rect 20855 16065 20864 16099
rect 20812 16056 20864 16065
rect 21364 16056 21416 16108
rect 22560 16124 22612 16176
rect 23204 16124 23256 16176
rect 22376 16056 22428 16108
rect 22744 16056 22796 16108
rect 23388 16056 23440 16108
rect 17960 15988 18012 16040
rect 23664 16056 23716 16108
rect 16856 15963 16908 15972
rect 16856 15929 16865 15963
rect 16865 15929 16899 15963
rect 16899 15929 16908 15963
rect 16856 15920 16908 15929
rect 27344 16124 27396 16176
rect 24584 16031 24636 16040
rect 23296 15920 23348 15972
rect 24584 15997 24593 16031
rect 24593 15997 24627 16031
rect 24627 15997 24636 16031
rect 24584 15988 24636 15997
rect 24860 15988 24912 16040
rect 27988 16056 28040 16108
rect 26148 16031 26200 16040
rect 26148 15997 26157 16031
rect 26157 15997 26191 16031
rect 26191 15997 26200 16031
rect 26148 15988 26200 15997
rect 28264 15920 28316 15972
rect 1400 15852 1452 15904
rect 23480 15895 23532 15904
rect 23480 15861 23489 15895
rect 23489 15861 23523 15895
rect 23523 15861 23532 15895
rect 23480 15852 23532 15861
rect 5582 15750 5634 15802
rect 5646 15750 5698 15802
rect 5710 15750 5762 15802
rect 5774 15750 5826 15802
rect 5838 15750 5890 15802
rect 14846 15750 14898 15802
rect 14910 15750 14962 15802
rect 14974 15750 15026 15802
rect 15038 15750 15090 15802
rect 15102 15750 15154 15802
rect 24110 15750 24162 15802
rect 24174 15750 24226 15802
rect 24238 15750 24290 15802
rect 24302 15750 24354 15802
rect 24366 15750 24418 15802
rect 17132 15691 17184 15700
rect 17132 15657 17141 15691
rect 17141 15657 17175 15691
rect 17175 15657 17184 15691
rect 17132 15648 17184 15657
rect 23664 15648 23716 15700
rect 27528 15648 27580 15700
rect 1400 15555 1452 15564
rect 1400 15521 1409 15555
rect 1409 15521 1443 15555
rect 1443 15521 1452 15555
rect 1400 15512 1452 15521
rect 2780 15555 2832 15564
rect 2780 15521 2789 15555
rect 2789 15521 2823 15555
rect 2823 15521 2832 15555
rect 2780 15512 2832 15521
rect 16948 15444 17000 15496
rect 17776 15444 17828 15496
rect 23480 15512 23532 15564
rect 24492 15580 24544 15632
rect 26332 15580 26384 15632
rect 25596 15444 25648 15496
rect 26332 15487 26384 15496
rect 26332 15453 26341 15487
rect 26341 15453 26375 15487
rect 26375 15453 26384 15487
rect 26332 15444 26384 15453
rect 1584 15419 1636 15428
rect 1584 15385 1593 15419
rect 1593 15385 1627 15419
rect 1627 15385 1636 15419
rect 1584 15376 1636 15385
rect 13820 15376 13872 15428
rect 23848 15376 23900 15428
rect 25136 15419 25188 15428
rect 25136 15385 25145 15419
rect 25145 15385 25179 15419
rect 25179 15385 25188 15419
rect 25136 15376 25188 15385
rect 23572 15308 23624 15360
rect 24860 15308 24912 15360
rect 25688 15376 25740 15428
rect 26516 15419 26568 15428
rect 26516 15385 26525 15419
rect 26525 15385 26559 15419
rect 26559 15385 26568 15419
rect 26516 15376 26568 15385
rect 28172 15419 28224 15428
rect 28172 15385 28181 15419
rect 28181 15385 28215 15419
rect 28215 15385 28224 15419
rect 28172 15376 28224 15385
rect 10214 15206 10266 15258
rect 10278 15206 10330 15258
rect 10342 15206 10394 15258
rect 10406 15206 10458 15258
rect 10470 15206 10522 15258
rect 19478 15206 19530 15258
rect 19542 15206 19594 15258
rect 19606 15206 19658 15258
rect 19670 15206 19722 15258
rect 19734 15206 19786 15258
rect 1584 15104 1636 15156
rect 23940 15104 23992 15156
rect 25044 15147 25096 15156
rect 25044 15113 25053 15147
rect 25053 15113 25087 15147
rect 25087 15113 25096 15147
rect 25044 15104 25096 15113
rect 26240 15104 26292 15156
rect 26516 15104 26568 15156
rect 27068 15104 27120 15156
rect 25228 15036 25280 15088
rect 1492 14968 1544 15020
rect 23388 14968 23440 15020
rect 24768 14968 24820 15020
rect 25136 14968 25188 15020
rect 25044 14900 25096 14952
rect 28540 15036 28592 15088
rect 27252 14968 27304 15020
rect 27804 14900 27856 14952
rect 14464 14832 14516 14884
rect 1400 14764 1452 14816
rect 27988 14764 28040 14816
rect 5582 14662 5634 14714
rect 5646 14662 5698 14714
rect 5710 14662 5762 14714
rect 5774 14662 5826 14714
rect 5838 14662 5890 14714
rect 14846 14662 14898 14714
rect 14910 14662 14962 14714
rect 14974 14662 15026 14714
rect 15038 14662 15090 14714
rect 15102 14662 15154 14714
rect 24110 14662 24162 14714
rect 24174 14662 24226 14714
rect 24238 14662 24290 14714
rect 24302 14662 24354 14714
rect 24366 14662 24418 14714
rect 24952 14603 25004 14612
rect 24952 14569 24961 14603
rect 24961 14569 24995 14603
rect 24995 14569 25004 14603
rect 24952 14560 25004 14569
rect 25872 14560 25924 14612
rect 25320 14492 25372 14544
rect 1400 14467 1452 14476
rect 1400 14433 1409 14467
rect 1409 14433 1443 14467
rect 1443 14433 1452 14467
rect 1400 14424 1452 14433
rect 1860 14467 1912 14476
rect 1860 14433 1869 14467
rect 1869 14433 1903 14467
rect 1903 14433 1912 14467
rect 1860 14424 1912 14433
rect 7656 14424 7708 14476
rect 9956 14424 10008 14476
rect 24860 14399 24912 14408
rect 24860 14365 24869 14399
rect 24869 14365 24903 14399
rect 24903 14365 24912 14399
rect 24860 14356 24912 14365
rect 26424 14492 26476 14544
rect 28080 14424 28132 14476
rect 1584 14331 1636 14340
rect 1584 14297 1593 14331
rect 1593 14297 1627 14331
rect 1627 14297 1636 14331
rect 1584 14288 1636 14297
rect 27804 14288 27856 14340
rect 28172 14331 28224 14340
rect 28172 14297 28181 14331
rect 28181 14297 28215 14331
rect 28215 14297 28224 14331
rect 28172 14288 28224 14297
rect 10214 14118 10266 14170
rect 10278 14118 10330 14170
rect 10342 14118 10394 14170
rect 10406 14118 10458 14170
rect 10470 14118 10522 14170
rect 19478 14118 19530 14170
rect 19542 14118 19594 14170
rect 19606 14118 19658 14170
rect 19670 14118 19722 14170
rect 19734 14118 19786 14170
rect 1584 14016 1636 14068
rect 25780 14059 25832 14068
rect 25780 14025 25789 14059
rect 25789 14025 25823 14059
rect 25823 14025 25832 14059
rect 25780 14016 25832 14025
rect 26884 14016 26936 14068
rect 27804 14059 27856 14068
rect 27804 14025 27813 14059
rect 27813 14025 27847 14059
rect 27847 14025 27856 14059
rect 27804 14016 27856 14025
rect 1860 13880 1912 13932
rect 25412 13880 25464 13932
rect 26976 13880 27028 13932
rect 12992 13812 13044 13864
rect 20628 13812 20680 13864
rect 25044 13812 25096 13864
rect 27252 13880 27304 13932
rect 27804 13812 27856 13864
rect 5582 13574 5634 13626
rect 5646 13574 5698 13626
rect 5710 13574 5762 13626
rect 5774 13574 5826 13626
rect 5838 13574 5890 13626
rect 14846 13574 14898 13626
rect 14910 13574 14962 13626
rect 14974 13574 15026 13626
rect 15038 13574 15090 13626
rect 15102 13574 15154 13626
rect 24110 13574 24162 13626
rect 24174 13574 24226 13626
rect 24238 13574 24290 13626
rect 24302 13574 24354 13626
rect 24366 13574 24418 13626
rect 24584 13472 24636 13524
rect 26056 13515 26108 13524
rect 26056 13481 26065 13515
rect 26065 13481 26099 13515
rect 26099 13481 26108 13515
rect 26056 13472 26108 13481
rect 27160 13515 27212 13524
rect 27160 13481 27169 13515
rect 27169 13481 27203 13515
rect 27203 13481 27212 13515
rect 27160 13472 27212 13481
rect 27344 13472 27396 13524
rect 1492 13268 1544 13320
rect 2412 13311 2464 13320
rect 2412 13277 2421 13311
rect 2421 13277 2455 13311
rect 2455 13277 2464 13311
rect 2412 13268 2464 13277
rect 27620 13336 27672 13388
rect 1400 13200 1452 13252
rect 26700 13268 26752 13320
rect 27804 13311 27856 13320
rect 25964 13200 26016 13252
rect 27804 13277 27813 13311
rect 27813 13277 27847 13311
rect 27847 13277 27856 13311
rect 27804 13268 27856 13277
rect 1584 13132 1636 13184
rect 10214 13030 10266 13082
rect 10278 13030 10330 13082
rect 10342 13030 10394 13082
rect 10406 13030 10458 13082
rect 10470 13030 10522 13082
rect 19478 13030 19530 13082
rect 19542 13030 19594 13082
rect 19606 13030 19658 13082
rect 19670 13030 19722 13082
rect 19734 13030 19786 13082
rect 1584 12903 1636 12912
rect 1584 12869 1593 12903
rect 1593 12869 1627 12903
rect 1627 12869 1636 12903
rect 1584 12860 1636 12869
rect 1400 12835 1452 12844
rect 1400 12801 1409 12835
rect 1409 12801 1443 12835
rect 1443 12801 1452 12835
rect 1400 12792 1452 12801
rect 26332 12792 26384 12844
rect 27436 12835 27488 12844
rect 27436 12801 27445 12835
rect 27445 12801 27479 12835
rect 27479 12801 27488 12835
rect 27436 12792 27488 12801
rect 2780 12767 2832 12776
rect 2780 12733 2789 12767
rect 2789 12733 2823 12767
rect 2823 12733 2832 12767
rect 2780 12724 2832 12733
rect 26792 12724 26844 12776
rect 5582 12486 5634 12538
rect 5646 12486 5698 12538
rect 5710 12486 5762 12538
rect 5774 12486 5826 12538
rect 5838 12486 5890 12538
rect 14846 12486 14898 12538
rect 14910 12486 14962 12538
rect 14974 12486 15026 12538
rect 15038 12486 15090 12538
rect 15102 12486 15154 12538
rect 24110 12486 24162 12538
rect 24174 12486 24226 12538
rect 24238 12486 24290 12538
rect 24302 12486 24354 12538
rect 24366 12486 24418 12538
rect 28080 12427 28132 12436
rect 28080 12393 28089 12427
rect 28089 12393 28123 12427
rect 28123 12393 28132 12427
rect 28080 12384 28132 12393
rect 2412 12248 2464 12300
rect 2780 12291 2832 12300
rect 2780 12257 2789 12291
rect 2789 12257 2823 12291
rect 2823 12257 2832 12291
rect 2780 12248 2832 12257
rect 26332 12180 26384 12232
rect 2504 12112 2556 12164
rect 10214 11942 10266 11994
rect 10278 11942 10330 11994
rect 10342 11942 10394 11994
rect 10406 11942 10458 11994
rect 10470 11942 10522 11994
rect 19478 11942 19530 11994
rect 19542 11942 19594 11994
rect 19606 11942 19658 11994
rect 19670 11942 19722 11994
rect 19734 11942 19786 11994
rect 2504 11883 2556 11892
rect 2504 11849 2513 11883
rect 2513 11849 2547 11883
rect 2547 11849 2556 11883
rect 2504 11840 2556 11849
rect 3700 11704 3752 11756
rect 7288 11704 7340 11756
rect 23756 11704 23808 11756
rect 27988 11747 28040 11756
rect 27988 11713 27997 11747
rect 27997 11713 28031 11747
rect 28031 11713 28040 11747
rect 27988 11704 28040 11713
rect 1860 11636 1912 11688
rect 12992 11636 13044 11688
rect 10140 11568 10192 11620
rect 1584 11500 1636 11552
rect 3240 11543 3292 11552
rect 3240 11509 3249 11543
rect 3249 11509 3283 11543
rect 3283 11509 3292 11543
rect 3240 11500 3292 11509
rect 26516 11500 26568 11552
rect 5582 11398 5634 11450
rect 5646 11398 5698 11450
rect 5710 11398 5762 11450
rect 5774 11398 5826 11450
rect 5838 11398 5890 11450
rect 14846 11398 14898 11450
rect 14910 11398 14962 11450
rect 14974 11398 15026 11450
rect 15038 11398 15090 11450
rect 15102 11398 15154 11450
rect 24110 11398 24162 11450
rect 24174 11398 24226 11450
rect 24238 11398 24290 11450
rect 24302 11398 24354 11450
rect 24366 11398 24418 11450
rect 3240 11228 3292 11280
rect 1584 11203 1636 11212
rect 1584 11169 1593 11203
rect 1593 11169 1627 11203
rect 1627 11169 1636 11203
rect 1584 11160 1636 11169
rect 1860 11203 1912 11212
rect 1860 11169 1869 11203
rect 1869 11169 1903 11203
rect 1903 11169 1912 11203
rect 1860 11160 1912 11169
rect 26332 11203 26384 11212
rect 26332 11169 26341 11203
rect 26341 11169 26375 11203
rect 26375 11169 26384 11203
rect 26332 11160 26384 11169
rect 26516 11203 26568 11212
rect 26516 11169 26525 11203
rect 26525 11169 26559 11203
rect 26559 11169 26568 11203
rect 26516 11160 26568 11169
rect 3976 11135 4028 11144
rect 3976 11101 3985 11135
rect 3985 11101 4019 11135
rect 4019 11101 4028 11135
rect 3976 11092 4028 11101
rect 28172 11067 28224 11076
rect 28172 11033 28181 11067
rect 28181 11033 28215 11067
rect 28215 11033 28224 11067
rect 28172 11024 28224 11033
rect 10214 10854 10266 10906
rect 10278 10854 10330 10906
rect 10342 10854 10394 10906
rect 10406 10854 10458 10906
rect 10470 10854 10522 10906
rect 19478 10854 19530 10906
rect 19542 10854 19594 10906
rect 19606 10854 19658 10906
rect 19670 10854 19722 10906
rect 19734 10854 19786 10906
rect 3976 10684 4028 10736
rect 17224 10616 17276 10668
rect 1952 10548 2004 10600
rect 2872 10591 2924 10600
rect 2872 10557 2881 10591
rect 2881 10557 2915 10591
rect 2915 10557 2924 10591
rect 2872 10548 2924 10557
rect 27344 10455 27396 10464
rect 27344 10421 27353 10455
rect 27353 10421 27387 10455
rect 27387 10421 27396 10455
rect 27344 10412 27396 10421
rect 27896 10455 27948 10464
rect 27896 10421 27905 10455
rect 27905 10421 27939 10455
rect 27939 10421 27948 10455
rect 27896 10412 27948 10421
rect 5582 10310 5634 10362
rect 5646 10310 5698 10362
rect 5710 10310 5762 10362
rect 5774 10310 5826 10362
rect 5838 10310 5890 10362
rect 14846 10310 14898 10362
rect 14910 10310 14962 10362
rect 14974 10310 15026 10362
rect 15038 10310 15090 10362
rect 15102 10310 15154 10362
rect 24110 10310 24162 10362
rect 24174 10310 24226 10362
rect 24238 10310 24290 10362
rect 24302 10310 24354 10362
rect 24366 10310 24418 10362
rect 1952 10251 2004 10260
rect 1952 10217 1961 10251
rect 1961 10217 1995 10251
rect 1995 10217 2004 10251
rect 1952 10208 2004 10217
rect 27896 10072 27948 10124
rect 2044 10004 2096 10056
rect 26332 10047 26384 10056
rect 26332 10013 26341 10047
rect 26341 10013 26375 10047
rect 26375 10013 26384 10047
rect 26332 10004 26384 10013
rect 27436 9936 27488 9988
rect 10214 9766 10266 9818
rect 10278 9766 10330 9818
rect 10342 9766 10394 9818
rect 10406 9766 10458 9818
rect 10470 9766 10522 9818
rect 19478 9766 19530 9818
rect 19542 9766 19594 9818
rect 19606 9766 19658 9818
rect 19670 9766 19722 9818
rect 19734 9766 19786 9818
rect 5448 9596 5500 9648
rect 24860 9596 24912 9648
rect 1492 9528 1544 9580
rect 26332 9528 26384 9580
rect 27712 9571 27764 9580
rect 27712 9537 27721 9571
rect 27721 9537 27755 9571
rect 27755 9537 27764 9571
rect 27712 9528 27764 9537
rect 1584 9324 1636 9376
rect 2412 9367 2464 9376
rect 2412 9333 2421 9367
rect 2421 9333 2455 9367
rect 2455 9333 2464 9367
rect 2412 9324 2464 9333
rect 27804 9367 27856 9376
rect 27804 9333 27813 9367
rect 27813 9333 27847 9367
rect 27847 9333 27856 9367
rect 27804 9324 27856 9333
rect 5582 9222 5634 9274
rect 5646 9222 5698 9274
rect 5710 9222 5762 9274
rect 5774 9222 5826 9274
rect 5838 9222 5890 9274
rect 14846 9222 14898 9274
rect 14910 9222 14962 9274
rect 14974 9222 15026 9274
rect 15038 9222 15090 9274
rect 15102 9222 15154 9274
rect 24110 9222 24162 9274
rect 24174 9222 24226 9274
rect 24238 9222 24290 9274
rect 24302 9222 24354 9274
rect 24366 9222 24418 9274
rect 2412 9052 2464 9104
rect 1584 9027 1636 9036
rect 1584 8993 1593 9027
rect 1593 8993 1627 9027
rect 1627 8993 1636 9027
rect 1584 8984 1636 8993
rect 2780 9027 2832 9036
rect 2780 8993 2789 9027
rect 2789 8993 2823 9027
rect 2823 8993 2832 9027
rect 27344 9052 27396 9104
rect 2780 8984 2832 8993
rect 27804 8984 27856 9036
rect 28172 9027 28224 9036
rect 28172 8993 28181 9027
rect 28181 8993 28215 9027
rect 28215 8993 28224 9027
rect 28172 8984 28224 8993
rect 10214 8678 10266 8730
rect 10278 8678 10330 8730
rect 10342 8678 10394 8730
rect 10406 8678 10458 8730
rect 10470 8678 10522 8730
rect 19478 8678 19530 8730
rect 19542 8678 19594 8730
rect 19606 8678 19658 8730
rect 19670 8678 19722 8730
rect 19734 8678 19786 8730
rect 1860 8483 1912 8492
rect 1860 8449 1869 8483
rect 1869 8449 1903 8483
rect 1903 8449 1912 8483
rect 1860 8440 1912 8449
rect 5448 8440 5500 8492
rect 21364 8372 21416 8424
rect 27988 8372 28040 8424
rect 27620 8304 27672 8356
rect 1584 8236 1636 8288
rect 2136 8236 2188 8288
rect 3332 8279 3384 8288
rect 3332 8245 3341 8279
rect 3341 8245 3375 8279
rect 3375 8245 3384 8279
rect 3332 8236 3384 8245
rect 27252 8279 27304 8288
rect 27252 8245 27261 8279
rect 27261 8245 27295 8279
rect 27295 8245 27304 8279
rect 27252 8236 27304 8245
rect 5582 8134 5634 8186
rect 5646 8134 5698 8186
rect 5710 8134 5762 8186
rect 5774 8134 5826 8186
rect 5838 8134 5890 8186
rect 14846 8134 14898 8186
rect 14910 8134 14962 8186
rect 14974 8134 15026 8186
rect 15038 8134 15090 8186
rect 15102 8134 15154 8186
rect 24110 8134 24162 8186
rect 24174 8134 24226 8186
rect 24238 8134 24290 8186
rect 24302 8134 24354 8186
rect 24366 8134 24418 8186
rect 3332 7964 3384 8016
rect 1584 7939 1636 7948
rect 1584 7905 1593 7939
rect 1593 7905 1627 7939
rect 1627 7905 1636 7939
rect 1584 7896 1636 7905
rect 2780 7939 2832 7948
rect 2780 7905 2789 7939
rect 2789 7905 2823 7939
rect 2823 7905 2832 7939
rect 2780 7896 2832 7905
rect 27252 7896 27304 7948
rect 1952 7760 2004 7812
rect 27804 7760 27856 7812
rect 28172 7803 28224 7812
rect 28172 7769 28181 7803
rect 28181 7769 28215 7803
rect 28215 7769 28224 7803
rect 28172 7760 28224 7769
rect 10214 7590 10266 7642
rect 10278 7590 10330 7642
rect 10342 7590 10394 7642
rect 10406 7590 10458 7642
rect 10470 7590 10522 7642
rect 19478 7590 19530 7642
rect 19542 7590 19594 7642
rect 19606 7590 19658 7642
rect 19670 7590 19722 7642
rect 19734 7590 19786 7642
rect 27804 7531 27856 7540
rect 27804 7497 27813 7531
rect 27813 7497 27847 7531
rect 27847 7497 27856 7531
rect 27804 7488 27856 7497
rect 2136 7463 2188 7472
rect 2136 7429 2145 7463
rect 2145 7429 2179 7463
rect 2179 7429 2188 7463
rect 2136 7420 2188 7429
rect 1952 7395 2004 7404
rect 1952 7361 1961 7395
rect 1961 7361 1995 7395
rect 1995 7361 2004 7395
rect 1952 7352 2004 7361
rect 27712 7395 27764 7404
rect 27712 7361 27721 7395
rect 27721 7361 27755 7395
rect 27755 7361 27764 7395
rect 27712 7352 27764 7361
rect 2964 7327 3016 7336
rect 2964 7293 2973 7327
rect 2973 7293 3007 7327
rect 3007 7293 3016 7327
rect 2964 7284 3016 7293
rect 4436 7191 4488 7200
rect 4436 7157 4445 7191
rect 4445 7157 4479 7191
rect 4479 7157 4488 7191
rect 4436 7148 4488 7157
rect 27252 7191 27304 7200
rect 27252 7157 27261 7191
rect 27261 7157 27295 7191
rect 27295 7157 27304 7191
rect 27252 7148 27304 7157
rect 5582 7046 5634 7098
rect 5646 7046 5698 7098
rect 5710 7046 5762 7098
rect 5774 7046 5826 7098
rect 5838 7046 5890 7098
rect 14846 7046 14898 7098
rect 14910 7046 14962 7098
rect 14974 7046 15026 7098
rect 15038 7046 15090 7098
rect 15102 7046 15154 7098
rect 24110 7046 24162 7098
rect 24174 7046 24226 7098
rect 24238 7046 24290 7098
rect 24302 7046 24354 7098
rect 24366 7046 24418 7098
rect 2596 6672 2648 6724
rect 2872 6851 2924 6860
rect 2872 6817 2881 6851
rect 2881 6817 2915 6851
rect 2915 6817 2924 6851
rect 2872 6808 2924 6817
rect 27252 6808 27304 6860
rect 28172 6851 28224 6860
rect 28172 6817 28181 6851
rect 28181 6817 28215 6851
rect 28215 6817 28224 6851
rect 28172 6808 28224 6817
rect 14004 6740 14056 6792
rect 27896 6672 27948 6724
rect 3608 6604 3660 6656
rect 10214 6502 10266 6554
rect 10278 6502 10330 6554
rect 10342 6502 10394 6554
rect 10406 6502 10458 6554
rect 10470 6502 10522 6554
rect 19478 6502 19530 6554
rect 19542 6502 19594 6554
rect 19606 6502 19658 6554
rect 19670 6502 19722 6554
rect 19734 6502 19786 6554
rect 1768 6400 1820 6452
rect 2596 6443 2648 6452
rect 2596 6409 2605 6443
rect 2605 6409 2639 6443
rect 2639 6409 2648 6443
rect 2596 6400 2648 6409
rect 4712 6400 4764 6452
rect 27896 6443 27948 6452
rect 27896 6409 27905 6443
rect 27905 6409 27939 6443
rect 27939 6409 27948 6443
rect 27896 6400 27948 6409
rect 3608 6375 3660 6384
rect 3608 6341 3617 6375
rect 3617 6341 3651 6375
rect 3651 6341 3660 6375
rect 3608 6332 3660 6341
rect 4160 6332 4212 6384
rect 2596 6264 2648 6316
rect 4436 6196 4488 6248
rect 4528 6239 4580 6248
rect 4528 6205 4537 6239
rect 4537 6205 4571 6239
rect 4571 6205 4580 6239
rect 24584 6239 24636 6248
rect 4528 6196 4580 6205
rect 24584 6205 24593 6239
rect 24593 6205 24627 6239
rect 24627 6205 24636 6239
rect 24584 6196 24636 6205
rect 24952 6196 25004 6248
rect 26056 6239 26108 6248
rect 26056 6205 26065 6239
rect 26065 6205 26099 6239
rect 26099 6205 26108 6239
rect 26056 6196 26108 6205
rect 2688 6128 2740 6180
rect 8668 6128 8720 6180
rect 27804 6128 27856 6180
rect 26516 6060 26568 6112
rect 5582 5958 5634 6010
rect 5646 5958 5698 6010
rect 5710 5958 5762 6010
rect 5774 5958 5826 6010
rect 5838 5958 5890 6010
rect 14846 5958 14898 6010
rect 14910 5958 14962 6010
rect 14974 5958 15026 6010
rect 15038 5958 15090 6010
rect 15102 5958 15154 6010
rect 24110 5958 24162 6010
rect 24174 5958 24226 6010
rect 24238 5958 24290 6010
rect 24302 5958 24354 6010
rect 24366 5958 24418 6010
rect 24584 5856 24636 5908
rect 1860 5763 1912 5772
rect 1860 5729 1869 5763
rect 1869 5729 1903 5763
rect 1903 5729 1912 5763
rect 1860 5720 1912 5729
rect 5356 5720 5408 5772
rect 27620 5788 27672 5840
rect 26516 5763 26568 5772
rect 26516 5729 26525 5763
rect 26525 5729 26559 5763
rect 26559 5729 26568 5763
rect 26516 5720 26568 5729
rect 28172 5763 28224 5772
rect 28172 5729 28181 5763
rect 28181 5729 28215 5763
rect 28215 5729 28224 5763
rect 28172 5720 28224 5729
rect 4160 5652 4212 5704
rect 4620 5695 4672 5704
rect 4620 5661 4629 5695
rect 4629 5661 4663 5695
rect 4663 5661 4672 5695
rect 4620 5652 4672 5661
rect 6368 5652 6420 5704
rect 6552 5695 6604 5704
rect 6552 5661 6561 5695
rect 6561 5661 6595 5695
rect 6595 5661 6604 5695
rect 6552 5652 6604 5661
rect 24860 5652 24912 5704
rect 1584 5627 1636 5636
rect 1584 5593 1593 5627
rect 1593 5593 1627 5627
rect 1627 5593 1636 5627
rect 1584 5584 1636 5593
rect 3884 5559 3936 5568
rect 3884 5525 3893 5559
rect 3893 5525 3927 5559
rect 3927 5525 3936 5559
rect 3884 5516 3936 5525
rect 10214 5414 10266 5466
rect 10278 5414 10330 5466
rect 10342 5414 10394 5466
rect 10406 5414 10458 5466
rect 10470 5414 10522 5466
rect 19478 5414 19530 5466
rect 19542 5414 19594 5466
rect 19606 5414 19658 5466
rect 19670 5414 19722 5466
rect 19734 5414 19786 5466
rect 1584 5312 1636 5364
rect 1676 5176 1728 5228
rect 6552 5312 6604 5364
rect 24952 5312 25004 5364
rect 3884 5244 3936 5296
rect 27160 5219 27212 5228
rect 27160 5185 27169 5219
rect 27169 5185 27203 5219
rect 27203 5185 27212 5219
rect 27160 5176 27212 5185
rect 27988 5176 28040 5228
rect 2780 5151 2832 5160
rect 2780 5117 2789 5151
rect 2789 5117 2823 5151
rect 2823 5117 2832 5151
rect 2780 5108 2832 5117
rect 24860 5108 24912 5160
rect 26148 5151 26200 5160
rect 26148 5117 26157 5151
rect 26157 5117 26191 5151
rect 26191 5117 26200 5151
rect 26148 5108 26200 5117
rect 2320 5040 2372 5092
rect 4436 5040 4488 5092
rect 5080 5040 5132 5092
rect 17132 5040 17184 5092
rect 17592 5040 17644 5092
rect 27712 5040 27764 5092
rect 4252 4972 4304 5024
rect 5172 5015 5224 5024
rect 5172 4981 5181 5015
rect 5181 4981 5215 5015
rect 5215 4981 5224 5015
rect 5172 4972 5224 4981
rect 5908 4972 5960 5024
rect 7196 5015 7248 5024
rect 7196 4981 7205 5015
rect 7205 4981 7239 5015
rect 7239 4981 7248 5015
rect 7196 4972 7248 4981
rect 5582 4870 5634 4922
rect 5646 4870 5698 4922
rect 5710 4870 5762 4922
rect 5774 4870 5826 4922
rect 5838 4870 5890 4922
rect 14846 4870 14898 4922
rect 14910 4870 14962 4922
rect 14974 4870 15026 4922
rect 15038 4870 15090 4922
rect 15102 4870 15154 4922
rect 24110 4870 24162 4922
rect 24174 4870 24226 4922
rect 24238 4870 24290 4922
rect 24302 4870 24354 4922
rect 24366 4870 24418 4922
rect 7196 4632 7248 4684
rect 2412 4607 2464 4616
rect 2412 4573 2421 4607
rect 2421 4573 2455 4607
rect 2455 4573 2464 4607
rect 2412 4564 2464 4573
rect 3056 4607 3108 4616
rect 3056 4573 3065 4607
rect 3065 4573 3099 4607
rect 3099 4573 3108 4607
rect 3056 4564 3108 4573
rect 6276 4607 6328 4616
rect 6276 4573 6285 4607
rect 6285 4573 6319 4607
rect 6319 4573 6328 4607
rect 6276 4564 6328 4573
rect 7288 4607 7340 4616
rect 7288 4573 7297 4607
rect 7297 4573 7331 4607
rect 7331 4573 7340 4607
rect 17132 4632 17184 4684
rect 8116 4607 8168 4616
rect 7288 4564 7340 4573
rect 8116 4573 8125 4607
rect 8125 4573 8159 4607
rect 8159 4573 8168 4607
rect 8116 4564 8168 4573
rect 9036 4564 9088 4616
rect 23848 4607 23900 4616
rect 23848 4573 23857 4607
rect 23857 4573 23891 4607
rect 23891 4573 23900 4607
rect 23848 4564 23900 4573
rect 4344 4496 4396 4548
rect 24860 4539 24912 4548
rect 24860 4505 24869 4539
rect 24869 4505 24903 4539
rect 24903 4505 24912 4539
rect 24860 4496 24912 4505
rect 27712 4496 27764 4548
rect 28356 4496 28408 4548
rect 1584 4428 1636 4480
rect 2504 4471 2556 4480
rect 2504 4437 2513 4471
rect 2513 4437 2547 4471
rect 2547 4437 2556 4471
rect 2504 4428 2556 4437
rect 7380 4471 7432 4480
rect 7380 4437 7389 4471
rect 7389 4437 7423 4471
rect 7423 4437 7432 4471
rect 7380 4428 7432 4437
rect 24952 4471 25004 4480
rect 24952 4437 24961 4471
rect 24961 4437 24995 4471
rect 24995 4437 25004 4471
rect 24952 4428 25004 4437
rect 10214 4326 10266 4378
rect 10278 4326 10330 4378
rect 10342 4326 10394 4378
rect 10406 4326 10458 4378
rect 10470 4326 10522 4378
rect 19478 4326 19530 4378
rect 19542 4326 19594 4378
rect 19606 4326 19658 4378
rect 19670 4326 19722 4378
rect 19734 4326 19786 4378
rect 2412 4224 2464 4276
rect 1584 4199 1636 4208
rect 1584 4165 1593 4199
rect 1593 4165 1627 4199
rect 1627 4165 1636 4199
rect 1584 4156 1636 4165
rect 1400 4131 1452 4140
rect 1400 4097 1409 4131
rect 1409 4097 1443 4131
rect 1443 4097 1452 4131
rect 1400 4088 1452 4097
rect 5080 4156 5132 4208
rect 7380 4199 7432 4208
rect 7380 4165 7389 4199
rect 7389 4165 7423 4199
rect 7423 4165 7432 4199
rect 7380 4156 7432 4165
rect 12900 4088 12952 4140
rect 24860 4088 24912 4140
rect 27160 4131 27212 4140
rect 27160 4097 27169 4131
rect 27169 4097 27203 4131
rect 27203 4097 27212 4131
rect 27160 4088 27212 4097
rect 28264 4088 28316 4140
rect 664 4020 716 4072
rect 4160 4063 4212 4072
rect 4160 4029 4169 4063
rect 4169 4029 4203 4063
rect 4203 4029 4212 4063
rect 4160 4020 4212 4029
rect 8116 4020 8168 4072
rect 1400 3884 1452 3936
rect 5172 3884 5224 3936
rect 6920 3884 6972 3936
rect 7748 3952 7800 4004
rect 12532 4020 12584 4072
rect 13176 4063 13228 4072
rect 13176 4029 13185 4063
rect 13185 4029 13219 4063
rect 13219 4029 13228 4063
rect 13176 4020 13228 4029
rect 13544 4063 13596 4072
rect 13544 4029 13553 4063
rect 13553 4029 13587 4063
rect 13587 4029 13596 4063
rect 13544 4020 13596 4029
rect 17684 4063 17736 4072
rect 17408 3952 17460 4004
rect 17684 4029 17693 4063
rect 17693 4029 17727 4063
rect 17727 4029 17736 4063
rect 17684 4020 17736 4029
rect 18052 4063 18104 4072
rect 18052 4029 18061 4063
rect 18061 4029 18095 4063
rect 18095 4029 18104 4063
rect 18052 4020 18104 4029
rect 23480 4063 23532 4072
rect 23480 4029 23489 4063
rect 23489 4029 23523 4063
rect 23523 4029 23532 4063
rect 23480 4020 23532 4029
rect 17960 3952 18012 4004
rect 23112 3952 23164 4004
rect 29000 3952 29052 4004
rect 9312 3884 9364 3936
rect 10324 3927 10376 3936
rect 10324 3893 10333 3927
rect 10333 3893 10367 3927
rect 10367 3893 10376 3927
rect 10324 3884 10376 3893
rect 15660 3884 15712 3936
rect 22192 3884 22244 3936
rect 25136 3884 25188 3936
rect 5582 3782 5634 3834
rect 5646 3782 5698 3834
rect 5710 3782 5762 3834
rect 5774 3782 5826 3834
rect 5838 3782 5890 3834
rect 14846 3782 14898 3834
rect 14910 3782 14962 3834
rect 14974 3782 15026 3834
rect 15038 3782 15090 3834
rect 15102 3782 15154 3834
rect 24110 3782 24162 3834
rect 24174 3782 24226 3834
rect 24238 3782 24290 3834
rect 24302 3782 24354 3834
rect 24366 3782 24418 3834
rect 5908 3680 5960 3732
rect 3332 3612 3384 3664
rect 4344 3612 4396 3664
rect 12348 3680 12400 3732
rect 12532 3723 12584 3732
rect 12532 3689 12541 3723
rect 12541 3689 12575 3723
rect 12575 3689 12584 3723
rect 12532 3680 12584 3689
rect 13176 3680 13228 3732
rect 17408 3680 17460 3732
rect 23112 3723 23164 3732
rect 23112 3689 23121 3723
rect 23121 3689 23155 3723
rect 23155 3689 23164 3723
rect 23112 3680 23164 3689
rect 23480 3680 23532 3732
rect 3056 3476 3108 3528
rect 5356 3587 5408 3596
rect 5356 3553 5365 3587
rect 5365 3553 5399 3587
rect 5399 3553 5408 3587
rect 5356 3544 5408 3553
rect 5908 3587 5960 3596
rect 5908 3553 5917 3587
rect 5917 3553 5951 3587
rect 5951 3553 5960 3587
rect 5908 3544 5960 3553
rect 10324 3612 10376 3664
rect 12900 3612 12952 3664
rect 16672 3612 16724 3664
rect 19984 3612 20036 3664
rect 24860 3612 24912 3664
rect 9312 3587 9364 3596
rect 9312 3553 9321 3587
rect 9321 3553 9355 3587
rect 9355 3553 9364 3587
rect 9312 3544 9364 3553
rect 9680 3587 9732 3596
rect 9680 3553 9689 3587
rect 9689 3553 9723 3587
rect 9723 3553 9732 3587
rect 9680 3544 9732 3553
rect 15660 3587 15712 3596
rect 15660 3553 15669 3587
rect 15669 3553 15703 3587
rect 15703 3553 15712 3587
rect 15660 3544 15712 3553
rect 16120 3587 16172 3596
rect 16120 3553 16129 3587
rect 16129 3553 16163 3587
rect 16163 3553 16172 3587
rect 16120 3544 16172 3553
rect 7656 3519 7708 3528
rect 3240 3451 3292 3460
rect 3240 3417 3249 3451
rect 3249 3417 3283 3451
rect 3283 3417 3292 3451
rect 3240 3408 3292 3417
rect 3884 3408 3936 3460
rect 4528 3408 4580 3460
rect 2228 3340 2280 3392
rect 7656 3485 7665 3519
rect 7665 3485 7699 3519
rect 7699 3485 7708 3519
rect 7656 3476 7708 3485
rect 11704 3476 11756 3528
rect 12992 3519 13044 3528
rect 12992 3485 13001 3519
rect 13001 3485 13035 3519
rect 13035 3485 13044 3519
rect 12992 3476 13044 3485
rect 14188 3476 14240 3528
rect 18880 3476 18932 3528
rect 20720 3544 20772 3596
rect 25136 3587 25188 3596
rect 19984 3519 20036 3528
rect 5540 3451 5592 3460
rect 5540 3417 5549 3451
rect 5549 3417 5583 3451
rect 5583 3417 5592 3451
rect 5540 3408 5592 3417
rect 15660 3408 15712 3460
rect 15844 3451 15896 3460
rect 15844 3417 15853 3451
rect 15853 3417 15887 3451
rect 15887 3417 15896 3451
rect 15844 3408 15896 3417
rect 18236 3408 18288 3460
rect 19984 3485 19993 3519
rect 19993 3485 20027 3519
rect 20027 3485 20036 3519
rect 19984 3476 20036 3485
rect 20168 3476 20220 3528
rect 21916 3476 21968 3528
rect 25136 3553 25145 3587
rect 25145 3553 25179 3587
rect 25179 3553 25188 3587
rect 25136 3544 25188 3553
rect 26148 3587 26200 3596
rect 26148 3553 26157 3587
rect 26157 3553 26191 3587
rect 26191 3553 26200 3587
rect 26148 3544 26200 3553
rect 23020 3519 23072 3528
rect 23020 3485 23029 3519
rect 23029 3485 23063 3519
rect 23063 3485 23072 3519
rect 23020 3476 23072 3485
rect 24952 3476 25004 3528
rect 27988 3476 28040 3528
rect 6552 3340 6604 3392
rect 7104 3340 7156 3392
rect 14096 3340 14148 3392
rect 20076 3383 20128 3392
rect 20076 3349 20085 3383
rect 20085 3349 20119 3383
rect 20119 3349 20128 3383
rect 20076 3340 20128 3349
rect 22100 3340 22152 3392
rect 23756 3340 23808 3392
rect 10214 3238 10266 3290
rect 10278 3238 10330 3290
rect 10342 3238 10394 3290
rect 10406 3238 10458 3290
rect 10470 3238 10522 3290
rect 19478 3238 19530 3290
rect 19542 3238 19594 3290
rect 19606 3238 19658 3290
rect 19670 3238 19722 3290
rect 19734 3238 19786 3290
rect 4252 3136 4304 3188
rect 5540 3136 5592 3188
rect 5632 3136 5684 3188
rect 27712 3179 27764 3188
rect 2504 3111 2556 3120
rect 2504 3077 2513 3111
rect 2513 3077 2547 3111
rect 2547 3077 2556 3111
rect 2504 3068 2556 3077
rect 2596 3068 2648 3120
rect 7104 3111 7156 3120
rect 4436 3000 4488 3052
rect 7104 3077 7113 3111
rect 7113 3077 7147 3111
rect 7147 3077 7156 3111
rect 7104 3068 7156 3077
rect 6920 3043 6972 3052
rect 2596 2932 2648 2984
rect 5632 2932 5684 2984
rect 3056 2864 3108 2916
rect 6920 3009 6929 3043
rect 6929 3009 6963 3043
rect 6963 3009 6972 3043
rect 6920 3000 6972 3009
rect 7380 2975 7432 2984
rect 7380 2941 7389 2975
rect 7389 2941 7423 2975
rect 7423 2941 7432 2975
rect 7380 2932 7432 2941
rect 14096 3068 14148 3120
rect 17684 3111 17736 3120
rect 17684 3077 17693 3111
rect 17693 3077 17727 3111
rect 17727 3077 17736 3111
rect 17684 3068 17736 3077
rect 22100 3111 22152 3120
rect 22100 3077 22109 3111
rect 22109 3077 22143 3111
rect 22143 3077 22152 3111
rect 22100 3068 22152 3077
rect 9772 3000 9824 3052
rect 11704 3043 11756 3052
rect 11704 3009 11713 3043
rect 11713 3009 11747 3043
rect 11747 3009 11756 3043
rect 11704 3000 11756 3009
rect 14188 3043 14240 3052
rect 14188 3009 14197 3043
rect 14197 3009 14231 3043
rect 14231 3009 14240 3043
rect 14188 3000 14240 3009
rect 11888 2975 11940 2984
rect 11888 2941 11897 2975
rect 11897 2941 11931 2975
rect 11931 2941 11940 2975
rect 11888 2932 11940 2941
rect 12256 2975 12308 2984
rect 12256 2941 12265 2975
rect 12265 2941 12299 2975
rect 12299 2941 12308 2975
rect 12256 2932 12308 2941
rect 14372 2975 14424 2984
rect 14372 2941 14381 2975
rect 14381 2941 14415 2975
rect 14415 2941 14424 2975
rect 14372 2932 14424 2941
rect 14740 2975 14792 2984
rect 14740 2941 14749 2975
rect 14749 2941 14783 2975
rect 14783 2941 14792 2975
rect 14740 2932 14792 2941
rect 8668 2864 8720 2916
rect 18236 3043 18288 3052
rect 1584 2796 1636 2848
rect 4160 2796 4212 2848
rect 9772 2839 9824 2848
rect 9772 2805 9781 2839
rect 9781 2805 9815 2839
rect 9815 2805 9824 2839
rect 9772 2796 9824 2805
rect 18236 3009 18245 3043
rect 18245 3009 18279 3043
rect 18279 3009 18288 3043
rect 18236 3000 18288 3009
rect 18880 3043 18932 3052
rect 18880 3009 18889 3043
rect 18889 3009 18923 3043
rect 18923 3009 18932 3043
rect 18880 3000 18932 3009
rect 21916 3043 21968 3052
rect 21916 3009 21925 3043
rect 21925 3009 21959 3043
rect 21959 3009 21968 3043
rect 21916 3000 21968 3009
rect 26056 3000 26108 3052
rect 19340 2975 19392 2984
rect 19340 2941 19349 2975
rect 19349 2941 19383 2975
rect 19383 2941 19392 2975
rect 19340 2932 19392 2941
rect 22560 2975 22612 2984
rect 22560 2941 22569 2975
rect 22569 2941 22603 2975
rect 22603 2941 22612 2975
rect 22560 2932 22612 2941
rect 24584 2975 24636 2984
rect 24584 2941 24593 2975
rect 24593 2941 24627 2975
rect 24627 2941 24636 2975
rect 24584 2932 24636 2941
rect 24768 2864 24820 2916
rect 25228 2864 25280 2916
rect 25504 2932 25556 2984
rect 26516 2932 26568 2984
rect 27712 3145 27721 3179
rect 27721 3145 27755 3179
rect 27755 3145 27764 3179
rect 27712 3136 27764 3145
rect 27804 3000 27856 3052
rect 25044 2796 25096 2848
rect 29644 2796 29696 2848
rect 5582 2694 5634 2746
rect 5646 2694 5698 2746
rect 5710 2694 5762 2746
rect 5774 2694 5826 2746
rect 5838 2694 5890 2746
rect 14846 2694 14898 2746
rect 14910 2694 14962 2746
rect 14974 2694 15026 2746
rect 15038 2694 15090 2746
rect 15102 2694 15154 2746
rect 24110 2694 24162 2746
rect 24174 2694 24226 2746
rect 24238 2694 24290 2746
rect 24302 2694 24354 2746
rect 24366 2694 24418 2746
rect 6276 2592 6328 2644
rect 11888 2592 11940 2644
rect 14372 2592 14424 2644
rect 15844 2635 15896 2644
rect 15844 2601 15853 2635
rect 15853 2601 15887 2635
rect 15887 2601 15896 2635
rect 15844 2592 15896 2601
rect 16304 2592 16356 2644
rect 17960 2635 18012 2644
rect 17960 2601 17969 2635
rect 17969 2601 18003 2635
rect 18003 2601 18012 2635
rect 17960 2592 18012 2601
rect 1584 2499 1636 2508
rect 1584 2465 1593 2499
rect 1593 2465 1627 2499
rect 1627 2465 1636 2499
rect 1584 2456 1636 2465
rect 2780 2499 2832 2508
rect 2780 2465 2789 2499
rect 2789 2465 2823 2499
rect 2823 2465 2832 2499
rect 2780 2456 2832 2465
rect 4620 2524 4672 2576
rect 5172 2524 5224 2576
rect 4160 2499 4212 2508
rect 4160 2465 4169 2499
rect 4169 2465 4203 2499
rect 4203 2465 4212 2499
rect 4160 2456 4212 2465
rect 4528 2499 4580 2508
rect 4528 2465 4537 2499
rect 4537 2465 4571 2499
rect 4571 2465 4580 2499
rect 4528 2456 4580 2465
rect 6368 2499 6420 2508
rect 6368 2465 6377 2499
rect 6377 2465 6411 2499
rect 6411 2465 6420 2499
rect 6368 2456 6420 2465
rect 6552 2499 6604 2508
rect 6552 2465 6561 2499
rect 6561 2465 6595 2499
rect 6595 2465 6604 2499
rect 6552 2456 6604 2465
rect 9128 2524 9180 2576
rect 9036 2499 9088 2508
rect 9036 2465 9045 2499
rect 9045 2465 9079 2499
rect 9079 2465 9088 2499
rect 9036 2456 9088 2465
rect 9772 2456 9824 2508
rect 12440 2388 12492 2440
rect 14096 2388 14148 2440
rect 15660 2388 15712 2440
rect 18696 2524 18748 2576
rect 26516 2592 26568 2644
rect 20076 2456 20128 2508
rect 27068 2524 27120 2576
rect 22192 2456 22244 2508
rect 23848 2456 23900 2508
rect 16764 2320 16816 2372
rect 27988 2388 28040 2440
rect 20168 2320 20220 2372
rect 23756 2320 23808 2372
rect 25044 2320 25096 2372
rect 26148 2320 26200 2372
rect 10214 2150 10266 2202
rect 10278 2150 10330 2202
rect 10342 2150 10394 2202
rect 10406 2150 10458 2202
rect 10470 2150 10522 2202
rect 19478 2150 19530 2202
rect 19542 2150 19594 2202
rect 19606 2150 19658 2202
rect 19670 2150 19722 2202
rect 19734 2150 19786 2202
rect 3056 1776 3108 1828
rect 7380 1776 7432 1828
<< metal2 >>
rect -10 41200 102 42000
rect 634 41200 746 42000
rect 1278 41200 1390 42000
rect 1922 41200 2034 42000
rect 2566 41200 2678 42000
rect 3210 41200 3322 42000
rect 3854 41200 3966 42000
rect 4498 41200 4610 42000
rect 5142 41200 5254 42000
rect 5786 41200 5898 42000
rect 7074 41200 7186 42000
rect 7718 41200 7830 42000
rect 8362 41200 8474 42000
rect 9006 41200 9118 42000
rect 9650 41200 9762 42000
rect 10294 41200 10406 42000
rect 10938 41200 11050 42000
rect 11582 41200 11694 42000
rect 12226 41200 12338 42000
rect 12870 41200 12982 42000
rect 13514 41200 13626 42000
rect 14158 41200 14270 42000
rect 14802 41200 14914 42000
rect 15446 41200 15558 42000
rect 16090 41200 16202 42000
rect 16734 41200 16846 42000
rect 17378 41200 17490 42000
rect 18022 41200 18134 42000
rect 18666 41200 18778 42000
rect 19310 41200 19422 42000
rect 19954 41200 20066 42000
rect 20598 41200 20710 42000
rect 21242 41200 21354 42000
rect 21886 41200 21998 42000
rect 22530 41200 22642 42000
rect 23174 41200 23286 42000
rect 23818 41200 23930 42000
rect 24462 41200 24574 42000
rect 25106 41200 25218 42000
rect 25750 41200 25862 42000
rect 26394 41200 26506 42000
rect 27038 41200 27150 42000
rect 27682 41200 27794 42000
rect 28326 41200 28438 42000
rect 28970 41200 29082 42000
rect 29614 41200 29726 42000
rect 32 38554 60 41200
rect 1766 39536 1822 39545
rect 1766 39471 1822 39480
rect 1780 39438 1808 39471
rect 1768 39432 1820 39438
rect 1768 39374 1820 39380
rect 1676 39296 1728 39302
rect 1676 39238 1728 39244
rect 1688 39030 1716 39238
rect 1676 39024 1728 39030
rect 1676 38966 1728 38972
rect 1492 38888 1544 38894
rect 1492 38830 1544 38836
rect 20 38548 72 38554
rect 20 38490 72 38496
rect 1400 38548 1452 38554
rect 1400 38490 1452 38496
rect 1412 35894 1440 38490
rect 1504 36378 1532 38830
rect 1676 38820 1728 38826
rect 1676 38762 1728 38768
rect 1584 37188 1636 37194
rect 1584 37130 1636 37136
rect 1596 36922 1624 37130
rect 1584 36916 1636 36922
rect 1584 36858 1636 36864
rect 1584 36780 1636 36786
rect 1584 36722 1636 36728
rect 1492 36372 1544 36378
rect 1492 36314 1544 36320
rect 1596 36242 1624 36722
rect 1584 36236 1636 36242
rect 1584 36178 1636 36184
rect 1412 35866 1532 35894
rect 1400 34400 1452 34406
rect 1400 34342 1452 34348
rect 1412 34066 1440 34342
rect 1400 34060 1452 34066
rect 1400 34002 1452 34008
rect 1400 33516 1452 33522
rect 1400 33458 1452 33464
rect 1412 33425 1440 33458
rect 1398 33416 1454 33425
rect 1398 33351 1454 33360
rect 1504 32910 1532 35866
rect 1492 32904 1544 32910
rect 1492 32846 1544 32852
rect 1688 32450 1716 38762
rect 1964 38282 1992 41200
rect 2778 40216 2834 40225
rect 2778 40151 2834 40160
rect 2412 39432 2464 39438
rect 2412 39374 2464 39380
rect 2424 38826 2452 39374
rect 2504 39296 2556 39302
rect 2504 39238 2556 39244
rect 2412 38820 2464 38826
rect 2412 38762 2464 38768
rect 2516 38418 2544 39238
rect 2792 38418 2820 40151
rect 2870 39400 2926 39409
rect 2870 39335 2926 39344
rect 2884 38894 2912 39335
rect 3148 39296 3200 39302
rect 3148 39238 3200 39244
rect 3160 39030 3188 39238
rect 3148 39024 3200 39030
rect 3148 38966 3200 38972
rect 2872 38888 2924 38894
rect 2872 38830 2924 38836
rect 3252 38554 3280 41200
rect 3896 39488 3924 41200
rect 4160 39500 4212 39506
rect 3896 39460 4160 39488
rect 4160 39442 4212 39448
rect 3976 39364 4028 39370
rect 3976 39306 4028 39312
rect 3240 38548 3292 38554
rect 3240 38490 3292 38496
rect 2504 38412 2556 38418
rect 2504 38354 2556 38360
rect 2780 38412 2832 38418
rect 2780 38354 2832 38360
rect 1952 38276 2004 38282
rect 1952 38218 2004 38224
rect 2872 38276 2924 38282
rect 2872 38218 2924 38224
rect 2778 38176 2834 38185
rect 2778 38111 2834 38120
rect 2792 37806 2820 38111
rect 2780 37800 2832 37806
rect 2780 37742 2832 37748
rect 1858 37496 1914 37505
rect 1858 37431 1914 37440
rect 1872 37330 1900 37431
rect 1860 37324 1912 37330
rect 1860 37266 1912 37272
rect 2596 36916 2648 36922
rect 2596 36858 2648 36864
rect 2044 36644 2096 36650
rect 2044 36586 2096 36592
rect 1768 35624 1820 35630
rect 1768 35566 1820 35572
rect 1780 35290 1808 35566
rect 1768 35284 1820 35290
rect 1768 35226 1820 35232
rect 1860 34944 1912 34950
rect 1860 34886 1912 34892
rect 1872 34678 1900 34886
rect 1860 34672 1912 34678
rect 1860 34614 1912 34620
rect 2056 33658 2084 36586
rect 2608 36174 2636 36858
rect 2596 36168 2648 36174
rect 2596 36110 2648 36116
rect 2884 35630 2912 38218
rect 3792 37936 3844 37942
rect 3792 37878 3844 37884
rect 3700 36712 3752 36718
rect 3700 36654 3752 36660
rect 3712 36174 3740 36654
rect 3700 36168 3752 36174
rect 3700 36110 3752 36116
rect 2872 35624 2924 35630
rect 2872 35566 2924 35572
rect 3424 35488 3476 35494
rect 3424 35430 3476 35436
rect 2412 35080 2464 35086
rect 2412 35022 2464 35028
rect 3240 35080 3292 35086
rect 3240 35022 3292 35028
rect 2136 35012 2188 35018
rect 2136 34954 2188 34960
rect 2044 33652 2096 33658
rect 2044 33594 2096 33600
rect 1952 33516 2004 33522
rect 1952 33458 2004 33464
rect 1688 32422 1900 32450
rect 1492 32360 1544 32366
rect 1492 32302 1544 32308
rect 1768 32360 1820 32366
rect 1768 32302 1820 32308
rect 1504 32026 1532 32302
rect 1492 32020 1544 32026
rect 1492 31962 1544 31968
rect 1676 31816 1728 31822
rect 1676 31758 1728 31764
rect 1688 31346 1716 31758
rect 1676 31340 1728 31346
rect 1676 31282 1728 31288
rect 1400 29640 1452 29646
rect 1400 29582 1452 29588
rect 1412 29170 1440 29582
rect 1400 29164 1452 29170
rect 1400 29106 1452 29112
rect 1584 29096 1636 29102
rect 1584 29038 1636 29044
rect 1596 28762 1624 29038
rect 1584 28756 1636 28762
rect 1584 28698 1636 28704
rect 1676 28552 1728 28558
rect 1676 28494 1728 28500
rect 1492 23724 1544 23730
rect 1492 23666 1544 23672
rect 1400 15904 1452 15910
rect 1400 15846 1452 15852
rect 1412 15570 1440 15846
rect 1400 15564 1452 15570
rect 1400 15506 1452 15512
rect 1504 15026 1532 23666
rect 1584 17128 1636 17134
rect 1584 17070 1636 17076
rect 1596 16794 1624 17070
rect 1584 16788 1636 16794
rect 1584 16730 1636 16736
rect 1688 16600 1716 28494
rect 1676 16594 1728 16600
rect 1676 16536 1728 16542
rect 1584 15428 1636 15434
rect 1584 15370 1636 15376
rect 1596 15162 1624 15370
rect 1584 15156 1636 15162
rect 1584 15098 1636 15104
rect 1492 15020 1544 15026
rect 1492 14962 1544 14968
rect 1400 14816 1452 14822
rect 1400 14758 1452 14764
rect 1412 14482 1440 14758
rect 1400 14476 1452 14482
rect 1400 14418 1452 14424
rect 1504 13326 1532 14962
rect 1584 14340 1636 14346
rect 1584 14282 1636 14288
rect 1596 14074 1624 14282
rect 1584 14068 1636 14074
rect 1584 14010 1636 14016
rect 1492 13320 1544 13326
rect 1492 13262 1544 13268
rect 1400 13252 1452 13258
rect 1400 13194 1452 13200
rect 1412 12850 1440 13194
rect 1400 12844 1452 12850
rect 1400 12786 1452 12792
rect 1504 9586 1532 13262
rect 1584 13184 1636 13190
rect 1584 13126 1636 13132
rect 1596 12918 1624 13126
rect 1584 12912 1636 12918
rect 1584 12854 1636 12860
rect 1584 11552 1636 11558
rect 1584 11494 1636 11500
rect 1596 11218 1624 11494
rect 1584 11212 1636 11218
rect 1584 11154 1636 11160
rect 1492 9580 1544 9586
rect 1492 9522 1544 9528
rect 1584 9376 1636 9382
rect 1584 9318 1636 9324
rect 1596 9042 1624 9318
rect 1584 9036 1636 9042
rect 1584 8978 1636 8984
rect 1584 8288 1636 8294
rect 1584 8230 1636 8236
rect 1596 7954 1624 8230
rect 1584 7948 1636 7954
rect 1584 7890 1636 7896
rect 1584 5636 1636 5642
rect 1584 5578 1636 5584
rect 1596 5370 1624 5578
rect 1584 5364 1636 5370
rect 1584 5306 1636 5312
rect 1688 5234 1716 16536
rect 1780 6458 1808 32302
rect 1872 21434 1900 32422
rect 1964 23610 1992 33458
rect 2148 26234 2176 34954
rect 2228 33924 2280 33930
rect 2228 33866 2280 33872
rect 2240 33658 2268 33866
rect 2228 33652 2280 33658
rect 2228 33594 2280 33600
rect 2228 31748 2280 31754
rect 2228 31690 2280 31696
rect 2240 30734 2268 31690
rect 2320 31272 2372 31278
rect 2320 31214 2372 31220
rect 2332 30938 2360 31214
rect 2320 30932 2372 30938
rect 2320 30874 2372 30880
rect 2228 30728 2280 30734
rect 2228 30670 2280 30676
rect 2056 26206 2176 26234
rect 2056 23730 2084 26206
rect 2044 23724 2096 23730
rect 2044 23666 2096 23672
rect 1964 23582 2084 23610
rect 1952 23520 2004 23526
rect 1952 23462 2004 23468
rect 1964 23186 1992 23462
rect 1952 23180 2004 23186
rect 1952 23122 2004 23128
rect 1872 21406 1992 21434
rect 1860 18080 1912 18086
rect 1860 18022 1912 18028
rect 1872 17746 1900 18022
rect 1860 17740 1912 17746
rect 1860 17682 1912 17688
rect 1860 17128 1912 17134
rect 1858 17096 1860 17105
rect 1912 17096 1914 17105
rect 1858 17031 1914 17040
rect 1860 14476 1912 14482
rect 1860 14418 1912 14424
rect 1872 14385 1900 14418
rect 1858 14376 1914 14385
rect 1858 14311 1914 14320
rect 1860 13932 1912 13938
rect 1860 13874 1912 13880
rect 1872 11694 1900 13874
rect 1860 11688 1912 11694
rect 1860 11630 1912 11636
rect 1860 11212 1912 11218
rect 1860 11154 1912 11160
rect 1872 10985 1900 11154
rect 1858 10976 1914 10985
rect 1858 10911 1914 10920
rect 1964 10826 1992 21406
rect 1872 10798 1992 10826
rect 1872 8498 1900 10798
rect 1952 10600 2004 10606
rect 1952 10542 2004 10548
rect 1964 10266 1992 10542
rect 1952 10260 2004 10266
rect 1952 10202 2004 10208
rect 2056 10062 2084 23582
rect 2044 10056 2096 10062
rect 2044 9998 2096 10004
rect 1860 8492 1912 8498
rect 1860 8434 1912 8440
rect 2136 8288 2188 8294
rect 2136 8230 2188 8236
rect 1952 7812 2004 7818
rect 1952 7754 2004 7760
rect 1964 7410 1992 7754
rect 2148 7478 2176 8230
rect 2136 7472 2188 7478
rect 2136 7414 2188 7420
rect 1952 7404 2004 7410
rect 1952 7346 2004 7352
rect 1768 6452 1820 6458
rect 1768 6394 1820 6400
rect 1860 5772 1912 5778
rect 1860 5714 1912 5720
rect 1872 5545 1900 5714
rect 1858 5536 1914 5545
rect 1858 5471 1914 5480
rect 1676 5228 1728 5234
rect 1676 5170 1728 5176
rect 1584 4480 1636 4486
rect 1584 4422 1636 4428
rect 1596 4214 1624 4422
rect 1584 4208 1636 4214
rect 1584 4150 1636 4156
rect 1400 4140 1452 4146
rect 1400 4082 1452 4088
rect 664 4072 716 4078
rect 664 4014 716 4020
rect 676 800 704 4014
rect 1412 3942 1440 4082
rect 1400 3936 1452 3942
rect 1400 3878 1452 3884
rect 2240 3398 2268 30670
rect 2424 26234 2452 35022
rect 2778 34776 2834 34785
rect 3252 34746 3280 35022
rect 2778 34711 2834 34720
rect 3240 34740 3292 34746
rect 2792 34542 2820 34711
rect 3240 34682 3292 34688
rect 2780 34536 2832 34542
rect 2780 34478 2832 34484
rect 2778 34096 2834 34105
rect 2778 34031 2780 34040
rect 2832 34031 2834 34040
rect 2780 34002 2832 34008
rect 3436 33114 3464 35430
rect 3424 33108 3476 33114
rect 3424 33050 3476 33056
rect 2870 32736 2926 32745
rect 2870 32671 2926 32680
rect 2884 32366 2912 32671
rect 2872 32360 2924 32366
rect 2872 32302 2924 32308
rect 2778 31376 2834 31385
rect 2778 31311 2834 31320
rect 2792 31278 2820 31311
rect 2780 31272 2832 31278
rect 2780 31214 2832 31220
rect 2778 29336 2834 29345
rect 2778 29271 2834 29280
rect 2792 29102 2820 29271
rect 2780 29096 2832 29102
rect 2780 29038 2832 29044
rect 2332 26206 2452 26234
rect 2332 5098 2360 26206
rect 2778 23216 2834 23225
rect 2778 23151 2780 23160
rect 2832 23151 2834 23160
rect 2780 23122 2832 23128
rect 2504 23044 2556 23050
rect 2504 22986 2556 22992
rect 2516 22778 2544 22986
rect 2504 22772 2556 22778
rect 2504 22714 2556 22720
rect 2596 22636 2648 22642
rect 2596 22578 2648 22584
rect 2412 18080 2464 18086
rect 2412 18022 2464 18028
rect 2424 17610 2452 18022
rect 2412 17604 2464 17610
rect 2412 17546 2464 17552
rect 2504 17060 2556 17066
rect 2504 17002 2556 17008
rect 2516 16794 2544 17002
rect 2504 16788 2556 16794
rect 2504 16730 2556 16736
rect 2608 16574 2636 22578
rect 2778 17776 2834 17785
rect 2778 17711 2780 17720
rect 2832 17711 2834 17720
rect 2780 17682 2832 17688
rect 2608 16546 2728 16574
rect 2412 13320 2464 13326
rect 2412 13262 2464 13268
rect 2424 12306 2452 13262
rect 2412 12300 2464 12306
rect 2412 12242 2464 12248
rect 2504 12164 2556 12170
rect 2504 12106 2556 12112
rect 2516 11898 2544 12106
rect 2504 11892 2556 11898
rect 2504 11834 2556 11840
rect 2412 9376 2464 9382
rect 2412 9318 2464 9324
rect 2424 9110 2452 9318
rect 2412 9104 2464 9110
rect 2412 9046 2464 9052
rect 2596 6724 2648 6730
rect 2596 6666 2648 6672
rect 2608 6458 2636 6666
rect 2596 6452 2648 6458
rect 2596 6394 2648 6400
rect 2596 6316 2648 6322
rect 2596 6258 2648 6264
rect 2320 5092 2372 5098
rect 2320 5034 2372 5040
rect 2412 4616 2464 4622
rect 2412 4558 2464 4564
rect 2424 4282 2452 4558
rect 2504 4480 2556 4486
rect 2504 4422 2556 4428
rect 2412 4276 2464 4282
rect 2412 4218 2464 4224
rect 2228 3392 2280 3398
rect 2228 3334 2280 3340
rect 2516 3126 2544 4422
rect 2608 3126 2636 6258
rect 2700 6186 2728 16546
rect 2778 15736 2834 15745
rect 2778 15671 2834 15680
rect 2792 15570 2820 15671
rect 2780 15564 2832 15570
rect 2780 15506 2832 15512
rect 2778 13016 2834 13025
rect 2778 12951 2834 12960
rect 2792 12782 2820 12951
rect 2780 12776 2832 12782
rect 2780 12718 2832 12724
rect 2778 12336 2834 12345
rect 2778 12271 2780 12280
rect 2832 12271 2834 12280
rect 2780 12242 2832 12248
rect 3712 11762 3740 36110
rect 3804 35834 3832 37878
rect 3884 37800 3936 37806
rect 3884 37742 3936 37748
rect 3896 37466 3924 37742
rect 3884 37460 3936 37466
rect 3884 37402 3936 37408
rect 3884 37120 3936 37126
rect 3884 37062 3936 37068
rect 3792 35828 3844 35834
rect 3792 35770 3844 35776
rect 3896 35290 3924 37062
rect 3988 36378 4016 39306
rect 4252 38344 4304 38350
rect 4252 38286 4304 38292
rect 4264 37194 4292 38286
rect 4540 37806 4568 41200
rect 4620 38888 4672 38894
rect 4620 38830 4672 38836
rect 4712 38888 4764 38894
rect 4712 38830 4764 38836
rect 4528 37800 4580 37806
rect 4528 37742 4580 37748
rect 4436 37732 4488 37738
rect 4436 37674 4488 37680
rect 4344 37256 4396 37262
rect 4344 37198 4396 37204
rect 4252 37188 4304 37194
rect 4252 37130 4304 37136
rect 4356 36786 4384 37198
rect 4344 36780 4396 36786
rect 4344 36722 4396 36728
rect 3976 36372 4028 36378
rect 3976 36314 4028 36320
rect 4066 36136 4122 36145
rect 4122 36094 4200 36122
rect 4066 36071 4122 36080
rect 3884 35284 3936 35290
rect 3884 35226 3936 35232
rect 4172 35086 4200 36094
rect 4448 35698 4476 37674
rect 4632 36378 4660 38830
rect 4724 38554 4752 38830
rect 4712 38548 4764 38554
rect 4712 38490 4764 38496
rect 5184 38418 5212 41200
rect 9036 40860 9088 40866
rect 9036 40802 9088 40808
rect 8852 40792 8904 40798
rect 8852 40734 8904 40740
rect 7564 40724 7616 40730
rect 7564 40666 7616 40672
rect 7472 40588 7524 40594
rect 7472 40530 7524 40536
rect 7380 40452 7432 40458
rect 7380 40394 7432 40400
rect 7196 40384 7248 40390
rect 7196 40326 7248 40332
rect 7102 39944 7158 39953
rect 7102 39879 7158 39888
rect 6644 39840 6696 39846
rect 6644 39782 6696 39788
rect 5582 39740 5890 39760
rect 5582 39738 5588 39740
rect 5644 39738 5668 39740
rect 5724 39738 5748 39740
rect 5804 39738 5828 39740
rect 5884 39738 5890 39740
rect 5644 39686 5646 39738
rect 5826 39686 5828 39738
rect 5582 39684 5588 39686
rect 5644 39684 5668 39686
rect 5724 39684 5748 39686
rect 5804 39684 5828 39686
rect 5884 39684 5890 39686
rect 5582 39664 5890 39684
rect 5448 39568 5500 39574
rect 5448 39510 5500 39516
rect 5264 39296 5316 39302
rect 5264 39238 5316 39244
rect 5172 38412 5224 38418
rect 5172 38354 5224 38360
rect 5172 38276 5224 38282
rect 5172 38218 5224 38224
rect 4712 37188 4764 37194
rect 4712 37130 4764 37136
rect 4620 36372 4672 36378
rect 4620 36314 4672 36320
rect 4436 35692 4488 35698
rect 4436 35634 4488 35640
rect 4528 35624 4580 35630
rect 4528 35566 4580 35572
rect 4540 35290 4568 35566
rect 4528 35284 4580 35290
rect 4528 35226 4580 35232
rect 4160 35080 4212 35086
rect 4160 35022 4212 35028
rect 3792 35012 3844 35018
rect 3792 34954 3844 34960
rect 3804 34746 3832 34954
rect 3792 34740 3844 34746
rect 3792 34682 3844 34688
rect 3882 30016 3938 30025
rect 3882 29951 3938 29960
rect 3896 29646 3924 29951
rect 3884 29640 3936 29646
rect 3884 29582 3936 29588
rect 3700 11756 3752 11762
rect 3700 11698 3752 11704
rect 3240 11552 3292 11558
rect 3240 11494 3292 11500
rect 3252 11286 3280 11494
rect 3240 11280 3292 11286
rect 3240 11222 3292 11228
rect 3976 11144 4028 11150
rect 3976 11086 4028 11092
rect 3988 10742 4016 11086
rect 3976 10736 4028 10742
rect 3976 10678 4028 10684
rect 2872 10600 2924 10606
rect 2872 10542 2924 10548
rect 2884 10305 2912 10542
rect 2870 10296 2926 10305
rect 2870 10231 2926 10240
rect 2780 9036 2832 9042
rect 2780 8978 2832 8984
rect 2792 8265 2820 8978
rect 3332 8288 3384 8294
rect 2778 8256 2834 8265
rect 3332 8230 3384 8236
rect 2778 8191 2834 8200
rect 3344 8022 3372 8230
rect 3332 8016 3384 8022
rect 3332 7958 3384 7964
rect 2780 7948 2832 7954
rect 2780 7890 2832 7896
rect 2792 7585 2820 7890
rect 2778 7576 2834 7585
rect 2778 7511 2834 7520
rect 2964 7336 3016 7342
rect 2964 7278 3016 7284
rect 2870 6896 2926 6905
rect 2870 6831 2872 6840
rect 2924 6831 2926 6840
rect 2872 6802 2924 6808
rect 2688 6180 2740 6186
rect 2688 6122 2740 6128
rect 2780 5160 2832 5166
rect 2780 5102 2832 5108
rect 2792 4865 2820 5102
rect 2778 4856 2834 4865
rect 2778 4791 2834 4800
rect 2976 3505 3004 7278
rect 4436 7200 4488 7206
rect 4436 7142 4488 7148
rect 3608 6656 3660 6662
rect 3608 6598 3660 6604
rect 3620 6390 3648 6598
rect 3608 6384 3660 6390
rect 3608 6326 3660 6332
rect 4160 6384 4212 6390
rect 4160 6326 4212 6332
rect 4172 5710 4200 6326
rect 4448 6254 4476 7142
rect 4724 6458 4752 37130
rect 4988 36848 5040 36854
rect 4988 36790 5040 36796
rect 5000 22642 5028 36790
rect 5184 36786 5212 38218
rect 5172 36780 5224 36786
rect 5172 36722 5224 36728
rect 5276 36378 5304 39238
rect 5356 38412 5408 38418
rect 5356 38354 5408 38360
rect 5368 36854 5396 38354
rect 5460 37330 5488 39510
rect 6552 38752 6604 38758
rect 6552 38694 6604 38700
rect 5582 38652 5890 38672
rect 5582 38650 5588 38652
rect 5644 38650 5668 38652
rect 5724 38650 5748 38652
rect 5804 38650 5828 38652
rect 5884 38650 5890 38652
rect 5644 38598 5646 38650
rect 5826 38598 5828 38650
rect 5582 38596 5588 38598
rect 5644 38596 5668 38598
rect 5724 38596 5748 38598
rect 5804 38596 5828 38598
rect 5884 38596 5890 38598
rect 5582 38576 5890 38596
rect 6564 38486 6592 38694
rect 6552 38480 6604 38486
rect 6552 38422 6604 38428
rect 6368 38276 6420 38282
rect 6368 38218 6420 38224
rect 6380 37874 6408 38218
rect 6368 37868 6420 37874
rect 6368 37810 6420 37816
rect 5582 37564 5890 37584
rect 5582 37562 5588 37564
rect 5644 37562 5668 37564
rect 5724 37562 5748 37564
rect 5804 37562 5828 37564
rect 5884 37562 5890 37564
rect 5644 37510 5646 37562
rect 5826 37510 5828 37562
rect 5582 37508 5588 37510
rect 5644 37508 5668 37510
rect 5724 37508 5748 37510
rect 5804 37508 5828 37510
rect 5884 37508 5890 37510
rect 5582 37488 5890 37508
rect 5448 37324 5500 37330
rect 5448 37266 5500 37272
rect 5356 36848 5408 36854
rect 5356 36790 5408 36796
rect 5264 36372 5316 36378
rect 5264 36314 5316 36320
rect 4988 22636 5040 22642
rect 4988 22578 5040 22584
rect 5460 9654 5488 37266
rect 5582 36476 5890 36496
rect 5582 36474 5588 36476
rect 5644 36474 5668 36476
rect 5724 36474 5748 36476
rect 5804 36474 5828 36476
rect 5884 36474 5890 36476
rect 5644 36422 5646 36474
rect 5826 36422 5828 36474
rect 5582 36420 5588 36422
rect 5644 36420 5668 36422
rect 5724 36420 5748 36422
rect 5804 36420 5828 36422
rect 5884 36420 5890 36422
rect 5582 36400 5890 36420
rect 6274 36408 6330 36417
rect 6274 36343 6330 36352
rect 5908 35556 5960 35562
rect 5908 35498 5960 35504
rect 5582 35388 5890 35408
rect 5582 35386 5588 35388
rect 5644 35386 5668 35388
rect 5724 35386 5748 35388
rect 5804 35386 5828 35388
rect 5884 35386 5890 35388
rect 5644 35334 5646 35386
rect 5826 35334 5828 35386
rect 5582 35332 5588 35334
rect 5644 35332 5668 35334
rect 5724 35332 5748 35334
rect 5804 35332 5828 35334
rect 5884 35332 5890 35334
rect 5582 35312 5890 35332
rect 5920 35222 5948 35498
rect 5998 35456 6054 35465
rect 5998 35391 6054 35400
rect 5908 35216 5960 35222
rect 5908 35158 5960 35164
rect 6012 35086 6040 35391
rect 6288 35290 6316 36343
rect 6380 36242 6408 37810
rect 6368 36236 6420 36242
rect 6368 36178 6420 36184
rect 6656 35698 6684 39782
rect 7116 39642 7144 39879
rect 7104 39636 7156 39642
rect 7104 39578 7156 39584
rect 7012 39568 7064 39574
rect 7012 39510 7064 39516
rect 6920 37800 6972 37806
rect 6920 37742 6972 37748
rect 6932 36378 6960 37742
rect 6920 36372 6972 36378
rect 6920 36314 6972 36320
rect 6736 36304 6788 36310
rect 6736 36246 6788 36252
rect 6644 35692 6696 35698
rect 6644 35634 6696 35640
rect 6276 35284 6328 35290
rect 6276 35226 6328 35232
rect 6748 35086 6776 36246
rect 6000 35080 6052 35086
rect 6000 35022 6052 35028
rect 6736 35080 6788 35086
rect 6736 35022 6788 35028
rect 5582 34300 5890 34320
rect 5582 34298 5588 34300
rect 5644 34298 5668 34300
rect 5724 34298 5748 34300
rect 5804 34298 5828 34300
rect 5884 34298 5890 34300
rect 5644 34246 5646 34298
rect 5826 34246 5828 34298
rect 5582 34244 5588 34246
rect 5644 34244 5668 34246
rect 5724 34244 5748 34246
rect 5804 34244 5828 34246
rect 5884 34244 5890 34246
rect 5582 34224 5890 34244
rect 5582 33212 5890 33232
rect 5582 33210 5588 33212
rect 5644 33210 5668 33212
rect 5724 33210 5748 33212
rect 5804 33210 5828 33212
rect 5884 33210 5890 33212
rect 5644 33158 5646 33210
rect 5826 33158 5828 33210
rect 5582 33156 5588 33158
rect 5644 33156 5668 33158
rect 5724 33156 5748 33158
rect 5804 33156 5828 33158
rect 5884 33156 5890 33158
rect 5582 33136 5890 33156
rect 5582 32124 5890 32144
rect 5582 32122 5588 32124
rect 5644 32122 5668 32124
rect 5724 32122 5748 32124
rect 5804 32122 5828 32124
rect 5884 32122 5890 32124
rect 5644 32070 5646 32122
rect 5826 32070 5828 32122
rect 5582 32068 5588 32070
rect 5644 32068 5668 32070
rect 5724 32068 5748 32070
rect 5804 32068 5828 32070
rect 5884 32068 5890 32070
rect 5582 32048 5890 32068
rect 6276 31816 6328 31822
rect 6276 31758 6328 31764
rect 5582 31036 5890 31056
rect 5582 31034 5588 31036
rect 5644 31034 5668 31036
rect 5724 31034 5748 31036
rect 5804 31034 5828 31036
rect 5884 31034 5890 31036
rect 5644 30982 5646 31034
rect 5826 30982 5828 31034
rect 5582 30980 5588 30982
rect 5644 30980 5668 30982
rect 5724 30980 5748 30982
rect 5804 30980 5828 30982
rect 5884 30980 5890 30982
rect 5582 30960 5890 30980
rect 5582 29948 5890 29968
rect 5582 29946 5588 29948
rect 5644 29946 5668 29948
rect 5724 29946 5748 29948
rect 5804 29946 5828 29948
rect 5884 29946 5890 29948
rect 5644 29894 5646 29946
rect 5826 29894 5828 29946
rect 5582 29892 5588 29894
rect 5644 29892 5668 29894
rect 5724 29892 5748 29894
rect 5804 29892 5828 29894
rect 5884 29892 5890 29894
rect 5582 29872 5890 29892
rect 5582 28860 5890 28880
rect 5582 28858 5588 28860
rect 5644 28858 5668 28860
rect 5724 28858 5748 28860
rect 5804 28858 5828 28860
rect 5884 28858 5890 28860
rect 5644 28806 5646 28858
rect 5826 28806 5828 28858
rect 5582 28804 5588 28806
rect 5644 28804 5668 28806
rect 5724 28804 5748 28806
rect 5804 28804 5828 28806
rect 5884 28804 5890 28806
rect 5582 28784 5890 28804
rect 5582 27772 5890 27792
rect 5582 27770 5588 27772
rect 5644 27770 5668 27772
rect 5724 27770 5748 27772
rect 5804 27770 5828 27772
rect 5884 27770 5890 27772
rect 5644 27718 5646 27770
rect 5826 27718 5828 27770
rect 5582 27716 5588 27718
rect 5644 27716 5668 27718
rect 5724 27716 5748 27718
rect 5804 27716 5828 27718
rect 5884 27716 5890 27718
rect 5582 27696 5890 27716
rect 5582 26684 5890 26704
rect 5582 26682 5588 26684
rect 5644 26682 5668 26684
rect 5724 26682 5748 26684
rect 5804 26682 5828 26684
rect 5884 26682 5890 26684
rect 5644 26630 5646 26682
rect 5826 26630 5828 26682
rect 5582 26628 5588 26630
rect 5644 26628 5668 26630
rect 5724 26628 5748 26630
rect 5804 26628 5828 26630
rect 5884 26628 5890 26630
rect 5582 26608 5890 26628
rect 5582 25596 5890 25616
rect 5582 25594 5588 25596
rect 5644 25594 5668 25596
rect 5724 25594 5748 25596
rect 5804 25594 5828 25596
rect 5884 25594 5890 25596
rect 5644 25542 5646 25594
rect 5826 25542 5828 25594
rect 5582 25540 5588 25542
rect 5644 25540 5668 25542
rect 5724 25540 5748 25542
rect 5804 25540 5828 25542
rect 5884 25540 5890 25542
rect 5582 25520 5890 25540
rect 5582 24508 5890 24528
rect 5582 24506 5588 24508
rect 5644 24506 5668 24508
rect 5724 24506 5748 24508
rect 5804 24506 5828 24508
rect 5884 24506 5890 24508
rect 5644 24454 5646 24506
rect 5826 24454 5828 24506
rect 5582 24452 5588 24454
rect 5644 24452 5668 24454
rect 5724 24452 5748 24454
rect 5804 24452 5828 24454
rect 5884 24452 5890 24454
rect 5582 24432 5890 24452
rect 5582 23420 5890 23440
rect 5582 23418 5588 23420
rect 5644 23418 5668 23420
rect 5724 23418 5748 23420
rect 5804 23418 5828 23420
rect 5884 23418 5890 23420
rect 5644 23366 5646 23418
rect 5826 23366 5828 23418
rect 5582 23364 5588 23366
rect 5644 23364 5668 23366
rect 5724 23364 5748 23366
rect 5804 23364 5828 23366
rect 5884 23364 5890 23366
rect 5582 23344 5890 23364
rect 5582 22332 5890 22352
rect 5582 22330 5588 22332
rect 5644 22330 5668 22332
rect 5724 22330 5748 22332
rect 5804 22330 5828 22332
rect 5884 22330 5890 22332
rect 5644 22278 5646 22330
rect 5826 22278 5828 22330
rect 5582 22276 5588 22278
rect 5644 22276 5668 22278
rect 5724 22276 5748 22278
rect 5804 22276 5828 22278
rect 5884 22276 5890 22278
rect 5582 22256 5890 22276
rect 5582 21244 5890 21264
rect 5582 21242 5588 21244
rect 5644 21242 5668 21244
rect 5724 21242 5748 21244
rect 5804 21242 5828 21244
rect 5884 21242 5890 21244
rect 5644 21190 5646 21242
rect 5826 21190 5828 21242
rect 5582 21188 5588 21190
rect 5644 21188 5668 21190
rect 5724 21188 5748 21190
rect 5804 21188 5828 21190
rect 5884 21188 5890 21190
rect 5582 21168 5890 21188
rect 5582 20156 5890 20176
rect 5582 20154 5588 20156
rect 5644 20154 5668 20156
rect 5724 20154 5748 20156
rect 5804 20154 5828 20156
rect 5884 20154 5890 20156
rect 5644 20102 5646 20154
rect 5826 20102 5828 20154
rect 5582 20100 5588 20102
rect 5644 20100 5668 20102
rect 5724 20100 5748 20102
rect 5804 20100 5828 20102
rect 5884 20100 5890 20102
rect 5582 20080 5890 20100
rect 5582 19068 5890 19088
rect 5582 19066 5588 19068
rect 5644 19066 5668 19068
rect 5724 19066 5748 19068
rect 5804 19066 5828 19068
rect 5884 19066 5890 19068
rect 5644 19014 5646 19066
rect 5826 19014 5828 19066
rect 5582 19012 5588 19014
rect 5644 19012 5668 19014
rect 5724 19012 5748 19014
rect 5804 19012 5828 19014
rect 5884 19012 5890 19014
rect 5582 18992 5890 19012
rect 5582 17980 5890 18000
rect 5582 17978 5588 17980
rect 5644 17978 5668 17980
rect 5724 17978 5748 17980
rect 5804 17978 5828 17980
rect 5884 17978 5890 17980
rect 5644 17926 5646 17978
rect 5826 17926 5828 17978
rect 5582 17924 5588 17926
rect 5644 17924 5668 17926
rect 5724 17924 5748 17926
rect 5804 17924 5828 17926
rect 5884 17924 5890 17926
rect 5582 17904 5890 17924
rect 6288 17882 6316 31758
rect 6736 31680 6788 31686
rect 6788 31628 6868 31634
rect 6736 31622 6868 31628
rect 6748 31606 6868 31622
rect 6736 30048 6788 30054
rect 6736 29990 6788 29996
rect 6748 29714 6776 29990
rect 6736 29708 6788 29714
rect 6736 29650 6788 29656
rect 6840 27334 6868 31606
rect 7024 30938 7052 39510
rect 7104 39296 7156 39302
rect 7104 39238 7156 39244
rect 7116 36378 7144 39238
rect 7208 37466 7236 40326
rect 7286 39808 7342 39817
rect 7286 39743 7342 39752
rect 7196 37460 7248 37466
rect 7196 37402 7248 37408
rect 7300 36786 7328 39743
rect 7392 38962 7420 40394
rect 7380 38956 7432 38962
rect 7380 38898 7432 38904
rect 7378 38312 7434 38321
rect 7378 38247 7434 38256
rect 7288 36780 7340 36786
rect 7288 36722 7340 36728
rect 7286 36680 7342 36689
rect 7286 36615 7342 36624
rect 7104 36372 7156 36378
rect 7104 36314 7156 36320
rect 7300 35154 7328 36615
rect 7392 35766 7420 38247
rect 7380 35760 7432 35766
rect 7380 35702 7432 35708
rect 7288 35148 7340 35154
rect 7288 35090 7340 35096
rect 7104 35080 7156 35086
rect 7104 35022 7156 35028
rect 7116 34649 7144 35022
rect 7102 34640 7158 34649
rect 7102 34575 7158 34584
rect 7484 34474 7512 40530
rect 7576 36310 7604 40666
rect 7656 40656 7708 40662
rect 7656 40598 7708 40604
rect 7564 36304 7616 36310
rect 7564 36246 7616 36252
rect 7562 35728 7618 35737
rect 7562 35663 7564 35672
rect 7616 35663 7618 35672
rect 7564 35634 7616 35640
rect 7564 34944 7616 34950
rect 7564 34886 7616 34892
rect 7576 34649 7604 34886
rect 7562 34640 7618 34649
rect 7562 34575 7618 34584
rect 7472 34468 7524 34474
rect 7472 34410 7524 34416
rect 7564 34400 7616 34406
rect 7564 34342 7616 34348
rect 7576 34105 7604 34342
rect 7562 34096 7618 34105
rect 7562 34031 7618 34040
rect 7668 33998 7696 40598
rect 8666 40488 8722 40497
rect 8666 40423 8722 40432
rect 8392 40112 8444 40118
rect 8392 40054 8444 40060
rect 7932 40044 7984 40050
rect 7932 39986 7984 39992
rect 7838 39400 7894 39409
rect 7838 39335 7894 39344
rect 7748 38480 7800 38486
rect 7746 38448 7748 38457
rect 7800 38448 7802 38457
rect 7746 38383 7802 38392
rect 7852 37466 7880 39335
rect 7840 37460 7892 37466
rect 7840 37402 7892 37408
rect 7944 37346 7972 39986
rect 8298 38992 8354 39001
rect 8298 38927 8354 38936
rect 8022 38856 8078 38865
rect 8022 38791 8024 38800
rect 8076 38791 8078 38800
rect 8024 38762 8076 38768
rect 8206 38040 8262 38049
rect 8206 37975 8262 37984
rect 8116 37664 8168 37670
rect 8116 37606 8168 37612
rect 8220 37618 8248 37975
rect 8312 37738 8340 38927
rect 8404 38554 8432 40054
rect 8484 39908 8536 39914
rect 8484 39850 8536 39856
rect 8392 38548 8444 38554
rect 8392 38490 8444 38496
rect 8496 38282 8524 39850
rect 8680 38962 8708 40423
rect 8668 38956 8720 38962
rect 8668 38898 8720 38904
rect 8576 38888 8628 38894
rect 8576 38830 8628 38836
rect 8588 38418 8616 38830
rect 8576 38412 8628 38418
rect 8576 38354 8628 38360
rect 8484 38276 8536 38282
rect 8484 38218 8536 38224
rect 8666 37768 8722 37777
rect 8300 37732 8352 37738
rect 8300 37674 8352 37680
rect 8484 37732 8536 37738
rect 8666 37703 8722 37712
rect 8484 37674 8536 37680
rect 8392 37664 8444 37670
rect 8022 37496 8078 37505
rect 8128 37466 8156 37606
rect 8220 37590 8340 37618
rect 8392 37606 8444 37612
rect 8022 37431 8078 37440
rect 8116 37460 8168 37466
rect 7852 37318 7972 37346
rect 7852 36174 7880 37318
rect 7932 36712 7984 36718
rect 7932 36654 7984 36660
rect 7840 36168 7892 36174
rect 7840 36110 7892 36116
rect 7840 35012 7892 35018
rect 7840 34954 7892 34960
rect 7748 34196 7800 34202
rect 7748 34138 7800 34144
rect 7760 33998 7788 34138
rect 7656 33992 7708 33998
rect 7656 33934 7708 33940
rect 7748 33992 7800 33998
rect 7748 33934 7800 33940
rect 7564 33856 7616 33862
rect 7564 33798 7616 33804
rect 7576 33289 7604 33798
rect 7852 33522 7880 34954
rect 7840 33516 7892 33522
rect 7840 33458 7892 33464
rect 7562 33280 7618 33289
rect 7562 33215 7618 33224
rect 7840 32904 7892 32910
rect 7840 32846 7892 32852
rect 7012 30932 7064 30938
rect 7012 30874 7064 30880
rect 7564 29640 7616 29646
rect 7564 29582 7616 29588
rect 6828 27328 6880 27334
rect 6828 27270 6880 27276
rect 6276 17876 6328 17882
rect 6276 17818 6328 17824
rect 7576 17785 7604 29582
rect 7748 29028 7800 29034
rect 7748 28970 7800 28976
rect 7562 17776 7618 17785
rect 7562 17711 7618 17720
rect 5582 16892 5890 16912
rect 5582 16890 5588 16892
rect 5644 16890 5668 16892
rect 5724 16890 5748 16892
rect 5804 16890 5828 16892
rect 5884 16890 5890 16892
rect 5644 16838 5646 16890
rect 5826 16838 5828 16890
rect 5582 16836 5588 16838
rect 5644 16836 5668 16838
rect 5724 16836 5748 16838
rect 5804 16836 5828 16838
rect 5884 16836 5890 16838
rect 5582 16816 5890 16836
rect 7760 16561 7788 28970
rect 7852 24857 7880 32846
rect 7944 31822 7972 36654
rect 8036 35834 8064 37431
rect 8116 37402 8168 37408
rect 8116 37256 8168 37262
rect 8116 37198 8168 37204
rect 8206 37224 8262 37233
rect 8128 36582 8156 37198
rect 8206 37159 8262 37168
rect 8220 36786 8248 37159
rect 8208 36780 8260 36786
rect 8208 36722 8260 36728
rect 8116 36576 8168 36582
rect 8116 36518 8168 36524
rect 8024 35828 8076 35834
rect 8024 35770 8076 35776
rect 8206 35728 8262 35737
rect 8206 35663 8208 35672
rect 8260 35663 8262 35672
rect 8208 35634 8260 35640
rect 8024 35216 8076 35222
rect 8024 35158 8076 35164
rect 7932 31816 7984 31822
rect 7932 31758 7984 31764
rect 8036 30734 8064 35158
rect 8114 33552 8170 33561
rect 8114 33487 8170 33496
rect 8128 32434 8156 33487
rect 8116 32428 8168 32434
rect 8116 32370 8168 32376
rect 8312 31668 8340 37590
rect 8404 36174 8432 37606
rect 8496 36786 8524 37674
rect 8484 36780 8536 36786
rect 8484 36722 8536 36728
rect 8392 36168 8444 36174
rect 8392 36110 8444 36116
rect 8390 35184 8446 35193
rect 8390 35119 8446 35128
rect 8404 35086 8432 35119
rect 8392 35080 8444 35086
rect 8392 35022 8444 35028
rect 8484 34944 8536 34950
rect 8390 34912 8446 34921
rect 8484 34886 8536 34892
rect 8390 34847 8446 34856
rect 8404 34610 8432 34847
rect 8392 34604 8444 34610
rect 8392 34546 8444 34552
rect 8496 34241 8524 34886
rect 8482 34232 8538 34241
rect 8482 34167 8538 34176
rect 8484 33992 8536 33998
rect 8482 33960 8484 33969
rect 8536 33960 8538 33969
rect 8482 33895 8538 33904
rect 8496 33522 8524 33895
rect 8484 33516 8536 33522
rect 8484 33458 8536 33464
rect 8392 31680 8444 31686
rect 8312 31640 8392 31668
rect 8392 31622 8444 31628
rect 8300 31340 8352 31346
rect 8300 31282 8352 31288
rect 8208 31272 8260 31278
rect 8114 31240 8170 31249
rect 8208 31214 8260 31220
rect 8114 31175 8116 31184
rect 8168 31175 8170 31184
rect 8116 31146 8168 31152
rect 8024 30728 8076 30734
rect 8024 30670 8076 30676
rect 8220 30569 8248 31214
rect 8312 30802 8340 31282
rect 8300 30796 8352 30802
rect 8300 30738 8352 30744
rect 8206 30560 8262 30569
rect 8206 30495 8262 30504
rect 8496 30258 8524 33458
rect 8680 32994 8708 37703
rect 8758 37360 8814 37369
rect 8758 37295 8814 37304
rect 8772 35562 8800 37295
rect 8864 36854 8892 40734
rect 8944 40520 8996 40526
rect 8944 40462 8996 40468
rect 8852 36848 8904 36854
rect 8852 36790 8904 36796
rect 8956 36786 8984 40462
rect 8944 36780 8996 36786
rect 8944 36722 8996 36728
rect 8850 36544 8906 36553
rect 8850 36479 8906 36488
rect 8760 35556 8812 35562
rect 8760 35498 8812 35504
rect 8760 34672 8812 34678
rect 8760 34614 8812 34620
rect 8772 34377 8800 34614
rect 8758 34368 8814 34377
rect 8758 34303 8814 34312
rect 8864 34134 8892 36479
rect 8944 36304 8996 36310
rect 8942 36272 8944 36281
rect 8996 36272 8998 36281
rect 8942 36207 8998 36216
rect 9048 35873 9076 40802
rect 9312 40316 9364 40322
rect 9312 40258 9364 40264
rect 9324 38962 9352 40258
rect 10324 40248 10376 40254
rect 10324 40190 10376 40196
rect 9864 40180 9916 40186
rect 9864 40122 9916 40128
rect 9680 39976 9732 39982
rect 9680 39918 9732 39924
rect 9692 39438 9720 39918
rect 9680 39432 9732 39438
rect 9680 39374 9732 39380
rect 9772 39364 9824 39370
rect 9772 39306 9824 39312
rect 9312 38956 9364 38962
rect 9312 38898 9364 38904
rect 9220 38888 9272 38894
rect 9220 38830 9272 38836
rect 9232 38758 9260 38830
rect 9128 38752 9180 38758
rect 9128 38694 9180 38700
rect 9220 38752 9272 38758
rect 9220 38694 9272 38700
rect 9140 38282 9168 38694
rect 9404 38548 9456 38554
rect 9404 38490 9456 38496
rect 9416 38418 9444 38490
rect 9784 38418 9812 39306
rect 9404 38412 9456 38418
rect 9404 38354 9456 38360
rect 9772 38412 9824 38418
rect 9772 38354 9824 38360
rect 9496 38344 9548 38350
rect 9494 38312 9496 38321
rect 9548 38312 9550 38321
rect 9128 38276 9180 38282
rect 9494 38247 9550 38256
rect 9678 38312 9734 38321
rect 9678 38247 9734 38256
rect 9128 38218 9180 38224
rect 9140 37806 9168 38218
rect 9218 37904 9274 37913
rect 9218 37839 9274 37848
rect 9128 37800 9180 37806
rect 9128 37742 9180 37748
rect 9128 37256 9180 37262
rect 9128 37198 9180 37204
rect 9140 36310 9168 37198
rect 9232 36786 9260 37839
rect 9312 37800 9364 37806
rect 9312 37742 9364 37748
rect 9220 36780 9272 36786
rect 9220 36722 9272 36728
rect 9324 36378 9352 37742
rect 9494 37632 9550 37641
rect 9494 37567 9550 37576
rect 9404 36712 9456 36718
rect 9404 36654 9456 36660
rect 9312 36372 9364 36378
rect 9312 36314 9364 36320
rect 9128 36304 9180 36310
rect 9416 36281 9444 36654
rect 9128 36246 9180 36252
rect 9402 36272 9458 36281
rect 9402 36207 9458 36216
rect 9310 36136 9366 36145
rect 9220 36100 9272 36106
rect 9310 36071 9366 36080
rect 9220 36042 9272 36048
rect 9126 36000 9182 36009
rect 9126 35935 9182 35944
rect 9034 35864 9090 35873
rect 9034 35799 9090 35808
rect 9036 35624 9088 35630
rect 9036 35566 9088 35572
rect 8944 35148 8996 35154
rect 8944 35090 8996 35096
rect 8852 34128 8904 34134
rect 8852 34070 8904 34076
rect 8956 33697 8984 35090
rect 9048 34746 9076 35566
rect 9140 35086 9168 35935
rect 9232 35834 9260 36042
rect 9220 35828 9272 35834
rect 9220 35770 9272 35776
rect 9324 35698 9352 36071
rect 9508 35894 9536 37567
rect 9588 37392 9640 37398
rect 9588 37334 9640 37340
rect 9600 36961 9628 37334
rect 9692 37262 9720 38247
rect 9772 37868 9824 37874
rect 9772 37810 9824 37816
rect 9784 37398 9812 37810
rect 9772 37392 9824 37398
rect 9772 37334 9824 37340
rect 9680 37256 9732 37262
rect 9680 37198 9732 37204
rect 9772 37256 9824 37262
rect 9772 37198 9824 37204
rect 9586 36952 9642 36961
rect 9692 36922 9720 37198
rect 9586 36887 9642 36896
rect 9680 36916 9732 36922
rect 9680 36858 9732 36864
rect 9586 36816 9642 36825
rect 9784 36786 9812 37198
rect 9876 37097 9904 40122
rect 10336 39506 10364 40190
rect 10876 39636 10928 39642
rect 10876 39578 10928 39584
rect 10140 39500 10192 39506
rect 10140 39442 10192 39448
rect 10324 39500 10376 39506
rect 10324 39442 10376 39448
rect 10692 39500 10744 39506
rect 10692 39442 10744 39448
rect 10048 39432 10100 39438
rect 10048 39374 10100 39380
rect 10060 38350 10088 39374
rect 10152 38418 10180 39442
rect 10704 39302 10732 39442
rect 10888 39438 10916 39578
rect 10784 39432 10836 39438
rect 10784 39374 10836 39380
rect 10876 39432 10928 39438
rect 10876 39374 10928 39380
rect 10692 39296 10744 39302
rect 10692 39238 10744 39244
rect 10214 39196 10522 39216
rect 10214 39194 10220 39196
rect 10276 39194 10300 39196
rect 10356 39194 10380 39196
rect 10436 39194 10460 39196
rect 10516 39194 10522 39196
rect 10276 39142 10278 39194
rect 10458 39142 10460 39194
rect 10214 39140 10220 39142
rect 10276 39140 10300 39142
rect 10356 39140 10380 39142
rect 10436 39140 10460 39142
rect 10516 39140 10522 39142
rect 10214 39120 10522 39140
rect 10232 38956 10284 38962
rect 10232 38898 10284 38904
rect 10140 38412 10192 38418
rect 10140 38354 10192 38360
rect 10048 38344 10100 38350
rect 10244 38298 10272 38898
rect 10324 38888 10376 38894
rect 10324 38830 10376 38836
rect 10336 38758 10364 38830
rect 10324 38752 10376 38758
rect 10324 38694 10376 38700
rect 10508 38752 10560 38758
rect 10508 38694 10560 38700
rect 10690 38720 10746 38729
rect 10520 38418 10548 38694
rect 10690 38655 10746 38664
rect 10508 38412 10560 38418
rect 10508 38354 10560 38360
rect 10048 38286 10100 38292
rect 10152 38270 10272 38298
rect 10048 38208 10100 38214
rect 10048 38150 10100 38156
rect 9954 38040 10010 38049
rect 9954 37975 10010 37984
rect 9968 37652 9996 37975
rect 10060 37806 10088 38150
rect 10152 37806 10180 38270
rect 10214 38108 10522 38128
rect 10214 38106 10220 38108
rect 10276 38106 10300 38108
rect 10356 38106 10380 38108
rect 10436 38106 10460 38108
rect 10516 38106 10522 38108
rect 10276 38054 10278 38106
rect 10458 38054 10460 38106
rect 10214 38052 10220 38054
rect 10276 38052 10300 38054
rect 10356 38052 10380 38054
rect 10436 38052 10460 38054
rect 10516 38052 10522 38054
rect 10214 38032 10522 38052
rect 10416 37868 10468 37874
rect 10416 37810 10468 37816
rect 10508 37868 10560 37874
rect 10508 37810 10560 37816
rect 10048 37800 10100 37806
rect 10048 37742 10100 37748
rect 10140 37800 10192 37806
rect 10140 37742 10192 37748
rect 10152 37652 10180 37742
rect 9968 37624 10180 37652
rect 10428 37262 10456 37810
rect 10416 37256 10468 37262
rect 10416 37198 10468 37204
rect 10520 37108 10548 37810
rect 10704 37312 10732 38655
rect 10796 38185 10824 39374
rect 10874 39128 10930 39137
rect 10874 39063 10930 39072
rect 10888 39030 10916 39063
rect 10876 39024 10928 39030
rect 10876 38966 10928 38972
rect 10980 38418 11008 41200
rect 11426 40352 11482 40361
rect 11426 40287 11482 40296
rect 11060 40112 11112 40118
rect 11060 40054 11112 40060
rect 11072 39642 11100 40054
rect 11060 39636 11112 39642
rect 11060 39578 11112 39584
rect 11336 38820 11388 38826
rect 11336 38762 11388 38768
rect 11244 38752 11296 38758
rect 11244 38694 11296 38700
rect 10968 38412 11020 38418
rect 10968 38354 11020 38360
rect 11256 38264 11284 38694
rect 11164 38236 11284 38264
rect 10782 38176 10838 38185
rect 10782 38111 10838 38120
rect 10874 38040 10930 38049
rect 10874 37975 10930 37984
rect 10704 37284 10824 37312
rect 10692 37188 10744 37194
rect 10692 37130 10744 37136
rect 9862 37088 9918 37097
rect 9862 37023 9918 37032
rect 9968 37080 10548 37108
rect 10704 37097 10732 37130
rect 10690 37088 10746 37097
rect 9586 36751 9642 36760
rect 9772 36780 9824 36786
rect 9600 36378 9628 36751
rect 9772 36722 9824 36728
rect 9588 36372 9640 36378
rect 9588 36314 9640 36320
rect 9770 36272 9826 36281
rect 9770 36207 9826 36216
rect 9784 36174 9812 36207
rect 9772 36168 9824 36174
rect 9772 36110 9824 36116
rect 9968 36038 9996 37080
rect 10214 37020 10522 37040
rect 10690 37023 10746 37032
rect 10214 37018 10220 37020
rect 10276 37018 10300 37020
rect 10356 37018 10380 37020
rect 10436 37018 10460 37020
rect 10516 37018 10522 37020
rect 10276 36966 10278 37018
rect 10458 36966 10460 37018
rect 10214 36964 10220 36966
rect 10276 36964 10300 36966
rect 10356 36964 10380 36966
rect 10436 36964 10460 36966
rect 10516 36964 10522 36966
rect 10046 36952 10102 36961
rect 10214 36944 10522 36964
rect 10046 36887 10102 36896
rect 10060 36786 10088 36887
rect 10796 36786 10824 37284
rect 10888 37194 10916 37975
rect 11060 37868 11112 37874
rect 11060 37810 11112 37816
rect 11072 37194 11100 37810
rect 10876 37188 10928 37194
rect 10876 37130 10928 37136
rect 11060 37188 11112 37194
rect 11060 37130 11112 37136
rect 11060 36848 11112 36854
rect 11164 36836 11192 38236
rect 11244 37868 11296 37874
rect 11244 37810 11296 37816
rect 11112 36808 11192 36836
rect 11060 36790 11112 36796
rect 10048 36780 10100 36786
rect 10416 36780 10468 36786
rect 10048 36722 10100 36728
rect 10152 36740 10416 36768
rect 9956 36032 10008 36038
rect 10048 36032 10100 36038
rect 9956 35974 10008 35980
rect 10046 36000 10048 36009
rect 10100 36000 10102 36009
rect 10046 35935 10102 35944
rect 10152 35894 10180 36740
rect 10416 36722 10468 36728
rect 10784 36780 10836 36786
rect 10784 36722 10836 36728
rect 10968 36780 11020 36786
rect 11256 36768 11284 37810
rect 10968 36722 11020 36728
rect 11164 36740 11284 36768
rect 10324 36576 10376 36582
rect 10980 36564 11008 36722
rect 10324 36518 10376 36524
rect 10612 36536 11008 36564
rect 10336 36281 10364 36518
rect 10612 36310 10640 36536
rect 10600 36304 10652 36310
rect 10322 36272 10378 36281
rect 10600 36246 10652 36252
rect 10322 36207 10378 36216
rect 10784 36236 10836 36242
rect 10784 36178 10836 36184
rect 10598 36000 10654 36009
rect 9416 35866 9536 35894
rect 9312 35692 9364 35698
rect 9312 35634 9364 35640
rect 9218 35320 9274 35329
rect 9218 35255 9220 35264
rect 9272 35255 9274 35264
rect 9220 35226 9272 35232
rect 9416 35086 9444 35866
rect 9862 35864 9918 35873
rect 9862 35799 9918 35808
rect 9968 35866 10180 35894
rect 10214 35932 10522 35952
rect 10598 35935 10654 35944
rect 10214 35930 10220 35932
rect 10276 35930 10300 35932
rect 10356 35930 10380 35932
rect 10436 35930 10460 35932
rect 10516 35930 10522 35932
rect 10276 35878 10278 35930
rect 10458 35878 10460 35930
rect 10214 35876 10220 35878
rect 10276 35876 10300 35878
rect 10356 35876 10380 35878
rect 10436 35876 10460 35878
rect 10516 35876 10522 35878
rect 9496 35692 9548 35698
rect 9496 35634 9548 35640
rect 9508 35601 9536 35634
rect 9876 35630 9904 35799
rect 9968 35698 9996 35866
rect 10214 35856 10522 35876
rect 10612 35816 10640 35935
rect 10612 35788 10732 35816
rect 10232 35760 10284 35766
rect 10060 35720 10232 35748
rect 9956 35692 10008 35698
rect 9956 35634 10008 35640
rect 9864 35624 9916 35630
rect 9494 35592 9550 35601
rect 9864 35566 9916 35572
rect 9494 35527 9550 35536
rect 9494 35320 9550 35329
rect 10060 35306 10088 35720
rect 10232 35702 10284 35708
rect 10704 35680 10732 35788
rect 10520 35652 10732 35680
rect 10520 35578 10548 35652
rect 10796 35612 10824 36178
rect 10968 36168 11020 36174
rect 10968 36110 11020 36116
rect 11060 36168 11112 36174
rect 11060 36110 11112 36116
rect 10980 36038 11008 36110
rect 10876 36032 10928 36038
rect 10876 35974 10928 35980
rect 10968 36032 11020 36038
rect 11072 36009 11100 36110
rect 10968 35974 11020 35980
rect 11058 36000 11114 36009
rect 10888 35873 10916 35974
rect 11058 35935 11114 35944
rect 10874 35864 10930 35873
rect 10874 35799 10930 35808
rect 11060 35760 11112 35766
rect 11060 35702 11112 35708
rect 10876 35624 10928 35630
rect 10796 35584 10876 35612
rect 10244 35550 10548 35578
rect 10876 35566 10928 35572
rect 10244 35494 10272 35550
rect 10232 35488 10284 35494
rect 10232 35430 10284 35436
rect 10324 35488 10376 35494
rect 10324 35430 10376 35436
rect 10336 35306 10364 35430
rect 9494 35255 9550 35264
rect 9588 35284 9640 35290
rect 9128 35080 9180 35086
rect 9128 35022 9180 35028
rect 9220 35080 9272 35086
rect 9220 35022 9272 35028
rect 9404 35080 9456 35086
rect 9404 35022 9456 35028
rect 9036 34740 9088 34746
rect 9036 34682 9088 34688
rect 8942 33688 8998 33697
rect 8942 33623 8998 33632
rect 9036 33040 9088 33046
rect 8680 32966 8892 32994
rect 9036 32982 9088 32988
rect 8760 32836 8812 32842
rect 8760 32778 8812 32784
rect 8772 32434 8800 32778
rect 8760 32428 8812 32434
rect 8760 32370 8812 32376
rect 8666 32328 8722 32337
rect 8666 32263 8668 32272
rect 8720 32263 8722 32272
rect 8668 32234 8720 32240
rect 8576 31136 8628 31142
rect 8576 31078 8628 31084
rect 8668 31136 8720 31142
rect 8668 31078 8720 31084
rect 8588 30841 8616 31078
rect 8574 30832 8630 30841
rect 8574 30767 8630 30776
rect 8680 30734 8708 31078
rect 8668 30728 8720 30734
rect 8668 30670 8720 30676
rect 8484 30252 8536 30258
rect 8484 30194 8536 30200
rect 8760 30252 8812 30258
rect 8760 30194 8812 30200
rect 8576 30048 8628 30054
rect 8576 29990 8628 29996
rect 8668 30048 8720 30054
rect 8668 29990 8720 29996
rect 8588 29889 8616 29990
rect 8574 29880 8630 29889
rect 8574 29815 8630 29824
rect 8680 29753 8708 29990
rect 8666 29744 8722 29753
rect 8666 29679 8722 29688
rect 8392 29640 8444 29646
rect 8390 29608 8392 29617
rect 8444 29608 8446 29617
rect 8390 29543 8446 29552
rect 8772 28558 8800 30194
rect 8864 28626 8892 32966
rect 8944 32904 8996 32910
rect 8944 32846 8996 32852
rect 8956 31521 8984 32846
rect 8942 31512 8998 31521
rect 8942 31447 8998 31456
rect 8944 31340 8996 31346
rect 9048 31328 9076 32982
rect 9128 32224 9180 32230
rect 9126 32192 9128 32201
rect 9180 32192 9182 32201
rect 9126 32127 9182 32136
rect 9126 32056 9182 32065
rect 9126 31991 9182 32000
rect 9140 31754 9168 31991
rect 9128 31748 9180 31754
rect 9128 31690 9180 31696
rect 9128 31340 9180 31346
rect 9048 31300 9128 31328
rect 8944 31282 8996 31288
rect 9128 31282 9180 31288
rect 8852 28620 8904 28626
rect 8852 28562 8904 28568
rect 8760 28552 8812 28558
rect 8760 28494 8812 28500
rect 8208 28416 8260 28422
rect 8208 28358 8260 28364
rect 8220 28014 8248 28358
rect 8300 28212 8352 28218
rect 8300 28154 8352 28160
rect 8312 28121 8340 28154
rect 8298 28112 8354 28121
rect 8298 28047 8354 28056
rect 8208 28008 8260 28014
rect 8208 27950 8260 27956
rect 8956 27577 8984 31282
rect 9140 30705 9168 31282
rect 9126 30696 9182 30705
rect 9126 30631 9182 30640
rect 9036 30592 9088 30598
rect 9036 30534 9088 30540
rect 9048 28529 9076 30534
rect 9232 30172 9260 35022
rect 9508 34746 9536 35255
rect 9588 35226 9640 35232
rect 9968 35278 10088 35306
rect 10152 35278 10364 35306
rect 10968 35284 11020 35290
rect 9600 35193 9628 35226
rect 9586 35184 9642 35193
rect 9586 35119 9642 35128
rect 9862 35048 9918 35057
rect 9862 34983 9918 34992
rect 9876 34950 9904 34983
rect 9864 34944 9916 34950
rect 9968 34921 9996 35278
rect 10152 35222 10180 35278
rect 10968 35226 11020 35232
rect 10140 35216 10192 35222
rect 10416 35216 10468 35222
rect 10140 35158 10192 35164
rect 10244 35164 10416 35170
rect 10244 35158 10468 35164
rect 10244 35142 10456 35158
rect 10244 35018 10272 35142
rect 10324 35080 10376 35086
rect 10376 35040 10640 35068
rect 10324 35022 10376 35028
rect 10232 35012 10284 35018
rect 10232 34954 10284 34960
rect 10140 34944 10192 34950
rect 9864 34886 9916 34892
rect 9954 34912 10010 34921
rect 10612 34921 10640 35040
rect 10980 34950 11008 35226
rect 10968 34944 11020 34950
rect 10140 34886 10192 34892
rect 10598 34912 10654 34921
rect 9954 34847 10010 34856
rect 10046 34776 10102 34785
rect 9496 34740 9548 34746
rect 10046 34711 10102 34720
rect 9496 34682 9548 34688
rect 10060 34610 10088 34711
rect 9588 34604 9640 34610
rect 9588 34546 9640 34552
rect 10048 34604 10100 34610
rect 10048 34546 10100 34552
rect 9310 34504 9366 34513
rect 9310 34439 9366 34448
rect 9324 33998 9352 34439
rect 9600 34406 9628 34546
rect 10152 34490 10180 34886
rect 10214 34844 10522 34864
rect 10598 34847 10654 34856
rect 10874 34912 10930 34921
rect 10968 34886 11020 34892
rect 10874 34847 10930 34856
rect 10214 34842 10220 34844
rect 10276 34842 10300 34844
rect 10356 34842 10380 34844
rect 10436 34842 10460 34844
rect 10516 34842 10522 34844
rect 10276 34790 10278 34842
rect 10458 34790 10460 34842
rect 10214 34788 10220 34790
rect 10276 34788 10300 34790
rect 10356 34788 10380 34790
rect 10436 34788 10460 34790
rect 10516 34788 10522 34790
rect 10214 34768 10522 34788
rect 10888 34660 10916 34847
rect 10796 34632 10916 34660
rect 10152 34462 10732 34490
rect 9876 34428 10088 34456
rect 9588 34400 9640 34406
rect 9588 34342 9640 34348
rect 9404 34128 9456 34134
rect 9876 34116 9904 34428
rect 10060 34354 10088 34428
rect 10600 34400 10652 34406
rect 10060 34326 10548 34354
rect 10600 34342 10652 34348
rect 10704 34354 10732 34462
rect 10796 34456 10824 34632
rect 11072 34610 11100 35702
rect 11164 35018 11192 36740
rect 11256 35222 11284 35253
rect 11244 35216 11296 35222
rect 11348 35170 11376 38762
rect 11440 37874 11468 40287
rect 12162 40216 12218 40225
rect 12162 40151 12218 40160
rect 11888 39908 11940 39914
rect 11888 39850 11940 39856
rect 11796 39500 11848 39506
rect 11532 39460 11796 39488
rect 11532 39370 11560 39460
rect 11796 39442 11848 39448
rect 11520 39364 11572 39370
rect 11520 39306 11572 39312
rect 11900 38962 11928 39850
rect 12176 39681 12204 40151
rect 12162 39672 12218 39681
rect 12162 39607 12218 39616
rect 12268 39506 12296 41200
rect 12530 40216 12586 40225
rect 12530 40151 12586 40160
rect 12624 40180 12676 40186
rect 12544 39953 12572 40151
rect 12624 40122 12676 40128
rect 12530 39944 12586 39953
rect 12440 39908 12492 39914
rect 12530 39879 12586 39888
rect 12440 39850 12492 39856
rect 12346 39672 12402 39681
rect 12346 39607 12402 39616
rect 12256 39500 12308 39506
rect 12256 39442 12308 39448
rect 12360 39386 12388 39607
rect 12452 39488 12480 39850
rect 12532 39500 12584 39506
rect 12452 39460 12532 39488
rect 12532 39442 12584 39448
rect 12268 39358 12388 39386
rect 11888 38956 11940 38962
rect 11888 38898 11940 38904
rect 12268 38654 12296 39358
rect 12348 39296 12400 39302
rect 12348 39238 12400 39244
rect 12084 38626 12296 38654
rect 11796 38344 11848 38350
rect 11796 38286 11848 38292
rect 11808 38214 11836 38286
rect 11796 38208 11848 38214
rect 11796 38150 11848 38156
rect 11980 38208 12032 38214
rect 11980 38150 12032 38156
rect 11992 38049 12020 38150
rect 11978 38040 12034 38049
rect 11978 37975 12034 37984
rect 11888 37936 11940 37942
rect 11888 37878 11940 37884
rect 11428 37868 11480 37874
rect 11428 37810 11480 37816
rect 11520 37868 11572 37874
rect 11520 37810 11572 37816
rect 11532 37398 11560 37810
rect 11612 37800 11664 37806
rect 11900 37788 11928 37878
rect 11664 37760 11928 37788
rect 11980 37800 12032 37806
rect 11612 37742 11664 37748
rect 12084 37777 12112 38626
rect 12164 38548 12216 38554
rect 12164 38490 12216 38496
rect 12176 38350 12204 38490
rect 12164 38344 12216 38350
rect 12164 38286 12216 38292
rect 12360 38196 12388 39238
rect 12636 38944 12664 40122
rect 12716 39976 12768 39982
rect 12716 39918 12768 39924
rect 12728 38962 12756 39918
rect 12808 39296 12860 39302
rect 12808 39238 12860 39244
rect 12176 38168 12388 38196
rect 12452 38916 12664 38944
rect 12716 38956 12768 38962
rect 12176 37806 12204 38168
rect 12452 37856 12480 38916
rect 12716 38898 12768 38904
rect 12820 38842 12848 39238
rect 12728 38814 12848 38842
rect 12532 38752 12584 38758
rect 12532 38694 12584 38700
rect 12544 38049 12572 38694
rect 12624 38412 12676 38418
rect 12624 38354 12676 38360
rect 12530 38040 12586 38049
rect 12530 37975 12586 37984
rect 12636 37942 12664 38354
rect 12624 37936 12676 37942
rect 12624 37878 12676 37884
rect 12268 37828 12480 37856
rect 12164 37800 12216 37806
rect 11980 37742 12032 37748
rect 12070 37768 12126 37777
rect 11992 37652 12020 37742
rect 12164 37742 12216 37748
rect 12070 37703 12126 37712
rect 12268 37652 12296 37828
rect 12728 37788 12756 38814
rect 12808 38344 12860 38350
rect 12808 38286 12860 38292
rect 12820 37942 12848 38286
rect 12808 37936 12860 37942
rect 12808 37878 12860 37884
rect 12912 37806 12940 41200
rect 13084 40112 13136 40118
rect 13084 40054 13136 40060
rect 12992 39908 13044 39914
rect 12992 39850 13044 39856
rect 13004 38962 13032 39850
rect 12992 38956 13044 38962
rect 12992 38898 13044 38904
rect 13096 38758 13124 40054
rect 13556 38894 13584 41200
rect 13912 40724 13964 40730
rect 13912 40666 13964 40672
rect 13176 38888 13228 38894
rect 13176 38830 13228 38836
rect 13544 38888 13596 38894
rect 13544 38830 13596 38836
rect 13084 38752 13136 38758
rect 13084 38694 13136 38700
rect 12990 38584 13046 38593
rect 13188 38554 13216 38830
rect 13268 38820 13320 38826
rect 13268 38762 13320 38768
rect 13360 38820 13412 38826
rect 13360 38762 13412 38768
rect 12990 38519 12992 38528
rect 13044 38519 13046 38528
rect 13176 38548 13228 38554
rect 12992 38490 13044 38496
rect 13176 38490 13228 38496
rect 13280 38350 13308 38762
rect 13176 38344 13228 38350
rect 13176 38286 13228 38292
rect 13268 38344 13320 38350
rect 13268 38286 13320 38292
rect 13188 38214 13216 38286
rect 13176 38208 13228 38214
rect 13176 38150 13228 38156
rect 12990 38040 13046 38049
rect 12990 37975 13046 37984
rect 13004 37806 13032 37975
rect 11992 37624 12296 37652
rect 12452 37760 12756 37788
rect 12900 37800 12952 37806
rect 11428 37392 11480 37398
rect 11428 37334 11480 37340
rect 11520 37392 11572 37398
rect 11520 37334 11572 37340
rect 11440 36904 11468 37334
rect 11532 37097 11560 37334
rect 11980 37324 12032 37330
rect 12452 37312 12480 37760
rect 12900 37742 12952 37748
rect 12992 37800 13044 37806
rect 12992 37742 13044 37748
rect 12544 37454 13308 37482
rect 12544 37330 12572 37454
rect 12716 37392 12768 37398
rect 12768 37352 12848 37380
rect 12716 37334 12768 37340
rect 12032 37284 12480 37312
rect 12532 37324 12584 37330
rect 11980 37266 12032 37272
rect 12256 37188 12308 37194
rect 12256 37130 12308 37136
rect 12268 37097 12296 37130
rect 11518 37088 11574 37097
rect 11518 37023 11574 37032
rect 12254 37088 12310 37097
rect 12254 37023 12310 37032
rect 11440 36876 12112 36904
rect 12084 36836 12112 36876
rect 12164 36848 12216 36854
rect 11532 36808 11928 36836
rect 12084 36808 12164 36836
rect 11532 36802 11560 36808
rect 11440 36786 11560 36802
rect 11428 36780 11560 36786
rect 11480 36774 11560 36780
rect 11428 36722 11480 36728
rect 11520 36712 11572 36718
rect 11520 36654 11572 36660
rect 11428 35692 11480 35698
rect 11428 35634 11480 35640
rect 11440 35222 11468 35634
rect 11532 35494 11560 36654
rect 11612 36644 11664 36650
rect 11612 36586 11664 36592
rect 11624 36106 11652 36586
rect 11796 36576 11848 36582
rect 11796 36518 11848 36524
rect 11808 36242 11836 36518
rect 11796 36236 11848 36242
rect 11716 36196 11796 36224
rect 11612 36100 11664 36106
rect 11612 36042 11664 36048
rect 11610 36000 11666 36009
rect 11610 35935 11666 35944
rect 11520 35488 11572 35494
rect 11520 35430 11572 35436
rect 11624 35290 11652 35935
rect 11612 35284 11664 35290
rect 11612 35226 11664 35232
rect 11296 35164 11376 35170
rect 11244 35158 11376 35164
rect 11428 35216 11480 35222
rect 11428 35158 11480 35164
rect 11256 35142 11376 35158
rect 11256 35086 11284 35142
rect 11716 35136 11744 36196
rect 11796 36178 11848 36184
rect 11900 36009 11928 36808
rect 12164 36790 12216 36796
rect 12070 36680 12126 36689
rect 12360 36666 12388 37284
rect 12532 37266 12584 37272
rect 12438 37088 12494 37097
rect 12438 37023 12494 37032
rect 12452 36922 12480 37023
rect 12440 36916 12492 36922
rect 12440 36858 12492 36864
rect 12532 36916 12584 36922
rect 12532 36858 12584 36864
rect 12126 36638 12388 36666
rect 12070 36615 12126 36624
rect 12070 36544 12126 36553
rect 12070 36479 12126 36488
rect 11886 36000 11942 36009
rect 11886 35935 11942 35944
rect 11980 35828 12032 35834
rect 11980 35770 12032 35776
rect 11796 35624 11848 35630
rect 11796 35566 11848 35572
rect 11532 35108 11744 35136
rect 11244 35080 11296 35086
rect 11244 35022 11296 35028
rect 11336 35080 11388 35086
rect 11336 35022 11388 35028
rect 11152 35012 11204 35018
rect 11152 34954 11204 34960
rect 11244 34740 11296 34746
rect 11244 34682 11296 34688
rect 11256 34649 11284 34682
rect 11242 34640 11298 34649
rect 11060 34604 11112 34610
rect 11242 34575 11298 34584
rect 11060 34546 11112 34552
rect 10876 34468 10928 34474
rect 10796 34428 10876 34456
rect 10876 34410 10928 34416
rect 9404 34070 9456 34076
rect 9692 34088 9904 34116
rect 9968 34190 10272 34218
rect 9416 33998 9444 34070
rect 9312 33992 9364 33998
rect 9312 33934 9364 33940
rect 9404 33992 9456 33998
rect 9692 33969 9720 34088
rect 9968 34066 9996 34190
rect 10244 34134 10272 34190
rect 10232 34128 10284 34134
rect 10232 34070 10284 34076
rect 9956 34060 10008 34066
rect 9956 34002 10008 34008
rect 10048 33992 10100 33998
rect 9404 33934 9456 33940
rect 9678 33960 9734 33969
rect 9496 33924 9548 33930
rect 10048 33934 10100 33940
rect 10232 33992 10284 33998
rect 10416 33992 10468 33998
rect 10232 33934 10284 33940
rect 10414 33960 10416 33969
rect 10468 33960 10470 33969
rect 9678 33895 9734 33904
rect 9956 33924 10008 33930
rect 9496 33866 9548 33872
rect 9956 33866 10008 33872
rect 9508 33640 9536 33866
rect 9770 33824 9826 33833
rect 9826 33782 9904 33810
rect 9770 33759 9826 33768
rect 9508 33612 9720 33640
rect 9404 33516 9456 33522
rect 9588 33516 9640 33522
rect 9404 33458 9456 33464
rect 9508 33476 9588 33504
rect 9416 33153 9444 33458
rect 9402 33144 9458 33153
rect 9402 33079 9458 33088
rect 9508 33046 9536 33476
rect 9588 33458 9640 33464
rect 9496 33040 9548 33046
rect 9496 32982 9548 32988
rect 9692 32881 9720 33612
rect 9770 33008 9826 33017
rect 9770 32943 9826 32952
rect 9784 32910 9812 32943
rect 9876 32910 9904 33782
rect 9968 33658 9996 33866
rect 10060 33844 10088 33934
rect 10244 33844 10272 33934
rect 10520 33946 10548 34326
rect 10612 34218 10640 34342
rect 10704 34326 11100 34354
rect 11072 34241 11100 34326
rect 11058 34232 11114 34241
rect 10612 34190 10824 34218
rect 10796 34066 10824 34190
rect 11058 34167 11114 34176
rect 10968 34128 11020 34134
rect 10874 34096 10930 34105
rect 10784 34060 10836 34066
rect 10968 34070 11020 34076
rect 10874 34031 10930 34040
rect 10784 34002 10836 34008
rect 10888 33946 10916 34031
rect 10520 33918 10916 33946
rect 10414 33895 10470 33904
rect 10060 33816 10094 33844
rect 10244 33833 10640 33844
rect 10980 33833 11008 34070
rect 11152 33992 11204 33998
rect 11348 33980 11376 35022
rect 11532 34592 11560 35108
rect 11612 35012 11664 35018
rect 11612 34954 11664 34960
rect 11512 34564 11560 34592
rect 11428 34468 11480 34474
rect 11512 34456 11540 34564
rect 11480 34428 11540 34456
rect 11428 34410 11480 34416
rect 11512 34388 11540 34428
rect 11512 34360 11560 34388
rect 11204 33952 11376 33980
rect 11152 33934 11204 33940
rect 10244 33824 10654 33833
rect 10244 33816 10598 33824
rect 10066 33697 10094 33816
rect 10214 33756 10522 33776
rect 10598 33759 10654 33768
rect 10966 33824 11022 33833
rect 10966 33759 11022 33768
rect 10214 33754 10220 33756
rect 10276 33754 10300 33756
rect 10356 33754 10380 33756
rect 10436 33754 10460 33756
rect 10516 33754 10522 33756
rect 10276 33702 10278 33754
rect 10458 33702 10460 33754
rect 10214 33700 10220 33702
rect 10276 33700 10300 33702
rect 10356 33700 10380 33702
rect 10436 33700 10460 33702
rect 10516 33700 10522 33702
rect 10046 33688 10102 33697
rect 9956 33652 10008 33658
rect 10214 33680 10522 33700
rect 10598 33688 10654 33697
rect 10046 33623 10102 33632
rect 10336 33632 10598 33640
rect 11428 33652 11480 33658
rect 10336 33623 10654 33632
rect 9956 33594 10008 33600
rect 10336 33612 10640 33623
rect 10796 33612 11284 33640
rect 10048 33516 10100 33522
rect 10048 33458 10100 33464
rect 10060 33425 10088 33458
rect 10046 33416 10102 33425
rect 10046 33351 10102 33360
rect 10048 33312 10100 33318
rect 10336 33289 10364 33612
rect 10414 33552 10470 33561
rect 10414 33487 10470 33496
rect 10600 33516 10652 33522
rect 10428 33454 10456 33487
rect 10600 33458 10652 33464
rect 10416 33448 10468 33454
rect 10416 33390 10468 33396
rect 10612 33386 10640 33458
rect 10508 33380 10560 33386
rect 10508 33322 10560 33328
rect 10600 33380 10652 33386
rect 10600 33322 10652 33328
rect 10048 33254 10100 33260
rect 10322 33280 10378 33289
rect 9772 32904 9824 32910
rect 9678 32872 9734 32881
rect 9772 32846 9824 32852
rect 9864 32904 9916 32910
rect 9916 32864 9996 32892
rect 9864 32846 9916 32852
rect 9678 32807 9734 32816
rect 9496 32768 9548 32774
rect 9496 32710 9548 32716
rect 9508 32502 9536 32710
rect 9496 32496 9548 32502
rect 9864 32496 9916 32502
rect 9496 32438 9548 32444
rect 9770 32464 9826 32473
rect 9864 32438 9916 32444
rect 9770 32399 9826 32408
rect 9680 32292 9732 32298
rect 9784 32280 9812 32399
rect 9732 32252 9812 32280
rect 9680 32234 9732 32240
rect 9312 32224 9364 32230
rect 9312 32166 9364 32172
rect 9324 31890 9352 32166
rect 9416 32014 9812 32042
rect 9416 31958 9444 32014
rect 9404 31952 9456 31958
rect 9404 31894 9456 31900
rect 9312 31884 9364 31890
rect 9312 31826 9364 31832
rect 9404 31816 9456 31822
rect 9404 31758 9456 31764
rect 9588 31816 9640 31822
rect 9588 31758 9640 31764
rect 9312 31748 9364 31754
rect 9312 31690 9364 31696
rect 9324 30870 9352 31690
rect 9416 31657 9444 31758
rect 9402 31648 9458 31657
rect 9402 31583 9458 31592
rect 9600 31278 9628 31758
rect 9680 31680 9732 31686
rect 9680 31622 9732 31628
rect 9784 31634 9812 32014
rect 9876 32008 9904 32438
rect 9968 32178 9996 32864
rect 10060 32756 10088 33254
rect 10520 33266 10548 33322
rect 10796 33266 10824 33612
rect 10876 33516 10928 33522
rect 10876 33458 10928 33464
rect 11060 33516 11112 33522
rect 11060 33458 11112 33464
rect 10520 33238 10824 33266
rect 10322 33215 10378 33224
rect 10888 33153 10916 33458
rect 11072 33289 11100 33458
rect 11256 33318 11284 33612
rect 11428 33594 11480 33600
rect 11440 33561 11468 33594
rect 11426 33552 11482 33561
rect 11426 33487 11482 33496
rect 11244 33312 11296 33318
rect 11058 33280 11114 33289
rect 11244 33254 11296 33260
rect 11058 33215 11114 33224
rect 10874 33144 10930 33153
rect 10600 33108 10652 33114
rect 10600 33050 10652 33056
rect 10692 33108 10744 33114
rect 10874 33079 10930 33088
rect 10692 33050 10744 33056
rect 10612 32910 10640 33050
rect 10140 32904 10192 32910
rect 10324 32904 10376 32910
rect 10192 32864 10324 32892
rect 10140 32846 10192 32852
rect 10324 32846 10376 32852
rect 10600 32904 10652 32910
rect 10600 32846 10652 32852
rect 10060 32728 10640 32756
rect 10214 32668 10522 32688
rect 10214 32666 10220 32668
rect 10276 32666 10300 32668
rect 10356 32666 10380 32668
rect 10436 32666 10460 32668
rect 10516 32666 10522 32668
rect 10276 32614 10278 32666
rect 10458 32614 10460 32666
rect 10214 32612 10220 32614
rect 10276 32612 10300 32614
rect 10356 32612 10380 32614
rect 10436 32612 10460 32614
rect 10516 32612 10522 32614
rect 10214 32592 10522 32612
rect 10048 32496 10100 32502
rect 10324 32496 10376 32502
rect 10100 32456 10272 32484
rect 10048 32438 10100 32444
rect 10244 32178 10272 32456
rect 10324 32438 10376 32444
rect 10336 32298 10364 32438
rect 10416 32360 10468 32366
rect 10416 32302 10468 32308
rect 10612 32314 10640 32728
rect 10704 32434 10732 33050
rect 10784 33040 10836 33046
rect 10784 32982 10836 32988
rect 10796 32824 10824 32982
rect 10876 32972 10928 32978
rect 10928 32932 11100 32960
rect 10876 32914 10928 32920
rect 11072 32881 11100 32932
rect 11532 32910 11560 34360
rect 11624 33114 11652 34954
rect 11704 34128 11756 34134
rect 11702 34096 11704 34105
rect 11756 34096 11758 34105
rect 11702 34031 11758 34040
rect 11612 33108 11664 33114
rect 11612 33050 11664 33056
rect 11520 32904 11572 32910
rect 11058 32872 11114 32881
rect 10796 32796 11008 32824
rect 11520 32846 11572 32852
rect 11336 32836 11388 32842
rect 11058 32807 11114 32816
rect 10692 32428 10744 32434
rect 10692 32370 10744 32376
rect 10784 32428 10836 32434
rect 10784 32370 10836 32376
rect 10796 32314 10824 32370
rect 10324 32292 10376 32298
rect 10324 32234 10376 32240
rect 9968 32150 10180 32178
rect 10244 32150 10364 32178
rect 9876 31980 10088 32008
rect 9954 31920 10010 31929
rect 9954 31855 10010 31864
rect 9968 31754 9996 31855
rect 10060 31754 10088 31980
rect 10152 31822 10180 32150
rect 10336 32026 10364 32150
rect 10232 32020 10284 32026
rect 10232 31962 10284 31968
rect 10324 32020 10376 32026
rect 10324 31962 10376 31968
rect 10244 31906 10272 31962
rect 10244 31878 10364 31906
rect 10336 31822 10364 31878
rect 10140 31816 10192 31822
rect 10140 31758 10192 31764
rect 10324 31816 10376 31822
rect 10324 31758 10376 31764
rect 9956 31748 10008 31754
rect 9956 31690 10008 31696
rect 10048 31748 10100 31754
rect 10048 31690 10100 31696
rect 10428 31668 10456 32302
rect 10612 32286 10824 32314
rect 10796 31872 10824 32286
rect 10980 32212 11008 32796
rect 11164 32796 11336 32824
rect 11164 32366 11192 32796
rect 11336 32778 11388 32784
rect 11242 32736 11298 32745
rect 11242 32671 11298 32680
rect 11152 32360 11204 32366
rect 11152 32302 11204 32308
rect 11060 32224 11112 32230
rect 10980 32184 11060 32212
rect 11060 32166 11112 32172
rect 11256 32042 11284 32671
rect 11532 32366 11560 32846
rect 11704 32836 11756 32842
rect 11624 32796 11704 32824
rect 11520 32360 11572 32366
rect 11520 32302 11572 32308
rect 11624 32178 11652 32796
rect 11704 32778 11756 32784
rect 11808 32745 11836 35566
rect 11992 35018 12020 35770
rect 12084 35630 12112 36479
rect 12544 36292 12572 36858
rect 12624 36848 12676 36854
rect 12624 36790 12676 36796
rect 12176 36264 12572 36292
rect 12176 36038 12204 36264
rect 12254 36136 12310 36145
rect 12636 36122 12664 36790
rect 12714 36408 12770 36417
rect 12714 36343 12770 36352
rect 12254 36071 12310 36080
rect 12360 36094 12664 36122
rect 12164 36032 12216 36038
rect 12164 35974 12216 35980
rect 12162 35864 12218 35873
rect 12162 35799 12218 35808
rect 12176 35630 12204 35799
rect 12268 35698 12296 36071
rect 12360 35834 12388 36094
rect 12440 36032 12492 36038
rect 12440 35974 12492 35980
rect 12348 35828 12400 35834
rect 12348 35770 12400 35776
rect 12256 35692 12308 35698
rect 12256 35634 12308 35640
rect 12348 35692 12400 35698
rect 12348 35634 12400 35640
rect 12072 35624 12124 35630
rect 12072 35566 12124 35572
rect 12164 35624 12216 35630
rect 12164 35566 12216 35572
rect 12162 35320 12218 35329
rect 12162 35255 12218 35264
rect 12176 35154 12204 35255
rect 12164 35148 12216 35154
rect 12164 35090 12216 35096
rect 12256 35080 12308 35086
rect 12256 35022 12308 35028
rect 11980 35012 12032 35018
rect 11980 34954 12032 34960
rect 11980 34740 12032 34746
rect 11980 34682 12032 34688
rect 11888 34672 11940 34678
rect 11888 34614 11940 34620
rect 11900 34134 11928 34614
rect 11992 34513 12020 34682
rect 12268 34513 12296 35022
rect 11978 34504 12034 34513
rect 11978 34439 12034 34448
rect 12254 34504 12310 34513
rect 12254 34439 12310 34448
rect 11888 34128 11940 34134
rect 11888 34070 11940 34076
rect 12072 34060 12124 34066
rect 12072 34002 12124 34008
rect 11980 33992 12032 33998
rect 11980 33934 12032 33940
rect 11888 33652 11940 33658
rect 11888 33594 11940 33600
rect 11900 33522 11928 33594
rect 11888 33516 11940 33522
rect 11888 33458 11940 33464
rect 11992 33134 12020 33934
rect 12084 33658 12112 34002
rect 12164 33992 12216 33998
rect 12164 33934 12216 33940
rect 12254 33960 12310 33969
rect 12072 33652 12124 33658
rect 12072 33594 12124 33600
rect 12176 33522 12204 33934
rect 12254 33895 12310 33904
rect 12164 33516 12216 33522
rect 12164 33458 12216 33464
rect 11992 33114 12112 33134
rect 11992 33108 12124 33114
rect 11992 33106 12072 33108
rect 12072 33050 12124 33056
rect 11980 33040 12032 33046
rect 11980 32982 12032 32988
rect 11794 32736 11850 32745
rect 11992 32722 12020 32982
rect 12084 32978 12112 33050
rect 12072 32972 12124 32978
rect 12072 32914 12124 32920
rect 11794 32671 11850 32680
rect 11900 32694 12020 32722
rect 10968 32020 11020 32026
rect 10968 31962 11020 31968
rect 11072 32014 11284 32042
rect 11348 32150 11652 32178
rect 10152 31640 10456 31668
rect 10704 31844 10824 31872
rect 9692 31414 9720 31622
rect 9784 31606 10088 31634
rect 9862 31512 9918 31521
rect 10060 31482 10088 31606
rect 9862 31447 9918 31456
rect 9956 31476 10008 31482
rect 9680 31408 9732 31414
rect 9680 31350 9732 31356
rect 9588 31272 9640 31278
rect 9876 31260 9904 31447
rect 9956 31418 10008 31424
rect 10048 31476 10100 31482
rect 10048 31418 10100 31424
rect 9968 31385 9996 31418
rect 9954 31376 10010 31385
rect 9954 31311 10010 31320
rect 10048 31272 10100 31278
rect 9876 31232 10048 31260
rect 9588 31214 9640 31220
rect 10048 31214 10100 31220
rect 9402 30968 9458 30977
rect 9402 30903 9458 30912
rect 9312 30864 9364 30870
rect 9312 30806 9364 30812
rect 9416 30734 9444 30903
rect 9404 30728 9456 30734
rect 9404 30670 9456 30676
rect 9404 30592 9456 30598
rect 9404 30534 9456 30540
rect 10046 30560 10102 30569
rect 9416 30326 9444 30534
rect 10046 30495 10102 30504
rect 9862 30424 9918 30433
rect 9680 30388 9732 30394
rect 9862 30359 9918 30368
rect 9680 30330 9732 30336
rect 9404 30320 9456 30326
rect 9404 30262 9456 30268
rect 9494 30288 9550 30297
rect 9494 30223 9550 30232
rect 9588 30252 9640 30258
rect 9232 30144 9444 30172
rect 9310 30016 9366 30025
rect 9310 29951 9366 29960
rect 9324 29850 9352 29951
rect 9416 29850 9444 30144
rect 9312 29844 9364 29850
rect 9312 29786 9364 29792
rect 9404 29844 9456 29850
rect 9404 29786 9456 29792
rect 9220 29572 9272 29578
rect 9220 29514 9272 29520
rect 9128 29504 9180 29510
rect 9128 29446 9180 29452
rect 9140 29073 9168 29446
rect 9232 29306 9260 29514
rect 9404 29504 9456 29510
rect 9404 29446 9456 29452
rect 9220 29300 9272 29306
rect 9220 29242 9272 29248
rect 9416 29209 9444 29446
rect 9402 29200 9458 29209
rect 9402 29135 9458 29144
rect 9126 29064 9182 29073
rect 9126 28999 9182 29008
rect 9508 28966 9536 30223
rect 9588 30194 9640 30200
rect 9128 28960 9180 28966
rect 9126 28928 9128 28937
rect 9496 28960 9548 28966
rect 9180 28928 9182 28937
rect 9496 28902 9548 28908
rect 9126 28863 9182 28872
rect 9034 28520 9090 28529
rect 9034 28455 9090 28464
rect 9220 28416 9272 28422
rect 9220 28358 9272 28364
rect 8942 27568 8998 27577
rect 8942 27503 8998 27512
rect 9232 27130 9260 28358
rect 9496 28076 9548 28082
rect 9600 28064 9628 30194
rect 9692 29578 9720 30330
rect 9680 29572 9732 29578
rect 9680 29514 9732 29520
rect 9770 29336 9826 29345
rect 9770 29271 9826 29280
rect 9680 28144 9732 28150
rect 9680 28086 9732 28092
rect 9548 28036 9628 28064
rect 9496 28018 9548 28024
rect 9508 27674 9536 28018
rect 9586 27704 9642 27713
rect 9496 27668 9548 27674
rect 9586 27639 9642 27648
rect 9496 27610 9548 27616
rect 9496 27464 9548 27470
rect 9494 27432 9496 27441
rect 9548 27432 9550 27441
rect 9494 27367 9550 27376
rect 9600 27334 9628 27639
rect 9692 27402 9720 28086
rect 9680 27396 9732 27402
rect 9680 27338 9732 27344
rect 9588 27328 9640 27334
rect 9588 27270 9640 27276
rect 9220 27124 9272 27130
rect 9220 27066 9272 27072
rect 9784 26926 9812 29271
rect 9772 26920 9824 26926
rect 9678 26888 9734 26897
rect 9772 26862 9824 26868
rect 9678 26823 9680 26832
rect 9732 26823 9734 26832
rect 9680 26794 9732 26800
rect 9036 26784 9088 26790
rect 9876 26772 9904 30359
rect 9954 30152 10010 30161
rect 9954 30087 10010 30096
rect 10060 30104 10088 30495
rect 10152 30326 10180 31640
rect 10214 31580 10522 31600
rect 10214 31578 10220 31580
rect 10276 31578 10300 31580
rect 10356 31578 10380 31580
rect 10436 31578 10460 31580
rect 10516 31578 10522 31580
rect 10276 31526 10278 31578
rect 10458 31526 10460 31578
rect 10214 31524 10220 31526
rect 10276 31524 10300 31526
rect 10356 31524 10380 31526
rect 10436 31524 10460 31526
rect 10516 31524 10522 31526
rect 10214 31504 10522 31524
rect 10232 31408 10284 31414
rect 10232 31350 10284 31356
rect 10244 31142 10272 31350
rect 10336 31334 10548 31362
rect 10704 31346 10732 31844
rect 10782 31784 10838 31793
rect 10782 31719 10784 31728
rect 10836 31719 10838 31728
rect 10784 31690 10836 31696
rect 10980 31346 11008 31962
rect 10336 31210 10364 31334
rect 10416 31272 10468 31278
rect 10416 31214 10468 31220
rect 10324 31204 10376 31210
rect 10324 31146 10376 31152
rect 10428 31142 10456 31214
rect 10520 31210 10548 31334
rect 10692 31340 10744 31346
rect 10692 31282 10744 31288
rect 10968 31340 11020 31346
rect 10968 31282 11020 31288
rect 10508 31204 10560 31210
rect 10508 31146 10560 31152
rect 10232 31136 10284 31142
rect 10232 31078 10284 31084
rect 10416 31136 10468 31142
rect 10874 31104 10930 31113
rect 10416 31078 10468 31084
rect 10704 31062 10874 31090
rect 10704 30802 10732 31062
rect 10874 31039 10930 31048
rect 10508 30796 10560 30802
rect 10508 30738 10560 30744
rect 10692 30796 10744 30802
rect 10692 30738 10744 30744
rect 10520 30682 10548 30738
rect 10876 30728 10928 30734
rect 10782 30696 10838 30705
rect 10520 30654 10782 30682
rect 10876 30670 10928 30676
rect 10782 30631 10838 30640
rect 10214 30492 10522 30512
rect 10214 30490 10220 30492
rect 10276 30490 10300 30492
rect 10356 30490 10380 30492
rect 10436 30490 10460 30492
rect 10516 30490 10522 30492
rect 10276 30438 10278 30490
rect 10458 30438 10460 30490
rect 10214 30436 10220 30438
rect 10276 30436 10300 30438
rect 10356 30436 10380 30438
rect 10436 30436 10460 30438
rect 10516 30436 10522 30438
rect 10214 30416 10522 30436
rect 10600 30388 10652 30394
rect 10888 30376 10916 30670
rect 10652 30348 10916 30376
rect 10600 30330 10652 30336
rect 10140 30320 10192 30326
rect 10140 30262 10192 30268
rect 10508 30320 10560 30326
rect 10508 30262 10560 30268
rect 10324 30116 10376 30122
rect 9968 30054 9996 30087
rect 10060 30076 10324 30104
rect 10324 30058 10376 30064
rect 9956 30048 10008 30054
rect 9956 29990 10008 29996
rect 10520 29850 10548 30262
rect 10416 29844 10468 29850
rect 10416 29786 10468 29792
rect 10508 29844 10560 29850
rect 10508 29786 10560 29792
rect 10428 29646 10456 29786
rect 10140 29640 10192 29646
rect 10140 29582 10192 29588
rect 10416 29640 10468 29646
rect 10784 29640 10836 29646
rect 10416 29582 10468 29588
rect 10704 29600 10784 29628
rect 10152 29492 10180 29582
rect 10152 29464 10640 29492
rect 10214 29404 10522 29424
rect 10214 29402 10220 29404
rect 10276 29402 10300 29404
rect 10356 29402 10380 29404
rect 10436 29402 10460 29404
rect 10516 29402 10522 29404
rect 10276 29350 10278 29402
rect 10458 29350 10460 29402
rect 10214 29348 10220 29350
rect 10276 29348 10300 29350
rect 10356 29348 10380 29350
rect 10436 29348 10460 29350
rect 10516 29348 10522 29350
rect 10214 29328 10522 29348
rect 10612 29345 10640 29464
rect 10598 29336 10654 29345
rect 10704 29306 10732 29600
rect 10784 29582 10836 29588
rect 10784 29504 10836 29510
rect 10784 29446 10836 29452
rect 10874 29472 10930 29481
rect 10796 29306 10824 29446
rect 10874 29407 10930 29416
rect 10598 29271 10654 29280
rect 10692 29300 10744 29306
rect 10692 29242 10744 29248
rect 10784 29300 10836 29306
rect 10784 29242 10836 29248
rect 10888 29238 10916 29407
rect 10876 29232 10928 29238
rect 10876 29174 10928 29180
rect 10048 29164 10100 29170
rect 10048 29106 10100 29112
rect 10232 29164 10284 29170
rect 10232 29106 10284 29112
rect 10416 29164 10468 29170
rect 10416 29106 10468 29112
rect 10508 29164 10560 29170
rect 10508 29106 10560 29112
rect 9954 28792 10010 28801
rect 9954 28727 10010 28736
rect 9968 28082 9996 28727
rect 10060 28665 10088 29106
rect 10140 28960 10192 28966
rect 10140 28902 10192 28908
rect 10046 28656 10102 28665
rect 10046 28591 10102 28600
rect 10048 28552 10100 28558
rect 10048 28494 10100 28500
rect 9956 28076 10008 28082
rect 9956 28018 10008 28024
rect 9968 27282 9996 28018
rect 10060 27985 10088 28494
rect 10046 27976 10102 27985
rect 10046 27911 10102 27920
rect 10152 27849 10180 28902
rect 10244 28626 10272 29106
rect 10232 28620 10284 28626
rect 10232 28562 10284 28568
rect 10428 28472 10456 29106
rect 10520 28801 10548 29106
rect 10506 28792 10562 28801
rect 10506 28727 10562 28736
rect 10600 28756 10652 28762
rect 10876 28756 10928 28762
rect 10652 28716 10876 28744
rect 10600 28698 10652 28704
rect 10876 28698 10928 28704
rect 10600 28620 10652 28626
rect 10652 28580 10916 28608
rect 10600 28562 10652 28568
rect 10692 28484 10744 28490
rect 10428 28444 10640 28472
rect 10612 28370 10640 28444
rect 10744 28444 10824 28472
rect 10692 28426 10744 28432
rect 10612 28342 10732 28370
rect 10214 28316 10522 28336
rect 10214 28314 10220 28316
rect 10276 28314 10300 28316
rect 10356 28314 10380 28316
rect 10436 28314 10460 28316
rect 10516 28314 10522 28316
rect 10276 28262 10278 28314
rect 10458 28262 10460 28314
rect 10214 28260 10220 28262
rect 10276 28260 10300 28262
rect 10356 28260 10380 28262
rect 10436 28260 10460 28262
rect 10516 28260 10522 28262
rect 10214 28240 10522 28260
rect 10598 27976 10654 27985
rect 10598 27911 10654 27920
rect 10138 27840 10194 27849
rect 10138 27775 10194 27784
rect 10140 27464 10192 27470
rect 10140 27406 10192 27412
rect 9968 27254 10088 27282
rect 9956 26920 10008 26926
rect 9956 26862 10008 26868
rect 9036 26726 9088 26732
rect 9784 26744 9904 26772
rect 9048 26353 9076 26726
rect 9588 26376 9640 26382
rect 9034 26344 9090 26353
rect 9588 26318 9640 26324
rect 9034 26279 9090 26288
rect 7838 24848 7894 24857
rect 7838 24783 7894 24792
rect 9496 23724 9548 23730
rect 9496 23666 9548 23672
rect 9508 23254 9536 23666
rect 9496 23248 9548 23254
rect 9496 23190 9548 23196
rect 7746 16552 7802 16561
rect 7746 16487 7802 16496
rect 9600 16153 9628 26318
rect 9784 24426 9812 26744
rect 9864 26376 9916 26382
rect 9864 26318 9916 26324
rect 9692 24398 9812 24426
rect 9692 22094 9720 24398
rect 9692 22066 9812 22094
rect 9586 16144 9642 16153
rect 9586 16079 9642 16088
rect 5582 15804 5890 15824
rect 5582 15802 5588 15804
rect 5644 15802 5668 15804
rect 5724 15802 5748 15804
rect 5804 15802 5828 15804
rect 5884 15802 5890 15804
rect 5644 15750 5646 15802
rect 5826 15750 5828 15802
rect 5582 15748 5588 15750
rect 5644 15748 5668 15750
rect 5724 15748 5748 15750
rect 5804 15748 5828 15750
rect 5884 15748 5890 15750
rect 5582 15728 5890 15748
rect 5582 14716 5890 14736
rect 5582 14714 5588 14716
rect 5644 14714 5668 14716
rect 5724 14714 5748 14716
rect 5804 14714 5828 14716
rect 5884 14714 5890 14716
rect 5644 14662 5646 14714
rect 5826 14662 5828 14714
rect 5582 14660 5588 14662
rect 5644 14660 5668 14662
rect 5724 14660 5748 14662
rect 5804 14660 5828 14662
rect 5884 14660 5890 14662
rect 5582 14640 5890 14660
rect 7656 14476 7708 14482
rect 7656 14418 7708 14424
rect 5582 13628 5890 13648
rect 5582 13626 5588 13628
rect 5644 13626 5668 13628
rect 5724 13626 5748 13628
rect 5804 13626 5828 13628
rect 5884 13626 5890 13628
rect 5644 13574 5646 13626
rect 5826 13574 5828 13626
rect 5582 13572 5588 13574
rect 5644 13572 5668 13574
rect 5724 13572 5748 13574
rect 5804 13572 5828 13574
rect 5884 13572 5890 13574
rect 5582 13552 5890 13572
rect 5582 12540 5890 12560
rect 5582 12538 5588 12540
rect 5644 12538 5668 12540
rect 5724 12538 5748 12540
rect 5804 12538 5828 12540
rect 5884 12538 5890 12540
rect 5644 12486 5646 12538
rect 5826 12486 5828 12538
rect 5582 12484 5588 12486
rect 5644 12484 5668 12486
rect 5724 12484 5748 12486
rect 5804 12484 5828 12486
rect 5884 12484 5890 12486
rect 5582 12464 5890 12484
rect 7288 11756 7340 11762
rect 7288 11698 7340 11704
rect 5582 11452 5890 11472
rect 5582 11450 5588 11452
rect 5644 11450 5668 11452
rect 5724 11450 5748 11452
rect 5804 11450 5828 11452
rect 5884 11450 5890 11452
rect 5644 11398 5646 11450
rect 5826 11398 5828 11450
rect 5582 11396 5588 11398
rect 5644 11396 5668 11398
rect 5724 11396 5748 11398
rect 5804 11396 5828 11398
rect 5884 11396 5890 11398
rect 5582 11376 5890 11396
rect 5582 10364 5890 10384
rect 5582 10362 5588 10364
rect 5644 10362 5668 10364
rect 5724 10362 5748 10364
rect 5804 10362 5828 10364
rect 5884 10362 5890 10364
rect 5644 10310 5646 10362
rect 5826 10310 5828 10362
rect 5582 10308 5588 10310
rect 5644 10308 5668 10310
rect 5724 10308 5748 10310
rect 5804 10308 5828 10310
rect 5884 10308 5890 10310
rect 5582 10288 5890 10308
rect 5448 9648 5500 9654
rect 5448 9590 5500 9596
rect 5460 8498 5488 9590
rect 5582 9276 5890 9296
rect 5582 9274 5588 9276
rect 5644 9274 5668 9276
rect 5724 9274 5748 9276
rect 5804 9274 5828 9276
rect 5884 9274 5890 9276
rect 5644 9222 5646 9274
rect 5826 9222 5828 9274
rect 5582 9220 5588 9222
rect 5644 9220 5668 9222
rect 5724 9220 5748 9222
rect 5804 9220 5828 9222
rect 5884 9220 5890 9222
rect 5582 9200 5890 9220
rect 5448 8492 5500 8498
rect 5448 8434 5500 8440
rect 5582 8188 5890 8208
rect 5582 8186 5588 8188
rect 5644 8186 5668 8188
rect 5724 8186 5748 8188
rect 5804 8186 5828 8188
rect 5884 8186 5890 8188
rect 5644 8134 5646 8186
rect 5826 8134 5828 8186
rect 5582 8132 5588 8134
rect 5644 8132 5668 8134
rect 5724 8132 5748 8134
rect 5804 8132 5828 8134
rect 5884 8132 5890 8134
rect 5582 8112 5890 8132
rect 5582 7100 5890 7120
rect 5582 7098 5588 7100
rect 5644 7098 5668 7100
rect 5724 7098 5748 7100
rect 5804 7098 5828 7100
rect 5884 7098 5890 7100
rect 5644 7046 5646 7098
rect 5826 7046 5828 7098
rect 5582 7044 5588 7046
rect 5644 7044 5668 7046
rect 5724 7044 5748 7046
rect 5804 7044 5828 7046
rect 5884 7044 5890 7046
rect 5582 7024 5890 7044
rect 4712 6452 4764 6458
rect 4712 6394 4764 6400
rect 4436 6248 4488 6254
rect 4436 6190 4488 6196
rect 4528 6248 4580 6254
rect 4528 6190 4580 6196
rect 4160 5704 4212 5710
rect 4160 5646 4212 5652
rect 3884 5568 3936 5574
rect 3884 5510 3936 5516
rect 3896 5302 3924 5510
rect 3884 5296 3936 5302
rect 3884 5238 3936 5244
rect 4436 5092 4488 5098
rect 4436 5034 4488 5040
rect 4252 5024 4304 5030
rect 4252 4966 4304 4972
rect 3056 4616 3108 4622
rect 3056 4558 3108 4564
rect 3068 3534 3096 4558
rect 4066 4176 4122 4185
rect 4122 4134 4200 4162
rect 4066 4111 4122 4120
rect 4172 4078 4200 4134
rect 4160 4072 4212 4078
rect 4160 4014 4212 4020
rect 3332 3664 3384 3670
rect 3332 3606 3384 3612
rect 3056 3528 3108 3534
rect 2962 3496 3018 3505
rect 3056 3470 3108 3476
rect 2962 3431 3018 3440
rect 2504 3120 2556 3126
rect 2504 3062 2556 3068
rect 2596 3120 2648 3126
rect 2596 3062 2648 3068
rect 2596 2984 2648 2990
rect 2596 2926 2648 2932
rect 1584 2848 1636 2854
rect 1584 2790 1636 2796
rect 1596 2514 1624 2790
rect 1584 2508 1636 2514
rect 1584 2450 1636 2456
rect 2608 800 2636 2926
rect 3068 2922 3096 3470
rect 3240 3460 3292 3466
rect 3240 3402 3292 3408
rect 3056 2916 3108 2922
rect 3056 2858 3108 2864
rect 2778 2816 2834 2825
rect 2778 2751 2834 2760
rect 2792 2514 2820 2751
rect 2780 2508 2832 2514
rect 2780 2450 2832 2456
rect 3252 2145 3280 3402
rect 3238 2136 3294 2145
rect 3238 2071 3294 2080
rect 3344 1986 3372 3606
rect 3884 3460 3936 3466
rect 3884 3402 3936 3408
rect 3252 1958 3372 1986
rect 3056 1828 3108 1834
rect 3056 1770 3108 1776
rect 3068 1465 3096 1770
rect 3054 1456 3110 1465
rect 3054 1391 3110 1400
rect 3252 800 3280 1958
rect 3896 800 3924 3402
rect 4264 3194 4292 4966
rect 4344 4548 4396 4554
rect 4344 4490 4396 4496
rect 4356 3670 4384 4490
rect 4344 3664 4396 3670
rect 4344 3606 4396 3612
rect 4252 3188 4304 3194
rect 4252 3130 4304 3136
rect 4448 3058 4476 5034
rect 4540 3466 4568 6190
rect 5582 6012 5890 6032
rect 5582 6010 5588 6012
rect 5644 6010 5668 6012
rect 5724 6010 5748 6012
rect 5804 6010 5828 6012
rect 5884 6010 5890 6012
rect 5644 5958 5646 6010
rect 5826 5958 5828 6010
rect 5582 5956 5588 5958
rect 5644 5956 5668 5958
rect 5724 5956 5748 5958
rect 5804 5956 5828 5958
rect 5884 5956 5890 5958
rect 5582 5936 5890 5956
rect 5356 5772 5408 5778
rect 5356 5714 5408 5720
rect 4620 5704 4672 5710
rect 4620 5646 4672 5652
rect 4528 3460 4580 3466
rect 4528 3402 4580 3408
rect 4436 3052 4488 3058
rect 4436 2994 4488 3000
rect 4160 2848 4212 2854
rect 4160 2790 4212 2796
rect 4172 2514 4200 2790
rect 4632 2582 4660 5646
rect 5080 5092 5132 5098
rect 5080 5034 5132 5040
rect 5092 4214 5120 5034
rect 5172 5024 5224 5030
rect 5172 4966 5224 4972
rect 5080 4208 5132 4214
rect 5080 4150 5132 4156
rect 5184 3942 5212 4966
rect 5172 3936 5224 3942
rect 5172 3878 5224 3884
rect 5368 3602 5396 5714
rect 6368 5704 6420 5710
rect 6368 5646 6420 5652
rect 6552 5704 6604 5710
rect 6552 5646 6604 5652
rect 5908 5024 5960 5030
rect 5908 4966 5960 4972
rect 5582 4924 5890 4944
rect 5582 4922 5588 4924
rect 5644 4922 5668 4924
rect 5724 4922 5748 4924
rect 5804 4922 5828 4924
rect 5884 4922 5890 4924
rect 5644 4870 5646 4922
rect 5826 4870 5828 4922
rect 5582 4868 5588 4870
rect 5644 4868 5668 4870
rect 5724 4868 5748 4870
rect 5804 4868 5828 4870
rect 5884 4868 5890 4870
rect 5582 4848 5890 4868
rect 5582 3836 5890 3856
rect 5582 3834 5588 3836
rect 5644 3834 5668 3836
rect 5724 3834 5748 3836
rect 5804 3834 5828 3836
rect 5884 3834 5890 3836
rect 5644 3782 5646 3834
rect 5826 3782 5828 3834
rect 5582 3780 5588 3782
rect 5644 3780 5668 3782
rect 5724 3780 5748 3782
rect 5804 3780 5828 3782
rect 5884 3780 5890 3782
rect 5582 3760 5890 3780
rect 5920 3738 5948 4966
rect 6276 4616 6328 4622
rect 6276 4558 6328 4564
rect 5908 3732 5960 3738
rect 5908 3674 5960 3680
rect 5356 3596 5408 3602
rect 5356 3538 5408 3544
rect 5908 3596 5960 3602
rect 5908 3538 5960 3544
rect 5540 3460 5592 3466
rect 5540 3402 5592 3408
rect 5552 3194 5580 3402
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 5632 3188 5684 3194
rect 5632 3130 5684 3136
rect 5644 2990 5672 3130
rect 5632 2984 5684 2990
rect 5632 2926 5684 2932
rect 5582 2748 5890 2768
rect 5582 2746 5588 2748
rect 5644 2746 5668 2748
rect 5724 2746 5748 2748
rect 5804 2746 5828 2748
rect 5884 2746 5890 2748
rect 5644 2694 5646 2746
rect 5826 2694 5828 2746
rect 5582 2692 5588 2694
rect 5644 2692 5668 2694
rect 5724 2692 5748 2694
rect 5804 2692 5828 2694
rect 5884 2692 5890 2694
rect 5582 2672 5890 2692
rect 4620 2576 4672 2582
rect 4620 2518 4672 2524
rect 5172 2576 5224 2582
rect 5172 2518 5224 2524
rect 4160 2508 4212 2514
rect 4160 2450 4212 2456
rect 4528 2508 4580 2514
rect 4528 2450 4580 2456
rect 4540 800 4568 2450
rect 5184 800 5212 2518
rect 5920 1850 5948 3538
rect 6288 2650 6316 4558
rect 6276 2644 6328 2650
rect 6276 2586 6328 2592
rect 6380 2514 6408 5646
rect 6564 5370 6592 5646
rect 6552 5364 6604 5370
rect 6552 5306 6604 5312
rect 7196 5024 7248 5030
rect 7196 4966 7248 4972
rect 7208 4690 7236 4966
rect 7196 4684 7248 4690
rect 7196 4626 7248 4632
rect 7300 4622 7328 11698
rect 7288 4616 7340 4622
rect 7288 4558 7340 4564
rect 7380 4480 7432 4486
rect 7380 4422 7432 4428
rect 7392 4214 7420 4422
rect 7380 4208 7432 4214
rect 7380 4150 7432 4156
rect 6920 3936 6972 3942
rect 6920 3878 6972 3884
rect 6552 3392 6604 3398
rect 6552 3334 6604 3340
rect 6564 2514 6592 3334
rect 6932 3058 6960 3878
rect 7668 3534 7696 14418
rect 8668 6180 8720 6186
rect 8668 6122 8720 6128
rect 8116 4616 8168 4622
rect 8116 4558 8168 4564
rect 8128 4078 8156 4558
rect 8116 4072 8168 4078
rect 8116 4014 8168 4020
rect 7748 4004 7800 4010
rect 7748 3946 7800 3952
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 7104 3392 7156 3398
rect 7104 3334 7156 3340
rect 7116 3126 7144 3334
rect 7104 3120 7156 3126
rect 7104 3062 7156 3068
rect 6920 3052 6972 3058
rect 6920 2994 6972 3000
rect 7380 2984 7432 2990
rect 7380 2926 7432 2932
rect 6368 2508 6420 2514
rect 6368 2450 6420 2456
rect 6552 2508 6604 2514
rect 6552 2450 6604 2456
rect 5828 1822 5948 1850
rect 7392 1834 7420 2926
rect 7380 1828 7432 1834
rect 5828 800 5856 1822
rect 7380 1770 7432 1776
rect 7760 800 7788 3946
rect 8680 2922 8708 6122
rect 9036 4616 9088 4622
rect 9036 4558 9088 4564
rect 8668 2916 8720 2922
rect 8668 2858 8720 2864
rect 9048 2514 9076 4558
rect 9312 3936 9364 3942
rect 9312 3878 9364 3884
rect 9324 3602 9352 3878
rect 9312 3596 9364 3602
rect 9312 3538 9364 3544
rect 9680 3596 9732 3602
rect 9680 3538 9732 3544
rect 9128 2576 9180 2582
rect 9128 2518 9180 2524
rect 9036 2508 9088 2514
rect 9036 2450 9088 2456
rect 9140 1170 9168 2518
rect 9048 1142 9168 1170
rect 9048 800 9076 1142
rect 9692 800 9720 3538
rect 9784 3058 9812 22066
rect 9876 20806 9904 26318
rect 9864 20800 9916 20806
rect 9864 20742 9916 20748
rect 9968 14482 9996 26862
rect 10060 26738 10088 27254
rect 10152 27062 10180 27406
rect 10214 27228 10522 27248
rect 10214 27226 10220 27228
rect 10276 27226 10300 27228
rect 10356 27226 10380 27228
rect 10436 27226 10460 27228
rect 10516 27226 10522 27228
rect 10276 27174 10278 27226
rect 10458 27174 10460 27226
rect 10214 27172 10220 27174
rect 10276 27172 10300 27174
rect 10356 27172 10380 27174
rect 10436 27172 10460 27174
rect 10516 27172 10522 27174
rect 10214 27152 10522 27172
rect 10140 27056 10192 27062
rect 10140 26998 10192 27004
rect 10232 26784 10284 26790
rect 10060 26710 10180 26738
rect 10232 26726 10284 26732
rect 9956 14476 10008 14482
rect 9956 14418 10008 14424
rect 10152 11626 10180 26710
rect 10244 26625 10272 26726
rect 10230 26616 10286 26625
rect 10230 26551 10286 26560
rect 10214 26140 10522 26160
rect 10214 26138 10220 26140
rect 10276 26138 10300 26140
rect 10356 26138 10380 26140
rect 10436 26138 10460 26140
rect 10516 26138 10522 26140
rect 10276 26086 10278 26138
rect 10458 26086 10460 26138
rect 10214 26084 10220 26086
rect 10276 26084 10300 26086
rect 10356 26084 10380 26086
rect 10436 26084 10460 26086
rect 10516 26084 10522 26086
rect 10214 26064 10522 26084
rect 10612 25401 10640 27911
rect 10704 27614 10732 28342
rect 10796 28257 10824 28444
rect 10782 28248 10838 28257
rect 10782 28183 10838 28192
rect 10796 27690 10824 28183
rect 10888 27985 10916 28580
rect 10874 27976 10930 27985
rect 10874 27911 10930 27920
rect 10796 27674 10916 27690
rect 10796 27668 10928 27674
rect 10796 27662 10876 27668
rect 10704 27586 10824 27614
rect 10876 27610 10928 27616
rect 10796 27470 10824 27586
rect 10692 27464 10744 27470
rect 10692 27406 10744 27412
rect 10784 27464 10836 27470
rect 10836 27424 10916 27452
rect 10784 27406 10836 27412
rect 10704 26081 10732 27406
rect 10782 27024 10838 27033
rect 10782 26959 10784 26968
rect 10836 26959 10838 26968
rect 10784 26930 10836 26936
rect 10690 26072 10746 26081
rect 10690 26007 10746 26016
rect 10784 25900 10836 25906
rect 10784 25842 10836 25848
rect 10796 25673 10824 25842
rect 10782 25664 10838 25673
rect 10782 25599 10838 25608
rect 10598 25392 10654 25401
rect 10598 25327 10654 25336
rect 10600 25288 10652 25294
rect 10784 25288 10836 25294
rect 10600 25230 10652 25236
rect 10782 25256 10784 25265
rect 10836 25256 10838 25265
rect 10214 25052 10522 25072
rect 10214 25050 10220 25052
rect 10276 25050 10300 25052
rect 10356 25050 10380 25052
rect 10436 25050 10460 25052
rect 10516 25050 10522 25052
rect 10276 24998 10278 25050
rect 10458 24998 10460 25050
rect 10214 24996 10220 24998
rect 10276 24996 10300 24998
rect 10356 24996 10380 24998
rect 10436 24996 10460 24998
rect 10516 24996 10522 24998
rect 10214 24976 10522 24996
rect 10612 24886 10640 25230
rect 10782 25191 10838 25200
rect 10888 25140 10916 27424
rect 10980 27305 11008 31282
rect 11072 28801 11100 32014
rect 11152 31680 11204 31686
rect 11348 31668 11376 32150
rect 11520 32020 11572 32026
rect 11520 31962 11572 31968
rect 11532 31822 11560 31962
rect 11704 31952 11756 31958
rect 11900 31940 11928 32694
rect 12176 32502 12204 33458
rect 12268 32745 12296 33895
rect 12254 32736 12310 32745
rect 12254 32671 12310 32680
rect 12164 32496 12216 32502
rect 12164 32438 12216 32444
rect 11756 31912 11928 31940
rect 11704 31894 11756 31900
rect 11520 31816 11572 31822
rect 11426 31784 11482 31793
rect 11520 31758 11572 31764
rect 11704 31816 11756 31822
rect 11756 31776 11836 31804
rect 11704 31758 11756 31764
rect 11426 31719 11482 31728
rect 11204 31640 11376 31668
rect 11152 31622 11204 31628
rect 11336 31136 11388 31142
rect 11336 31078 11388 31084
rect 11348 30802 11376 31078
rect 11440 30977 11468 31719
rect 11704 31340 11756 31346
rect 11532 31300 11704 31328
rect 11426 30968 11482 30977
rect 11426 30903 11482 30912
rect 11336 30796 11388 30802
rect 11336 30738 11388 30744
rect 11532 30326 11560 31300
rect 11704 31282 11756 31288
rect 11702 31104 11758 31113
rect 11702 31039 11758 31048
rect 11612 30932 11664 30938
rect 11612 30874 11664 30880
rect 11624 30326 11652 30874
rect 11716 30433 11744 31039
rect 11702 30424 11758 30433
rect 11702 30359 11758 30368
rect 11520 30320 11572 30326
rect 11164 30246 11468 30274
rect 11520 30262 11572 30268
rect 11612 30320 11664 30326
rect 11612 30262 11664 30268
rect 11164 29646 11192 30246
rect 11244 30184 11296 30190
rect 11440 30172 11468 30246
rect 11440 30144 11744 30172
rect 11244 30126 11296 30132
rect 11152 29640 11204 29646
rect 11152 29582 11204 29588
rect 11058 28792 11114 28801
rect 11058 28727 11114 28736
rect 11072 28694 11100 28727
rect 11060 28688 11112 28694
rect 11060 28630 11112 28636
rect 11256 28626 11284 30126
rect 11336 30116 11388 30122
rect 11336 30058 11388 30064
rect 11348 29034 11376 30058
rect 11518 29744 11574 29753
rect 11518 29679 11574 29688
rect 11532 29646 11560 29679
rect 11716 29646 11744 30144
rect 11808 29646 11836 31776
rect 11978 31784 12034 31793
rect 12360 31754 12388 35634
rect 12452 34066 12480 35974
rect 12624 35760 12676 35766
rect 12624 35702 12676 35708
rect 12532 35080 12584 35086
rect 12532 35022 12584 35028
rect 12440 34060 12492 34066
rect 12440 34002 12492 34008
rect 12452 33844 12480 34002
rect 12544 33998 12572 35022
rect 12532 33992 12584 33998
rect 12532 33934 12584 33940
rect 12452 33816 12572 33844
rect 12440 33448 12492 33454
rect 12440 33390 12492 33396
rect 12452 32842 12480 33390
rect 12544 32892 12572 33816
rect 12636 33522 12664 35702
rect 12728 35494 12756 36343
rect 12820 35766 12848 37352
rect 12992 37324 13044 37330
rect 12992 37266 13044 37272
rect 12898 37088 12954 37097
rect 12898 37023 12954 37032
rect 12912 36394 12940 37023
rect 13004 36553 13032 37266
rect 13280 37126 13308 37454
rect 13084 37120 13136 37126
rect 13082 37088 13084 37097
rect 13268 37120 13320 37126
rect 13136 37088 13138 37097
rect 13268 37062 13320 37068
rect 13082 37023 13138 37032
rect 13372 36938 13400 38762
rect 13452 37800 13504 37806
rect 13452 37742 13504 37748
rect 13280 36910 13400 36938
rect 13280 36854 13308 36910
rect 13268 36848 13320 36854
rect 13268 36790 13320 36796
rect 13084 36644 13136 36650
rect 13084 36586 13136 36592
rect 12990 36544 13046 36553
rect 12990 36479 13046 36488
rect 12912 36366 13032 36394
rect 13004 36310 13032 36366
rect 12992 36304 13044 36310
rect 12992 36246 13044 36252
rect 12992 36168 13044 36174
rect 12992 36110 13044 36116
rect 12898 36000 12954 36009
rect 12898 35935 12954 35944
rect 12808 35760 12860 35766
rect 12808 35702 12860 35708
rect 12716 35488 12768 35494
rect 12808 35488 12860 35494
rect 12716 35430 12768 35436
rect 12806 35456 12808 35465
rect 12860 35456 12862 35465
rect 12806 35391 12862 35400
rect 12912 35170 12940 35935
rect 13004 35766 13032 36110
rect 12992 35760 13044 35766
rect 12992 35702 13044 35708
rect 13096 35698 13124 36586
rect 13464 36582 13492 37742
rect 13726 37496 13782 37505
rect 13726 37431 13782 37440
rect 13636 37256 13688 37262
rect 13636 37198 13688 37204
rect 13542 37088 13598 37097
rect 13542 37023 13598 37032
rect 13556 36786 13584 37023
rect 13544 36780 13596 36786
rect 13544 36722 13596 36728
rect 13648 36718 13676 37198
rect 13740 37194 13768 37431
rect 13728 37188 13780 37194
rect 13728 37130 13780 37136
rect 13636 36712 13688 36718
rect 13636 36654 13688 36660
rect 13452 36576 13504 36582
rect 13452 36518 13504 36524
rect 13542 36544 13598 36553
rect 13542 36479 13598 36488
rect 13556 36394 13584 36479
rect 13372 36366 13584 36394
rect 13636 36372 13688 36378
rect 13372 36156 13400 36366
rect 13636 36314 13688 36320
rect 13728 36372 13780 36378
rect 13728 36314 13780 36320
rect 13188 36128 13400 36156
rect 13084 35692 13136 35698
rect 13084 35634 13136 35640
rect 13082 35592 13138 35601
rect 13188 35578 13216 36128
rect 13648 36106 13676 36314
rect 13636 36100 13688 36106
rect 13636 36042 13688 36048
rect 13268 35760 13320 35766
rect 13636 35760 13688 35766
rect 13320 35720 13400 35748
rect 13268 35702 13320 35708
rect 13138 35550 13216 35578
rect 13266 35592 13322 35601
rect 13082 35527 13138 35536
rect 13266 35527 13268 35536
rect 13320 35527 13322 35536
rect 13268 35498 13320 35504
rect 13266 35456 13322 35465
rect 13266 35391 13322 35400
rect 12820 35142 12940 35170
rect 12992 35148 13044 35154
rect 12716 34196 12768 34202
rect 12716 34138 12768 34144
rect 12624 33516 12676 33522
rect 12624 33458 12676 33464
rect 12728 33454 12756 34138
rect 12820 33930 12848 35142
rect 12992 35090 13044 35096
rect 12900 35080 12952 35086
rect 12900 35022 12952 35028
rect 12912 34406 12940 35022
rect 13004 34950 13032 35090
rect 13280 35057 13308 35391
rect 13266 35048 13322 35057
rect 13266 34983 13322 34992
rect 12992 34944 13044 34950
rect 12992 34886 13044 34892
rect 13084 34944 13136 34950
rect 13084 34886 13136 34892
rect 13096 34678 13124 34886
rect 13084 34672 13136 34678
rect 13084 34614 13136 34620
rect 13372 34542 13400 35720
rect 13740 35748 13768 36314
rect 13924 36038 13952 40666
rect 14004 39908 14056 39914
rect 14004 39850 14056 39856
rect 14016 39370 14044 39850
rect 14096 39500 14148 39506
rect 14096 39442 14148 39448
rect 14004 39364 14056 39370
rect 14004 39306 14056 39312
rect 14108 38894 14136 39442
rect 14096 38888 14148 38894
rect 14096 38830 14148 38836
rect 14200 38593 14228 41200
rect 15382 40488 15438 40497
rect 15382 40423 15438 40432
rect 15290 40080 15346 40089
rect 15290 40015 15346 40024
rect 14280 39840 14332 39846
rect 15304 39817 15332 40015
rect 14280 39782 14332 39788
rect 14646 39808 14702 39817
rect 14292 39438 14320 39782
rect 15290 39808 15346 39817
rect 14646 39743 14702 39752
rect 14554 39672 14610 39681
rect 14554 39607 14610 39616
rect 14280 39432 14332 39438
rect 14280 39374 14332 39380
rect 14568 39370 14596 39607
rect 14464 39364 14516 39370
rect 14464 39306 14516 39312
rect 14556 39364 14608 39370
rect 14556 39306 14608 39312
rect 14370 39128 14426 39137
rect 14476 39098 14504 39306
rect 14660 39137 14688 39743
rect 14846 39740 15154 39760
rect 15290 39743 15346 39752
rect 14846 39738 14852 39740
rect 14908 39738 14932 39740
rect 14988 39738 15012 39740
rect 15068 39738 15092 39740
rect 15148 39738 15154 39740
rect 14908 39686 14910 39738
rect 15090 39686 15092 39738
rect 14846 39684 14852 39686
rect 14908 39684 14932 39686
rect 14988 39684 15012 39686
rect 15068 39684 15092 39686
rect 15148 39684 15154 39686
rect 14846 39664 15154 39684
rect 14646 39128 14702 39137
rect 14370 39063 14426 39072
rect 14464 39092 14516 39098
rect 14384 38978 14412 39063
rect 14464 39034 14516 39040
rect 14556 39092 14608 39098
rect 14646 39063 14702 39072
rect 15292 39092 15344 39098
rect 14556 39034 14608 39040
rect 15292 39034 15344 39040
rect 14568 38978 14596 39034
rect 14384 38950 14596 38978
rect 14648 38956 14700 38962
rect 14648 38898 14700 38904
rect 14660 38729 14688 38898
rect 15304 38729 15332 39034
rect 14646 38720 14702 38729
rect 15290 38720 15346 38729
rect 14646 38655 14702 38664
rect 14846 38652 15154 38672
rect 15290 38655 15346 38664
rect 14846 38650 14852 38652
rect 14908 38650 14932 38652
rect 14988 38650 15012 38652
rect 15068 38650 15092 38652
rect 15148 38650 15154 38652
rect 14908 38598 14910 38650
rect 15090 38598 15092 38650
rect 15396 38654 15424 40423
rect 15488 39506 15516 41200
rect 15936 40792 15988 40798
rect 15936 40734 15988 40740
rect 15568 39840 15620 39846
rect 15568 39782 15620 39788
rect 15476 39500 15528 39506
rect 15476 39442 15528 39448
rect 15476 39092 15528 39098
rect 15476 39034 15528 39040
rect 15488 38758 15516 39034
rect 15580 38962 15608 39782
rect 15660 39500 15712 39506
rect 15660 39442 15712 39448
rect 15672 39030 15700 39442
rect 15660 39024 15712 39030
rect 15660 38966 15712 38972
rect 15568 38956 15620 38962
rect 15568 38898 15620 38904
rect 15476 38752 15528 38758
rect 15476 38694 15528 38700
rect 15752 38752 15804 38758
rect 15752 38694 15804 38700
rect 15396 38626 15608 38654
rect 14846 38596 14852 38598
rect 14908 38596 14932 38598
rect 14988 38596 15012 38598
rect 15068 38596 15092 38598
rect 15148 38596 15154 38598
rect 14186 38584 14242 38593
rect 14846 38576 15154 38596
rect 15290 38584 15346 38593
rect 14186 38519 14242 38528
rect 15212 38542 15290 38570
rect 14740 38480 14792 38486
rect 14740 38422 14792 38428
rect 14752 38282 14780 38422
rect 15212 38400 15240 38542
rect 15290 38519 15346 38528
rect 15580 38418 15608 38626
rect 15764 38418 15792 38694
rect 15028 38372 15240 38400
rect 15384 38412 15436 38418
rect 14832 38344 14884 38350
rect 15028 38332 15056 38372
rect 15384 38354 15436 38360
rect 15568 38412 15620 38418
rect 15568 38354 15620 38360
rect 15752 38412 15804 38418
rect 15752 38354 15804 38360
rect 14884 38304 15056 38332
rect 14832 38286 14884 38292
rect 14740 38276 14792 38282
rect 14740 38218 14792 38224
rect 14372 37868 14424 37874
rect 14372 37810 14424 37816
rect 14188 37324 14240 37330
rect 14188 37266 14240 37272
rect 14096 37256 14148 37262
rect 14096 37198 14148 37204
rect 14004 36304 14056 36310
rect 14002 36272 14004 36281
rect 14056 36272 14058 36281
rect 14108 36242 14136 37198
rect 14002 36207 14058 36216
rect 14096 36236 14148 36242
rect 14096 36178 14148 36184
rect 14200 36174 14228 37266
rect 14384 36689 14412 37810
rect 14648 37800 14700 37806
rect 15396 37777 15424 38354
rect 15476 38344 15528 38350
rect 15476 38286 15528 38292
rect 14648 37742 14700 37748
rect 15198 37768 15254 37777
rect 14660 36922 14688 37742
rect 15198 37703 15254 37712
rect 15382 37768 15438 37777
rect 15382 37703 15438 37712
rect 15212 37670 15240 37703
rect 15200 37664 15252 37670
rect 15200 37606 15252 37612
rect 14846 37564 15154 37584
rect 14846 37562 14852 37564
rect 14908 37562 14932 37564
rect 14988 37562 15012 37564
rect 15068 37562 15092 37564
rect 15148 37562 15154 37564
rect 14908 37510 14910 37562
rect 15090 37510 15092 37562
rect 14846 37508 14852 37510
rect 14908 37508 14932 37510
rect 14988 37508 15012 37510
rect 15068 37508 15092 37510
rect 15148 37508 15154 37510
rect 14846 37488 15154 37508
rect 15488 37505 15516 38286
rect 15752 37800 15804 37806
rect 15752 37742 15804 37748
rect 15474 37496 15530 37505
rect 15474 37431 15530 37440
rect 15764 37126 15792 37742
rect 15752 37120 15804 37126
rect 15752 37062 15804 37068
rect 14648 36916 14700 36922
rect 14648 36858 14700 36864
rect 15016 36916 15068 36922
rect 15016 36858 15068 36864
rect 15476 36916 15528 36922
rect 15476 36858 15528 36864
rect 15028 36786 15056 36858
rect 15016 36780 15068 36786
rect 15016 36722 15068 36728
rect 14370 36680 14426 36689
rect 14370 36615 14426 36624
rect 14384 36378 14412 36615
rect 14462 36544 14518 36553
rect 14462 36479 14518 36488
rect 14476 36378 14504 36479
rect 14846 36476 15154 36496
rect 14846 36474 14852 36476
rect 14908 36474 14932 36476
rect 14988 36474 15012 36476
rect 15068 36474 15092 36476
rect 15148 36474 15154 36476
rect 14908 36422 14910 36474
rect 15090 36422 15092 36474
rect 14846 36420 14852 36422
rect 14908 36420 14932 36422
rect 14988 36420 15012 36422
rect 15068 36420 15092 36422
rect 15148 36420 15154 36422
rect 14646 36408 14702 36417
rect 14372 36372 14424 36378
rect 14372 36314 14424 36320
rect 14464 36372 14516 36378
rect 14846 36400 15154 36420
rect 15382 36408 15438 36417
rect 14646 36343 14702 36352
rect 15382 36343 15384 36352
rect 14464 36314 14516 36320
rect 14188 36168 14240 36174
rect 14188 36110 14240 36116
rect 13820 36032 13872 36038
rect 13820 35974 13872 35980
rect 13912 36032 13964 36038
rect 13912 35974 13964 35980
rect 13688 35720 13768 35748
rect 13636 35702 13688 35708
rect 13452 35692 13504 35698
rect 13504 35652 13584 35680
rect 13452 35634 13504 35640
rect 13452 35556 13504 35562
rect 13556 35544 13584 35652
rect 13636 35556 13688 35562
rect 13556 35516 13636 35544
rect 13452 35498 13504 35504
rect 13636 35498 13688 35504
rect 13464 35222 13492 35498
rect 13728 35488 13780 35494
rect 13728 35430 13780 35436
rect 13452 35216 13504 35222
rect 13452 35158 13504 35164
rect 13740 35057 13768 35430
rect 13726 35048 13782 35057
rect 13726 34983 13782 34992
rect 13832 34950 13860 35974
rect 13912 35828 13964 35834
rect 13912 35770 13964 35776
rect 13924 35465 13952 35770
rect 14200 35686 14320 35714
rect 14384 35698 14412 36314
rect 14556 36032 14608 36038
rect 14556 35974 14608 35980
rect 14200 35630 14228 35686
rect 14188 35624 14240 35630
rect 14188 35566 14240 35572
rect 14004 35488 14056 35494
rect 13910 35456 13966 35465
rect 14004 35430 14056 35436
rect 13910 35391 13966 35400
rect 13912 35080 13964 35086
rect 13910 35048 13912 35057
rect 13964 35048 13966 35057
rect 13910 34983 13966 34992
rect 13728 34944 13780 34950
rect 13728 34886 13780 34892
rect 13820 34944 13872 34950
rect 13820 34886 13872 34892
rect 13360 34536 13412 34542
rect 13360 34478 13412 34484
rect 12900 34400 12952 34406
rect 12900 34342 12952 34348
rect 12992 34400 13044 34406
rect 12992 34342 13044 34348
rect 12912 34202 12940 34342
rect 12900 34196 12952 34202
rect 12900 34138 12952 34144
rect 13004 34066 13032 34342
rect 12992 34060 13044 34066
rect 12992 34002 13044 34008
rect 12808 33924 12860 33930
rect 12808 33866 12860 33872
rect 12990 33688 13046 33697
rect 12990 33623 13046 33632
rect 13004 33590 13032 33623
rect 12992 33584 13044 33590
rect 12992 33526 13044 33532
rect 13372 33522 13400 34478
rect 13360 33516 13412 33522
rect 13412 33476 13676 33504
rect 13360 33458 13412 33464
rect 12716 33448 12768 33454
rect 12716 33390 12768 33396
rect 12900 33448 12952 33454
rect 12900 33390 12952 33396
rect 12992 33448 13044 33454
rect 12992 33390 13044 33396
rect 12912 33130 12940 33390
rect 13004 33289 13032 33390
rect 13360 33380 13412 33386
rect 13360 33322 13412 33328
rect 12990 33280 13046 33289
rect 12990 33215 13046 33224
rect 13266 33280 13322 33289
rect 13266 33215 13322 33224
rect 12912 33102 13124 33130
rect 13280 33114 13308 33215
rect 13372 33114 13400 33322
rect 13096 33046 13124 33102
rect 13268 33108 13320 33114
rect 13268 33050 13320 33056
rect 13360 33108 13412 33114
rect 13360 33050 13412 33056
rect 13084 33040 13136 33046
rect 12714 33008 12770 33017
rect 13084 32982 13136 32988
rect 12714 32943 12770 32952
rect 13648 32960 13676 33476
rect 13740 33402 13768 34886
rect 13912 34604 13964 34610
rect 13912 34546 13964 34552
rect 13924 34354 13952 34546
rect 14016 34377 14044 35430
rect 14096 35080 14148 35086
rect 14096 35022 14148 35028
rect 13832 34326 13952 34354
rect 14002 34368 14058 34377
rect 13832 33561 13860 34326
rect 14002 34303 14058 34312
rect 14108 34241 14136 35022
rect 13910 34232 13966 34241
rect 14094 34232 14150 34241
rect 13966 34190 14044 34218
rect 13910 34167 13966 34176
rect 13912 34128 13964 34134
rect 13912 34070 13964 34076
rect 13924 33998 13952 34070
rect 13912 33992 13964 33998
rect 13912 33934 13964 33940
rect 13818 33552 13874 33561
rect 14016 33522 14044 34190
rect 14094 34167 14150 34176
rect 14188 34196 14240 34202
rect 14108 34134 14136 34167
rect 14188 34138 14240 34144
rect 14096 34128 14148 34134
rect 14096 34070 14148 34076
rect 14200 33998 14228 34138
rect 14188 33992 14240 33998
rect 14188 33934 14240 33940
rect 14292 33980 14320 35686
rect 14372 35692 14424 35698
rect 14372 35634 14424 35640
rect 14384 35086 14412 35634
rect 14568 35601 14596 35974
rect 14554 35592 14610 35601
rect 14554 35527 14610 35536
rect 14660 35494 14688 36343
rect 15436 36343 15438 36352
rect 15384 36314 15436 36320
rect 15292 36304 15344 36310
rect 15292 36246 15344 36252
rect 15200 35828 15252 35834
rect 15200 35770 15252 35776
rect 14738 35592 14794 35601
rect 14738 35527 14794 35536
rect 14648 35488 14700 35494
rect 14648 35430 14700 35436
rect 14646 35320 14702 35329
rect 14752 35306 14780 35527
rect 14846 35388 15154 35408
rect 14846 35386 14852 35388
rect 14908 35386 14932 35388
rect 14988 35386 15012 35388
rect 15068 35386 15092 35388
rect 15148 35386 15154 35388
rect 14908 35334 14910 35386
rect 15090 35334 15092 35386
rect 14846 35332 14852 35334
rect 14908 35332 14932 35334
rect 14988 35332 15012 35334
rect 15068 35332 15092 35334
rect 15148 35332 15154 35334
rect 14846 35312 15154 35332
rect 14702 35278 14780 35306
rect 15212 35306 15240 35770
rect 15304 35698 15332 36246
rect 15292 35692 15344 35698
rect 15292 35634 15344 35640
rect 15488 35494 15516 36858
rect 15764 36786 15792 37062
rect 15568 36780 15620 36786
rect 15568 36722 15620 36728
rect 15752 36780 15804 36786
rect 15752 36722 15804 36728
rect 15844 36780 15896 36786
rect 15844 36722 15896 36728
rect 15580 35698 15608 36722
rect 15660 36236 15712 36242
rect 15660 36178 15712 36184
rect 15568 35692 15620 35698
rect 15568 35634 15620 35640
rect 15568 35556 15620 35562
rect 15568 35498 15620 35504
rect 15292 35488 15344 35494
rect 15290 35456 15292 35465
rect 15476 35488 15528 35494
rect 15344 35456 15346 35465
rect 15476 35430 15528 35436
rect 15290 35391 15346 35400
rect 15290 35320 15346 35329
rect 15212 35278 15290 35306
rect 14646 35255 14702 35264
rect 15290 35255 15346 35264
rect 15580 35222 15608 35498
rect 15568 35216 15620 35222
rect 14752 35142 15240 35170
rect 15568 35158 15620 35164
rect 15672 35154 15700 36178
rect 15764 35766 15792 36722
rect 15856 36310 15884 36722
rect 15948 36378 15976 40734
rect 16132 38418 16160 41200
rect 18064 40118 18092 41200
rect 19062 40352 19118 40361
rect 19062 40287 19118 40296
rect 16580 40112 16632 40118
rect 16580 40054 16632 40060
rect 18052 40112 18104 40118
rect 18052 40054 18104 40060
rect 18880 40112 18932 40118
rect 18880 40054 18932 40060
rect 16592 39914 16620 40054
rect 16948 40044 17000 40050
rect 16948 39986 17000 39992
rect 16580 39908 16632 39914
rect 16580 39850 16632 39856
rect 16672 39908 16724 39914
rect 16672 39850 16724 39856
rect 16684 39438 16712 39850
rect 16672 39432 16724 39438
rect 16672 39374 16724 39380
rect 16960 39030 16988 39986
rect 17038 39672 17094 39681
rect 17038 39607 17094 39616
rect 17500 39636 17552 39642
rect 17052 39409 17080 39607
rect 17500 39578 17552 39584
rect 17038 39400 17094 39409
rect 17038 39335 17094 39344
rect 17316 39296 17368 39302
rect 17314 39264 17316 39273
rect 17368 39264 17370 39273
rect 17314 39199 17370 39208
rect 16764 39024 16816 39030
rect 16948 39024 17000 39030
rect 16816 38972 16896 38978
rect 16764 38966 16896 38972
rect 16948 38966 17000 38972
rect 16488 38956 16540 38962
rect 16776 38950 16896 38966
rect 17512 38962 17540 39578
rect 17592 39432 17644 39438
rect 17592 39374 17644 39380
rect 16488 38898 16540 38904
rect 16212 38820 16264 38826
rect 16212 38762 16264 38768
rect 16120 38412 16172 38418
rect 16120 38354 16172 38360
rect 16224 37874 16252 38762
rect 16304 38752 16356 38758
rect 16304 38694 16356 38700
rect 16212 37868 16264 37874
rect 16212 37810 16264 37816
rect 16118 37360 16174 37369
rect 16118 37295 16174 37304
rect 16028 37120 16080 37126
rect 16028 37062 16080 37068
rect 16040 36718 16068 37062
rect 16028 36712 16080 36718
rect 16028 36654 16080 36660
rect 15936 36372 15988 36378
rect 15936 36314 15988 36320
rect 15844 36304 15896 36310
rect 15844 36246 15896 36252
rect 15934 36272 15990 36281
rect 15934 36207 15990 36216
rect 15948 35766 15976 36207
rect 16132 36174 16160 37295
rect 16212 36712 16264 36718
rect 16210 36680 16212 36689
rect 16264 36680 16266 36689
rect 16210 36615 16266 36624
rect 16120 36168 16172 36174
rect 16120 36110 16172 36116
rect 16212 36168 16264 36174
rect 16212 36110 16264 36116
rect 16224 35834 16252 36110
rect 16212 35828 16264 35834
rect 16212 35770 16264 35776
rect 15752 35760 15804 35766
rect 15752 35702 15804 35708
rect 15936 35760 15988 35766
rect 15936 35702 15988 35708
rect 16316 35494 16344 38694
rect 16500 38418 16528 38898
rect 16488 38412 16540 38418
rect 16488 38354 16540 38360
rect 16500 37806 16528 38354
rect 16488 37800 16540 37806
rect 16488 37742 16540 37748
rect 16396 37732 16448 37738
rect 16396 37674 16448 37680
rect 16408 37330 16436 37674
rect 16396 37324 16448 37330
rect 16396 37266 16448 37272
rect 16408 36650 16436 37266
rect 16396 36644 16448 36650
rect 16396 36586 16448 36592
rect 16408 36242 16436 36586
rect 16396 36236 16448 36242
rect 16396 36178 16448 36184
rect 16500 36122 16528 37742
rect 16408 36094 16528 36122
rect 16304 35488 16356 35494
rect 16304 35430 16356 35436
rect 16408 35306 16436 36094
rect 16672 36032 16724 36038
rect 16672 35974 16724 35980
rect 16684 35698 16712 35974
rect 16764 35828 16816 35834
rect 16764 35770 16816 35776
rect 16672 35692 16724 35698
rect 16672 35634 16724 35640
rect 16486 35456 16542 35465
rect 16486 35391 16542 35400
rect 16316 35278 16436 35306
rect 14372 35080 14424 35086
rect 14372 35022 14424 35028
rect 14752 35018 14780 35142
rect 15212 35086 15240 35142
rect 15660 35148 15712 35154
rect 15660 35090 15712 35096
rect 14924 35080 14976 35086
rect 14924 35022 14976 35028
rect 15108 35080 15160 35086
rect 15108 35022 15160 35028
rect 15200 35080 15252 35086
rect 15200 35022 15252 35028
rect 14740 35012 14792 35018
rect 14740 34954 14792 34960
rect 14936 34950 14964 35022
rect 14924 34944 14976 34950
rect 14924 34886 14976 34892
rect 15120 34649 15148 35022
rect 15106 34640 15162 34649
rect 15106 34575 15162 34584
rect 14556 34536 14608 34542
rect 14556 34478 14608 34484
rect 14464 34196 14516 34202
rect 14464 34138 14516 34144
rect 14372 33992 14424 33998
rect 14292 33952 14372 33980
rect 14292 33862 14320 33952
rect 14372 33934 14424 33940
rect 14280 33856 14332 33862
rect 14280 33798 14332 33804
rect 14476 33674 14504 34138
rect 14568 33969 14596 34478
rect 14648 34400 14700 34406
rect 14648 34342 14700 34348
rect 14660 34241 14688 34342
rect 14846 34300 15154 34320
rect 14846 34298 14852 34300
rect 14908 34298 14932 34300
rect 14988 34298 15012 34300
rect 15068 34298 15092 34300
rect 15148 34298 15154 34300
rect 14908 34246 14910 34298
rect 15090 34246 15092 34298
rect 14846 34244 14852 34246
rect 14908 34244 14932 34246
rect 14988 34244 15012 34246
rect 15068 34244 15092 34246
rect 15148 34244 15154 34246
rect 14646 34232 14702 34241
rect 14846 34224 15154 34244
rect 14646 34167 14702 34176
rect 15212 34105 15240 35022
rect 15476 34468 15528 34474
rect 15476 34410 15528 34416
rect 15382 34368 15438 34377
rect 15382 34303 15438 34312
rect 15198 34096 15254 34105
rect 15198 34031 15254 34040
rect 14648 33992 14700 33998
rect 14554 33960 14610 33969
rect 14648 33934 14700 33940
rect 14924 33992 14976 33998
rect 14924 33934 14976 33940
rect 14554 33895 14610 33904
rect 14292 33646 14504 33674
rect 13818 33487 13874 33496
rect 14004 33516 14056 33522
rect 14004 33458 14056 33464
rect 13910 33416 13966 33425
rect 13740 33374 13910 33402
rect 13910 33351 13966 33360
rect 14188 32972 14240 32978
rect 12624 32904 12676 32910
rect 12544 32864 12624 32892
rect 12624 32846 12676 32852
rect 12440 32836 12492 32842
rect 12440 32778 12492 32784
rect 12728 32774 12756 32943
rect 13648 32932 13860 32960
rect 13084 32904 13136 32910
rect 13084 32846 13136 32852
rect 13542 32872 13598 32881
rect 12808 32836 12860 32842
rect 12808 32778 12860 32784
rect 12716 32768 12768 32774
rect 12716 32710 12768 32716
rect 12820 32502 12848 32778
rect 12900 32564 12952 32570
rect 12900 32506 12952 32512
rect 12808 32496 12860 32502
rect 12808 32438 12860 32444
rect 12532 32292 12584 32298
rect 12532 32234 12584 32240
rect 12544 32201 12572 32234
rect 12820 32230 12848 32438
rect 12716 32224 12768 32230
rect 12530 32192 12586 32201
rect 12716 32166 12768 32172
rect 12808 32224 12860 32230
rect 12808 32166 12860 32172
rect 12530 32127 12586 32136
rect 12728 31958 12756 32166
rect 12716 31952 12768 31958
rect 12716 31894 12768 31900
rect 12912 31822 12940 32506
rect 13096 32366 13124 32846
rect 13452 32836 13504 32842
rect 13542 32807 13544 32816
rect 13452 32778 13504 32784
rect 13596 32807 13598 32816
rect 13726 32872 13782 32881
rect 13726 32807 13782 32816
rect 13544 32778 13596 32784
rect 13176 32768 13228 32774
rect 13176 32710 13228 32716
rect 13188 32434 13216 32710
rect 13358 32600 13414 32609
rect 13358 32535 13360 32544
rect 13412 32535 13414 32544
rect 13360 32506 13412 32512
rect 13176 32428 13228 32434
rect 13176 32370 13228 32376
rect 13084 32360 13136 32366
rect 13084 32302 13136 32308
rect 12900 31816 12952 31822
rect 12900 31758 12952 31764
rect 11978 31719 12034 31728
rect 12084 31726 12388 31754
rect 11992 31142 12020 31719
rect 12084 31346 12112 31726
rect 13188 31686 13216 32370
rect 13464 32230 13492 32778
rect 13740 32722 13768 32807
rect 13556 32694 13768 32722
rect 13452 32224 13504 32230
rect 13452 32166 13504 32172
rect 13556 31958 13584 32694
rect 13728 32496 13780 32502
rect 13648 32456 13728 32484
rect 13544 31952 13596 31958
rect 13450 31920 13506 31929
rect 13544 31894 13596 31900
rect 13450 31855 13506 31864
rect 12348 31680 12400 31686
rect 12176 31640 12348 31668
rect 12072 31340 12124 31346
rect 12072 31282 12124 31288
rect 12176 31278 12204 31640
rect 12348 31622 12400 31628
rect 13176 31680 13228 31686
rect 13176 31622 13228 31628
rect 12268 31470 13124 31498
rect 12268 31414 12296 31470
rect 12256 31408 12308 31414
rect 12256 31350 12308 31356
rect 12348 31408 12400 31414
rect 12348 31350 12400 31356
rect 12164 31272 12216 31278
rect 12164 31214 12216 31220
rect 11980 31136 12032 31142
rect 11886 31104 11942 31113
rect 12360 31090 12388 31350
rect 11980 31078 12032 31084
rect 11886 31039 11942 31048
rect 12084 31062 12388 31090
rect 12452 31334 12940 31362
rect 11900 30569 11928 31039
rect 11980 30932 12032 30938
rect 11980 30874 12032 30880
rect 11886 30560 11942 30569
rect 11886 30495 11942 30504
rect 11520 29640 11572 29646
rect 11520 29582 11572 29588
rect 11704 29640 11756 29646
rect 11704 29582 11756 29588
rect 11796 29640 11848 29646
rect 11992 29617 12020 30874
rect 12084 30161 12112 31062
rect 12452 30954 12480 31334
rect 12808 31272 12860 31278
rect 12808 31214 12860 31220
rect 12624 31136 12676 31142
rect 12624 31078 12676 31084
rect 12176 30926 12480 30954
rect 12636 30938 12664 31078
rect 12714 30968 12770 30977
rect 12624 30932 12676 30938
rect 12176 30870 12204 30926
rect 12714 30903 12716 30912
rect 12624 30874 12676 30880
rect 12768 30903 12770 30912
rect 12716 30874 12768 30880
rect 12164 30864 12216 30870
rect 12164 30806 12216 30812
rect 12256 30864 12308 30870
rect 12820 30852 12848 31214
rect 12912 30977 12940 31334
rect 12898 30968 12954 30977
rect 12898 30903 12954 30912
rect 12820 30824 12940 30852
rect 12256 30806 12308 30812
rect 12268 30734 12296 30806
rect 12716 30796 12768 30802
rect 12716 30738 12768 30744
rect 12256 30728 12308 30734
rect 12256 30670 12308 30676
rect 12348 30728 12400 30734
rect 12624 30728 12676 30734
rect 12400 30676 12572 30682
rect 12348 30670 12572 30676
rect 12728 30705 12756 30738
rect 12624 30670 12676 30676
rect 12714 30696 12770 30705
rect 12360 30654 12572 30670
rect 12348 30592 12400 30598
rect 12346 30560 12348 30569
rect 12440 30592 12492 30598
rect 12400 30560 12402 30569
rect 12440 30534 12492 30540
rect 12346 30495 12402 30504
rect 12348 30388 12400 30394
rect 12348 30330 12400 30336
rect 12360 30258 12388 30330
rect 12348 30252 12400 30258
rect 12348 30194 12400 30200
rect 12452 30161 12480 30534
rect 12544 30394 12572 30654
rect 12532 30388 12584 30394
rect 12532 30330 12584 30336
rect 12070 30152 12126 30161
rect 12070 30087 12126 30096
rect 12438 30152 12494 30161
rect 12438 30087 12494 30096
rect 12164 29776 12216 29782
rect 12216 29736 12572 29764
rect 12636 29753 12664 30670
rect 12714 30631 12770 30640
rect 12816 30592 12868 30598
rect 12728 30552 12816 30580
rect 12728 30326 12756 30552
rect 12816 30534 12868 30540
rect 12716 30320 12768 30326
rect 12716 30262 12768 30268
rect 12714 30152 12770 30161
rect 12714 30087 12716 30096
rect 12768 30087 12770 30096
rect 12716 30058 12768 30064
rect 12808 30048 12860 30054
rect 12728 29996 12808 30002
rect 12912 30036 12940 30824
rect 13096 30705 13124 31470
rect 13464 31346 13492 31855
rect 13176 31340 13228 31346
rect 13176 31282 13228 31288
rect 13452 31340 13504 31346
rect 13452 31282 13504 31288
rect 13188 30734 13216 31282
rect 13648 31260 13676 32456
rect 13728 32438 13780 32444
rect 13832 32434 13860 32932
rect 14188 32914 14240 32920
rect 14096 32768 14148 32774
rect 14096 32710 14148 32716
rect 13820 32428 13872 32434
rect 13820 32370 13872 32376
rect 13728 32292 13780 32298
rect 13728 32234 13780 32240
rect 13740 31890 13768 32234
rect 13820 32224 13872 32230
rect 14004 32224 14056 32230
rect 13820 32166 13872 32172
rect 14002 32192 14004 32201
rect 14056 32192 14058 32201
rect 13832 32026 13860 32166
rect 14002 32127 14058 32136
rect 13820 32020 13872 32026
rect 13820 31962 13872 31968
rect 14108 31958 14136 32710
rect 14200 32502 14228 32914
rect 14292 32722 14320 33646
rect 14660 33572 14688 33934
rect 14832 33924 14884 33930
rect 14832 33866 14884 33872
rect 14384 33544 14688 33572
rect 14384 32842 14412 33544
rect 14844 33504 14872 33866
rect 14660 33476 14872 33504
rect 14464 33448 14516 33454
rect 14464 33390 14516 33396
rect 14476 33153 14504 33390
rect 14660 33289 14688 33476
rect 14832 33380 14884 33386
rect 14936 33368 14964 33934
rect 15200 33856 15252 33862
rect 15252 33816 15332 33844
rect 15200 33798 15252 33804
rect 15200 33516 15252 33522
rect 15200 33458 15252 33464
rect 15108 33448 15160 33454
rect 14884 33340 14964 33368
rect 15106 33416 15108 33425
rect 15160 33416 15162 33425
rect 15106 33351 15162 33360
rect 14832 33322 14884 33328
rect 15212 33318 15240 33458
rect 14740 33312 14792 33318
rect 14646 33280 14702 33289
rect 14740 33254 14792 33260
rect 15200 33312 15252 33318
rect 15200 33254 15252 33260
rect 14646 33215 14702 33224
rect 14462 33144 14518 33153
rect 14462 33079 14518 33088
rect 14752 32842 14780 33254
rect 14846 33212 15154 33232
rect 14846 33210 14852 33212
rect 14908 33210 14932 33212
rect 14988 33210 15012 33212
rect 15068 33210 15092 33212
rect 15148 33210 15154 33212
rect 14908 33158 14910 33210
rect 15090 33158 15092 33210
rect 14846 33156 14852 33158
rect 14908 33156 14932 33158
rect 14988 33156 15012 33158
rect 15068 33156 15092 33158
rect 15148 33156 15154 33158
rect 14846 33136 15154 33156
rect 14832 32972 14884 32978
rect 14832 32914 14884 32920
rect 14372 32836 14424 32842
rect 14372 32778 14424 32784
rect 14556 32836 14608 32842
rect 14556 32778 14608 32784
rect 14740 32836 14792 32842
rect 14740 32778 14792 32784
rect 14292 32694 14504 32722
rect 14188 32496 14240 32502
rect 14372 32496 14424 32502
rect 14188 32438 14240 32444
rect 14292 32456 14372 32484
rect 14292 32298 14320 32456
rect 14372 32438 14424 32444
rect 14476 32348 14504 32694
rect 14384 32320 14504 32348
rect 14280 32292 14332 32298
rect 14280 32234 14332 32240
rect 14278 32192 14334 32201
rect 14278 32127 14334 32136
rect 14096 31952 14148 31958
rect 13818 31920 13874 31929
rect 13728 31884 13780 31890
rect 14292 31929 14320 32127
rect 14096 31894 14148 31900
rect 14278 31920 14334 31929
rect 13818 31855 13874 31864
rect 14278 31855 14334 31864
rect 13728 31826 13780 31832
rect 13832 31657 13860 31855
rect 14096 31816 14148 31822
rect 14096 31758 14148 31764
rect 13912 31680 13964 31686
rect 13818 31648 13874 31657
rect 13912 31622 13964 31628
rect 14002 31648 14058 31657
rect 13818 31583 13874 31592
rect 13728 31408 13780 31414
rect 13726 31376 13728 31385
rect 13780 31376 13782 31385
rect 13726 31311 13782 31320
rect 13924 31278 13952 31622
rect 14002 31583 14058 31592
rect 13912 31272 13964 31278
rect 13648 31232 13768 31260
rect 13176 30728 13228 30734
rect 13082 30696 13138 30705
rect 12992 30660 13044 30666
rect 13452 30728 13504 30734
rect 13228 30688 13452 30716
rect 13176 30670 13228 30676
rect 13452 30670 13504 30676
rect 13636 30728 13688 30734
rect 13636 30670 13688 30676
rect 13082 30631 13138 30640
rect 12992 30602 13044 30608
rect 13004 30546 13032 30602
rect 13648 30546 13676 30670
rect 13004 30518 13676 30546
rect 13174 30424 13230 30433
rect 13174 30359 13230 30368
rect 13358 30424 13414 30433
rect 13740 30410 13768 31232
rect 13912 31214 13964 31220
rect 13358 30359 13414 30368
rect 13648 30382 13768 30410
rect 12992 30184 13044 30190
rect 12992 30126 13044 30132
rect 12860 30008 12940 30036
rect 12728 29990 12860 29996
rect 12728 29974 12848 29990
rect 12164 29718 12216 29724
rect 12164 29640 12216 29646
rect 11796 29582 11848 29588
rect 11978 29608 12034 29617
rect 12164 29582 12216 29588
rect 12254 29608 12310 29617
rect 11978 29543 12034 29552
rect 11794 29472 11850 29481
rect 11794 29407 11850 29416
rect 11808 29238 11836 29407
rect 11796 29232 11848 29238
rect 11796 29174 11848 29180
rect 12176 29170 12204 29582
rect 12544 29578 12572 29736
rect 12622 29744 12678 29753
rect 12622 29679 12678 29688
rect 12254 29543 12256 29552
rect 12308 29543 12310 29552
rect 12532 29572 12584 29578
rect 12256 29514 12308 29520
rect 12532 29514 12584 29520
rect 12624 29572 12676 29578
rect 12624 29514 12676 29520
rect 12438 29472 12494 29481
rect 12438 29407 12494 29416
rect 12256 29232 12308 29238
rect 12452 29220 12480 29407
rect 12636 29288 12664 29514
rect 12308 29192 12480 29220
rect 12544 29260 12664 29288
rect 12256 29174 12308 29180
rect 11428 29164 11480 29170
rect 12164 29164 12216 29170
rect 11428 29106 11480 29112
rect 12084 29124 12164 29152
rect 11336 29028 11388 29034
rect 11336 28970 11388 28976
rect 11440 28966 11468 29106
rect 11520 29096 11572 29102
rect 11612 29096 11664 29102
rect 11520 29038 11572 29044
rect 11610 29064 11612 29073
rect 11664 29064 11666 29073
rect 11978 29064 12034 29073
rect 11428 28960 11480 28966
rect 11428 28902 11480 28908
rect 11532 28914 11560 29038
rect 11610 28999 11666 29008
rect 11900 29022 11978 29050
rect 11900 28914 11928 29022
rect 11978 28999 12034 29008
rect 11532 28886 11928 28914
rect 11244 28620 11296 28626
rect 11244 28562 11296 28568
rect 11058 28520 11114 28529
rect 11058 28455 11114 28464
rect 11072 28422 11100 28455
rect 11060 28416 11112 28422
rect 11060 28358 11112 28364
rect 11256 28150 11284 28562
rect 11336 28552 11388 28558
rect 11336 28494 11388 28500
rect 11244 28144 11296 28150
rect 11348 28121 11376 28494
rect 11612 28484 11664 28490
rect 11440 28444 11612 28472
rect 11244 28086 11296 28092
rect 11334 28112 11390 28121
rect 11256 27470 11284 28086
rect 11334 28047 11390 28056
rect 11244 27464 11296 27470
rect 11244 27406 11296 27412
rect 11060 27396 11112 27402
rect 11060 27338 11112 27344
rect 10966 27296 11022 27305
rect 10966 27231 11022 27240
rect 10968 26240 11020 26246
rect 10968 26182 11020 26188
rect 10796 25112 10916 25140
rect 10600 24880 10652 24886
rect 10600 24822 10652 24828
rect 10324 24812 10376 24818
rect 10324 24754 10376 24760
rect 10336 24410 10364 24754
rect 10324 24404 10376 24410
rect 10324 24346 10376 24352
rect 10600 24200 10652 24206
rect 10600 24142 10652 24148
rect 10692 24200 10744 24206
rect 10692 24142 10744 24148
rect 10214 23964 10522 23984
rect 10214 23962 10220 23964
rect 10276 23962 10300 23964
rect 10356 23962 10380 23964
rect 10436 23962 10460 23964
rect 10516 23962 10522 23964
rect 10276 23910 10278 23962
rect 10458 23910 10460 23962
rect 10214 23908 10220 23910
rect 10276 23908 10300 23910
rect 10356 23908 10380 23910
rect 10436 23908 10460 23910
rect 10516 23908 10522 23910
rect 10214 23888 10522 23908
rect 10232 23724 10284 23730
rect 10232 23666 10284 23672
rect 10324 23724 10376 23730
rect 10324 23666 10376 23672
rect 10244 23225 10272 23666
rect 10336 23361 10364 23666
rect 10322 23352 10378 23361
rect 10322 23287 10378 23296
rect 10230 23216 10286 23225
rect 10230 23151 10286 23160
rect 10214 22876 10522 22896
rect 10214 22874 10220 22876
rect 10276 22874 10300 22876
rect 10356 22874 10380 22876
rect 10436 22874 10460 22876
rect 10516 22874 10522 22876
rect 10276 22822 10278 22874
rect 10458 22822 10460 22874
rect 10214 22820 10220 22822
rect 10276 22820 10300 22822
rect 10356 22820 10380 22822
rect 10436 22820 10460 22822
rect 10516 22820 10522 22822
rect 10214 22800 10522 22820
rect 10214 21788 10522 21808
rect 10214 21786 10220 21788
rect 10276 21786 10300 21788
rect 10356 21786 10380 21788
rect 10436 21786 10460 21788
rect 10516 21786 10522 21788
rect 10276 21734 10278 21786
rect 10458 21734 10460 21786
rect 10214 21732 10220 21734
rect 10276 21732 10300 21734
rect 10356 21732 10380 21734
rect 10436 21732 10460 21734
rect 10516 21732 10522 21734
rect 10214 21712 10522 21732
rect 10214 20700 10522 20720
rect 10214 20698 10220 20700
rect 10276 20698 10300 20700
rect 10356 20698 10380 20700
rect 10436 20698 10460 20700
rect 10516 20698 10522 20700
rect 10276 20646 10278 20698
rect 10458 20646 10460 20698
rect 10214 20644 10220 20646
rect 10276 20644 10300 20646
rect 10356 20644 10380 20646
rect 10436 20644 10460 20646
rect 10516 20644 10522 20646
rect 10214 20624 10522 20644
rect 10214 19612 10522 19632
rect 10214 19610 10220 19612
rect 10276 19610 10300 19612
rect 10356 19610 10380 19612
rect 10436 19610 10460 19612
rect 10516 19610 10522 19612
rect 10276 19558 10278 19610
rect 10458 19558 10460 19610
rect 10214 19556 10220 19558
rect 10276 19556 10300 19558
rect 10356 19556 10380 19558
rect 10436 19556 10460 19558
rect 10516 19556 10522 19558
rect 10214 19536 10522 19556
rect 10214 18524 10522 18544
rect 10214 18522 10220 18524
rect 10276 18522 10300 18524
rect 10356 18522 10380 18524
rect 10436 18522 10460 18524
rect 10516 18522 10522 18524
rect 10276 18470 10278 18522
rect 10458 18470 10460 18522
rect 10214 18468 10220 18470
rect 10276 18468 10300 18470
rect 10356 18468 10380 18470
rect 10436 18468 10460 18470
rect 10516 18468 10522 18470
rect 10214 18448 10522 18468
rect 10612 17649 10640 24142
rect 10704 24041 10732 24142
rect 10796 24052 10824 25112
rect 10876 24608 10928 24614
rect 10876 24550 10928 24556
rect 10888 24206 10916 24550
rect 10980 24410 11008 26182
rect 11072 25945 11100 27338
rect 11440 27130 11468 28444
rect 11612 28426 11664 28432
rect 11704 28484 11756 28490
rect 11704 28426 11756 28432
rect 11520 28076 11572 28082
rect 11520 28018 11572 28024
rect 11428 27124 11480 27130
rect 11428 27066 11480 27072
rect 11334 26480 11390 26489
rect 11334 26415 11390 26424
rect 11348 26382 11376 26415
rect 11532 26382 11560 28018
rect 11610 27976 11666 27985
rect 11610 27911 11666 27920
rect 11624 27402 11652 27911
rect 11612 27396 11664 27402
rect 11612 27338 11664 27344
rect 11716 27282 11744 28426
rect 11980 28144 12032 28150
rect 11794 28112 11850 28121
rect 12084 28132 12112 29124
rect 12544 29152 12572 29260
rect 12164 29106 12216 29112
rect 12452 29124 12572 29152
rect 12622 29200 12678 29209
rect 12622 29135 12678 29144
rect 12452 28937 12480 29124
rect 12532 29028 12584 29034
rect 12636 29016 12664 29135
rect 12584 28988 12664 29016
rect 12532 28970 12584 28976
rect 12438 28928 12494 28937
rect 12438 28863 12494 28872
rect 12348 28756 12400 28762
rect 12348 28698 12400 28704
rect 12360 28422 12388 28698
rect 12440 28688 12492 28694
rect 12438 28656 12440 28665
rect 12492 28656 12494 28665
rect 12622 28656 12678 28665
rect 12438 28591 12494 28600
rect 12544 28614 12622 28642
rect 12348 28416 12400 28422
rect 12348 28358 12400 28364
rect 12440 28416 12492 28422
rect 12440 28358 12492 28364
rect 12032 28104 12112 28132
rect 12452 28121 12480 28358
rect 11980 28086 12032 28092
rect 11794 28047 11850 28056
rect 11808 28014 11836 28047
rect 11796 28008 11848 28014
rect 11796 27950 11848 27956
rect 11886 27976 11942 27985
rect 11886 27911 11888 27920
rect 11940 27911 11942 27920
rect 11888 27882 11940 27888
rect 11980 27464 12032 27470
rect 11980 27406 12032 27412
rect 11624 27254 11744 27282
rect 11624 27062 11652 27254
rect 11702 27160 11758 27169
rect 11702 27095 11758 27104
rect 11612 27056 11664 27062
rect 11612 26998 11664 27004
rect 11716 26994 11744 27095
rect 11704 26988 11756 26994
rect 11704 26930 11756 26936
rect 11796 26920 11848 26926
rect 11796 26862 11848 26868
rect 11808 26761 11836 26862
rect 11992 26790 12020 27406
rect 11980 26784 12032 26790
rect 11794 26752 11850 26761
rect 11980 26726 12032 26732
rect 12084 26738 12112 28104
rect 12438 28112 12494 28121
rect 12438 28047 12494 28056
rect 12164 27872 12216 27878
rect 12164 27814 12216 27820
rect 12176 26858 12204 27814
rect 12452 27470 12480 28047
rect 12544 27985 12572 28614
rect 12622 28591 12678 28600
rect 12622 28520 12678 28529
rect 12622 28455 12678 28464
rect 12636 28218 12664 28455
rect 12624 28212 12676 28218
rect 12624 28154 12676 28160
rect 12622 28112 12678 28121
rect 12622 28047 12678 28056
rect 12530 27976 12586 27985
rect 12636 27946 12664 28047
rect 12530 27911 12586 27920
rect 12624 27940 12676 27946
rect 12624 27882 12676 27888
rect 12728 27674 12756 29974
rect 13004 29889 13032 30126
rect 12990 29880 13046 29889
rect 12990 29815 13046 29824
rect 13188 29714 13216 30359
rect 13266 29880 13322 29889
rect 13266 29815 13322 29824
rect 13176 29708 13228 29714
rect 13176 29650 13228 29656
rect 12990 29608 13046 29617
rect 12990 29543 13046 29552
rect 12900 28552 12952 28558
rect 12898 28520 12900 28529
rect 12952 28520 12954 28529
rect 12898 28455 12954 28464
rect 12808 28212 12860 28218
rect 12808 28154 12860 28160
rect 12820 28082 12848 28154
rect 12808 28076 12860 28082
rect 12808 28018 12860 28024
rect 13004 28014 13032 29543
rect 13084 29164 13136 29170
rect 13084 29106 13136 29112
rect 13096 29073 13124 29106
rect 13082 29064 13138 29073
rect 13082 28999 13138 29008
rect 13084 28552 13136 28558
rect 13084 28494 13136 28500
rect 12992 28008 13044 28014
rect 12992 27950 13044 27956
rect 13096 27826 13124 28494
rect 13280 28472 13308 29815
rect 13372 28626 13400 30359
rect 13452 30252 13504 30258
rect 13452 30194 13504 30200
rect 13464 29889 13492 30194
rect 13450 29880 13506 29889
rect 13450 29815 13506 29824
rect 13452 29776 13504 29782
rect 13452 29718 13504 29724
rect 13464 29617 13492 29718
rect 13450 29608 13506 29617
rect 13450 29543 13506 29552
rect 13648 29492 13676 30382
rect 14016 30376 14044 31583
rect 13924 30348 14044 30376
rect 13924 30122 13952 30348
rect 14004 30252 14056 30258
rect 14108 30240 14136 31758
rect 14188 31272 14240 31278
rect 14188 31214 14240 31220
rect 14200 30734 14228 31214
rect 14188 30728 14240 30734
rect 14188 30670 14240 30676
rect 14186 30560 14242 30569
rect 14186 30495 14242 30504
rect 14056 30212 14136 30240
rect 14004 30194 14056 30200
rect 13912 30116 13964 30122
rect 13912 30058 13964 30064
rect 13728 30048 13780 30054
rect 13728 29990 13780 29996
rect 13464 29464 13676 29492
rect 13360 28620 13412 28626
rect 13360 28562 13412 28568
rect 13280 28444 13400 28472
rect 13176 28416 13228 28422
rect 13228 28376 13308 28404
rect 13176 28358 13228 28364
rect 13176 28212 13228 28218
rect 13176 28154 13228 28160
rect 12820 27798 13124 27826
rect 12716 27668 12768 27674
rect 12544 27628 12716 27656
rect 12440 27464 12492 27470
rect 12440 27406 12492 27412
rect 12440 27328 12492 27334
rect 12254 27296 12310 27305
rect 12254 27231 12310 27240
rect 12438 27296 12440 27305
rect 12492 27296 12494 27305
rect 12438 27231 12494 27240
rect 12268 27130 12296 27231
rect 12256 27124 12308 27130
rect 12256 27066 12308 27072
rect 12544 26994 12572 27628
rect 12716 27610 12768 27616
rect 12716 27328 12768 27334
rect 12716 27270 12768 27276
rect 12728 26994 12756 27270
rect 12532 26988 12584 26994
rect 12532 26930 12584 26936
rect 12716 26988 12768 26994
rect 12716 26930 12768 26936
rect 12348 26920 12400 26926
rect 12348 26862 12400 26868
rect 12164 26852 12216 26858
rect 12164 26794 12216 26800
rect 12256 26784 12308 26790
rect 12084 26710 12204 26738
rect 12256 26726 12308 26732
rect 11794 26687 11850 26696
rect 12072 26512 12124 26518
rect 12072 26454 12124 26460
rect 11336 26376 11388 26382
rect 11336 26318 11388 26324
rect 11520 26376 11572 26382
rect 11888 26376 11940 26382
rect 11520 26318 11572 26324
rect 11808 26324 11888 26330
rect 11808 26318 11940 26324
rect 11058 25936 11114 25945
rect 11058 25871 11114 25880
rect 11336 25900 11388 25906
rect 11336 25842 11388 25848
rect 11428 25900 11480 25906
rect 11428 25842 11480 25848
rect 11150 25800 11206 25809
rect 11150 25735 11206 25744
rect 11058 25528 11114 25537
rect 11058 25463 11060 25472
rect 11112 25463 11114 25472
rect 11060 25434 11112 25440
rect 11164 25294 11192 25735
rect 11244 25696 11296 25702
rect 11244 25638 11296 25644
rect 11152 25288 11204 25294
rect 11152 25230 11204 25236
rect 11060 25220 11112 25226
rect 11060 25162 11112 25168
rect 11072 24993 11100 25162
rect 11058 24984 11114 24993
rect 11058 24919 11114 24928
rect 11256 24410 11284 25638
rect 11348 25498 11376 25842
rect 11336 25492 11388 25498
rect 11336 25434 11388 25440
rect 11440 25362 11468 25842
rect 11428 25356 11480 25362
rect 11532 25344 11560 26318
rect 11612 26308 11664 26314
rect 11808 26302 11928 26318
rect 11980 26308 12032 26314
rect 11808 26296 11836 26302
rect 11664 26268 11836 26296
rect 11612 26250 11664 26256
rect 11980 26250 12032 26256
rect 11532 25316 11652 25344
rect 11428 25298 11480 25304
rect 11520 25220 11572 25226
rect 11520 25162 11572 25168
rect 11532 24970 11560 25162
rect 11348 24942 11560 24970
rect 11624 24954 11652 25316
rect 11612 24948 11664 24954
rect 11348 24682 11376 24942
rect 11612 24890 11664 24896
rect 11428 24744 11480 24750
rect 11428 24686 11480 24692
rect 11888 24744 11940 24750
rect 11992 24732 12020 26250
rect 12084 26217 12112 26454
rect 12176 26450 12204 26710
rect 12164 26444 12216 26450
rect 12164 26386 12216 26392
rect 12268 26314 12296 26726
rect 12256 26308 12308 26314
rect 12256 26250 12308 26256
rect 12360 26246 12388 26862
rect 12624 26852 12676 26858
rect 12624 26794 12676 26800
rect 12636 26489 12664 26794
rect 12728 26790 12756 26930
rect 12716 26784 12768 26790
rect 12716 26726 12768 26732
rect 12622 26480 12678 26489
rect 12622 26415 12678 26424
rect 12636 26314 12664 26415
rect 12532 26308 12584 26314
rect 12532 26250 12584 26256
rect 12624 26308 12676 26314
rect 12624 26250 12676 26256
rect 12348 26240 12400 26246
rect 12070 26208 12126 26217
rect 12348 26182 12400 26188
rect 12070 26143 12126 26152
rect 12164 25900 12216 25906
rect 12164 25842 12216 25848
rect 12072 24948 12124 24954
rect 12072 24890 12124 24896
rect 12084 24818 12112 24890
rect 12072 24812 12124 24818
rect 12072 24754 12124 24760
rect 11940 24704 12020 24732
rect 12070 24712 12126 24721
rect 11888 24686 11940 24692
rect 11336 24676 11388 24682
rect 11336 24618 11388 24624
rect 10968 24404 11020 24410
rect 10968 24346 11020 24352
rect 11244 24404 11296 24410
rect 11244 24346 11296 24352
rect 11440 24206 11468 24686
rect 12070 24647 12126 24656
rect 11796 24608 11848 24614
rect 11518 24576 11574 24585
rect 11796 24550 11848 24556
rect 11518 24511 11574 24520
rect 10876 24200 10928 24206
rect 10876 24142 10928 24148
rect 11428 24200 11480 24206
rect 11428 24142 11480 24148
rect 10690 24032 10746 24041
rect 10796 24024 10916 24052
rect 10690 23967 10746 23976
rect 10782 23896 10838 23905
rect 10782 23831 10838 23840
rect 10796 23730 10824 23831
rect 10784 23724 10836 23730
rect 10784 23666 10836 23672
rect 10784 22636 10836 22642
rect 10784 22578 10836 22584
rect 10796 22234 10824 22578
rect 10784 22228 10836 22234
rect 10784 22170 10836 22176
rect 10888 20505 10916 24024
rect 11440 23769 11468 24142
rect 11426 23760 11482 23769
rect 11336 23724 11388 23730
rect 11426 23695 11482 23704
rect 11336 23666 11388 23672
rect 11348 23322 11376 23666
rect 11336 23316 11388 23322
rect 11336 23258 11388 23264
rect 11532 23118 11560 24511
rect 11808 24410 11836 24550
rect 11796 24404 11848 24410
rect 11796 24346 11848 24352
rect 12084 24342 12112 24647
rect 12176 24410 12204 25842
rect 12544 25537 12572 26250
rect 12636 25770 12664 26250
rect 12820 25945 12848 27798
rect 13188 27690 13216 28154
rect 13280 28082 13308 28376
rect 13268 28076 13320 28082
rect 13268 28018 13320 28024
rect 12912 27662 13216 27690
rect 12912 27402 12940 27662
rect 13266 27432 13322 27441
rect 12900 27396 12952 27402
rect 12900 27338 12952 27344
rect 13004 27390 13266 27418
rect 13004 27305 13032 27390
rect 13266 27367 13322 27376
rect 12990 27296 13046 27305
rect 12990 27231 13046 27240
rect 12992 26988 13044 26994
rect 12992 26930 13044 26936
rect 12806 25936 12862 25945
rect 12806 25871 12862 25880
rect 12624 25764 12676 25770
rect 12624 25706 12676 25712
rect 12530 25528 12586 25537
rect 12530 25463 12586 25472
rect 13004 25430 13032 26930
rect 13268 26852 13320 26858
rect 13268 26794 13320 26800
rect 13280 26738 13308 26794
rect 13096 26710 13308 26738
rect 13096 26246 13124 26710
rect 13372 26602 13400 28444
rect 13464 28082 13492 29464
rect 13740 29306 13768 29990
rect 14016 29714 14044 30194
rect 14094 30016 14150 30025
rect 14094 29951 14150 29960
rect 14004 29708 14056 29714
rect 14004 29650 14056 29656
rect 13820 29640 13872 29646
rect 13820 29582 13872 29588
rect 13832 29306 13860 29582
rect 14016 29492 14044 29650
rect 14108 29646 14136 29951
rect 14096 29640 14148 29646
rect 14096 29582 14148 29588
rect 14016 29464 14136 29492
rect 13728 29300 13780 29306
rect 13728 29242 13780 29248
rect 13820 29300 13872 29306
rect 13820 29242 13872 29248
rect 14108 29238 14136 29464
rect 14200 29238 14228 30495
rect 14096 29232 14148 29238
rect 14096 29174 14148 29180
rect 14188 29232 14240 29238
rect 14188 29174 14240 29180
rect 13636 29028 13688 29034
rect 13636 28970 13688 28976
rect 13544 28552 13596 28558
rect 13544 28494 13596 28500
rect 13452 28076 13504 28082
rect 13452 28018 13504 28024
rect 13556 27690 13584 28494
rect 13464 27674 13584 27690
rect 13452 27668 13584 27674
rect 13504 27662 13584 27668
rect 13452 27610 13504 27616
rect 13648 27614 13676 28970
rect 13912 28960 13964 28966
rect 13912 28902 13964 28908
rect 13728 28620 13780 28626
rect 13728 28562 13780 28568
rect 13556 27586 13676 27614
rect 13450 27296 13506 27305
rect 13556 27282 13584 27586
rect 13506 27254 13584 27282
rect 13634 27296 13690 27305
rect 13450 27231 13506 27240
rect 13634 27231 13690 27240
rect 13452 27124 13504 27130
rect 13452 27066 13504 27072
rect 13188 26574 13400 26602
rect 13084 26240 13136 26246
rect 13084 26182 13136 26188
rect 12716 25424 12768 25430
rect 12716 25366 12768 25372
rect 12992 25424 13044 25430
rect 12992 25366 13044 25372
rect 12532 25220 12584 25226
rect 12532 25162 12584 25168
rect 12440 24608 12492 24614
rect 12440 24550 12492 24556
rect 12164 24404 12216 24410
rect 12164 24346 12216 24352
rect 12072 24336 12124 24342
rect 12072 24278 12124 24284
rect 11980 24200 12032 24206
rect 11980 24142 12032 24148
rect 11992 23610 12020 24142
rect 12452 24138 12480 24550
rect 12440 24132 12492 24138
rect 12440 24074 12492 24080
rect 12438 23760 12494 23769
rect 12438 23695 12440 23704
rect 12492 23695 12494 23704
rect 12440 23666 12492 23672
rect 11992 23582 12112 23610
rect 11704 23520 11756 23526
rect 11704 23462 11756 23468
rect 11980 23520 12032 23526
rect 11980 23462 12032 23468
rect 11716 23186 11744 23462
rect 11704 23180 11756 23186
rect 11704 23122 11756 23128
rect 11992 23118 12020 23462
rect 11060 23112 11112 23118
rect 11060 23054 11112 23060
rect 11336 23112 11388 23118
rect 11336 23054 11388 23060
rect 11520 23112 11572 23118
rect 11520 23054 11572 23060
rect 11980 23112 12032 23118
rect 11980 23054 12032 23060
rect 10968 22976 11020 22982
rect 10968 22918 11020 22924
rect 10980 22642 11008 22918
rect 11072 22642 11100 23054
rect 11348 22817 11376 23054
rect 11334 22808 11390 22817
rect 11334 22743 11390 22752
rect 11978 22672 12034 22681
rect 10968 22636 11020 22642
rect 10968 22578 11020 22584
rect 11060 22636 11112 22642
rect 11978 22607 11980 22616
rect 11060 22578 11112 22584
rect 12032 22607 12034 22616
rect 11980 22578 12032 22584
rect 12084 22522 12112 23582
rect 12164 23112 12216 23118
rect 12162 23080 12164 23089
rect 12440 23112 12492 23118
rect 12216 23080 12218 23089
rect 12440 23054 12492 23060
rect 12162 23015 12218 23024
rect 12084 22494 12204 22522
rect 12072 22432 12124 22438
rect 12072 22374 12124 22380
rect 12084 22166 12112 22374
rect 12072 22160 12124 22166
rect 12072 22102 12124 22108
rect 11244 22024 11296 22030
rect 11244 21966 11296 21972
rect 11888 22024 11940 22030
rect 11888 21966 11940 21972
rect 11256 21729 11284 21966
rect 11242 21720 11298 21729
rect 11900 21690 11928 21966
rect 11242 21655 11298 21664
rect 11888 21684 11940 21690
rect 11888 21626 11940 21632
rect 11796 21548 11848 21554
rect 11796 21490 11848 21496
rect 11808 21010 11836 21490
rect 12072 21072 12124 21078
rect 12072 21014 12124 21020
rect 11796 21004 11848 21010
rect 11796 20946 11848 20952
rect 12084 20913 12112 21014
rect 12070 20904 12126 20913
rect 12070 20839 12126 20848
rect 10874 20496 10930 20505
rect 10874 20431 10930 20440
rect 12176 20369 12204 22494
rect 12254 22128 12310 22137
rect 12254 22063 12310 22072
rect 12268 21486 12296 22063
rect 12452 21706 12480 23054
rect 12360 21678 12480 21706
rect 12360 21622 12388 21678
rect 12348 21616 12400 21622
rect 12348 21558 12400 21564
rect 12256 21480 12308 21486
rect 12256 21422 12308 21428
rect 12440 20868 12492 20874
rect 12440 20810 12492 20816
rect 12162 20360 12218 20369
rect 12162 20295 12218 20304
rect 12452 19417 12480 20810
rect 12438 19408 12494 19417
rect 12438 19343 12494 19352
rect 10598 17640 10654 17649
rect 10598 17575 10654 17584
rect 10214 17436 10522 17456
rect 10214 17434 10220 17436
rect 10276 17434 10300 17436
rect 10356 17434 10380 17436
rect 10436 17434 10460 17436
rect 10516 17434 10522 17436
rect 10276 17382 10278 17434
rect 10458 17382 10460 17434
rect 10214 17380 10220 17382
rect 10276 17380 10300 17382
rect 10356 17380 10380 17382
rect 10436 17380 10460 17382
rect 10516 17380 10522 17382
rect 10214 17360 10522 17380
rect 10214 16348 10522 16368
rect 10214 16346 10220 16348
rect 10276 16346 10300 16348
rect 10356 16346 10380 16348
rect 10436 16346 10460 16348
rect 10516 16346 10522 16348
rect 10276 16294 10278 16346
rect 10458 16294 10460 16346
rect 10214 16292 10220 16294
rect 10276 16292 10300 16294
rect 10356 16292 10380 16294
rect 10436 16292 10460 16294
rect 10516 16292 10522 16294
rect 10214 16272 10522 16292
rect 10214 15260 10522 15280
rect 10214 15258 10220 15260
rect 10276 15258 10300 15260
rect 10356 15258 10380 15260
rect 10436 15258 10460 15260
rect 10516 15258 10522 15260
rect 10276 15206 10278 15258
rect 10458 15206 10460 15258
rect 10214 15204 10220 15206
rect 10276 15204 10300 15206
rect 10356 15204 10380 15206
rect 10436 15204 10460 15206
rect 10516 15204 10522 15206
rect 10214 15184 10522 15204
rect 10214 14172 10522 14192
rect 10214 14170 10220 14172
rect 10276 14170 10300 14172
rect 10356 14170 10380 14172
rect 10436 14170 10460 14172
rect 10516 14170 10522 14172
rect 10276 14118 10278 14170
rect 10458 14118 10460 14170
rect 10214 14116 10220 14118
rect 10276 14116 10300 14118
rect 10356 14116 10380 14118
rect 10436 14116 10460 14118
rect 10516 14116 10522 14118
rect 10214 14096 10522 14116
rect 10214 13084 10522 13104
rect 10214 13082 10220 13084
rect 10276 13082 10300 13084
rect 10356 13082 10380 13084
rect 10436 13082 10460 13084
rect 10516 13082 10522 13084
rect 10276 13030 10278 13082
rect 10458 13030 10460 13082
rect 10214 13028 10220 13030
rect 10276 13028 10300 13030
rect 10356 13028 10380 13030
rect 10436 13028 10460 13030
rect 10516 13028 10522 13030
rect 10214 13008 10522 13028
rect 10214 11996 10522 12016
rect 10214 11994 10220 11996
rect 10276 11994 10300 11996
rect 10356 11994 10380 11996
rect 10436 11994 10460 11996
rect 10516 11994 10522 11996
rect 10276 11942 10278 11994
rect 10458 11942 10460 11994
rect 10214 11940 10220 11942
rect 10276 11940 10300 11942
rect 10356 11940 10380 11942
rect 10436 11940 10460 11942
rect 10516 11940 10522 11942
rect 10214 11920 10522 11940
rect 10140 11620 10192 11626
rect 10140 11562 10192 11568
rect 10214 10908 10522 10928
rect 10214 10906 10220 10908
rect 10276 10906 10300 10908
rect 10356 10906 10380 10908
rect 10436 10906 10460 10908
rect 10516 10906 10522 10908
rect 10276 10854 10278 10906
rect 10458 10854 10460 10906
rect 10214 10852 10220 10854
rect 10276 10852 10300 10854
rect 10356 10852 10380 10854
rect 10436 10852 10460 10854
rect 10516 10852 10522 10854
rect 10214 10832 10522 10852
rect 10214 9820 10522 9840
rect 10214 9818 10220 9820
rect 10276 9818 10300 9820
rect 10356 9818 10380 9820
rect 10436 9818 10460 9820
rect 10516 9818 10522 9820
rect 10276 9766 10278 9818
rect 10458 9766 10460 9818
rect 10214 9764 10220 9766
rect 10276 9764 10300 9766
rect 10356 9764 10380 9766
rect 10436 9764 10460 9766
rect 10516 9764 10522 9766
rect 10214 9744 10522 9764
rect 10214 8732 10522 8752
rect 10214 8730 10220 8732
rect 10276 8730 10300 8732
rect 10356 8730 10380 8732
rect 10436 8730 10460 8732
rect 10516 8730 10522 8732
rect 10276 8678 10278 8730
rect 10458 8678 10460 8730
rect 10214 8676 10220 8678
rect 10276 8676 10300 8678
rect 10356 8676 10380 8678
rect 10436 8676 10460 8678
rect 10516 8676 10522 8678
rect 10214 8656 10522 8676
rect 10214 7644 10522 7664
rect 10214 7642 10220 7644
rect 10276 7642 10300 7644
rect 10356 7642 10380 7644
rect 10436 7642 10460 7644
rect 10516 7642 10522 7644
rect 10276 7590 10278 7642
rect 10458 7590 10460 7642
rect 10214 7588 10220 7590
rect 10276 7588 10300 7590
rect 10356 7588 10380 7590
rect 10436 7588 10460 7590
rect 10516 7588 10522 7590
rect 10214 7568 10522 7588
rect 12544 6914 12572 25162
rect 12622 25120 12678 25129
rect 12622 25055 12678 25064
rect 12636 24410 12664 25055
rect 12728 24750 12756 25366
rect 13188 25226 13216 26574
rect 13360 26444 13412 26450
rect 13360 26386 13412 26392
rect 13268 26240 13320 26246
rect 13268 26182 13320 26188
rect 13280 25906 13308 26182
rect 13268 25900 13320 25906
rect 13268 25842 13320 25848
rect 13372 25412 13400 26386
rect 13280 25384 13400 25412
rect 13176 25220 13228 25226
rect 13176 25162 13228 25168
rect 12990 24984 13046 24993
rect 12990 24919 12992 24928
rect 13044 24919 13046 24928
rect 13174 24984 13230 24993
rect 13174 24919 13230 24928
rect 12992 24890 13044 24896
rect 12716 24744 12768 24750
rect 12716 24686 12768 24692
rect 12808 24744 12860 24750
rect 12808 24686 12860 24692
rect 12624 24404 12676 24410
rect 12624 24346 12676 24352
rect 12716 23724 12768 23730
rect 12716 23666 12768 23672
rect 12622 23080 12678 23089
rect 12622 23015 12678 23024
rect 12636 22642 12664 23015
rect 12624 22636 12676 22642
rect 12624 22578 12676 22584
rect 12622 21448 12678 21457
rect 12622 21383 12678 21392
rect 12636 20806 12664 21383
rect 12624 20800 12676 20806
rect 12624 20742 12676 20748
rect 12728 18902 12756 23666
rect 12820 21962 12848 24686
rect 13082 24440 13138 24449
rect 13082 24375 13138 24384
rect 12898 24304 12954 24313
rect 12898 24239 12954 24248
rect 12992 24268 13044 24274
rect 12912 24206 12940 24239
rect 12992 24210 13044 24216
rect 12900 24200 12952 24206
rect 12900 24142 12952 24148
rect 12808 21956 12860 21962
rect 12808 21898 12860 21904
rect 12716 18896 12768 18902
rect 12716 18838 12768 18844
rect 12820 18698 12848 21898
rect 12900 21480 12952 21486
rect 12900 21422 12952 21428
rect 12912 20058 12940 21422
rect 13004 20777 13032 24210
rect 13096 23730 13124 24375
rect 13188 23798 13216 24919
rect 13280 24682 13308 25384
rect 13360 25220 13412 25226
rect 13360 25162 13412 25168
rect 13268 24676 13320 24682
rect 13268 24618 13320 24624
rect 13266 24168 13322 24177
rect 13266 24103 13322 24112
rect 13176 23792 13228 23798
rect 13176 23734 13228 23740
rect 13280 23730 13308 24103
rect 13084 23724 13136 23730
rect 13084 23666 13136 23672
rect 13268 23724 13320 23730
rect 13268 23666 13320 23672
rect 13372 23322 13400 25162
rect 13360 23316 13412 23322
rect 13360 23258 13412 23264
rect 13464 23118 13492 27066
rect 13544 26920 13596 26926
rect 13544 26862 13596 26868
rect 13556 26586 13584 26862
rect 13544 26580 13596 26586
rect 13544 26522 13596 26528
rect 13544 25968 13596 25974
rect 13544 25910 13596 25916
rect 13556 25838 13584 25910
rect 13544 25832 13596 25838
rect 13544 25774 13596 25780
rect 13544 24268 13596 24274
rect 13648 24256 13676 27231
rect 13740 26790 13768 28562
rect 13924 28218 13952 28902
rect 13912 28212 13964 28218
rect 13912 28154 13964 28160
rect 14004 28212 14056 28218
rect 14004 28154 14056 28160
rect 14016 28098 14044 28154
rect 13924 28070 14044 28098
rect 13820 28008 13872 28014
rect 13820 27950 13872 27956
rect 13832 27470 13860 27950
rect 13820 27464 13872 27470
rect 13820 27406 13872 27412
rect 13820 26988 13872 26994
rect 13820 26930 13872 26936
rect 13728 26784 13780 26790
rect 13728 26726 13780 26732
rect 13832 26314 13860 26930
rect 13924 26450 13952 28070
rect 14108 28014 14136 29174
rect 14186 28792 14242 28801
rect 14186 28727 14242 28736
rect 14200 28626 14228 28727
rect 14188 28620 14240 28626
rect 14188 28562 14240 28568
rect 14292 28150 14320 31855
rect 14384 31346 14412 32320
rect 14568 31754 14596 32778
rect 14844 32722 14872 32914
rect 14660 32694 14872 32722
rect 14660 32201 14688 32694
rect 15304 32230 15332 33816
rect 15396 32910 15424 34303
rect 15488 33386 15516 34410
rect 15672 33998 15700 35090
rect 16118 34776 16174 34785
rect 16118 34711 16174 34720
rect 16132 34678 16160 34711
rect 16120 34672 16172 34678
rect 16120 34614 16172 34620
rect 15936 34604 15988 34610
rect 15936 34546 15988 34552
rect 15948 34456 15976 34546
rect 16212 34468 16264 34474
rect 15948 34428 16212 34456
rect 15948 34202 15976 34428
rect 16212 34410 16264 34416
rect 15936 34196 15988 34202
rect 15936 34138 15988 34144
rect 15660 33992 15712 33998
rect 15660 33934 15712 33940
rect 15568 33652 15620 33658
rect 15568 33594 15620 33600
rect 15580 33425 15608 33594
rect 15672 33522 15700 33934
rect 15660 33516 15712 33522
rect 15660 33458 15712 33464
rect 15566 33416 15622 33425
rect 15476 33380 15528 33386
rect 15566 33351 15622 33360
rect 15476 33322 15528 33328
rect 15672 32978 15700 33458
rect 16316 33386 16344 35278
rect 16396 35012 16448 35018
rect 16396 34954 16448 34960
rect 16304 33380 16356 33386
rect 16304 33322 16356 33328
rect 15660 32972 15712 32978
rect 15660 32914 15712 32920
rect 15384 32904 15436 32910
rect 15384 32846 15436 32852
rect 15292 32224 15344 32230
rect 14646 32192 14702 32201
rect 15292 32166 15344 32172
rect 14646 32127 14702 32136
rect 14846 32124 15154 32144
rect 14846 32122 14852 32124
rect 14908 32122 14932 32124
rect 14988 32122 15012 32124
rect 15068 32122 15092 32124
rect 15148 32122 15154 32124
rect 14908 32070 14910 32122
rect 15090 32070 15092 32122
rect 14846 32068 14852 32070
rect 14908 32068 14932 32070
rect 14988 32068 15012 32070
rect 15068 32068 15092 32070
rect 15148 32068 15154 32070
rect 14846 32048 15154 32068
rect 15290 32056 15346 32065
rect 15200 32020 15252 32026
rect 15290 31991 15346 32000
rect 15200 31962 15252 31968
rect 15212 31906 15240 31962
rect 14660 31878 15240 31906
rect 14556 31748 14608 31754
rect 14556 31690 14608 31696
rect 14464 31476 14516 31482
rect 14464 31418 14516 31424
rect 14372 31340 14424 31346
rect 14372 31282 14424 31288
rect 14384 30734 14412 31282
rect 14476 31278 14504 31418
rect 14464 31272 14516 31278
rect 14464 31214 14516 31220
rect 14660 31192 14688 31878
rect 14740 31816 14792 31822
rect 14740 31758 14792 31764
rect 14830 31784 14886 31793
rect 14752 31346 14780 31758
rect 15198 31784 15254 31793
rect 14830 31719 14832 31728
rect 14884 31719 14886 31728
rect 15120 31728 15198 31754
rect 15120 31726 15254 31728
rect 14832 31690 14884 31696
rect 15120 31385 15148 31726
rect 15198 31719 15254 31726
rect 15200 31476 15252 31482
rect 15200 31418 15252 31424
rect 15106 31376 15162 31385
rect 14740 31340 14792 31346
rect 15106 31311 15162 31320
rect 14740 31282 14792 31288
rect 15212 31249 15240 31418
rect 14568 31164 14688 31192
rect 15198 31240 15254 31249
rect 15198 31175 15254 31184
rect 14462 30968 14518 30977
rect 14462 30903 14518 30912
rect 14372 30728 14424 30734
rect 14372 30670 14424 30676
rect 14476 30569 14504 30903
rect 14568 30802 14596 31164
rect 15304 31124 15332 31991
rect 14660 31113 15332 31124
rect 14646 31104 15332 31113
rect 14702 31096 15332 31104
rect 14646 31039 14702 31048
rect 14846 31036 15154 31056
rect 14846 31034 14852 31036
rect 14908 31034 14932 31036
rect 14988 31034 15012 31036
rect 15068 31034 15092 31036
rect 15148 31034 15154 31036
rect 14908 30982 14910 31034
rect 15090 30982 15092 31034
rect 14846 30980 14852 30982
rect 14908 30980 14932 30982
rect 14988 30980 15012 30982
rect 15068 30980 15092 30982
rect 15148 30980 15154 30982
rect 14846 30960 15154 30980
rect 15396 30938 15424 32846
rect 15672 31890 15700 32914
rect 16304 32768 16356 32774
rect 16304 32710 16356 32716
rect 16212 32292 16264 32298
rect 16212 32234 16264 32240
rect 15936 32224 15988 32230
rect 15936 32166 15988 32172
rect 15660 31884 15712 31890
rect 15660 31826 15712 31832
rect 15844 31340 15896 31346
rect 15844 31282 15896 31288
rect 15474 30968 15530 30977
rect 15384 30932 15436 30938
rect 15474 30903 15530 30912
rect 15384 30874 15436 30880
rect 14556 30796 14608 30802
rect 14556 30738 14608 30744
rect 14462 30560 14518 30569
rect 14462 30495 14518 30504
rect 14372 30320 14424 30326
rect 14372 30262 14424 30268
rect 14384 29889 14412 30262
rect 14370 29880 14426 29889
rect 14370 29815 14426 29824
rect 14462 29608 14518 29617
rect 14462 29543 14518 29552
rect 14372 28552 14424 28558
rect 14372 28494 14424 28500
rect 14280 28144 14332 28150
rect 14280 28086 14332 28092
rect 14096 28008 14148 28014
rect 14096 27950 14148 27956
rect 14004 27872 14056 27878
rect 14004 27814 14056 27820
rect 14016 27402 14044 27814
rect 14108 27470 14136 27950
rect 14186 27840 14242 27849
rect 14186 27775 14242 27784
rect 14096 27464 14148 27470
rect 14096 27406 14148 27412
rect 14004 27396 14056 27402
rect 14004 27338 14056 27344
rect 14200 27062 14228 27775
rect 14188 27056 14240 27062
rect 14188 26998 14240 27004
rect 14096 26988 14148 26994
rect 14096 26930 14148 26936
rect 14004 26852 14056 26858
rect 14004 26794 14056 26800
rect 13912 26444 13964 26450
rect 13912 26386 13964 26392
rect 14016 26314 14044 26794
rect 13820 26308 13872 26314
rect 13820 26250 13872 26256
rect 14004 26308 14056 26314
rect 14004 26250 14056 26256
rect 13818 25936 13874 25945
rect 13818 25871 13820 25880
rect 13872 25871 13874 25880
rect 13820 25842 13872 25848
rect 13728 25696 13780 25702
rect 13728 25638 13780 25644
rect 13740 24954 13768 25638
rect 14004 25424 14056 25430
rect 14004 25366 14056 25372
rect 14016 25158 14044 25366
rect 14004 25152 14056 25158
rect 14004 25094 14056 25100
rect 13728 24948 13780 24954
rect 13780 24908 13860 24936
rect 13728 24890 13780 24896
rect 13728 24336 13780 24342
rect 13728 24278 13780 24284
rect 13596 24228 13676 24256
rect 13544 24210 13596 24216
rect 13740 24154 13768 24278
rect 13648 24126 13768 24154
rect 13648 23866 13676 24126
rect 13728 24064 13780 24070
rect 13728 24006 13780 24012
rect 13636 23860 13688 23866
rect 13636 23802 13688 23808
rect 13740 23730 13768 24006
rect 13728 23724 13780 23730
rect 13728 23666 13780 23672
rect 13636 23316 13688 23322
rect 13688 23276 13768 23304
rect 13636 23258 13688 23264
rect 13268 23112 13320 23118
rect 13268 23054 13320 23060
rect 13452 23112 13504 23118
rect 13452 23054 13504 23060
rect 13740 23066 13768 23276
rect 13832 23186 13860 24908
rect 14004 24880 14056 24886
rect 14002 24848 14004 24857
rect 14056 24848 14058 24857
rect 13912 24812 13964 24818
rect 14002 24783 14058 24792
rect 13912 24754 13964 24760
rect 13924 24154 13952 24754
rect 13924 24126 14044 24154
rect 14016 23746 14044 24126
rect 14108 23866 14136 26930
rect 14280 26376 14332 26382
rect 14200 26336 14280 26364
rect 14200 24954 14228 26336
rect 14280 26318 14332 26324
rect 14280 25288 14332 25294
rect 14280 25230 14332 25236
rect 14188 24948 14240 24954
rect 14188 24890 14240 24896
rect 14200 24721 14228 24890
rect 14292 24750 14320 25230
rect 14280 24744 14332 24750
rect 14186 24712 14242 24721
rect 14280 24686 14332 24692
rect 14186 24647 14242 24656
rect 14384 24562 14412 28494
rect 14476 27713 14504 29543
rect 14462 27704 14518 27713
rect 14462 27639 14518 27648
rect 14568 26790 14596 30738
rect 15488 30734 15516 30903
rect 15856 30734 15884 31282
rect 14740 30728 14792 30734
rect 14740 30670 14792 30676
rect 15200 30728 15252 30734
rect 15200 30670 15252 30676
rect 15476 30728 15528 30734
rect 15476 30670 15528 30676
rect 15844 30728 15896 30734
rect 15844 30670 15896 30676
rect 14752 29832 14780 30670
rect 14846 29948 15154 29968
rect 14846 29946 14852 29948
rect 14908 29946 14932 29948
rect 14988 29946 15012 29948
rect 15068 29946 15092 29948
rect 15148 29946 15154 29948
rect 14908 29894 14910 29946
rect 15090 29894 15092 29946
rect 14846 29892 14852 29894
rect 14908 29892 14932 29894
rect 14988 29892 15012 29894
rect 15068 29892 15092 29894
rect 15148 29892 15154 29894
rect 14846 29872 15154 29892
rect 14752 29804 15056 29832
rect 14648 29776 14700 29782
rect 14648 29718 14700 29724
rect 14660 28948 14688 29718
rect 15028 29170 15056 29804
rect 15212 29209 15240 30670
rect 15292 30660 15344 30666
rect 15292 30602 15344 30608
rect 15304 30394 15332 30602
rect 15856 30394 15884 30670
rect 15292 30388 15344 30394
rect 15292 30330 15344 30336
rect 15844 30388 15896 30394
rect 15844 30330 15896 30336
rect 15292 30252 15344 30258
rect 15292 30194 15344 30200
rect 15384 30252 15436 30258
rect 15384 30194 15436 30200
rect 15844 30252 15896 30258
rect 15844 30194 15896 30200
rect 15304 29889 15332 30194
rect 15290 29880 15346 29889
rect 15290 29815 15346 29824
rect 15198 29200 15254 29209
rect 15016 29164 15068 29170
rect 15198 29135 15254 29144
rect 15016 29106 15068 29112
rect 14660 28937 15332 28948
rect 14660 28928 15346 28937
rect 14660 28920 15290 28928
rect 14846 28860 15154 28880
rect 15290 28863 15346 28872
rect 14846 28858 14852 28860
rect 14908 28858 14932 28860
rect 14988 28858 15012 28860
rect 15068 28858 15092 28860
rect 15148 28858 15154 28860
rect 14908 28806 14910 28858
rect 15090 28806 15092 28858
rect 14846 28804 14852 28806
rect 14908 28804 14932 28806
rect 14988 28804 15012 28806
rect 15068 28804 15092 28806
rect 15148 28804 15154 28806
rect 14846 28784 15154 28804
rect 15290 28792 15346 28801
rect 15290 28727 15346 28736
rect 15304 28642 15332 28727
rect 14660 28614 15332 28642
rect 14660 28558 14688 28614
rect 14648 28552 14700 28558
rect 14648 28494 14700 28500
rect 14740 28552 14792 28558
rect 14740 28494 14792 28500
rect 14648 28212 14700 28218
rect 14648 28154 14700 28160
rect 14660 26994 14688 28154
rect 14752 27334 14780 28494
rect 15292 28144 15344 28150
rect 15292 28086 15344 28092
rect 14846 27772 15154 27792
rect 14846 27770 14852 27772
rect 14908 27770 14932 27772
rect 14988 27770 15012 27772
rect 15068 27770 15092 27772
rect 15148 27770 15154 27772
rect 14908 27718 14910 27770
rect 15090 27718 15092 27770
rect 14846 27716 14852 27718
rect 14908 27716 14932 27718
rect 14988 27716 15012 27718
rect 15068 27716 15092 27718
rect 15148 27716 15154 27718
rect 14846 27696 15154 27716
rect 15108 27600 15160 27606
rect 14936 27560 15108 27588
rect 14740 27328 14792 27334
rect 14740 27270 14792 27276
rect 14752 26994 14780 27270
rect 14648 26988 14700 26994
rect 14648 26930 14700 26936
rect 14740 26988 14792 26994
rect 14740 26930 14792 26936
rect 14556 26784 14608 26790
rect 14936 26772 14964 27560
rect 15108 27542 15160 27548
rect 15200 27328 15252 27334
rect 15200 27270 15252 27276
rect 15016 26988 15068 26994
rect 15016 26930 15068 26936
rect 15028 26858 15056 26930
rect 15016 26852 15068 26858
rect 15016 26794 15068 26800
rect 14556 26726 14608 26732
rect 14660 26744 14964 26772
rect 14568 26450 14596 26726
rect 14556 26444 14608 26450
rect 14556 26386 14608 26392
rect 14554 25800 14610 25809
rect 14554 25735 14610 25744
rect 14568 25702 14596 25735
rect 14556 25696 14608 25702
rect 14660 25673 14688 26744
rect 14846 26684 15154 26704
rect 14846 26682 14852 26684
rect 14908 26682 14932 26684
rect 14988 26682 15012 26684
rect 15068 26682 15092 26684
rect 15148 26682 15154 26684
rect 14908 26630 14910 26682
rect 15090 26630 15092 26682
rect 14846 26628 14852 26630
rect 14908 26628 14932 26630
rect 14988 26628 15012 26630
rect 15068 26628 15092 26630
rect 15148 26628 15154 26630
rect 14846 26608 15154 26628
rect 15212 26518 15240 27270
rect 15200 26512 15252 26518
rect 15120 26472 15200 26500
rect 14740 26444 14792 26450
rect 14924 26444 14976 26450
rect 14740 26386 14792 26392
rect 14844 26404 14924 26432
rect 14752 25752 14780 26386
rect 14844 25906 14872 26404
rect 14924 26386 14976 26392
rect 15120 26296 15148 26472
rect 15200 26454 15252 26460
rect 15304 26364 15332 28086
rect 15396 27985 15424 30194
rect 15856 30025 15884 30194
rect 15842 30016 15898 30025
rect 15842 29951 15898 29960
rect 15752 29776 15804 29782
rect 15752 29718 15804 29724
rect 15660 29572 15712 29578
rect 15660 29514 15712 29520
rect 15568 29232 15620 29238
rect 15474 29200 15530 29209
rect 15568 29174 15620 29180
rect 15474 29135 15530 29144
rect 15488 28218 15516 29135
rect 15580 28966 15608 29174
rect 15672 29034 15700 29514
rect 15764 29238 15792 29718
rect 15948 29345 15976 32166
rect 16224 31249 16252 32234
rect 16316 31686 16344 32710
rect 16304 31680 16356 31686
rect 16304 31622 16356 31628
rect 16316 31385 16344 31622
rect 16302 31376 16358 31385
rect 16302 31311 16358 31320
rect 16210 31240 16266 31249
rect 16210 31175 16266 31184
rect 16028 31136 16080 31142
rect 16028 31078 16080 31084
rect 16040 30598 16068 31078
rect 16212 30660 16264 30666
rect 16212 30602 16264 30608
rect 16028 30592 16080 30598
rect 16028 30534 16080 30540
rect 16120 30592 16172 30598
rect 16120 30534 16172 30540
rect 15934 29336 15990 29345
rect 15934 29271 15990 29280
rect 15752 29232 15804 29238
rect 15752 29174 15804 29180
rect 15660 29028 15712 29034
rect 15660 28970 15712 28976
rect 16040 28966 16068 30534
rect 16132 29238 16160 30534
rect 16224 29782 16252 30602
rect 16304 30388 16356 30394
rect 16304 30330 16356 30336
rect 16212 29776 16264 29782
rect 16212 29718 16264 29724
rect 16120 29232 16172 29238
rect 16120 29174 16172 29180
rect 16316 29170 16344 30330
rect 16304 29164 16356 29170
rect 16304 29106 16356 29112
rect 15568 28960 15620 28966
rect 15568 28902 15620 28908
rect 16028 28960 16080 28966
rect 16028 28902 16080 28908
rect 16304 28552 16356 28558
rect 16304 28494 16356 28500
rect 16120 28416 16172 28422
rect 16120 28358 16172 28364
rect 16132 28218 16160 28358
rect 15476 28212 15528 28218
rect 15476 28154 15528 28160
rect 15844 28212 15896 28218
rect 15844 28154 15896 28160
rect 16120 28212 16172 28218
rect 16120 28154 16172 28160
rect 15382 27976 15438 27985
rect 15382 27911 15384 27920
rect 15436 27911 15438 27920
rect 15384 27882 15436 27888
rect 15396 27851 15424 27882
rect 15752 27532 15804 27538
rect 15752 27474 15804 27480
rect 15660 26988 15712 26994
rect 15660 26930 15712 26936
rect 15568 26920 15620 26926
rect 15568 26862 15620 26868
rect 15476 26784 15528 26790
rect 15476 26726 15528 26732
rect 15304 26353 15424 26364
rect 15304 26344 15438 26353
rect 15304 26336 15382 26344
rect 14936 26268 15148 26296
rect 15382 26279 15438 26288
rect 14936 26058 14964 26268
rect 15200 26240 15252 26246
rect 15488 26234 15516 26726
rect 15580 26602 15608 26862
rect 15672 26761 15700 26930
rect 15658 26752 15714 26761
rect 15658 26687 15714 26696
rect 15580 26574 15700 26602
rect 15568 26444 15620 26450
rect 15568 26386 15620 26392
rect 15580 26353 15608 26386
rect 15566 26344 15622 26353
rect 15566 26279 15622 26288
rect 15488 26206 15608 26234
rect 15200 26182 15252 26188
rect 14936 26030 15056 26058
rect 15028 26024 15056 26030
rect 15028 25996 15148 26024
rect 15120 25906 15148 25996
rect 15212 25956 15240 26182
rect 15212 25928 15333 25956
rect 15305 25922 15333 25928
rect 14832 25900 14884 25906
rect 14832 25842 14884 25848
rect 15016 25900 15068 25906
rect 15016 25842 15068 25848
rect 15108 25900 15160 25906
rect 15305 25894 15424 25922
rect 15108 25842 15160 25848
rect 15028 25752 15056 25842
rect 14752 25724 15056 25752
rect 15396 25752 15424 25894
rect 15580 25888 15608 26206
rect 15672 25956 15700 26574
rect 15764 26450 15792 27474
rect 15856 26994 15884 28154
rect 16210 27840 16266 27849
rect 16210 27775 16266 27784
rect 15936 27668 15988 27674
rect 15936 27610 15988 27616
rect 15948 27402 15976 27610
rect 16224 27606 16252 27775
rect 16212 27600 16264 27606
rect 16212 27542 16264 27548
rect 15936 27396 15988 27402
rect 15936 27338 15988 27344
rect 15844 26988 15896 26994
rect 15844 26930 15896 26936
rect 15752 26444 15804 26450
rect 15752 26386 15804 26392
rect 15672 25928 15711 25956
rect 15580 25860 15655 25888
rect 15474 25800 15530 25809
rect 15396 25744 15474 25752
rect 15627 25786 15655 25860
rect 15396 25735 15530 25744
rect 15562 25758 15655 25786
rect 15396 25724 15516 25735
rect 15562 25684 15590 25758
rect 15683 25702 15711 25928
rect 15752 25832 15804 25838
rect 15856 25820 15884 26930
rect 16120 26784 16172 26790
rect 16120 26726 16172 26732
rect 15936 26240 15988 26246
rect 15936 26182 15988 26188
rect 15804 25792 15884 25820
rect 15752 25774 15804 25780
rect 14556 25638 14608 25644
rect 14646 25664 14702 25673
rect 15290 25664 15346 25673
rect 15212 25622 15290 25650
rect 14646 25599 14702 25608
rect 14846 25596 15154 25616
rect 14846 25594 14852 25596
rect 14908 25594 14932 25596
rect 14988 25594 15012 25596
rect 15068 25594 15092 25596
rect 15148 25594 15154 25596
rect 14908 25542 14910 25594
rect 15090 25542 15092 25594
rect 14846 25540 14852 25542
rect 14908 25540 14932 25542
rect 14988 25540 15012 25542
rect 15068 25540 15092 25542
rect 15148 25540 15154 25542
rect 14846 25520 15154 25540
rect 15212 25378 15240 25622
rect 15290 25599 15346 25608
rect 15488 25656 15590 25684
rect 15660 25696 15712 25702
rect 14476 25350 14780 25378
rect 14476 25294 14504 25350
rect 14464 25288 14516 25294
rect 14464 25230 14516 25236
rect 14648 25288 14700 25294
rect 14648 25230 14700 25236
rect 14556 24948 14608 24954
rect 14556 24890 14608 24896
rect 14292 24534 14412 24562
rect 14464 24608 14516 24614
rect 14464 24550 14516 24556
rect 14096 23860 14148 23866
rect 14096 23802 14148 23808
rect 14188 23860 14240 23866
rect 14188 23802 14240 23808
rect 13912 23724 13964 23730
rect 14016 23718 14136 23746
rect 13912 23666 13964 23672
rect 13924 23633 13952 23666
rect 13910 23624 13966 23633
rect 13966 23582 14044 23610
rect 13910 23559 13966 23568
rect 13820 23180 13872 23186
rect 13820 23122 13872 23128
rect 13176 22636 13228 22642
rect 13176 22578 13228 22584
rect 13188 21876 13216 22578
rect 13280 22545 13308 23054
rect 13266 22536 13322 22545
rect 13266 22471 13322 22480
rect 13360 22024 13412 22030
rect 13358 21992 13360 22001
rect 13412 21992 13414 22001
rect 13464 21962 13492 23054
rect 13740 23038 13860 23066
rect 13726 22808 13782 22817
rect 13544 22772 13596 22778
rect 13726 22743 13782 22752
rect 13544 22714 13596 22720
rect 13358 21927 13414 21936
rect 13452 21956 13504 21962
rect 13452 21898 13504 21904
rect 13188 21848 13400 21876
rect 13176 21140 13228 21146
rect 13176 21082 13228 21088
rect 13084 20936 13136 20942
rect 13084 20878 13136 20884
rect 12990 20768 13046 20777
rect 12990 20703 13046 20712
rect 12900 20052 12952 20058
rect 12900 19994 12952 20000
rect 13096 19446 13124 20878
rect 13188 20262 13216 21082
rect 13268 20936 13320 20942
rect 13268 20878 13320 20884
rect 13280 20641 13308 20878
rect 13266 20632 13322 20641
rect 13266 20567 13322 20576
rect 13176 20256 13228 20262
rect 13176 20198 13228 20204
rect 13372 19514 13400 21848
rect 13556 20380 13584 22714
rect 13636 21956 13688 21962
rect 13636 21898 13688 21904
rect 13648 21865 13676 21898
rect 13634 21856 13690 21865
rect 13634 21791 13690 21800
rect 13648 21554 13676 21791
rect 13740 21622 13768 22743
rect 13728 21616 13780 21622
rect 13728 21558 13780 21564
rect 13636 21548 13688 21554
rect 13636 21490 13688 21496
rect 13636 21004 13688 21010
rect 13636 20946 13688 20952
rect 13648 20505 13676 20946
rect 13634 20496 13690 20505
rect 13634 20431 13690 20440
rect 13556 20352 13676 20380
rect 13544 19848 13596 19854
rect 13544 19790 13596 19796
rect 13360 19508 13412 19514
rect 13360 19450 13412 19456
rect 13084 19440 13136 19446
rect 13084 19382 13136 19388
rect 13556 19310 13584 19790
rect 13544 19304 13596 19310
rect 13544 19246 13596 19252
rect 12808 18692 12860 18698
rect 12808 18634 12860 18640
rect 13648 18290 13676 20352
rect 13636 18284 13688 18290
rect 13636 18226 13688 18232
rect 13832 15434 13860 23038
rect 13912 22568 13964 22574
rect 13912 22510 13964 22516
rect 13924 21554 13952 22510
rect 14016 22030 14044 23582
rect 14108 22642 14136 23718
rect 14200 23225 14228 23802
rect 14186 23216 14242 23225
rect 14186 23151 14242 23160
rect 14188 22976 14240 22982
rect 14186 22944 14188 22953
rect 14240 22944 14242 22953
rect 14186 22879 14242 22888
rect 14096 22636 14148 22642
rect 14096 22578 14148 22584
rect 14004 22024 14056 22030
rect 14004 21966 14056 21972
rect 14186 21992 14242 22001
rect 14186 21927 14242 21936
rect 13912 21548 13964 21554
rect 13912 21490 13964 21496
rect 13924 21146 13952 21490
rect 13912 21140 13964 21146
rect 13912 21082 13964 21088
rect 14096 21072 14148 21078
rect 13910 21040 13966 21049
rect 14096 21014 14148 21020
rect 13910 20975 13966 20984
rect 14004 21004 14056 21010
rect 13924 20806 13952 20975
rect 14004 20946 14056 20952
rect 13912 20800 13964 20806
rect 13912 20742 13964 20748
rect 14016 20466 14044 20946
rect 14108 20602 14136 21014
rect 14096 20596 14148 20602
rect 14096 20538 14148 20544
rect 14004 20460 14056 20466
rect 14004 20402 14056 20408
rect 14200 19854 14228 21927
rect 14188 19848 14240 19854
rect 14188 19790 14240 19796
rect 14200 18834 14228 19790
rect 14188 18828 14240 18834
rect 14188 18770 14240 18776
rect 14188 18352 14240 18358
rect 14186 18320 14188 18329
rect 14240 18320 14242 18329
rect 14186 18255 14242 18264
rect 13820 15428 13872 15434
rect 13820 15370 13872 15376
rect 12992 13864 13044 13870
rect 12992 13806 13044 13812
rect 13004 11694 13032 13806
rect 12992 11688 13044 11694
rect 12992 11630 13044 11636
rect 12452 6886 12572 6914
rect 10214 6556 10522 6576
rect 10214 6554 10220 6556
rect 10276 6554 10300 6556
rect 10356 6554 10380 6556
rect 10436 6554 10460 6556
rect 10516 6554 10522 6556
rect 10276 6502 10278 6554
rect 10458 6502 10460 6554
rect 10214 6500 10220 6502
rect 10276 6500 10300 6502
rect 10356 6500 10380 6502
rect 10436 6500 10460 6502
rect 10516 6500 10522 6502
rect 10214 6480 10522 6500
rect 10214 5468 10522 5488
rect 10214 5466 10220 5468
rect 10276 5466 10300 5468
rect 10356 5466 10380 5468
rect 10436 5466 10460 5468
rect 10516 5466 10522 5468
rect 10276 5414 10278 5466
rect 10458 5414 10460 5466
rect 10214 5412 10220 5414
rect 10276 5412 10300 5414
rect 10356 5412 10380 5414
rect 10436 5412 10460 5414
rect 10516 5412 10522 5414
rect 10214 5392 10522 5412
rect 10214 4380 10522 4400
rect 10214 4378 10220 4380
rect 10276 4378 10300 4380
rect 10356 4378 10380 4380
rect 10436 4378 10460 4380
rect 10516 4378 10522 4380
rect 10276 4326 10278 4378
rect 10458 4326 10460 4378
rect 10214 4324 10220 4326
rect 10276 4324 10300 4326
rect 10356 4324 10380 4326
rect 10436 4324 10460 4326
rect 10516 4324 10522 4326
rect 10214 4304 10522 4324
rect 10324 3936 10376 3942
rect 10324 3878 10376 3884
rect 10336 3670 10364 3878
rect 12452 3754 12480 6886
rect 12900 4140 12952 4146
rect 12900 4082 12952 4088
rect 12532 4072 12584 4078
rect 12532 4014 12584 4020
rect 12360 3738 12480 3754
rect 12544 3738 12572 4014
rect 12348 3732 12480 3738
rect 12400 3726 12480 3732
rect 12348 3674 12400 3680
rect 10324 3664 10376 3670
rect 10324 3606 10376 3612
rect 11704 3528 11756 3534
rect 11704 3470 11756 3476
rect 10214 3292 10522 3312
rect 10214 3290 10220 3292
rect 10276 3290 10300 3292
rect 10356 3290 10380 3292
rect 10436 3290 10460 3292
rect 10516 3290 10522 3292
rect 10276 3238 10278 3290
rect 10458 3238 10460 3290
rect 10214 3236 10220 3238
rect 10276 3236 10300 3238
rect 10356 3236 10380 3238
rect 10436 3236 10460 3238
rect 10516 3236 10522 3238
rect 10214 3216 10522 3236
rect 11716 3058 11744 3470
rect 9772 3052 9824 3058
rect 9772 2994 9824 3000
rect 11704 3052 11756 3058
rect 11704 2994 11756 3000
rect 11888 2984 11940 2990
rect 11888 2926 11940 2932
rect 12256 2984 12308 2990
rect 12256 2926 12308 2932
rect 9772 2848 9824 2854
rect 9772 2790 9824 2796
rect 9784 2514 9812 2790
rect 11900 2650 11928 2926
rect 11888 2644 11940 2650
rect 11888 2586 11940 2592
rect 9772 2508 9824 2514
rect 9772 2450 9824 2456
rect 10214 2204 10522 2224
rect 10214 2202 10220 2204
rect 10276 2202 10300 2204
rect 10356 2202 10380 2204
rect 10436 2202 10460 2204
rect 10516 2202 10522 2204
rect 10276 2150 10278 2202
rect 10458 2150 10460 2202
rect 10214 2148 10220 2150
rect 10276 2148 10300 2150
rect 10356 2148 10380 2150
rect 10436 2148 10460 2150
rect 10516 2148 10522 2150
rect 10214 2128 10522 2148
rect 12268 800 12296 2926
rect 12452 2446 12480 3726
rect 12532 3732 12584 3738
rect 12532 3674 12584 3680
rect 12912 3670 12940 4082
rect 12900 3664 12952 3670
rect 12900 3606 12952 3612
rect 13004 3534 13032 11630
rect 14292 6914 14320 24534
rect 14370 24168 14426 24177
rect 14370 24103 14426 24112
rect 14384 24070 14412 24103
rect 14372 24064 14424 24070
rect 14372 24006 14424 24012
rect 14476 23225 14504 24550
rect 14568 24188 14596 24890
rect 14660 24585 14688 25230
rect 14752 24954 14780 25350
rect 15016 25356 15068 25362
rect 15120 25350 15240 25378
rect 15400 25356 15452 25362
rect 15120 25344 15148 25350
rect 15068 25316 15148 25344
rect 15016 25298 15068 25304
rect 15488 25344 15516 25656
rect 15660 25638 15712 25644
rect 15452 25316 15516 25344
rect 15566 25392 15622 25401
rect 15566 25327 15622 25336
rect 15400 25298 15452 25304
rect 15200 25288 15252 25294
rect 14844 25236 15200 25242
rect 14844 25230 15252 25236
rect 14844 25214 15240 25230
rect 14740 24948 14792 24954
rect 14740 24890 14792 24896
rect 14844 24750 14872 25214
rect 14924 25152 14976 25158
rect 14924 25094 14976 25100
rect 14832 24744 14884 24750
rect 14738 24712 14794 24721
rect 14832 24686 14884 24692
rect 14738 24647 14794 24656
rect 14646 24576 14702 24585
rect 14646 24511 14702 24520
rect 14646 24440 14702 24449
rect 14752 24410 14780 24647
rect 14936 24596 14964 25094
rect 15016 24948 15068 24954
rect 15068 24908 15240 24936
rect 15016 24890 15068 24896
rect 15212 24800 15240 24908
rect 15384 24812 15436 24818
rect 15212 24772 15384 24800
rect 15384 24754 15436 24760
rect 15488 24732 15516 25316
rect 15580 25158 15608 25327
rect 15764 25265 15792 25774
rect 15948 25294 15976 26182
rect 16028 25764 16080 25770
rect 16028 25706 16080 25712
rect 16040 25673 16068 25706
rect 16026 25664 16082 25673
rect 16026 25599 16082 25608
rect 16132 25362 16160 26726
rect 16212 25900 16264 25906
rect 16212 25842 16264 25848
rect 16120 25356 16172 25362
rect 16040 25316 16120 25344
rect 15936 25288 15988 25294
rect 15750 25256 15806 25265
rect 15936 25230 15988 25236
rect 15750 25191 15806 25200
rect 15568 25152 15620 25158
rect 15568 25094 15620 25100
rect 15844 25152 15896 25158
rect 15844 25094 15896 25100
rect 15752 24948 15804 24954
rect 15752 24890 15804 24896
rect 15488 24704 15700 24732
rect 15304 24636 15516 24664
rect 15304 24596 15332 24636
rect 14936 24568 15332 24596
rect 15382 24576 15438 24585
rect 14846 24508 15154 24528
rect 15382 24511 15438 24520
rect 14846 24506 14852 24508
rect 14908 24506 14932 24508
rect 14988 24506 15012 24508
rect 15068 24506 15092 24508
rect 15148 24506 15154 24508
rect 14908 24454 14910 24506
rect 15090 24454 15092 24506
rect 14846 24452 14852 24454
rect 14908 24452 14932 24454
rect 14988 24452 15012 24454
rect 15068 24452 15092 24454
rect 15148 24452 15154 24454
rect 14846 24432 15154 24452
rect 15290 24440 15346 24449
rect 14646 24375 14702 24384
rect 14740 24404 14792 24410
rect 14660 24290 14688 24375
rect 14740 24346 14792 24352
rect 15120 24384 15290 24392
rect 15120 24375 15346 24384
rect 15120 24364 15332 24375
rect 15120 24290 15148 24364
rect 14660 24262 15148 24290
rect 15016 24200 15068 24206
rect 14568 24160 14872 24188
rect 14556 24064 14608 24070
rect 14556 24006 14608 24012
rect 14568 23730 14596 24006
rect 14738 23760 14794 23769
rect 14556 23724 14608 23730
rect 14844 23746 14872 24160
rect 15016 24142 15068 24148
rect 15292 24200 15344 24206
rect 15396 24188 15424 24511
rect 15488 24206 15516 24636
rect 15672 24614 15700 24704
rect 15764 24614 15792 24890
rect 15660 24608 15712 24614
rect 15660 24550 15712 24556
rect 15752 24608 15804 24614
rect 15856 24585 15884 25094
rect 15948 24954 15976 25230
rect 15936 24948 15988 24954
rect 15936 24890 15988 24896
rect 15948 24818 15976 24890
rect 16040 24886 16068 25316
rect 16120 25298 16172 25304
rect 16224 25226 16252 25842
rect 16212 25220 16264 25226
rect 16212 25162 16264 25168
rect 16028 24880 16080 24886
rect 16120 24880 16172 24886
rect 16028 24822 16080 24828
rect 16118 24848 16120 24857
rect 16172 24848 16174 24857
rect 15936 24812 15988 24818
rect 16118 24783 16174 24792
rect 15936 24754 15988 24760
rect 16120 24608 16172 24614
rect 15752 24550 15804 24556
rect 15842 24576 15898 24585
rect 16026 24576 16082 24585
rect 15842 24511 15898 24520
rect 15948 24534 16026 24562
rect 15948 24449 15976 24534
rect 16120 24550 16172 24556
rect 16026 24511 16082 24520
rect 16132 24449 16160 24550
rect 15934 24440 15990 24449
rect 15934 24375 15990 24384
rect 16118 24440 16174 24449
rect 16118 24375 16174 24384
rect 15844 24336 15896 24342
rect 15844 24278 15896 24284
rect 15344 24160 15424 24188
rect 15456 24200 15516 24206
rect 15292 24142 15344 24148
rect 15508 24160 15516 24200
rect 15456 24142 15508 24148
rect 15028 23905 15056 24142
rect 15476 24064 15528 24070
rect 15476 24006 15528 24012
rect 15014 23896 15070 23905
rect 15198 23896 15254 23905
rect 15014 23831 15070 23840
rect 15120 23854 15198 23882
rect 15120 23780 15148 23854
rect 15198 23831 15254 23840
rect 14922 23760 14978 23769
rect 14844 23718 14922 23746
rect 14738 23695 14740 23704
rect 14556 23666 14608 23672
rect 14792 23695 14794 23704
rect 14922 23695 14978 23704
rect 15028 23752 15148 23780
rect 15488 23780 15516 24006
rect 15856 23905 15884 24278
rect 16028 24132 16080 24138
rect 15948 24092 16028 24120
rect 15842 23896 15898 23905
rect 15842 23831 15898 23840
rect 15488 23752 15562 23780
rect 14740 23666 14792 23672
rect 14462 23216 14518 23225
rect 14462 23151 14518 23160
rect 14568 23100 14596 23666
rect 15028 23662 15056 23752
rect 15200 23724 15252 23730
rect 15384 23724 15436 23730
rect 15252 23684 15332 23712
rect 15200 23666 15252 23672
rect 15016 23656 15068 23662
rect 15016 23598 15068 23604
rect 15304 23474 15332 23684
rect 15534 23712 15562 23752
rect 15436 23684 15562 23712
rect 15844 23724 15896 23730
rect 15384 23666 15436 23672
rect 15304 23446 15433 23474
rect 14846 23420 15154 23440
rect 14846 23418 14852 23420
rect 14908 23418 14932 23420
rect 14988 23418 15012 23420
rect 15068 23418 15092 23420
rect 15148 23418 15154 23420
rect 14908 23366 14910 23418
rect 15090 23366 15092 23418
rect 14846 23364 14852 23366
rect 14908 23364 14932 23366
rect 14988 23364 15012 23366
rect 15068 23364 15092 23366
rect 15148 23364 15154 23366
rect 14646 23352 14702 23361
rect 14846 23344 15154 23364
rect 15278 23352 15334 23361
rect 14702 23296 15278 23304
rect 15405 23338 15433 23446
rect 14646 23287 15334 23296
rect 15396 23310 15433 23338
rect 14660 23276 15320 23287
rect 15396 23186 15424 23310
rect 15488 23254 15516 23684
rect 15844 23666 15896 23672
rect 15660 23656 15712 23662
rect 15580 23604 15660 23610
rect 15580 23598 15712 23604
rect 15580 23582 15700 23598
rect 15476 23248 15528 23254
rect 15476 23190 15528 23196
rect 15384 23180 15436 23186
rect 15384 23122 15436 23128
rect 14648 23112 14700 23118
rect 14568 23072 14648 23100
rect 14648 23054 14700 23060
rect 14464 23044 14516 23050
rect 14464 22986 14516 22992
rect 14476 22574 14504 22986
rect 15292 22772 15344 22778
rect 15212 22732 15292 22760
rect 14832 22636 14884 22642
rect 14832 22578 14884 22584
rect 14464 22568 14516 22574
rect 14464 22510 14516 22516
rect 14844 22488 14872 22578
rect 15016 22500 15068 22506
rect 14844 22460 15016 22488
rect 15016 22442 15068 22448
rect 14648 22432 14700 22438
rect 14648 22374 14700 22380
rect 14372 22092 14424 22098
rect 14660 22094 14688 22374
rect 14846 22332 15154 22352
rect 14846 22330 14852 22332
rect 14908 22330 14932 22332
rect 14988 22330 15012 22332
rect 15068 22330 15092 22332
rect 15148 22330 15154 22332
rect 14908 22278 14910 22330
rect 15090 22278 15092 22330
rect 14846 22276 14852 22278
rect 14908 22276 14932 22278
rect 14988 22276 15012 22278
rect 15068 22276 15092 22278
rect 15148 22276 15154 22278
rect 14846 22256 15154 22276
rect 14740 22228 14792 22234
rect 15212 22216 15240 22732
rect 15292 22714 15344 22720
rect 15488 22710 15516 23190
rect 15476 22704 15528 22710
rect 15476 22646 15528 22652
rect 15580 22506 15608 23582
rect 15856 23254 15884 23666
rect 15844 23248 15896 23254
rect 15844 23190 15896 23196
rect 15752 23180 15804 23186
rect 15672 23140 15752 23168
rect 15568 22500 15620 22506
rect 15568 22442 15620 22448
rect 15672 22438 15700 23140
rect 15752 23122 15804 23128
rect 15844 23112 15896 23118
rect 15844 23054 15896 23060
rect 15750 22672 15806 22681
rect 15750 22607 15752 22616
rect 15804 22607 15806 22616
rect 15752 22578 15804 22584
rect 15856 22438 15884 23054
rect 15384 22432 15436 22438
rect 15290 22400 15346 22409
rect 15384 22374 15436 22380
rect 15660 22432 15712 22438
rect 15660 22374 15712 22380
rect 15844 22432 15896 22438
rect 15844 22374 15896 22380
rect 15290 22335 15346 22344
rect 14792 22188 15240 22216
rect 14740 22170 14792 22176
rect 15304 22148 15332 22335
rect 15028 22120 15332 22148
rect 14660 22066 14964 22094
rect 14372 22034 14424 22040
rect 14384 21593 14412 22034
rect 14464 21956 14516 21962
rect 14464 21898 14516 21904
rect 14370 21584 14426 21593
rect 14370 21519 14426 21528
rect 14372 18760 14424 18766
rect 14372 18702 14424 18708
rect 14384 18630 14412 18702
rect 14372 18624 14424 18630
rect 14372 18566 14424 18572
rect 14476 14890 14504 21898
rect 14660 21814 14872 21842
rect 14660 21418 14688 21814
rect 14738 21720 14794 21729
rect 14738 21655 14794 21664
rect 14752 21434 14780 21655
rect 14844 21604 14872 21814
rect 14936 21729 14964 22066
rect 15028 22030 15056 22120
rect 15016 22024 15068 22030
rect 15396 21978 15424 22374
rect 15474 22264 15530 22273
rect 15474 22199 15530 22208
rect 15660 22228 15712 22234
rect 15488 22001 15516 22199
rect 15660 22170 15712 22176
rect 15016 21966 15068 21972
rect 15120 21950 15424 21978
rect 15474 21992 15530 22001
rect 15016 21888 15068 21894
rect 15016 21830 15068 21836
rect 14922 21720 14978 21729
rect 14922 21655 14978 21664
rect 15028 21604 15056 21830
rect 15120 21622 15148 21950
rect 15474 21927 15530 21936
rect 15384 21888 15436 21894
rect 15304 21848 15384 21876
rect 14844 21576 15056 21604
rect 15108 21616 15160 21622
rect 15108 21558 15160 21564
rect 14752 21418 14964 21434
rect 14648 21412 14700 21418
rect 14752 21412 14976 21418
rect 14752 21406 14924 21412
rect 14648 21354 14700 21360
rect 14924 21354 14976 21360
rect 14556 21344 14608 21350
rect 14556 21286 14608 21292
rect 14568 21010 14596 21286
rect 14556 21004 14608 21010
rect 14556 20946 14608 20952
rect 14660 20874 14688 21354
rect 14740 21344 14792 21350
rect 14740 21286 14792 21292
rect 15200 21344 15252 21350
rect 15200 21286 15252 21292
rect 14648 20868 14700 20874
rect 14648 20810 14700 20816
rect 14556 20800 14608 20806
rect 14556 20742 14608 20748
rect 14568 19258 14596 20742
rect 14648 20392 14700 20398
rect 14648 20334 14700 20340
rect 14660 19854 14688 20334
rect 14752 20330 14780 21286
rect 14846 21244 15154 21264
rect 14846 21242 14852 21244
rect 14908 21242 14932 21244
rect 14988 21242 15012 21244
rect 15068 21242 15092 21244
rect 15148 21242 15154 21244
rect 14908 21190 14910 21242
rect 15090 21190 15092 21242
rect 14846 21188 14852 21190
rect 14908 21188 14932 21190
rect 14988 21188 15012 21190
rect 15068 21188 15092 21190
rect 15148 21188 15154 21190
rect 14846 21168 15154 21188
rect 15212 21010 15240 21286
rect 15200 21004 15252 21010
rect 15200 20946 15252 20952
rect 14830 20904 14886 20913
rect 15304 20874 15332 21848
rect 15384 21830 15436 21836
rect 15568 21888 15620 21894
rect 15568 21830 15620 21836
rect 15384 21616 15436 21622
rect 15384 21558 15436 21564
rect 15396 21049 15424 21558
rect 15476 21480 15528 21486
rect 15476 21422 15528 21428
rect 15488 21146 15516 21422
rect 15476 21140 15528 21146
rect 15476 21082 15528 21088
rect 15382 21040 15438 21049
rect 15382 20975 15438 20984
rect 15396 20874 15424 20975
rect 14830 20839 14886 20848
rect 15292 20868 15344 20874
rect 14844 20806 14872 20839
rect 15292 20810 15344 20816
rect 15384 20868 15436 20874
rect 15384 20810 15436 20816
rect 14832 20800 14884 20806
rect 14832 20742 14884 20748
rect 15384 20596 15436 20602
rect 15384 20538 15436 20544
rect 15200 20528 15252 20534
rect 15200 20470 15252 20476
rect 14740 20324 14792 20330
rect 14740 20266 14792 20272
rect 14752 20058 14780 20266
rect 14846 20156 15154 20176
rect 14846 20154 14852 20156
rect 14908 20154 14932 20156
rect 14988 20154 15012 20156
rect 15068 20154 15092 20156
rect 15148 20154 15154 20156
rect 14908 20102 14910 20154
rect 15090 20102 15092 20154
rect 14846 20100 14852 20102
rect 14908 20100 14932 20102
rect 14988 20100 15012 20102
rect 15068 20100 15092 20102
rect 15148 20100 15154 20102
rect 14846 20080 15154 20100
rect 14740 20052 14792 20058
rect 14740 19994 14792 20000
rect 14648 19848 14700 19854
rect 14648 19790 14700 19796
rect 14752 19378 14780 19994
rect 15106 19952 15162 19961
rect 15106 19887 15162 19896
rect 15120 19854 15148 19887
rect 15108 19848 15160 19854
rect 15108 19790 15160 19796
rect 15106 19680 15162 19689
rect 15106 19615 15162 19624
rect 14740 19372 14792 19378
rect 14740 19314 14792 19320
rect 15120 19310 15148 19615
rect 15108 19304 15160 19310
rect 14568 19242 14688 19258
rect 15108 19246 15160 19252
rect 14568 19236 14700 19242
rect 14568 19230 14648 19236
rect 14648 19178 14700 19184
rect 14556 19168 14608 19174
rect 14556 19110 14608 19116
rect 14568 18086 14596 19110
rect 14846 19068 15154 19088
rect 14846 19066 14852 19068
rect 14908 19066 14932 19068
rect 14988 19066 15012 19068
rect 15068 19066 15092 19068
rect 15148 19066 15154 19068
rect 14908 19014 14910 19066
rect 15090 19014 15092 19066
rect 14846 19012 14852 19014
rect 14908 19012 14932 19014
rect 14988 19012 15012 19014
rect 15068 19012 15092 19014
rect 15148 19012 15154 19014
rect 14846 18992 15154 19012
rect 15212 18970 15240 20470
rect 15292 20256 15344 20262
rect 15292 20198 15344 20204
rect 15200 18964 15252 18970
rect 15200 18906 15252 18912
rect 14740 18828 14792 18834
rect 14740 18770 14792 18776
rect 14556 18080 14608 18086
rect 14556 18022 14608 18028
rect 14568 17678 14596 18022
rect 14752 17746 14780 18770
rect 15212 18358 15240 18906
rect 15200 18352 15252 18358
rect 15200 18294 15252 18300
rect 14846 17980 15154 18000
rect 14846 17978 14852 17980
rect 14908 17978 14932 17980
rect 14988 17978 15012 17980
rect 15068 17978 15092 17980
rect 15148 17978 15154 17980
rect 14908 17926 14910 17978
rect 15090 17926 15092 17978
rect 14846 17924 14852 17926
rect 14908 17924 14932 17926
rect 14988 17924 15012 17926
rect 15068 17924 15092 17926
rect 15148 17924 15154 17926
rect 14846 17904 15154 17924
rect 15212 17746 15240 18294
rect 15304 18290 15332 20198
rect 15396 19938 15424 20538
rect 15476 20052 15528 20058
rect 15580 20040 15608 21830
rect 15672 21146 15700 22170
rect 15844 22092 15896 22098
rect 15844 22034 15896 22040
rect 15752 22024 15804 22030
rect 15752 21966 15804 21972
rect 15660 21140 15712 21146
rect 15660 21082 15712 21088
rect 15764 21049 15792 21966
rect 15856 21146 15884 22034
rect 15948 21622 15976 24092
rect 16028 24074 16080 24080
rect 16120 24132 16172 24138
rect 16120 24074 16172 24080
rect 16028 23860 16080 23866
rect 16028 23802 16080 23808
rect 16040 22982 16068 23802
rect 16132 23254 16160 24074
rect 16120 23248 16172 23254
rect 16120 23190 16172 23196
rect 16120 23044 16172 23050
rect 16120 22986 16172 22992
rect 16212 23044 16264 23050
rect 16212 22986 16264 22992
rect 16028 22976 16080 22982
rect 16028 22918 16080 22924
rect 16132 22574 16160 22986
rect 16028 22568 16080 22574
rect 16028 22510 16080 22516
rect 16120 22568 16172 22574
rect 16120 22510 16172 22516
rect 16040 22001 16068 22510
rect 16026 21992 16082 22001
rect 16026 21927 16082 21936
rect 16120 21888 16172 21894
rect 16120 21830 16172 21836
rect 16132 21729 16160 21830
rect 16118 21720 16174 21729
rect 16028 21684 16080 21690
rect 16118 21655 16174 21664
rect 16028 21626 16080 21632
rect 15936 21616 15988 21622
rect 15936 21558 15988 21564
rect 15844 21140 15896 21146
rect 15844 21082 15896 21088
rect 15750 21040 15806 21049
rect 15750 20975 15806 20984
rect 15660 20868 15712 20874
rect 15660 20810 15712 20816
rect 15528 20012 15608 20040
rect 15476 19994 15528 20000
rect 15396 19910 15516 19938
rect 15488 19854 15516 19910
rect 15476 19848 15528 19854
rect 15476 19790 15528 19796
rect 15384 19780 15436 19786
rect 15384 19722 15436 19728
rect 15396 18630 15424 19722
rect 15568 19712 15620 19718
rect 15568 19654 15620 19660
rect 15580 19310 15608 19654
rect 15568 19304 15620 19310
rect 15568 19246 15620 19252
rect 15672 19242 15700 20810
rect 15752 20460 15804 20466
rect 15752 20402 15804 20408
rect 15764 20058 15792 20402
rect 15752 20052 15804 20058
rect 15752 19994 15804 20000
rect 15948 19378 15976 21558
rect 16040 21321 16068 21626
rect 16120 21548 16172 21554
rect 16120 21490 16172 21496
rect 16026 21312 16082 21321
rect 16026 21247 16082 21256
rect 16132 21078 16160 21490
rect 16120 21072 16172 21078
rect 16120 21014 16172 21020
rect 16028 21004 16080 21010
rect 16028 20946 16080 20952
rect 16040 20534 16068 20946
rect 16028 20528 16080 20534
rect 16028 20470 16080 20476
rect 16132 20466 16160 21014
rect 16224 21010 16252 22986
rect 16316 22692 16344 28494
rect 16408 27614 16436 34954
rect 16500 34785 16528 35391
rect 16672 35216 16724 35222
rect 16776 35193 16804 35770
rect 16672 35158 16724 35164
rect 16762 35184 16818 35193
rect 16486 34776 16542 34785
rect 16486 34711 16542 34720
rect 16684 34610 16712 35158
rect 16762 35119 16818 35128
rect 16488 34604 16540 34610
rect 16488 34546 16540 34552
rect 16672 34604 16724 34610
rect 16672 34546 16724 34552
rect 16500 34202 16528 34546
rect 16580 34536 16632 34542
rect 16580 34478 16632 34484
rect 16592 34202 16620 34478
rect 16488 34196 16540 34202
rect 16488 34138 16540 34144
rect 16580 34196 16632 34202
rect 16580 34138 16632 34144
rect 16592 32434 16620 34138
rect 16580 32428 16632 32434
rect 16580 32370 16632 32376
rect 16486 31920 16542 31929
rect 16486 31855 16542 31864
rect 16500 31754 16528 31855
rect 16488 31748 16540 31754
rect 16488 31690 16540 31696
rect 16592 31414 16620 32370
rect 16868 31754 16896 38950
rect 17500 38956 17552 38962
rect 17500 38898 17552 38904
rect 17604 38758 17632 39374
rect 17868 39364 17920 39370
rect 17868 39306 17920 39312
rect 17684 39296 17736 39302
rect 17684 39238 17736 39244
rect 17696 39030 17724 39238
rect 17684 39024 17736 39030
rect 17684 38966 17736 38972
rect 17592 38752 17644 38758
rect 17880 38740 17908 39306
rect 18604 39296 18656 39302
rect 18418 39264 18474 39273
rect 18604 39238 18656 39244
rect 18418 39199 18474 39208
rect 18432 39098 18460 39199
rect 18420 39092 18472 39098
rect 18420 39034 18472 39040
rect 18328 39024 18380 39030
rect 18328 38966 18380 38972
rect 18340 38826 18368 38966
rect 18328 38820 18380 38826
rect 18328 38762 18380 38768
rect 18420 38752 18472 38758
rect 17880 38712 18000 38740
rect 17592 38694 17644 38700
rect 17868 38412 17920 38418
rect 17868 38354 17920 38360
rect 17130 38040 17186 38049
rect 17130 37975 17186 37984
rect 16948 37256 17000 37262
rect 16948 37198 17000 37204
rect 16960 37097 16988 37198
rect 16946 37088 17002 37097
rect 16946 37023 17002 37032
rect 17040 36712 17092 36718
rect 17040 36654 17092 36660
rect 16946 36000 17002 36009
rect 16946 35935 17002 35944
rect 16960 33998 16988 35935
rect 17052 35737 17080 36654
rect 17144 36417 17172 37975
rect 17316 37868 17368 37874
rect 17316 37810 17368 37816
rect 17328 37466 17356 37810
rect 17880 37466 17908 38354
rect 17316 37460 17368 37466
rect 17316 37402 17368 37408
rect 17868 37460 17920 37466
rect 17868 37402 17920 37408
rect 17880 37369 17908 37402
rect 17866 37360 17922 37369
rect 17866 37295 17922 37304
rect 17972 37126 18000 38712
rect 18156 38700 18420 38706
rect 18156 38694 18472 38700
rect 18156 38678 18460 38694
rect 18052 37664 18104 37670
rect 18052 37606 18104 37612
rect 18064 37330 18092 37606
rect 18052 37324 18104 37330
rect 18052 37266 18104 37272
rect 18156 37262 18184 38678
rect 18420 38548 18472 38554
rect 18420 38490 18472 38496
rect 18236 38208 18288 38214
rect 18236 38150 18288 38156
rect 18328 38208 18380 38214
rect 18328 38150 18380 38156
rect 18248 37448 18276 38150
rect 18340 38010 18368 38150
rect 18328 38004 18380 38010
rect 18328 37946 18380 37952
rect 18432 37738 18460 38490
rect 18420 37732 18472 37738
rect 18420 37674 18472 37680
rect 18328 37460 18380 37466
rect 18248 37420 18328 37448
rect 18328 37402 18380 37408
rect 18144 37256 18196 37262
rect 18144 37198 18196 37204
rect 18328 37256 18380 37262
rect 18328 37198 18380 37204
rect 17960 37120 18012 37126
rect 17960 37062 18012 37068
rect 18144 36916 18196 36922
rect 18144 36858 18196 36864
rect 18052 36780 18104 36786
rect 18052 36722 18104 36728
rect 17130 36408 17186 36417
rect 17130 36343 17186 36352
rect 17868 36372 17920 36378
rect 17038 35728 17094 35737
rect 17038 35663 17094 35672
rect 17040 35216 17092 35222
rect 17040 35158 17092 35164
rect 16948 33992 17000 33998
rect 16948 33934 17000 33940
rect 16948 32428 17000 32434
rect 17052 32416 17080 35158
rect 17144 35154 17172 36343
rect 17868 36314 17920 36320
rect 17590 36272 17646 36281
rect 17590 36207 17646 36216
rect 17774 36272 17830 36281
rect 17774 36207 17830 36216
rect 17224 36100 17276 36106
rect 17224 36042 17276 36048
rect 17236 35766 17264 36042
rect 17604 36009 17632 36207
rect 17788 36038 17816 36207
rect 17776 36032 17828 36038
rect 17590 36000 17646 36009
rect 17776 35974 17828 35980
rect 17590 35935 17646 35944
rect 17224 35760 17276 35766
rect 17224 35702 17276 35708
rect 17684 35692 17736 35698
rect 17684 35634 17736 35640
rect 17224 35556 17276 35562
rect 17224 35498 17276 35504
rect 17132 35148 17184 35154
rect 17132 35090 17184 35096
rect 17144 33930 17172 35090
rect 17236 34762 17264 35498
rect 17498 35456 17554 35465
rect 17498 35391 17554 35400
rect 17316 35080 17368 35086
rect 17316 35022 17368 35028
rect 17328 34921 17356 35022
rect 17314 34912 17370 34921
rect 17314 34847 17370 34856
rect 17236 34734 17356 34762
rect 17224 34468 17276 34474
rect 17224 34410 17276 34416
rect 17236 34134 17264 34410
rect 17224 34128 17276 34134
rect 17224 34070 17276 34076
rect 17132 33924 17184 33930
rect 17132 33866 17184 33872
rect 17328 33289 17356 34734
rect 17512 34610 17540 35391
rect 17590 35184 17646 35193
rect 17590 35119 17646 35128
rect 17500 34604 17552 34610
rect 17500 34546 17552 34552
rect 17500 34196 17552 34202
rect 17500 34138 17552 34144
rect 17314 33280 17370 33289
rect 17314 33215 17370 33224
rect 17512 32910 17540 34138
rect 17500 32904 17552 32910
rect 17420 32864 17500 32892
rect 17132 32768 17184 32774
rect 17132 32710 17184 32716
rect 17144 32434 17172 32710
rect 17314 32600 17370 32609
rect 17314 32535 17370 32544
rect 17224 32496 17276 32502
rect 17224 32438 17276 32444
rect 17000 32388 17080 32416
rect 17132 32428 17184 32434
rect 16948 32370 17000 32376
rect 17132 32370 17184 32376
rect 16684 31726 16896 31754
rect 16580 31408 16632 31414
rect 16486 31376 16542 31385
rect 16580 31350 16632 31356
rect 16486 31311 16488 31320
rect 16540 31311 16542 31320
rect 16488 31282 16540 31288
rect 16488 28416 16540 28422
rect 16488 28358 16540 28364
rect 16500 27946 16528 28358
rect 16488 27940 16540 27946
rect 16488 27882 16540 27888
rect 16408 27586 16620 27614
rect 16592 26353 16620 27586
rect 16394 26344 16450 26353
rect 16394 26279 16450 26288
rect 16578 26344 16634 26353
rect 16578 26279 16634 26288
rect 16408 25906 16436 26279
rect 16578 26072 16634 26081
rect 16578 26007 16580 26016
rect 16632 26007 16634 26016
rect 16580 25978 16632 25984
rect 16396 25900 16448 25906
rect 16396 25842 16448 25848
rect 16408 25362 16436 25842
rect 16396 25356 16448 25362
rect 16396 25298 16448 25304
rect 16408 24410 16436 25298
rect 16488 24608 16540 24614
rect 16488 24550 16540 24556
rect 16396 24404 16448 24410
rect 16396 24346 16448 24352
rect 16316 22664 16436 22692
rect 16304 22228 16356 22234
rect 16304 22170 16356 22176
rect 16316 21894 16344 22170
rect 16304 21888 16356 21894
rect 16304 21830 16356 21836
rect 16304 21344 16356 21350
rect 16304 21286 16356 21292
rect 16212 21004 16264 21010
rect 16212 20946 16264 20952
rect 16316 20874 16344 21286
rect 16304 20868 16356 20874
rect 16304 20810 16356 20816
rect 16212 20800 16264 20806
rect 16212 20742 16264 20748
rect 16120 20460 16172 20466
rect 16120 20402 16172 20408
rect 16028 19916 16080 19922
rect 16028 19858 16080 19864
rect 15936 19372 15988 19378
rect 15936 19314 15988 19320
rect 15660 19236 15712 19242
rect 15660 19178 15712 19184
rect 15568 19168 15620 19174
rect 15568 19110 15620 19116
rect 15580 18902 15608 19110
rect 15568 18896 15620 18902
rect 15568 18838 15620 18844
rect 15384 18624 15436 18630
rect 15384 18566 15436 18572
rect 15292 18284 15344 18290
rect 15292 18226 15344 18232
rect 15396 18154 15424 18566
rect 15384 18148 15436 18154
rect 15384 18090 15436 18096
rect 15672 17814 15700 19178
rect 16040 19174 16068 19858
rect 16224 19854 16252 20742
rect 16304 20460 16356 20466
rect 16304 20402 16356 20408
rect 16316 19922 16344 20402
rect 16304 19916 16356 19922
rect 16304 19858 16356 19864
rect 16212 19848 16264 19854
rect 16212 19790 16264 19796
rect 16120 19712 16172 19718
rect 16120 19654 16172 19660
rect 16028 19168 16080 19174
rect 16028 19110 16080 19116
rect 16132 18834 16160 19654
rect 16316 18970 16344 19858
rect 16304 18964 16356 18970
rect 16304 18906 16356 18912
rect 16120 18828 16172 18834
rect 16120 18770 16172 18776
rect 15660 17808 15712 17814
rect 15660 17750 15712 17756
rect 14740 17740 14792 17746
rect 14740 17682 14792 17688
rect 15200 17740 15252 17746
rect 15200 17682 15252 17688
rect 15844 17740 15896 17746
rect 15844 17682 15896 17688
rect 14556 17672 14608 17678
rect 14556 17614 14608 17620
rect 15660 17604 15712 17610
rect 15660 17546 15712 17552
rect 15672 17338 15700 17546
rect 15660 17332 15712 17338
rect 15660 17274 15712 17280
rect 15856 17184 15884 17682
rect 16028 17264 16080 17270
rect 16028 17206 16080 17212
rect 15936 17196 15988 17202
rect 15856 17156 15936 17184
rect 14846 16892 15154 16912
rect 14846 16890 14852 16892
rect 14908 16890 14932 16892
rect 14988 16890 15012 16892
rect 15068 16890 15092 16892
rect 15148 16890 15154 16892
rect 14908 16838 14910 16890
rect 15090 16838 15092 16890
rect 14846 16836 14852 16838
rect 14908 16836 14932 16838
rect 14988 16836 15012 16838
rect 15068 16836 15092 16838
rect 15148 16836 15154 16838
rect 14846 16816 15154 16836
rect 15856 16658 15884 17156
rect 15936 17138 15988 17144
rect 15844 16652 15896 16658
rect 15844 16594 15896 16600
rect 16040 16590 16068 17206
rect 16028 16584 16080 16590
rect 16028 16526 16080 16532
rect 14846 15804 15154 15824
rect 14846 15802 14852 15804
rect 14908 15802 14932 15804
rect 14988 15802 15012 15804
rect 15068 15802 15092 15804
rect 15148 15802 15154 15804
rect 14908 15750 14910 15802
rect 15090 15750 15092 15802
rect 14846 15748 14852 15750
rect 14908 15748 14932 15750
rect 14988 15748 15012 15750
rect 15068 15748 15092 15750
rect 15148 15748 15154 15750
rect 14846 15728 15154 15748
rect 14464 14884 14516 14890
rect 14464 14826 14516 14832
rect 14846 14716 15154 14736
rect 14846 14714 14852 14716
rect 14908 14714 14932 14716
rect 14988 14714 15012 14716
rect 15068 14714 15092 14716
rect 15148 14714 15154 14716
rect 14908 14662 14910 14714
rect 15090 14662 15092 14714
rect 14846 14660 14852 14662
rect 14908 14660 14932 14662
rect 14988 14660 15012 14662
rect 15068 14660 15092 14662
rect 15148 14660 15154 14662
rect 14846 14640 15154 14660
rect 14846 13628 15154 13648
rect 14846 13626 14852 13628
rect 14908 13626 14932 13628
rect 14988 13626 15012 13628
rect 15068 13626 15092 13628
rect 15148 13626 15154 13628
rect 14908 13574 14910 13626
rect 15090 13574 15092 13626
rect 14846 13572 14852 13574
rect 14908 13572 14932 13574
rect 14988 13572 15012 13574
rect 15068 13572 15092 13574
rect 15148 13572 15154 13574
rect 14846 13552 15154 13572
rect 14846 12540 15154 12560
rect 14846 12538 14852 12540
rect 14908 12538 14932 12540
rect 14988 12538 15012 12540
rect 15068 12538 15092 12540
rect 15148 12538 15154 12540
rect 14908 12486 14910 12538
rect 15090 12486 15092 12538
rect 14846 12484 14852 12486
rect 14908 12484 14932 12486
rect 14988 12484 15012 12486
rect 15068 12484 15092 12486
rect 15148 12484 15154 12486
rect 14846 12464 15154 12484
rect 16408 12434 16436 22664
rect 16500 22273 16528 24550
rect 16684 22642 16712 31726
rect 16764 31680 16816 31686
rect 16960 31668 16988 32370
rect 17040 32224 17092 32230
rect 17040 32166 17092 32172
rect 16764 31622 16816 31628
rect 16868 31640 16988 31668
rect 16776 31278 16804 31622
rect 16764 31272 16816 31278
rect 16764 31214 16816 31220
rect 16868 31142 16896 31640
rect 16856 31136 16908 31142
rect 16856 31078 16908 31084
rect 16948 31136 17000 31142
rect 16948 31078 17000 31084
rect 16960 30870 16988 31078
rect 16948 30864 17000 30870
rect 16948 30806 17000 30812
rect 17052 30734 17080 32166
rect 17236 31686 17264 32438
rect 17328 31890 17356 32535
rect 17316 31884 17368 31890
rect 17316 31826 17368 31832
rect 17420 31754 17448 32864
rect 17500 32846 17552 32852
rect 17500 32496 17552 32502
rect 17498 32464 17500 32473
rect 17552 32464 17554 32473
rect 17498 32399 17554 32408
rect 17500 31816 17552 31822
rect 17500 31758 17552 31764
rect 17408 31748 17460 31754
rect 17408 31690 17460 31696
rect 17224 31680 17276 31686
rect 17512 31657 17540 31758
rect 17224 31622 17276 31628
rect 17498 31648 17554 31657
rect 17498 31583 17554 31592
rect 17132 31340 17184 31346
rect 17132 31282 17184 31288
rect 17040 30728 17092 30734
rect 17040 30670 17092 30676
rect 16856 30592 16908 30598
rect 16856 30534 16908 30540
rect 16948 30592 17000 30598
rect 16948 30534 17000 30540
rect 16868 30326 16896 30534
rect 16960 30433 16988 30534
rect 16946 30424 17002 30433
rect 16946 30359 17002 30368
rect 16856 30320 16908 30326
rect 16762 30288 16818 30297
rect 16856 30262 16908 30268
rect 16762 30223 16818 30232
rect 16776 29170 16804 30223
rect 16856 30184 16908 30190
rect 16856 30126 16908 30132
rect 17040 30184 17092 30190
rect 17144 30161 17172 31282
rect 17604 30954 17632 35119
rect 17696 31362 17724 35634
rect 17880 35494 17908 36314
rect 18064 35834 18092 36722
rect 18052 35828 18104 35834
rect 18052 35770 18104 35776
rect 18156 35698 18184 36858
rect 18340 36038 18368 37198
rect 18512 36644 18564 36650
rect 18512 36586 18564 36592
rect 18524 36242 18552 36586
rect 18512 36236 18564 36242
rect 18512 36178 18564 36184
rect 18328 36032 18380 36038
rect 18234 36000 18290 36009
rect 18328 35974 18380 35980
rect 18418 36000 18474 36009
rect 18234 35935 18290 35944
rect 18418 35935 18474 35944
rect 18144 35692 18196 35698
rect 18144 35634 18196 35640
rect 18248 35601 18276 35935
rect 18432 35850 18460 35935
rect 18340 35834 18460 35850
rect 18328 35828 18460 35834
rect 18380 35822 18460 35828
rect 18328 35770 18380 35776
rect 18420 35760 18472 35766
rect 18616 35748 18644 39238
rect 18892 39030 18920 40054
rect 18972 39364 19024 39370
rect 18972 39306 19024 39312
rect 18880 39024 18932 39030
rect 18880 38966 18932 38972
rect 18696 38412 18748 38418
rect 18696 38354 18748 38360
rect 18708 37262 18736 38354
rect 18696 37256 18748 37262
rect 18696 37198 18748 37204
rect 18708 36106 18736 37198
rect 18878 36952 18934 36961
rect 18878 36887 18934 36896
rect 18786 36680 18842 36689
rect 18786 36615 18842 36624
rect 18696 36100 18748 36106
rect 18696 36042 18748 36048
rect 18800 35894 18828 36615
rect 18892 36310 18920 36887
rect 18880 36304 18932 36310
rect 18880 36246 18932 36252
rect 18800 35866 18920 35894
rect 18892 35834 18920 35866
rect 18880 35828 18932 35834
rect 18880 35770 18932 35776
rect 18696 35760 18748 35766
rect 18616 35720 18696 35748
rect 18420 35702 18472 35708
rect 18696 35702 18748 35708
rect 18432 35612 18460 35702
rect 18234 35592 18290 35601
rect 18432 35584 18644 35612
rect 18234 35527 18290 35536
rect 17868 35488 17920 35494
rect 17868 35430 17920 35436
rect 18248 35222 18276 35527
rect 18420 35284 18472 35290
rect 18420 35226 18472 35232
rect 17960 35216 18012 35222
rect 17774 35184 17830 35193
rect 17960 35158 18012 35164
rect 18236 35216 18288 35222
rect 18236 35158 18288 35164
rect 17774 35119 17830 35128
rect 17788 34610 17816 35119
rect 17868 34944 17920 34950
rect 17868 34886 17920 34892
rect 17776 34604 17828 34610
rect 17776 34546 17828 34552
rect 17880 34241 17908 34886
rect 17972 34746 18000 35158
rect 18328 35148 18380 35154
rect 18328 35090 18380 35096
rect 18144 35080 18196 35086
rect 18144 35022 18196 35028
rect 17960 34740 18012 34746
rect 17960 34682 18012 34688
rect 18050 34504 18106 34513
rect 18050 34439 18106 34448
rect 18156 34490 18184 35022
rect 18340 34610 18368 35090
rect 18432 34921 18460 35226
rect 18616 35222 18644 35584
rect 18604 35216 18656 35222
rect 18604 35158 18656 35164
rect 18984 35086 19012 39306
rect 19076 38894 19104 40287
rect 19996 39506 20024 41200
rect 20352 40656 20404 40662
rect 20352 40598 20404 40604
rect 20074 39672 20130 39681
rect 20074 39607 20130 39616
rect 19984 39500 20036 39506
rect 19984 39442 20036 39448
rect 19340 39432 19392 39438
rect 20088 39409 20116 39607
rect 20168 39568 20220 39574
rect 20168 39510 20220 39516
rect 19340 39374 19392 39380
rect 20074 39400 20130 39409
rect 19352 39137 19380 39374
rect 20074 39335 20130 39344
rect 19892 39296 19944 39302
rect 19892 39238 19944 39244
rect 19478 39196 19786 39216
rect 19478 39194 19484 39196
rect 19540 39194 19564 39196
rect 19620 39194 19644 39196
rect 19700 39194 19724 39196
rect 19780 39194 19786 39196
rect 19540 39142 19542 39194
rect 19722 39142 19724 39194
rect 19478 39140 19484 39142
rect 19540 39140 19564 39142
rect 19620 39140 19644 39142
rect 19700 39140 19724 39142
rect 19780 39140 19786 39142
rect 19338 39128 19394 39137
rect 19478 39120 19786 39140
rect 19338 39063 19394 39072
rect 19064 38888 19116 38894
rect 19064 38830 19116 38836
rect 19800 38888 19852 38894
rect 19904 38876 19932 39238
rect 20076 39024 20128 39030
rect 20076 38966 20128 38972
rect 19852 38848 19932 38876
rect 19800 38830 19852 38836
rect 19892 38752 19944 38758
rect 19892 38694 19944 38700
rect 19982 38720 20038 38729
rect 19168 38542 19380 38570
rect 19062 38176 19118 38185
rect 19062 38111 19118 38120
rect 19076 37874 19104 38111
rect 19064 37868 19116 37874
rect 19064 37810 19116 37816
rect 19168 37754 19196 38542
rect 19076 37726 19196 37754
rect 19076 37505 19104 37726
rect 19156 37664 19208 37670
rect 19156 37606 19208 37612
rect 19062 37496 19118 37505
rect 19062 37431 19118 37440
rect 19168 37126 19196 37606
rect 19352 37210 19380 38542
rect 19478 38108 19786 38128
rect 19478 38106 19484 38108
rect 19540 38106 19564 38108
rect 19620 38106 19644 38108
rect 19700 38106 19724 38108
rect 19780 38106 19786 38108
rect 19540 38054 19542 38106
rect 19722 38054 19724 38106
rect 19478 38052 19484 38054
rect 19540 38052 19564 38054
rect 19620 38052 19644 38054
rect 19700 38052 19724 38054
rect 19780 38052 19786 38054
rect 19478 38032 19786 38052
rect 19904 38010 19932 38694
rect 19982 38655 20038 38664
rect 19892 38004 19944 38010
rect 19892 37946 19944 37952
rect 19614 37768 19670 37777
rect 19614 37703 19616 37712
rect 19668 37703 19670 37712
rect 19616 37674 19668 37680
rect 19614 37224 19670 37233
rect 19352 37182 19614 37210
rect 19614 37159 19616 37168
rect 19668 37159 19670 37168
rect 19616 37130 19668 37136
rect 19156 37120 19208 37126
rect 19156 37062 19208 37068
rect 19064 36780 19116 36786
rect 19064 36722 19116 36728
rect 19076 36689 19104 36722
rect 19168 36718 19196 37062
rect 19478 37020 19786 37040
rect 19478 37018 19484 37020
rect 19540 37018 19564 37020
rect 19620 37018 19644 37020
rect 19700 37018 19724 37020
rect 19780 37018 19786 37020
rect 19540 36966 19542 37018
rect 19722 36966 19724 37018
rect 19478 36964 19484 36966
rect 19540 36964 19564 36966
rect 19620 36964 19644 36966
rect 19700 36964 19724 36966
rect 19780 36964 19786 36966
rect 19338 36952 19394 36961
rect 19478 36944 19786 36964
rect 19338 36887 19394 36896
rect 19156 36712 19208 36718
rect 19062 36680 19118 36689
rect 19156 36654 19208 36660
rect 19246 36680 19302 36689
rect 19062 36615 19118 36624
rect 19168 36360 19196 36654
rect 19246 36615 19248 36624
rect 19300 36615 19302 36624
rect 19248 36586 19300 36592
rect 19352 36530 19380 36887
rect 19352 36502 19656 36530
rect 19076 36332 19196 36360
rect 19524 36372 19576 36378
rect 19076 35766 19104 36332
rect 19524 36314 19576 36320
rect 19536 36242 19564 36314
rect 19628 36242 19656 36502
rect 19524 36236 19576 36242
rect 19524 36178 19576 36184
rect 19616 36236 19668 36242
rect 19616 36178 19668 36184
rect 19154 36136 19210 36145
rect 19904 36106 19932 37946
rect 19996 37806 20024 38655
rect 19984 37800 20036 37806
rect 19984 37742 20036 37748
rect 19154 36071 19210 36080
rect 19340 36100 19392 36106
rect 19064 35760 19116 35766
rect 19064 35702 19116 35708
rect 19168 35442 19196 36071
rect 19340 36042 19392 36048
rect 19892 36100 19944 36106
rect 19892 36042 19944 36048
rect 19984 36100 20036 36106
rect 19984 36042 20036 36048
rect 19352 36009 19380 36042
rect 19338 36000 19394 36009
rect 19890 36000 19946 36009
rect 19338 35935 19394 35944
rect 19478 35932 19786 35952
rect 19890 35935 19946 35944
rect 19478 35930 19484 35932
rect 19540 35930 19564 35932
rect 19620 35930 19644 35932
rect 19700 35930 19724 35932
rect 19780 35930 19786 35932
rect 19540 35878 19542 35930
rect 19722 35878 19724 35930
rect 19478 35876 19484 35878
rect 19540 35876 19564 35878
rect 19620 35876 19644 35878
rect 19700 35876 19724 35878
rect 19780 35876 19786 35878
rect 19338 35864 19394 35873
rect 19478 35856 19786 35876
rect 19338 35799 19394 35808
rect 19248 35760 19300 35766
rect 19248 35702 19300 35708
rect 19076 35414 19196 35442
rect 18972 35080 19024 35086
rect 18972 35022 19024 35028
rect 18418 34912 18474 34921
rect 18418 34847 18474 34856
rect 18786 34776 18842 34785
rect 18786 34711 18842 34720
rect 18696 34672 18748 34678
rect 18616 34632 18696 34660
rect 18328 34604 18380 34610
rect 18328 34546 18380 34552
rect 18234 34504 18290 34513
rect 18156 34462 18234 34490
rect 17866 34232 17922 34241
rect 17866 34167 17922 34176
rect 18064 34134 18092 34439
rect 18052 34128 18104 34134
rect 18052 34070 18104 34076
rect 18064 33590 18092 34070
rect 18156 33862 18184 34462
rect 18234 34439 18290 34448
rect 18340 34066 18368 34546
rect 18512 34400 18564 34406
rect 18512 34342 18564 34348
rect 18328 34060 18380 34066
rect 18328 34002 18380 34008
rect 18236 33924 18288 33930
rect 18236 33866 18288 33872
rect 18144 33856 18196 33862
rect 18144 33798 18196 33804
rect 18052 33584 18104 33590
rect 18052 33526 18104 33532
rect 18050 33144 18106 33153
rect 18248 33114 18276 33866
rect 18050 33079 18052 33088
rect 18104 33079 18106 33088
rect 18236 33108 18288 33114
rect 18052 33050 18104 33056
rect 18236 33050 18288 33056
rect 17696 31334 17816 31362
rect 17684 31272 17736 31278
rect 17684 31214 17736 31220
rect 17224 30932 17276 30938
rect 17224 30874 17276 30880
rect 17328 30926 17632 30954
rect 17236 30734 17264 30874
rect 17224 30728 17276 30734
rect 17224 30670 17276 30676
rect 17040 30126 17092 30132
rect 17130 30152 17186 30161
rect 16868 29345 16896 30126
rect 16948 30116 17000 30122
rect 16948 30058 17000 30064
rect 16960 29889 16988 30058
rect 16946 29880 17002 29889
rect 16946 29815 17002 29824
rect 16854 29336 16910 29345
rect 16854 29271 16910 29280
rect 16764 29164 16816 29170
rect 16764 29106 16816 29112
rect 17052 29102 17080 30126
rect 17130 30087 17186 30096
rect 17328 30036 17356 30926
rect 17408 30864 17460 30870
rect 17408 30806 17460 30812
rect 17144 30008 17356 30036
rect 16856 29096 16908 29102
rect 16856 29038 16908 29044
rect 17040 29096 17092 29102
rect 17040 29038 17092 29044
rect 16762 28656 16818 28665
rect 16762 28591 16818 28600
rect 16776 26926 16804 28591
rect 16868 28121 16896 29038
rect 16948 28960 17000 28966
rect 16948 28902 17000 28908
rect 16960 28665 16988 28902
rect 16946 28656 17002 28665
rect 16946 28591 17002 28600
rect 16854 28112 16910 28121
rect 16854 28047 16910 28056
rect 16868 27713 16896 28047
rect 17052 28014 17080 29038
rect 17144 28966 17172 30008
rect 17224 29028 17276 29034
rect 17224 28970 17276 28976
rect 17132 28960 17184 28966
rect 17132 28902 17184 28908
rect 17144 28626 17172 28902
rect 17132 28620 17184 28626
rect 17132 28562 17184 28568
rect 17236 28558 17264 28970
rect 17224 28552 17276 28558
rect 17276 28512 17356 28540
rect 17224 28494 17276 28500
rect 17132 28484 17184 28490
rect 17132 28426 17184 28432
rect 17144 28257 17172 28426
rect 17130 28248 17186 28257
rect 17130 28183 17186 28192
rect 17224 28076 17276 28082
rect 17224 28018 17276 28024
rect 17040 28008 17092 28014
rect 17040 27950 17092 27956
rect 16854 27704 16910 27713
rect 17052 27674 17080 27950
rect 16854 27639 16910 27648
rect 17040 27668 17092 27674
rect 17040 27610 17092 27616
rect 16856 27396 16908 27402
rect 16856 27338 16908 27344
rect 16868 27062 16896 27338
rect 16856 27056 16908 27062
rect 16856 26998 16908 27004
rect 16948 26988 17000 26994
rect 16948 26930 17000 26936
rect 16764 26920 16816 26926
rect 16764 26862 16816 26868
rect 16960 26625 16988 26930
rect 16946 26616 17002 26625
rect 16946 26551 17002 26560
rect 16856 25696 16908 25702
rect 17236 25673 17264 28018
rect 17328 27577 17356 28512
rect 17420 28393 17448 30806
rect 17500 30728 17552 30734
rect 17500 30670 17552 30676
rect 17512 29753 17540 30670
rect 17696 30258 17724 31214
rect 17788 30977 17816 31334
rect 17774 30968 17830 30977
rect 17774 30903 17830 30912
rect 17788 30802 17816 30903
rect 17776 30796 17828 30802
rect 17776 30738 17828 30744
rect 18064 30394 18092 33050
rect 18236 32904 18288 32910
rect 18236 32846 18288 32852
rect 18248 32774 18276 32846
rect 18236 32768 18288 32774
rect 18236 32710 18288 32716
rect 18236 32428 18288 32434
rect 18340 32416 18368 34002
rect 18524 33862 18552 34342
rect 18616 34202 18644 34632
rect 18696 34614 18748 34620
rect 18604 34196 18656 34202
rect 18604 34138 18656 34144
rect 18800 33862 18828 34711
rect 19076 34377 19104 35414
rect 19260 35222 19288 35702
rect 19352 35698 19380 35799
rect 19432 35760 19484 35766
rect 19432 35702 19484 35708
rect 19616 35760 19668 35766
rect 19616 35702 19668 35708
rect 19800 35760 19852 35766
rect 19800 35702 19852 35708
rect 19340 35692 19392 35698
rect 19340 35634 19392 35640
rect 19156 35216 19208 35222
rect 19156 35158 19208 35164
rect 19248 35216 19300 35222
rect 19248 35158 19300 35164
rect 19168 35034 19196 35158
rect 19444 35034 19472 35702
rect 19524 35624 19576 35630
rect 19524 35566 19576 35572
rect 19536 35465 19564 35566
rect 19522 35456 19578 35465
rect 19522 35391 19578 35400
rect 19168 35006 19472 35034
rect 19628 35018 19656 35702
rect 19812 35222 19840 35702
rect 19904 35494 19932 35935
rect 19996 35562 20024 36042
rect 19984 35556 20036 35562
rect 19984 35498 20036 35504
rect 19892 35488 19944 35494
rect 19892 35430 19944 35436
rect 19800 35216 19852 35222
rect 19800 35158 19852 35164
rect 19616 35012 19668 35018
rect 19616 34954 19668 34960
rect 19478 34844 19786 34864
rect 19478 34842 19484 34844
rect 19540 34842 19564 34844
rect 19620 34842 19644 34844
rect 19700 34842 19724 34844
rect 19780 34842 19786 34844
rect 19540 34790 19542 34842
rect 19722 34790 19724 34842
rect 19478 34788 19484 34790
rect 19540 34788 19564 34790
rect 19620 34788 19644 34790
rect 19700 34788 19724 34790
rect 19780 34788 19786 34790
rect 19478 34768 19786 34788
rect 19984 34604 20036 34610
rect 19984 34546 20036 34552
rect 19892 34400 19944 34406
rect 19168 34377 19380 34388
rect 19062 34368 19118 34377
rect 19062 34303 19118 34312
rect 19168 34368 19394 34377
rect 19168 34360 19338 34368
rect 18972 33924 19024 33930
rect 18972 33866 19024 33872
rect 18420 33856 18472 33862
rect 18420 33798 18472 33804
rect 18512 33856 18564 33862
rect 18512 33798 18564 33804
rect 18788 33856 18840 33862
rect 18788 33798 18840 33804
rect 18432 33658 18460 33798
rect 18420 33652 18472 33658
rect 18420 33594 18472 33600
rect 18432 33017 18460 33594
rect 18418 33008 18474 33017
rect 18418 32943 18474 32952
rect 18432 32910 18460 32943
rect 18420 32904 18472 32910
rect 18420 32846 18472 32852
rect 18524 32774 18552 33798
rect 18694 33688 18750 33697
rect 18694 33623 18750 33632
rect 18604 33584 18656 33590
rect 18604 33526 18656 33532
rect 18616 33386 18644 33526
rect 18604 33380 18656 33386
rect 18604 33322 18656 33328
rect 18616 32910 18644 33322
rect 18708 33017 18736 33623
rect 18694 33008 18750 33017
rect 18694 32943 18750 32952
rect 18604 32904 18656 32910
rect 18604 32846 18656 32852
rect 18512 32768 18564 32774
rect 18512 32710 18564 32716
rect 18696 32768 18748 32774
rect 18696 32710 18748 32716
rect 18708 32502 18736 32710
rect 18696 32496 18748 32502
rect 18696 32438 18748 32444
rect 18288 32388 18368 32416
rect 18236 32370 18288 32376
rect 18604 32020 18656 32026
rect 18604 31962 18656 31968
rect 18236 31748 18288 31754
rect 18236 31690 18288 31696
rect 18052 30388 18104 30394
rect 18052 30330 18104 30336
rect 17684 30252 17736 30258
rect 17684 30194 17736 30200
rect 17696 29850 17724 30194
rect 17774 30016 17830 30025
rect 17774 29951 17830 29960
rect 17684 29844 17736 29850
rect 17684 29786 17736 29792
rect 17592 29776 17644 29782
rect 17498 29744 17554 29753
rect 17592 29718 17644 29724
rect 17498 29679 17554 29688
rect 17604 28937 17632 29718
rect 17590 28928 17646 28937
rect 17590 28863 17646 28872
rect 17500 28620 17552 28626
rect 17500 28562 17552 28568
rect 17406 28384 17462 28393
rect 17406 28319 17462 28328
rect 17408 27668 17460 27674
rect 17408 27610 17460 27616
rect 17314 27568 17370 27577
rect 17314 27503 17370 27512
rect 17328 26518 17356 27503
rect 17420 27305 17448 27610
rect 17406 27296 17462 27305
rect 17406 27231 17462 27240
rect 17408 26920 17460 26926
rect 17408 26862 17460 26868
rect 17316 26512 17368 26518
rect 17316 26454 17368 26460
rect 16856 25638 16908 25644
rect 17222 25664 17278 25673
rect 16868 24818 16896 25638
rect 17222 25599 17278 25608
rect 17040 25288 17092 25294
rect 17040 25230 17092 25236
rect 16948 25220 17000 25226
rect 16948 25162 17000 25168
rect 16960 25129 16988 25162
rect 16946 25120 17002 25129
rect 16946 25055 17002 25064
rect 16856 24812 16908 24818
rect 16856 24754 16908 24760
rect 16764 24676 16816 24682
rect 16764 24618 16816 24624
rect 16776 24410 16804 24618
rect 17052 24614 17080 25230
rect 17224 25152 17276 25158
rect 17224 25094 17276 25100
rect 17130 24984 17186 24993
rect 17130 24919 17132 24928
rect 17184 24919 17186 24928
rect 17132 24890 17184 24896
rect 17040 24608 17092 24614
rect 17040 24550 17092 24556
rect 16764 24404 16816 24410
rect 16764 24346 16816 24352
rect 17236 24342 17264 25094
rect 17420 24818 17448 26862
rect 17512 26858 17540 28562
rect 17696 28082 17724 29786
rect 17684 28076 17736 28082
rect 17684 28018 17736 28024
rect 17788 27928 17816 29951
rect 17958 29744 18014 29753
rect 17868 29708 17920 29714
rect 18014 29702 18184 29730
rect 17958 29679 18014 29688
rect 17868 29650 17920 29656
rect 17880 29578 17908 29650
rect 17868 29572 17920 29578
rect 17868 29514 17920 29520
rect 17960 29504 18012 29510
rect 17960 29446 18012 29452
rect 17972 29238 18000 29446
rect 17960 29232 18012 29238
rect 17960 29174 18012 29180
rect 18052 29232 18104 29238
rect 18052 29174 18104 29180
rect 18064 29073 18092 29174
rect 18156 29170 18184 29702
rect 18144 29164 18196 29170
rect 18144 29106 18196 29112
rect 18050 29064 18106 29073
rect 18050 28999 18106 29008
rect 17868 28756 17920 28762
rect 17868 28698 17920 28704
rect 17604 27900 17816 27928
rect 17500 26852 17552 26858
rect 17500 26794 17552 26800
rect 17604 26518 17632 27900
rect 17880 27826 17908 28698
rect 18248 28608 18276 31690
rect 18512 31680 18564 31686
rect 18512 31622 18564 31628
rect 18420 30796 18472 30802
rect 18420 30738 18472 30744
rect 18432 30161 18460 30738
rect 18418 30152 18474 30161
rect 18418 30087 18474 30096
rect 18420 30048 18472 30054
rect 18420 29990 18472 29996
rect 18432 29782 18460 29990
rect 18420 29776 18472 29782
rect 18420 29718 18472 29724
rect 18328 29504 18380 29510
rect 18328 29446 18380 29452
rect 18340 28966 18368 29446
rect 18418 29336 18474 29345
rect 18418 29271 18474 29280
rect 18432 29102 18460 29271
rect 18420 29096 18472 29102
rect 18420 29038 18472 29044
rect 18328 28960 18380 28966
rect 18328 28902 18380 28908
rect 18340 28762 18368 28902
rect 18328 28756 18380 28762
rect 18328 28698 18380 28704
rect 18328 28620 18380 28626
rect 18248 28580 18328 28608
rect 18328 28562 18380 28568
rect 18052 28552 18104 28558
rect 18052 28494 18104 28500
rect 18418 28520 18474 28529
rect 17788 27798 17908 27826
rect 17788 26994 17816 27798
rect 18064 27606 18092 28494
rect 18418 28455 18474 28464
rect 18236 28416 18288 28422
rect 18236 28358 18288 28364
rect 18248 28150 18276 28358
rect 18236 28144 18288 28150
rect 18236 28086 18288 28092
rect 18236 28008 18288 28014
rect 18236 27950 18288 27956
rect 17868 27600 17920 27606
rect 17868 27542 17920 27548
rect 18052 27600 18104 27606
rect 18052 27542 18104 27548
rect 18142 27568 18198 27577
rect 17880 27044 17908 27542
rect 18248 27538 18276 27950
rect 18328 27940 18380 27946
rect 18328 27882 18380 27888
rect 18142 27503 18198 27512
rect 18236 27532 18288 27538
rect 18052 27464 18104 27470
rect 18052 27406 18104 27412
rect 17960 27328 18012 27334
rect 17958 27296 17960 27305
rect 18012 27296 18014 27305
rect 17958 27231 18014 27240
rect 17960 27056 18012 27062
rect 17880 27016 17960 27044
rect 17960 26998 18012 27004
rect 17684 26988 17736 26994
rect 17684 26930 17736 26936
rect 17776 26988 17828 26994
rect 17776 26930 17828 26936
rect 17592 26512 17644 26518
rect 17592 26454 17644 26460
rect 17592 26376 17644 26382
rect 17592 26318 17644 26324
rect 17408 24812 17460 24818
rect 17408 24754 17460 24760
rect 17224 24336 17276 24342
rect 17224 24278 17276 24284
rect 16764 23792 16816 23798
rect 16764 23734 16816 23740
rect 16776 23594 16804 23734
rect 16856 23656 16908 23662
rect 16856 23598 16908 23604
rect 16948 23656 17000 23662
rect 16948 23598 17000 23604
rect 16764 23588 16816 23594
rect 16764 23530 16816 23536
rect 16762 22944 16818 22953
rect 16762 22879 16818 22888
rect 16776 22642 16804 22879
rect 16672 22636 16724 22642
rect 16672 22578 16724 22584
rect 16764 22636 16816 22642
rect 16764 22578 16816 22584
rect 16486 22264 16542 22273
rect 16486 22199 16542 22208
rect 16580 22024 16632 22030
rect 16580 21966 16632 21972
rect 16488 21956 16540 21962
rect 16488 21898 16540 21904
rect 16500 21554 16528 21898
rect 16592 21865 16620 21966
rect 16578 21856 16634 21865
rect 16578 21791 16634 21800
rect 16578 21720 16634 21729
rect 16578 21655 16634 21664
rect 16488 21548 16540 21554
rect 16488 21490 16540 21496
rect 16500 19174 16528 21490
rect 16592 21185 16620 21655
rect 16578 21176 16634 21185
rect 16578 21111 16634 21120
rect 16684 21026 16712 22578
rect 16764 22432 16816 22438
rect 16764 22374 16816 22380
rect 16776 22234 16804 22374
rect 16764 22228 16816 22234
rect 16764 22170 16816 22176
rect 16762 21720 16818 21729
rect 16762 21655 16818 21664
rect 16776 21418 16804 21655
rect 16764 21412 16816 21418
rect 16764 21354 16816 21360
rect 16592 20998 16712 21026
rect 16488 19168 16540 19174
rect 16488 19110 16540 19116
rect 16488 17604 16540 17610
rect 16488 17546 16540 17552
rect 16500 17134 16528 17546
rect 16488 17128 16540 17134
rect 16488 17070 16540 17076
rect 16500 16250 16528 17070
rect 16488 16244 16540 16250
rect 16488 16186 16540 16192
rect 16316 12406 16436 12434
rect 14846 11452 15154 11472
rect 14846 11450 14852 11452
rect 14908 11450 14932 11452
rect 14988 11450 15012 11452
rect 15068 11450 15092 11452
rect 15148 11450 15154 11452
rect 14908 11398 14910 11450
rect 15090 11398 15092 11450
rect 14846 11396 14852 11398
rect 14908 11396 14932 11398
rect 14988 11396 15012 11398
rect 15068 11396 15092 11398
rect 15148 11396 15154 11398
rect 14846 11376 15154 11396
rect 14846 10364 15154 10384
rect 14846 10362 14852 10364
rect 14908 10362 14932 10364
rect 14988 10362 15012 10364
rect 15068 10362 15092 10364
rect 15148 10362 15154 10364
rect 14908 10310 14910 10362
rect 15090 10310 15092 10362
rect 14846 10308 14852 10310
rect 14908 10308 14932 10310
rect 14988 10308 15012 10310
rect 15068 10308 15092 10310
rect 15148 10308 15154 10310
rect 14846 10288 15154 10308
rect 14846 9276 15154 9296
rect 14846 9274 14852 9276
rect 14908 9274 14932 9276
rect 14988 9274 15012 9276
rect 15068 9274 15092 9276
rect 15148 9274 15154 9276
rect 14908 9222 14910 9274
rect 15090 9222 15092 9274
rect 14846 9220 14852 9222
rect 14908 9220 14932 9222
rect 14988 9220 15012 9222
rect 15068 9220 15092 9222
rect 15148 9220 15154 9222
rect 14846 9200 15154 9220
rect 14846 8188 15154 8208
rect 14846 8186 14852 8188
rect 14908 8186 14932 8188
rect 14988 8186 15012 8188
rect 15068 8186 15092 8188
rect 15148 8186 15154 8188
rect 14908 8134 14910 8186
rect 15090 8134 15092 8186
rect 14846 8132 14852 8134
rect 14908 8132 14932 8134
rect 14988 8132 15012 8134
rect 15068 8132 15092 8134
rect 15148 8132 15154 8134
rect 14846 8112 15154 8132
rect 14846 7100 15154 7120
rect 14846 7098 14852 7100
rect 14908 7098 14932 7100
rect 14988 7098 15012 7100
rect 15068 7098 15092 7100
rect 15148 7098 15154 7100
rect 14908 7046 14910 7098
rect 15090 7046 15092 7098
rect 14846 7044 14852 7046
rect 14908 7044 14932 7046
rect 14988 7044 15012 7046
rect 15068 7044 15092 7046
rect 15148 7044 15154 7046
rect 14846 7024 15154 7044
rect 14016 6886 14320 6914
rect 14016 6798 14044 6886
rect 14004 6792 14056 6798
rect 14004 6734 14056 6740
rect 14846 6012 15154 6032
rect 14846 6010 14852 6012
rect 14908 6010 14932 6012
rect 14988 6010 15012 6012
rect 15068 6010 15092 6012
rect 15148 6010 15154 6012
rect 14908 5958 14910 6010
rect 15090 5958 15092 6010
rect 14846 5956 14852 5958
rect 14908 5956 14932 5958
rect 14988 5956 15012 5958
rect 15068 5956 15092 5958
rect 15148 5956 15154 5958
rect 14846 5936 15154 5956
rect 14846 4924 15154 4944
rect 14846 4922 14852 4924
rect 14908 4922 14932 4924
rect 14988 4922 15012 4924
rect 15068 4922 15092 4924
rect 15148 4922 15154 4924
rect 14908 4870 14910 4922
rect 15090 4870 15092 4922
rect 14846 4868 14852 4870
rect 14908 4868 14932 4870
rect 14988 4868 15012 4870
rect 15068 4868 15092 4870
rect 15148 4868 15154 4870
rect 14846 4848 15154 4868
rect 13176 4072 13228 4078
rect 13176 4014 13228 4020
rect 13544 4072 13596 4078
rect 13544 4014 13596 4020
rect 13188 3738 13216 4014
rect 13176 3732 13228 3738
rect 13176 3674 13228 3680
rect 12992 3528 13044 3534
rect 12992 3470 13044 3476
rect 12440 2440 12492 2446
rect 12440 2382 12492 2388
rect 13556 800 13584 4014
rect 15660 3936 15712 3942
rect 15660 3878 15712 3884
rect 14846 3836 15154 3856
rect 14846 3834 14852 3836
rect 14908 3834 14932 3836
rect 14988 3834 15012 3836
rect 15068 3834 15092 3836
rect 15148 3834 15154 3836
rect 14908 3782 14910 3834
rect 15090 3782 15092 3834
rect 14846 3780 14852 3782
rect 14908 3780 14932 3782
rect 14988 3780 15012 3782
rect 15068 3780 15092 3782
rect 15148 3780 15154 3782
rect 14846 3760 15154 3780
rect 15672 3602 15700 3878
rect 15660 3596 15712 3602
rect 15660 3538 15712 3544
rect 16120 3596 16172 3602
rect 16120 3538 16172 3544
rect 14188 3528 14240 3534
rect 14188 3470 14240 3476
rect 14096 3392 14148 3398
rect 14096 3334 14148 3340
rect 14108 3126 14136 3334
rect 14096 3120 14148 3126
rect 14096 3062 14148 3068
rect 14108 2446 14136 3062
rect 14200 3058 14228 3470
rect 15660 3460 15712 3466
rect 15660 3402 15712 3408
rect 15844 3460 15896 3466
rect 15844 3402 15896 3408
rect 14188 3052 14240 3058
rect 14188 2994 14240 3000
rect 14372 2984 14424 2990
rect 14372 2926 14424 2932
rect 14740 2984 14792 2990
rect 14740 2926 14792 2932
rect 14384 2650 14412 2926
rect 14372 2644 14424 2650
rect 14372 2586 14424 2592
rect 14096 2440 14148 2446
rect 14096 2382 14148 2388
rect 14752 1578 14780 2926
rect 14846 2748 15154 2768
rect 14846 2746 14852 2748
rect 14908 2746 14932 2748
rect 14988 2746 15012 2748
rect 15068 2746 15092 2748
rect 15148 2746 15154 2748
rect 14908 2694 14910 2746
rect 15090 2694 15092 2746
rect 14846 2692 14852 2694
rect 14908 2692 14932 2694
rect 14988 2692 15012 2694
rect 15068 2692 15092 2694
rect 15148 2692 15154 2694
rect 14846 2672 15154 2692
rect 15672 2446 15700 3402
rect 15856 2650 15884 3402
rect 15844 2644 15896 2650
rect 15844 2586 15896 2592
rect 15660 2440 15712 2446
rect 15660 2382 15712 2388
rect 14752 1550 14872 1578
rect 14844 800 14872 1550
rect 16132 800 16160 3538
rect 16316 2650 16344 12406
rect 16592 6914 16620 20998
rect 16672 20914 16724 20920
rect 16672 20856 16724 20862
rect 16684 20602 16712 20856
rect 16672 20596 16724 20602
rect 16672 20538 16724 20544
rect 16868 20398 16896 23598
rect 16960 23361 16988 23598
rect 16946 23352 17002 23361
rect 16946 23287 17002 23296
rect 16946 23216 17002 23225
rect 17236 23202 17264 24278
rect 17052 23186 17264 23202
rect 16946 23151 17002 23160
rect 17040 23180 17264 23186
rect 16960 23118 16988 23151
rect 17092 23174 17264 23180
rect 17040 23122 17092 23128
rect 16948 23112 17000 23118
rect 16948 23054 17000 23060
rect 17132 23112 17184 23118
rect 17132 23054 17184 23060
rect 17040 23044 17092 23050
rect 17040 22986 17092 22992
rect 16948 22772 17000 22778
rect 16948 22714 17000 22720
rect 16960 22506 16988 22714
rect 17052 22574 17080 22986
rect 17144 22710 17172 23054
rect 17132 22704 17184 22710
rect 17132 22646 17184 22652
rect 17040 22568 17092 22574
rect 17040 22510 17092 22516
rect 16948 22500 17000 22506
rect 16948 22442 17000 22448
rect 16948 21956 17000 21962
rect 17132 21956 17184 21962
rect 16948 21898 17000 21904
rect 17052 21916 17132 21944
rect 16960 21010 16988 21898
rect 16948 21004 17000 21010
rect 16948 20946 17000 20952
rect 16856 20392 16908 20398
rect 16856 20334 16908 20340
rect 16868 19961 16896 20334
rect 16854 19952 16910 19961
rect 16960 19938 16988 20946
rect 17052 20398 17080 21916
rect 17132 21898 17184 21904
rect 17132 20800 17184 20806
rect 17132 20742 17184 20748
rect 17144 20398 17172 20742
rect 17040 20392 17092 20398
rect 17040 20334 17092 20340
rect 17132 20392 17184 20398
rect 17132 20334 17184 20340
rect 17040 20052 17092 20058
rect 17144 20040 17172 20334
rect 17092 20012 17172 20040
rect 17040 19994 17092 20000
rect 16960 19910 17080 19938
rect 16854 19887 16910 19896
rect 16948 19848 17000 19854
rect 16948 19790 17000 19796
rect 16764 19440 16816 19446
rect 16764 19382 16816 19388
rect 16854 19408 16910 19417
rect 16672 18692 16724 18698
rect 16672 18634 16724 18640
rect 16684 17134 16712 18634
rect 16672 17128 16724 17134
rect 16672 17070 16724 17076
rect 16684 16454 16712 17070
rect 16672 16448 16724 16454
rect 16672 16390 16724 16396
rect 16776 16182 16804 19382
rect 16854 19343 16910 19352
rect 16868 19242 16896 19343
rect 16960 19310 16988 19790
rect 17052 19689 17080 19910
rect 17038 19680 17094 19689
rect 17038 19615 17094 19624
rect 17040 19372 17092 19378
rect 17040 19314 17092 19320
rect 16948 19304 17000 19310
rect 16948 19246 17000 19252
rect 16856 19236 16908 19242
rect 16856 19178 16908 19184
rect 16868 18290 16896 19178
rect 16856 18284 16908 18290
rect 16856 18226 16908 18232
rect 16856 17060 16908 17066
rect 16856 17002 16908 17008
rect 16764 16176 16816 16182
rect 16764 16118 16816 16124
rect 16868 15978 16896 17002
rect 16948 16992 17000 16998
rect 16948 16934 17000 16940
rect 16960 16114 16988 16934
rect 17052 16674 17080 19314
rect 17132 18760 17184 18766
rect 17132 18702 17184 18708
rect 17144 17882 17172 18702
rect 17132 17876 17184 17882
rect 17132 17818 17184 17824
rect 17236 16776 17264 23174
rect 17316 23180 17368 23186
rect 17316 23122 17368 23128
rect 17328 21690 17356 23122
rect 17316 21684 17368 21690
rect 17316 21626 17368 21632
rect 17316 21480 17368 21486
rect 17316 21422 17368 21428
rect 17328 21010 17356 21422
rect 17316 21004 17368 21010
rect 17316 20946 17368 20952
rect 17316 18624 17368 18630
rect 17316 18566 17368 18572
rect 17328 18290 17356 18566
rect 17316 18284 17368 18290
rect 17316 18226 17368 18232
rect 17316 16788 17368 16794
rect 17236 16748 17316 16776
rect 17316 16730 17368 16736
rect 17052 16646 17264 16674
rect 17236 16590 17264 16646
rect 17224 16584 17276 16590
rect 17224 16526 17276 16532
rect 17132 16516 17184 16522
rect 17132 16458 17184 16464
rect 16948 16108 17000 16114
rect 16948 16050 17000 16056
rect 16856 15972 16908 15978
rect 16856 15914 16908 15920
rect 16960 15502 16988 16050
rect 17144 15706 17172 16458
rect 17132 15700 17184 15706
rect 17132 15642 17184 15648
rect 16948 15496 17000 15502
rect 16948 15438 17000 15444
rect 17420 12434 17448 24754
rect 17500 24336 17552 24342
rect 17500 24278 17552 24284
rect 17512 23730 17540 24278
rect 17500 23724 17552 23730
rect 17500 23666 17552 23672
rect 17500 23316 17552 23322
rect 17500 23258 17552 23264
rect 17512 22273 17540 23258
rect 17498 22264 17554 22273
rect 17498 22199 17554 22208
rect 17500 22160 17552 22166
rect 17500 22102 17552 22108
rect 17512 21690 17540 22102
rect 17500 21684 17552 21690
rect 17500 21626 17552 21632
rect 17500 18760 17552 18766
rect 17500 18702 17552 18708
rect 17512 18426 17540 18702
rect 17500 18420 17552 18426
rect 17500 18362 17552 18368
rect 17500 18284 17552 18290
rect 17500 18226 17552 18232
rect 17512 17610 17540 18226
rect 17500 17604 17552 17610
rect 17500 17546 17552 17552
rect 17236 12406 17448 12434
rect 17236 10674 17264 12406
rect 17224 10668 17276 10674
rect 17224 10610 17276 10616
rect 16592 6886 16712 6914
rect 16684 3670 16712 6886
rect 17604 5098 17632 26318
rect 17696 25906 17724 26930
rect 17684 25900 17736 25906
rect 17684 25842 17736 25848
rect 17788 25158 17816 26930
rect 18064 26908 18092 27406
rect 18156 27062 18184 27503
rect 18236 27474 18288 27480
rect 18236 27328 18288 27334
rect 18236 27270 18288 27276
rect 18248 27130 18276 27270
rect 18236 27124 18288 27130
rect 18236 27066 18288 27072
rect 18144 27056 18196 27062
rect 18144 26998 18196 27004
rect 18064 26880 18276 26908
rect 18052 26784 18104 26790
rect 18144 26784 18196 26790
rect 18052 26726 18104 26732
rect 18142 26752 18144 26761
rect 18196 26752 18198 26761
rect 17868 26512 17920 26518
rect 17868 26454 17920 26460
rect 17776 25152 17828 25158
rect 17776 25094 17828 25100
rect 17684 23860 17736 23866
rect 17684 23802 17736 23808
rect 17696 22953 17724 23802
rect 17880 23050 17908 26454
rect 17958 26208 18014 26217
rect 17958 26143 18014 26152
rect 17972 25430 18000 26143
rect 18064 25702 18092 26726
rect 18142 26687 18198 26696
rect 18144 26444 18196 26450
rect 18144 26386 18196 26392
rect 18052 25696 18104 25702
rect 18052 25638 18104 25644
rect 17960 25424 18012 25430
rect 17960 25366 18012 25372
rect 18064 24750 18092 25638
rect 18156 25362 18184 26386
rect 18248 26314 18276 26880
rect 18340 26450 18368 27882
rect 18432 27538 18460 28455
rect 18420 27532 18472 27538
rect 18420 27474 18472 27480
rect 18418 27296 18474 27305
rect 18418 27231 18474 27240
rect 18432 27062 18460 27231
rect 18524 27130 18552 31622
rect 18616 27946 18644 31962
rect 18696 31680 18748 31686
rect 18696 31622 18748 31628
rect 18708 28014 18736 31622
rect 18788 30660 18840 30666
rect 18788 30602 18840 30608
rect 18880 30660 18932 30666
rect 18880 30602 18932 30608
rect 18800 29034 18828 30602
rect 18892 30569 18920 30602
rect 18984 30598 19012 33866
rect 19168 33522 19196 34360
rect 19892 34342 19944 34348
rect 19338 34303 19394 34312
rect 19248 34060 19300 34066
rect 19248 34002 19300 34008
rect 19156 33516 19208 33522
rect 19260 33504 19288 34002
rect 19340 33924 19392 33930
rect 19340 33866 19392 33872
rect 19352 33833 19380 33866
rect 19338 33824 19394 33833
rect 19338 33759 19394 33768
rect 19478 33756 19786 33776
rect 19478 33754 19484 33756
rect 19540 33754 19564 33756
rect 19620 33754 19644 33756
rect 19700 33754 19724 33756
rect 19780 33754 19786 33756
rect 19540 33702 19542 33754
rect 19722 33702 19724 33754
rect 19478 33700 19484 33702
rect 19540 33700 19564 33702
rect 19620 33700 19644 33702
rect 19700 33700 19724 33702
rect 19780 33700 19786 33702
rect 19478 33680 19786 33700
rect 19904 33590 19932 34342
rect 19996 34202 20024 34546
rect 20088 34474 20116 38966
rect 20180 38418 20208 39510
rect 20364 39030 20392 40598
rect 20352 39024 20404 39030
rect 20352 38966 20404 38972
rect 20260 38956 20312 38962
rect 20640 38944 20668 41200
rect 21272 40044 21324 40050
rect 21272 39986 21324 39992
rect 20812 39908 20864 39914
rect 20812 39850 20864 39856
rect 20260 38898 20312 38904
rect 20548 38916 20668 38944
rect 20720 38956 20772 38962
rect 20168 38412 20220 38418
rect 20168 38354 20220 38360
rect 20168 36916 20220 36922
rect 20168 36858 20220 36864
rect 20180 36009 20208 36858
rect 20166 36000 20222 36009
rect 20166 35935 20222 35944
rect 20272 35612 20300 38898
rect 20548 38418 20576 38916
rect 20720 38898 20772 38904
rect 20628 38752 20680 38758
rect 20628 38694 20680 38700
rect 20536 38412 20588 38418
rect 20536 38354 20588 38360
rect 20352 37868 20404 37874
rect 20352 37810 20404 37816
rect 20364 37262 20392 37810
rect 20444 37664 20496 37670
rect 20444 37606 20496 37612
rect 20352 37256 20404 37262
rect 20352 37198 20404 37204
rect 20364 36174 20392 37198
rect 20352 36168 20404 36174
rect 20352 36110 20404 36116
rect 20350 35864 20406 35873
rect 20350 35799 20406 35808
rect 20364 35630 20392 35799
rect 20180 35584 20300 35612
rect 20352 35624 20404 35630
rect 20180 35000 20208 35584
rect 20352 35566 20404 35572
rect 20456 35136 20484 37606
rect 20534 37360 20590 37369
rect 20534 37295 20590 37304
rect 20548 35766 20576 37295
rect 20536 35760 20588 35766
rect 20536 35702 20588 35708
rect 20364 35108 20484 35136
rect 20534 35184 20590 35193
rect 20534 35119 20590 35128
rect 20180 34972 20300 35000
rect 20166 34912 20222 34921
rect 20166 34847 20222 34856
rect 20180 34746 20208 34847
rect 20168 34740 20220 34746
rect 20168 34682 20220 34688
rect 20168 34536 20220 34542
rect 20168 34478 20220 34484
rect 20076 34468 20128 34474
rect 20076 34410 20128 34416
rect 20180 34202 20208 34478
rect 19984 34196 20036 34202
rect 19984 34138 20036 34144
rect 20168 34196 20220 34202
rect 20168 34138 20220 34144
rect 20168 33856 20220 33862
rect 20168 33798 20220 33804
rect 20180 33658 20208 33798
rect 20168 33652 20220 33658
rect 20168 33594 20220 33600
rect 19432 33584 19484 33590
rect 19432 33526 19484 33532
rect 19892 33584 19944 33590
rect 20272 33538 20300 34972
rect 19892 33526 19944 33532
rect 19340 33516 19392 33522
rect 19260 33476 19340 33504
rect 19156 33458 19208 33464
rect 19340 33458 19392 33464
rect 19444 33318 19472 33526
rect 19616 33516 19668 33522
rect 19616 33458 19668 33464
rect 20180 33510 20300 33538
rect 19432 33312 19484 33318
rect 19432 33254 19484 33260
rect 19444 32910 19472 33254
rect 19628 32978 19656 33458
rect 19800 33380 19852 33386
rect 19800 33322 19852 33328
rect 19616 32972 19668 32978
rect 19616 32914 19668 32920
rect 19812 32910 19840 33322
rect 19248 32904 19300 32910
rect 19248 32846 19300 32852
rect 19432 32904 19484 32910
rect 19432 32846 19484 32852
rect 19708 32904 19760 32910
rect 19708 32846 19760 32852
rect 19800 32904 19852 32910
rect 19800 32846 19852 32852
rect 19260 32366 19288 32846
rect 19340 32768 19392 32774
rect 19338 32736 19340 32745
rect 19720 32756 19748 32846
rect 19892 32768 19944 32774
rect 19392 32736 19394 32745
rect 19720 32728 19892 32756
rect 19892 32710 19944 32716
rect 19338 32671 19394 32680
rect 19352 32473 19380 32671
rect 19478 32668 19786 32688
rect 19478 32666 19484 32668
rect 19540 32666 19564 32668
rect 19620 32666 19644 32668
rect 19700 32666 19724 32668
rect 19780 32666 19786 32668
rect 19540 32614 19542 32666
rect 19722 32614 19724 32666
rect 19478 32612 19484 32614
rect 19540 32612 19564 32614
rect 19620 32612 19644 32614
rect 19700 32612 19724 32614
rect 19780 32612 19786 32614
rect 19478 32592 19786 32612
rect 19338 32464 19394 32473
rect 19338 32399 19394 32408
rect 19984 32428 20036 32434
rect 19984 32370 20036 32376
rect 19248 32360 19300 32366
rect 19248 32302 19300 32308
rect 19260 32065 19288 32302
rect 19996 32230 20024 32370
rect 19984 32224 20036 32230
rect 19522 32192 19578 32201
rect 19984 32166 20036 32172
rect 19522 32127 19578 32136
rect 19246 32056 19302 32065
rect 19246 31991 19302 32000
rect 19536 31890 19564 32127
rect 19708 32020 19760 32026
rect 19708 31962 19760 31968
rect 19524 31884 19576 31890
rect 19524 31826 19576 31832
rect 19720 31822 19748 31962
rect 19892 31884 19944 31890
rect 19892 31826 19944 31832
rect 19708 31816 19760 31822
rect 19708 31758 19760 31764
rect 19340 31748 19392 31754
rect 19340 31690 19392 31696
rect 19154 31240 19210 31249
rect 19154 31175 19210 31184
rect 19064 31136 19116 31142
rect 19064 31078 19116 31084
rect 19076 30802 19104 31078
rect 19064 30796 19116 30802
rect 19064 30738 19116 30744
rect 19076 30705 19104 30738
rect 19062 30696 19118 30705
rect 19062 30631 19118 30640
rect 18972 30592 19024 30598
rect 18878 30560 18934 30569
rect 18972 30534 19024 30540
rect 18878 30495 18934 30504
rect 18972 30388 19024 30394
rect 18972 30330 19024 30336
rect 18880 30320 18932 30326
rect 18880 30262 18932 30268
rect 18892 29850 18920 30262
rect 18880 29844 18932 29850
rect 18880 29786 18932 29792
rect 18880 29504 18932 29510
rect 18880 29446 18932 29452
rect 18892 29306 18920 29446
rect 18880 29300 18932 29306
rect 18880 29242 18932 29248
rect 18788 29028 18840 29034
rect 18788 28970 18840 28976
rect 18696 28008 18748 28014
rect 18696 27950 18748 27956
rect 18604 27940 18656 27946
rect 18604 27882 18656 27888
rect 18602 27704 18658 27713
rect 18602 27639 18658 27648
rect 18616 27554 18644 27639
rect 18616 27526 18736 27554
rect 18604 27464 18656 27470
rect 18604 27406 18656 27412
rect 18512 27124 18564 27130
rect 18512 27066 18564 27072
rect 18420 27056 18472 27062
rect 18420 26998 18472 27004
rect 18512 26920 18564 26926
rect 18512 26862 18564 26868
rect 18418 26616 18474 26625
rect 18418 26551 18420 26560
rect 18472 26551 18474 26560
rect 18420 26522 18472 26528
rect 18328 26444 18380 26450
rect 18328 26386 18380 26392
rect 18236 26308 18288 26314
rect 18236 26250 18288 26256
rect 18248 25702 18276 26250
rect 18524 25906 18552 26862
rect 18616 26586 18644 27406
rect 18604 26580 18656 26586
rect 18604 26522 18656 26528
rect 18604 26240 18656 26246
rect 18604 26182 18656 26188
rect 18616 25974 18644 26182
rect 18604 25968 18656 25974
rect 18604 25910 18656 25916
rect 18328 25900 18380 25906
rect 18328 25842 18380 25848
rect 18512 25900 18564 25906
rect 18512 25842 18564 25848
rect 18236 25696 18288 25702
rect 18236 25638 18288 25644
rect 18144 25356 18196 25362
rect 18144 25298 18196 25304
rect 18142 24848 18198 24857
rect 18248 24818 18276 25638
rect 18340 25276 18368 25842
rect 18708 25294 18736 27526
rect 18800 26450 18828 28970
rect 18880 27600 18932 27606
rect 18880 27542 18932 27548
rect 18892 27441 18920 27542
rect 18878 27432 18934 27441
rect 18878 27367 18934 27376
rect 18880 26988 18932 26994
rect 18880 26930 18932 26936
rect 18892 26489 18920 26930
rect 18878 26480 18934 26489
rect 18788 26444 18840 26450
rect 18878 26415 18934 26424
rect 18788 26386 18840 26392
rect 18880 26376 18932 26382
rect 18880 26318 18932 26324
rect 18892 26246 18920 26318
rect 18880 26240 18932 26246
rect 18880 26182 18932 26188
rect 18604 25288 18656 25294
rect 18340 25248 18604 25276
rect 18340 24936 18368 25248
rect 18604 25230 18656 25236
rect 18696 25288 18748 25294
rect 18696 25230 18748 25236
rect 18340 24908 18460 24936
rect 18432 24818 18460 24908
rect 18142 24783 18198 24792
rect 18236 24812 18288 24818
rect 18052 24744 18104 24750
rect 18052 24686 18104 24692
rect 18156 24206 18184 24783
rect 18236 24754 18288 24760
rect 18420 24812 18472 24818
rect 18472 24772 18552 24800
rect 18420 24754 18472 24760
rect 18144 24200 18196 24206
rect 17972 24160 18144 24188
rect 17868 23044 17920 23050
rect 17868 22986 17920 22992
rect 17682 22944 17738 22953
rect 17682 22879 17738 22888
rect 17774 22808 17830 22817
rect 17774 22743 17830 22752
rect 17788 22574 17816 22743
rect 17972 22681 18000 24160
rect 18144 24142 18196 24148
rect 18236 24132 18288 24138
rect 18288 24092 18368 24120
rect 18236 24074 18288 24080
rect 18234 24032 18290 24041
rect 18340 24018 18368 24092
rect 18418 24032 18474 24041
rect 18340 23990 18418 24018
rect 18234 23967 18290 23976
rect 18418 23967 18474 23976
rect 18144 23724 18196 23730
rect 18144 23666 18196 23672
rect 18052 23656 18104 23662
rect 18052 23598 18104 23604
rect 18064 22778 18092 23598
rect 18156 23322 18184 23666
rect 18144 23316 18196 23322
rect 18144 23258 18196 23264
rect 18142 23216 18198 23225
rect 18248 23202 18276 23967
rect 18420 23724 18472 23730
rect 18420 23666 18472 23672
rect 18328 23588 18380 23594
rect 18328 23530 18380 23536
rect 18340 23361 18368 23530
rect 18326 23352 18382 23361
rect 18326 23287 18382 23296
rect 18432 23254 18460 23666
rect 18420 23248 18472 23254
rect 18326 23216 18382 23225
rect 18248 23174 18326 23202
rect 18142 23151 18198 23160
rect 18420 23190 18472 23196
rect 18326 23151 18382 23160
rect 18156 22778 18184 23151
rect 18420 23112 18472 23118
rect 18420 23054 18472 23060
rect 18328 23044 18380 23050
rect 18328 22986 18380 22992
rect 18052 22772 18104 22778
rect 18052 22714 18104 22720
rect 18144 22772 18196 22778
rect 18144 22714 18196 22720
rect 17958 22672 18014 22681
rect 17958 22607 18014 22616
rect 17776 22568 17828 22574
rect 17776 22510 17828 22516
rect 17684 22024 17736 22030
rect 17684 21966 17736 21972
rect 17696 21554 17724 21966
rect 17684 21548 17736 21554
rect 17684 21490 17736 21496
rect 17788 21010 17816 22510
rect 18050 22400 18106 22409
rect 18050 22335 18106 22344
rect 17868 22160 17920 22166
rect 17868 22102 17920 22108
rect 17776 21004 17828 21010
rect 17776 20946 17828 20952
rect 17880 20942 17908 22102
rect 17960 21480 18012 21486
rect 17960 21422 18012 21428
rect 17972 20942 18000 21422
rect 18064 21078 18092 22335
rect 18340 22094 18368 22986
rect 18432 22506 18460 23054
rect 18524 22794 18552 24772
rect 18696 24608 18748 24614
rect 18696 24550 18748 24556
rect 18708 24342 18736 24550
rect 18696 24336 18748 24342
rect 18696 24278 18748 24284
rect 18984 24206 19012 30330
rect 19064 30252 19116 30258
rect 19064 30194 19116 30200
rect 19076 29628 19104 30194
rect 19168 30054 19196 31175
rect 19352 30802 19380 31690
rect 19478 31580 19786 31600
rect 19478 31578 19484 31580
rect 19540 31578 19564 31580
rect 19620 31578 19644 31580
rect 19700 31578 19724 31580
rect 19780 31578 19786 31580
rect 19540 31526 19542 31578
rect 19722 31526 19724 31578
rect 19478 31524 19484 31526
rect 19540 31524 19564 31526
rect 19620 31524 19644 31526
rect 19700 31524 19724 31526
rect 19780 31524 19786 31526
rect 19478 31504 19786 31524
rect 19904 31362 19932 31826
rect 19996 31754 20024 32166
rect 20076 31816 20128 31822
rect 20076 31758 20128 31764
rect 19984 31748 20036 31754
rect 19984 31690 20036 31696
rect 19812 31334 19932 31362
rect 19340 30796 19392 30802
rect 19340 30738 19392 30744
rect 19616 30728 19668 30734
rect 19614 30696 19616 30705
rect 19668 30696 19670 30705
rect 19812 30666 19840 31334
rect 19892 31272 19944 31278
rect 19892 31214 19944 31220
rect 19904 30682 19932 31214
rect 19996 30938 20024 31690
rect 20088 31482 20116 31758
rect 20076 31476 20128 31482
rect 20076 31418 20128 31424
rect 19984 30932 20036 30938
rect 19984 30874 20036 30880
rect 20088 30802 20116 31418
rect 20180 30938 20208 33510
rect 20364 32842 20392 35108
rect 20548 34785 20576 35119
rect 20534 34776 20590 34785
rect 20534 34711 20590 34720
rect 20640 34610 20668 38694
rect 20628 34604 20680 34610
rect 20628 34546 20680 34552
rect 20444 34536 20496 34542
rect 20444 34478 20496 34484
rect 20352 32836 20404 32842
rect 20352 32778 20404 32784
rect 20364 32065 20392 32778
rect 20350 32056 20406 32065
rect 20260 32020 20312 32026
rect 20456 32026 20484 34478
rect 20536 34400 20588 34406
rect 20536 34342 20588 34348
rect 20628 34400 20680 34406
rect 20628 34342 20680 34348
rect 20350 31991 20406 32000
rect 20444 32020 20496 32026
rect 20260 31962 20312 31968
rect 20444 31962 20496 31968
rect 20272 31890 20300 31962
rect 20260 31884 20312 31890
rect 20548 31872 20576 34342
rect 20640 34202 20668 34342
rect 20628 34196 20680 34202
rect 20628 34138 20680 34144
rect 20628 33992 20680 33998
rect 20628 33934 20680 33940
rect 20640 32910 20668 33934
rect 20628 32904 20680 32910
rect 20628 32846 20680 32852
rect 20640 32434 20668 32846
rect 20732 32502 20760 38898
rect 20824 37874 20852 39850
rect 20996 39296 21048 39302
rect 20996 39238 21048 39244
rect 20904 38208 20956 38214
rect 20904 38150 20956 38156
rect 20916 37913 20944 38150
rect 20902 37904 20958 37913
rect 20812 37868 20864 37874
rect 20902 37839 20958 37848
rect 20812 37810 20864 37816
rect 20824 37670 20852 37810
rect 20812 37664 20864 37670
rect 20812 37606 20864 37612
rect 20904 37188 20956 37194
rect 20904 37130 20956 37136
rect 20916 36786 20944 37130
rect 20904 36780 20956 36786
rect 20904 36722 20956 36728
rect 20812 36712 20864 36718
rect 20810 36680 20812 36689
rect 20864 36680 20866 36689
rect 20810 36615 20866 36624
rect 20812 36576 20864 36582
rect 20810 36544 20812 36553
rect 20864 36544 20866 36553
rect 20810 36479 20866 36488
rect 20824 36156 20852 36479
rect 20916 36281 20944 36722
rect 20902 36272 20958 36281
rect 20902 36207 20958 36216
rect 20824 36128 20944 36156
rect 20812 36032 20864 36038
rect 20812 35974 20864 35980
rect 20824 35834 20852 35974
rect 20812 35828 20864 35834
rect 20812 35770 20864 35776
rect 20810 35728 20866 35737
rect 20916 35698 20944 36128
rect 21008 35737 21036 39238
rect 21178 38584 21234 38593
rect 21178 38519 21234 38528
rect 21192 36106 21220 38519
rect 21180 36100 21232 36106
rect 21180 36042 21232 36048
rect 20994 35728 21050 35737
rect 20810 35663 20866 35672
rect 20904 35692 20956 35698
rect 20824 35630 20852 35663
rect 20994 35663 21050 35672
rect 20904 35634 20956 35640
rect 20812 35624 20864 35630
rect 20812 35566 20864 35572
rect 20916 35193 20944 35634
rect 21088 35624 21140 35630
rect 21088 35566 21140 35572
rect 21100 35465 21128 35566
rect 21086 35456 21142 35465
rect 21086 35391 21142 35400
rect 20902 35184 20958 35193
rect 20902 35119 20958 35128
rect 20996 35012 21048 35018
rect 20996 34954 21048 34960
rect 20904 34944 20956 34950
rect 20810 34912 20866 34921
rect 20904 34886 20956 34892
rect 20810 34847 20866 34856
rect 20824 34746 20852 34847
rect 20812 34740 20864 34746
rect 20812 34682 20864 34688
rect 20810 34640 20866 34649
rect 20810 34575 20866 34584
rect 20824 33862 20852 34575
rect 20916 34542 20944 34886
rect 21008 34610 21036 34954
rect 20996 34604 21048 34610
rect 20996 34546 21048 34552
rect 20904 34536 20956 34542
rect 20904 34478 20956 34484
rect 20996 34468 21048 34474
rect 20996 34410 21048 34416
rect 20902 34368 20958 34377
rect 20902 34303 20958 34312
rect 20812 33856 20864 33862
rect 20812 33798 20864 33804
rect 20916 33402 20944 34303
rect 21008 33538 21036 34410
rect 21100 34134 21128 35391
rect 21192 34474 21220 36042
rect 21284 36009 21312 39986
rect 21822 39808 21878 39817
rect 21822 39743 21878 39752
rect 21548 38344 21600 38350
rect 21548 38286 21600 38292
rect 21364 37392 21416 37398
rect 21364 37334 21416 37340
rect 21270 36000 21326 36009
rect 21270 35935 21326 35944
rect 21272 35556 21324 35562
rect 21272 35498 21324 35504
rect 21284 34950 21312 35498
rect 21272 34944 21324 34950
rect 21270 34912 21272 34921
rect 21324 34912 21326 34921
rect 21270 34847 21326 34856
rect 21180 34468 21232 34474
rect 21180 34410 21232 34416
rect 21178 34368 21234 34377
rect 21178 34303 21234 34312
rect 21088 34128 21140 34134
rect 21192 34105 21220 34303
rect 21376 34184 21404 37334
rect 21456 37256 21508 37262
rect 21456 37198 21508 37204
rect 21468 36922 21496 37198
rect 21456 36916 21508 36922
rect 21456 36858 21508 36864
rect 21456 36780 21508 36786
rect 21456 36722 21508 36728
rect 21284 34156 21404 34184
rect 21088 34070 21140 34076
rect 21178 34096 21234 34105
rect 21100 33658 21128 34070
rect 21178 34031 21234 34040
rect 21088 33652 21140 33658
rect 21088 33594 21140 33600
rect 21008 33510 21220 33538
rect 20916 33374 21036 33402
rect 20902 33008 20958 33017
rect 20902 32943 20958 32952
rect 20720 32496 20772 32502
rect 20720 32438 20772 32444
rect 20628 32428 20680 32434
rect 20628 32370 20680 32376
rect 20640 32178 20668 32370
rect 20640 32150 20760 32178
rect 20732 31906 20760 32150
rect 20732 31878 20852 31906
rect 20260 31826 20312 31832
rect 20456 31844 20576 31872
rect 20352 31680 20404 31686
rect 20352 31622 20404 31628
rect 20260 31136 20312 31142
rect 20260 31078 20312 31084
rect 20272 30938 20300 31078
rect 20168 30932 20220 30938
rect 20168 30874 20220 30880
rect 20260 30932 20312 30938
rect 20260 30874 20312 30880
rect 20076 30796 20128 30802
rect 20076 30738 20128 30744
rect 20168 30728 20220 30734
rect 19904 30676 20168 30682
rect 19904 30670 20220 30676
rect 19614 30631 19670 30640
rect 19800 30660 19852 30666
rect 19800 30602 19852 30608
rect 19904 30654 20208 30670
rect 20260 30660 20312 30666
rect 19478 30492 19786 30512
rect 19478 30490 19484 30492
rect 19540 30490 19564 30492
rect 19620 30490 19644 30492
rect 19700 30490 19724 30492
rect 19780 30490 19786 30492
rect 19540 30438 19542 30490
rect 19722 30438 19724 30490
rect 19478 30436 19484 30438
rect 19540 30436 19564 30438
rect 19620 30436 19644 30438
rect 19700 30436 19724 30438
rect 19780 30436 19786 30438
rect 19478 30416 19786 30436
rect 19904 30394 19932 30654
rect 20260 30602 20312 30608
rect 19892 30388 19944 30394
rect 19892 30330 19944 30336
rect 20076 30388 20128 30394
rect 20076 30330 20128 30336
rect 19248 30320 19300 30326
rect 19248 30262 19300 30268
rect 19156 30048 19208 30054
rect 19156 29990 19208 29996
rect 19260 29753 19288 30262
rect 19430 30152 19486 30161
rect 19430 30087 19486 30096
rect 19246 29744 19302 29753
rect 19246 29679 19302 29688
rect 19444 29646 19472 30087
rect 19248 29640 19300 29646
rect 19076 29600 19248 29628
rect 19432 29640 19484 29646
rect 19248 29582 19300 29588
rect 19338 29608 19394 29617
rect 19432 29582 19484 29588
rect 19338 29543 19394 29552
rect 19062 29472 19118 29481
rect 19062 29407 19118 29416
rect 19076 29306 19104 29407
rect 19064 29300 19116 29306
rect 19064 29242 19116 29248
rect 19352 28801 19380 29543
rect 19478 29404 19786 29424
rect 19478 29402 19484 29404
rect 19540 29402 19564 29404
rect 19620 29402 19644 29404
rect 19700 29402 19724 29404
rect 19780 29402 19786 29404
rect 19540 29350 19542 29402
rect 19722 29350 19724 29402
rect 19478 29348 19484 29350
rect 19540 29348 19564 29350
rect 19620 29348 19644 29350
rect 19700 29348 19724 29350
rect 19780 29348 19786 29350
rect 19478 29328 19786 29348
rect 19708 29096 19760 29102
rect 19904 29084 19932 30330
rect 19982 30152 20038 30161
rect 19982 30087 20038 30096
rect 19996 29850 20024 30087
rect 19984 29844 20036 29850
rect 19984 29786 20036 29792
rect 19984 29572 20036 29578
rect 19984 29514 20036 29520
rect 19760 29056 19932 29084
rect 19708 29038 19760 29044
rect 19338 28792 19394 28801
rect 19338 28727 19394 28736
rect 19890 28792 19946 28801
rect 19890 28727 19946 28736
rect 19904 28694 19932 28727
rect 19892 28688 19944 28694
rect 19798 28656 19854 28665
rect 19156 28620 19208 28626
rect 19156 28562 19208 28568
rect 19708 28620 19760 28626
rect 19892 28630 19944 28636
rect 19798 28591 19854 28600
rect 19708 28562 19760 28568
rect 19062 28520 19118 28529
rect 19062 28455 19118 28464
rect 19076 28082 19104 28455
rect 19064 28076 19116 28082
rect 19064 28018 19116 28024
rect 19064 27396 19116 27402
rect 19064 27338 19116 27344
rect 19076 26761 19104 27338
rect 19062 26752 19118 26761
rect 19168 26738 19196 28562
rect 19720 28529 19748 28562
rect 19706 28520 19762 28529
rect 19340 28484 19392 28490
rect 19812 28490 19840 28591
rect 19706 28455 19762 28464
rect 19800 28484 19852 28490
rect 19340 28426 19392 28432
rect 19800 28426 19852 28432
rect 19246 27840 19302 27849
rect 19246 27775 19302 27784
rect 19260 27402 19288 27775
rect 19352 27402 19380 28426
rect 19892 28416 19944 28422
rect 19892 28358 19944 28364
rect 19478 28316 19786 28336
rect 19478 28314 19484 28316
rect 19540 28314 19564 28316
rect 19620 28314 19644 28316
rect 19700 28314 19724 28316
rect 19780 28314 19786 28316
rect 19540 28262 19542 28314
rect 19722 28262 19724 28314
rect 19478 28260 19484 28262
rect 19540 28260 19564 28262
rect 19620 28260 19644 28262
rect 19700 28260 19724 28262
rect 19780 28260 19786 28262
rect 19478 28240 19786 28260
rect 19248 27396 19300 27402
rect 19248 27338 19300 27344
rect 19340 27396 19392 27402
rect 19340 27338 19392 27344
rect 19478 27228 19786 27248
rect 19478 27226 19484 27228
rect 19540 27226 19564 27228
rect 19620 27226 19644 27228
rect 19700 27226 19724 27228
rect 19780 27226 19786 27228
rect 19540 27174 19542 27226
rect 19722 27174 19724 27226
rect 19478 27172 19484 27174
rect 19540 27172 19564 27174
rect 19620 27172 19644 27174
rect 19700 27172 19724 27174
rect 19780 27172 19786 27174
rect 19478 27152 19786 27172
rect 19260 26858 19380 26874
rect 19248 26852 19380 26858
rect 19300 26846 19380 26852
rect 19248 26794 19300 26800
rect 19168 26710 19288 26738
rect 19062 26687 19118 26696
rect 18696 24200 18748 24206
rect 18696 24142 18748 24148
rect 18972 24200 19024 24206
rect 18972 24142 19024 24148
rect 18604 24132 18656 24138
rect 18604 24074 18656 24080
rect 18616 23798 18644 24074
rect 18604 23792 18656 23798
rect 18604 23734 18656 23740
rect 18604 23656 18656 23662
rect 18604 23598 18656 23604
rect 18616 23225 18644 23598
rect 18602 23216 18658 23225
rect 18602 23151 18658 23160
rect 18524 22766 18644 22794
rect 18510 22672 18566 22681
rect 18510 22607 18512 22616
rect 18564 22607 18566 22616
rect 18512 22578 18564 22584
rect 18420 22500 18472 22506
rect 18420 22442 18472 22448
rect 18340 22066 18460 22094
rect 18236 22024 18288 22030
rect 18328 22024 18380 22030
rect 18236 21966 18288 21972
rect 18326 21992 18328 22001
rect 18380 21992 18382 22001
rect 18144 21548 18196 21554
rect 18144 21490 18196 21496
rect 18052 21072 18104 21078
rect 18052 21014 18104 21020
rect 17684 20936 17736 20942
rect 17868 20936 17920 20942
rect 17684 20878 17736 20884
rect 17774 20904 17830 20913
rect 17696 20058 17724 20878
rect 17868 20878 17920 20884
rect 17960 20936 18012 20942
rect 17960 20878 18012 20884
rect 17774 20839 17830 20848
rect 17684 20052 17736 20058
rect 17684 19994 17736 20000
rect 17696 17270 17724 19994
rect 17684 17264 17736 17270
rect 17684 17206 17736 17212
rect 17788 16998 17816 20839
rect 17868 20596 17920 20602
rect 17868 20538 17920 20544
rect 17880 19242 17908 20538
rect 18156 20058 18184 21490
rect 18248 20602 18276 21966
rect 18326 21927 18382 21936
rect 18236 20596 18288 20602
rect 18236 20538 18288 20544
rect 18144 20052 18196 20058
rect 18144 19994 18196 20000
rect 18340 19990 18368 21927
rect 18328 19984 18380 19990
rect 18328 19926 18380 19932
rect 17960 19848 18012 19854
rect 17960 19790 18012 19796
rect 17868 19236 17920 19242
rect 17868 19178 17920 19184
rect 17972 18986 18000 19790
rect 18432 19446 18460 22066
rect 18616 22030 18644 22766
rect 18604 22024 18656 22030
rect 18604 21966 18656 21972
rect 18510 21720 18566 21729
rect 18510 21655 18566 21664
rect 18524 21418 18552 21655
rect 18512 21412 18564 21418
rect 18512 21354 18564 21360
rect 18708 21010 18736 24142
rect 18788 24132 18840 24138
rect 18788 24074 18840 24080
rect 18800 24041 18828 24074
rect 18786 24032 18842 24041
rect 18786 23967 18842 23976
rect 18786 23896 18842 23905
rect 19076 23882 19104 26687
rect 19156 25900 19208 25906
rect 19156 25842 19208 25848
rect 19168 25809 19196 25842
rect 19154 25800 19210 25809
rect 19154 25735 19210 25744
rect 19154 25392 19210 25401
rect 19154 25327 19156 25336
rect 19208 25327 19210 25336
rect 19156 25298 19208 25304
rect 19168 24206 19196 25298
rect 19260 25242 19288 26710
rect 19352 26568 19380 26846
rect 19616 26580 19668 26586
rect 19352 26540 19616 26568
rect 19616 26522 19668 26528
rect 19706 26344 19762 26353
rect 19706 26279 19708 26288
rect 19760 26279 19762 26288
rect 19708 26250 19760 26256
rect 19904 26246 19932 28358
rect 19996 27130 20024 29514
rect 19984 27124 20036 27130
rect 19984 27066 20036 27072
rect 20088 27010 20116 30330
rect 20168 30184 20220 30190
rect 20168 30126 20220 30132
rect 19996 26982 20116 27010
rect 19892 26240 19944 26246
rect 19892 26182 19944 26188
rect 19478 26140 19786 26160
rect 19478 26138 19484 26140
rect 19540 26138 19564 26140
rect 19620 26138 19644 26140
rect 19700 26138 19724 26140
rect 19780 26138 19786 26140
rect 19540 26086 19542 26138
rect 19722 26086 19724 26138
rect 19478 26084 19484 26086
rect 19540 26084 19564 26086
rect 19620 26084 19644 26086
rect 19700 26084 19724 26086
rect 19780 26084 19786 26086
rect 19478 26064 19786 26084
rect 19892 25492 19944 25498
rect 19892 25434 19944 25440
rect 19904 25401 19932 25434
rect 19890 25392 19946 25401
rect 19890 25327 19946 25336
rect 19260 25214 19380 25242
rect 19248 25152 19300 25158
rect 19248 25094 19300 25100
rect 19156 24200 19208 24206
rect 19156 24142 19208 24148
rect 18786 23831 18788 23840
rect 18840 23831 18842 23840
rect 18984 23854 19104 23882
rect 18788 23802 18840 23808
rect 18880 23724 18932 23730
rect 18880 23666 18932 23672
rect 18788 23520 18840 23526
rect 18788 23462 18840 23468
rect 18800 23322 18828 23462
rect 18788 23316 18840 23322
rect 18788 23258 18840 23264
rect 18892 21690 18920 23666
rect 18880 21684 18932 21690
rect 18880 21626 18932 21632
rect 18696 21004 18748 21010
rect 18696 20946 18748 20952
rect 18984 20942 19012 23854
rect 19064 23792 19116 23798
rect 19064 23734 19116 23740
rect 19076 23322 19104 23734
rect 19064 23316 19116 23322
rect 19064 23258 19116 23264
rect 19168 23186 19196 24142
rect 19156 23180 19208 23186
rect 19156 23122 19208 23128
rect 19064 23112 19116 23118
rect 19064 23054 19116 23060
rect 19076 22953 19104 23054
rect 19062 22944 19118 22953
rect 19062 22879 19118 22888
rect 19168 22710 19196 23122
rect 19156 22704 19208 22710
rect 19156 22646 19208 22652
rect 19260 22098 19288 25094
rect 19352 24818 19380 25214
rect 19892 25152 19944 25158
rect 19890 25120 19892 25129
rect 19944 25120 19946 25129
rect 19478 25052 19786 25072
rect 19890 25055 19946 25064
rect 19478 25050 19484 25052
rect 19540 25050 19564 25052
rect 19620 25050 19644 25052
rect 19700 25050 19724 25052
rect 19780 25050 19786 25052
rect 19540 24998 19542 25050
rect 19722 24998 19724 25050
rect 19478 24996 19484 24998
rect 19540 24996 19564 24998
rect 19620 24996 19644 24998
rect 19700 24996 19724 24998
rect 19780 24996 19786 24998
rect 19478 24976 19786 24996
rect 19340 24812 19392 24818
rect 19340 24754 19392 24760
rect 19352 24449 19380 24754
rect 19338 24440 19394 24449
rect 19338 24375 19394 24384
rect 19478 23964 19786 23984
rect 19478 23962 19484 23964
rect 19540 23962 19564 23964
rect 19620 23962 19644 23964
rect 19700 23962 19724 23964
rect 19780 23962 19786 23964
rect 19540 23910 19542 23962
rect 19722 23910 19724 23962
rect 19478 23908 19484 23910
rect 19540 23908 19564 23910
rect 19620 23908 19644 23910
rect 19700 23908 19724 23910
rect 19780 23908 19786 23910
rect 19478 23888 19786 23908
rect 19904 23662 19932 25055
rect 19892 23656 19944 23662
rect 19892 23598 19944 23604
rect 19708 23588 19760 23594
rect 19708 23530 19760 23536
rect 19616 23520 19668 23526
rect 19352 23480 19616 23508
rect 19352 22642 19380 23480
rect 19616 23462 19668 23468
rect 19720 23361 19748 23530
rect 19706 23352 19762 23361
rect 19432 23316 19484 23322
rect 19706 23287 19762 23296
rect 19432 23258 19484 23264
rect 19444 23118 19472 23258
rect 19798 23216 19854 23225
rect 19798 23151 19800 23160
rect 19852 23151 19854 23160
rect 19800 23122 19852 23128
rect 19432 23112 19484 23118
rect 19432 23054 19484 23060
rect 19478 22876 19786 22896
rect 19478 22874 19484 22876
rect 19540 22874 19564 22876
rect 19620 22874 19644 22876
rect 19700 22874 19724 22876
rect 19780 22874 19786 22876
rect 19540 22822 19542 22874
rect 19722 22822 19724 22874
rect 19478 22820 19484 22822
rect 19540 22820 19564 22822
rect 19620 22820 19644 22822
rect 19700 22820 19724 22822
rect 19780 22820 19786 22822
rect 19478 22800 19786 22820
rect 19340 22636 19392 22642
rect 19340 22578 19392 22584
rect 19432 22636 19484 22642
rect 19432 22578 19484 22584
rect 19248 22092 19300 22098
rect 19248 22034 19300 22040
rect 19156 21888 19208 21894
rect 19444 21876 19472 22578
rect 19614 22536 19670 22545
rect 19614 22471 19670 22480
rect 19798 22536 19854 22545
rect 19798 22471 19854 22480
rect 19628 22438 19656 22471
rect 19616 22432 19668 22438
rect 19616 22374 19668 22380
rect 19614 22128 19670 22137
rect 19614 22063 19616 22072
rect 19668 22063 19670 22072
rect 19616 22034 19668 22040
rect 19208 21848 19288 21876
rect 19156 21830 19208 21836
rect 19156 21684 19208 21690
rect 19156 21626 19208 21632
rect 19168 21321 19196 21626
rect 19260 21468 19288 21848
rect 19352 21848 19472 21876
rect 19812 21876 19840 22471
rect 19904 22030 19932 23598
rect 19892 22024 19944 22030
rect 19892 21966 19944 21972
rect 19812 21848 19932 21876
rect 19352 21468 19380 21848
rect 19478 21788 19786 21808
rect 19478 21786 19484 21788
rect 19540 21786 19564 21788
rect 19620 21786 19644 21788
rect 19700 21786 19724 21788
rect 19780 21786 19786 21788
rect 19540 21734 19542 21786
rect 19722 21734 19724 21786
rect 19478 21732 19484 21734
rect 19540 21732 19564 21734
rect 19620 21732 19644 21734
rect 19700 21732 19724 21734
rect 19780 21732 19786 21734
rect 19478 21712 19786 21732
rect 19260 21440 19380 21468
rect 19154 21312 19210 21321
rect 19154 21247 19210 21256
rect 19260 21010 19288 21440
rect 19340 21344 19392 21350
rect 19340 21286 19392 21292
rect 19248 21004 19300 21010
rect 19248 20946 19300 20952
rect 18972 20936 19024 20942
rect 18972 20878 19024 20884
rect 18512 20800 18564 20806
rect 18510 20768 18512 20777
rect 18564 20768 18566 20777
rect 18510 20703 18566 20712
rect 18878 20632 18934 20641
rect 18878 20567 18934 20576
rect 18696 20052 18748 20058
rect 18696 19994 18748 20000
rect 18708 19718 18736 19994
rect 18892 19786 18920 20567
rect 19352 20466 19380 21286
rect 19904 21146 19932 21848
rect 19892 21140 19944 21146
rect 19892 21082 19944 21088
rect 19616 20936 19668 20942
rect 19668 20896 19932 20924
rect 19616 20878 19668 20884
rect 19478 20700 19786 20720
rect 19478 20698 19484 20700
rect 19540 20698 19564 20700
rect 19620 20698 19644 20700
rect 19700 20698 19724 20700
rect 19780 20698 19786 20700
rect 19540 20646 19542 20698
rect 19722 20646 19724 20698
rect 19478 20644 19484 20646
rect 19540 20644 19564 20646
rect 19620 20644 19644 20646
rect 19700 20644 19724 20646
rect 19780 20644 19786 20646
rect 19478 20624 19786 20644
rect 19432 20528 19484 20534
rect 19432 20470 19484 20476
rect 19340 20460 19392 20466
rect 19340 20402 19392 20408
rect 19444 19922 19472 20470
rect 19432 19916 19484 19922
rect 19432 19858 19484 19864
rect 19248 19848 19300 19854
rect 19248 19790 19300 19796
rect 18880 19780 18932 19786
rect 18880 19722 18932 19728
rect 18696 19712 18748 19718
rect 18696 19654 18748 19660
rect 18800 19514 19012 19530
rect 18788 19508 19024 19514
rect 18840 19502 18972 19508
rect 18788 19450 18840 19456
rect 18972 19450 19024 19456
rect 19260 19446 19288 19790
rect 19444 19700 19472 19858
rect 19524 19848 19576 19854
rect 19904 19836 19932 20896
rect 19576 19808 19932 19836
rect 19524 19790 19576 19796
rect 19352 19672 19472 19700
rect 19892 19712 19944 19718
rect 18420 19440 18472 19446
rect 18420 19382 18472 19388
rect 19248 19440 19300 19446
rect 19248 19382 19300 19388
rect 18052 19372 18104 19378
rect 18052 19314 18104 19320
rect 18328 19372 18380 19378
rect 18328 19314 18380 19320
rect 17880 18958 18000 18986
rect 17880 18426 17908 18958
rect 18064 18902 18092 19314
rect 17960 18896 18012 18902
rect 17960 18838 18012 18844
rect 18052 18896 18104 18902
rect 18052 18838 18104 18844
rect 17868 18420 17920 18426
rect 17868 18362 17920 18368
rect 17868 18284 17920 18290
rect 17868 18226 17920 18232
rect 17880 18086 17908 18226
rect 17868 18080 17920 18086
rect 17868 18022 17920 18028
rect 17776 16992 17828 16998
rect 17776 16934 17828 16940
rect 17788 15502 17816 16934
rect 17972 16046 18000 18838
rect 18144 18828 18196 18834
rect 18144 18770 18196 18776
rect 18052 18692 18104 18698
rect 18052 18634 18104 18640
rect 18064 18426 18092 18634
rect 18052 18420 18104 18426
rect 18052 18362 18104 18368
rect 18156 18222 18184 18770
rect 18236 18624 18288 18630
rect 18236 18566 18288 18572
rect 18144 18216 18196 18222
rect 18144 18158 18196 18164
rect 18156 16522 18184 18158
rect 18248 17882 18276 18566
rect 18340 18426 18368 19314
rect 18880 18964 18932 18970
rect 18880 18906 18932 18912
rect 18892 18766 18920 18906
rect 18420 18760 18472 18766
rect 18420 18702 18472 18708
rect 18880 18760 18932 18766
rect 18880 18702 18932 18708
rect 18328 18420 18380 18426
rect 18328 18362 18380 18368
rect 18326 18320 18382 18329
rect 18326 18255 18382 18264
rect 18340 18086 18368 18255
rect 18328 18080 18380 18086
rect 18328 18022 18380 18028
rect 18236 17876 18288 17882
rect 18236 17818 18288 17824
rect 18248 17678 18276 17818
rect 18432 17678 18460 18702
rect 18892 18290 18920 18702
rect 19248 18352 19300 18358
rect 19248 18294 19300 18300
rect 18880 18284 18932 18290
rect 18880 18226 18932 18232
rect 18236 17672 18288 17678
rect 18236 17614 18288 17620
rect 18420 17672 18472 17678
rect 18420 17614 18472 17620
rect 18432 17270 18460 17614
rect 19260 17610 19288 18294
rect 19352 18290 19380 19672
rect 19892 19654 19944 19660
rect 19478 19612 19786 19632
rect 19478 19610 19484 19612
rect 19540 19610 19564 19612
rect 19620 19610 19644 19612
rect 19700 19610 19724 19612
rect 19780 19610 19786 19612
rect 19540 19558 19542 19610
rect 19722 19558 19724 19610
rect 19478 19556 19484 19558
rect 19540 19556 19564 19558
rect 19620 19556 19644 19558
rect 19700 19556 19724 19558
rect 19780 19556 19786 19558
rect 19478 19536 19786 19556
rect 19800 19372 19852 19378
rect 19904 19360 19932 19654
rect 19852 19332 19932 19360
rect 19800 19314 19852 19320
rect 19432 19304 19484 19310
rect 19432 19246 19484 19252
rect 19444 18970 19472 19246
rect 19524 19236 19576 19242
rect 19524 19178 19576 19184
rect 19432 18964 19484 18970
rect 19432 18906 19484 18912
rect 19536 18698 19564 19178
rect 19892 18964 19944 18970
rect 19892 18906 19944 18912
rect 19524 18692 19576 18698
rect 19524 18634 19576 18640
rect 19904 18630 19932 18906
rect 19892 18624 19944 18630
rect 19892 18566 19944 18572
rect 19478 18524 19786 18544
rect 19478 18522 19484 18524
rect 19540 18522 19564 18524
rect 19620 18522 19644 18524
rect 19700 18522 19724 18524
rect 19780 18522 19786 18524
rect 19540 18470 19542 18522
rect 19722 18470 19724 18522
rect 19478 18468 19484 18470
rect 19540 18468 19564 18470
rect 19620 18468 19644 18470
rect 19700 18468 19724 18470
rect 19780 18468 19786 18470
rect 19478 18448 19786 18468
rect 19904 18290 19932 18566
rect 19340 18284 19392 18290
rect 19340 18226 19392 18232
rect 19892 18284 19944 18290
rect 19892 18226 19944 18232
rect 19340 17808 19392 17814
rect 19340 17750 19392 17756
rect 19248 17604 19300 17610
rect 19248 17546 19300 17552
rect 19260 17338 19288 17546
rect 19248 17332 19300 17338
rect 19248 17274 19300 17280
rect 18420 17264 18472 17270
rect 18420 17206 18472 17212
rect 18236 17196 18288 17202
rect 18236 17138 18288 17144
rect 18144 16516 18196 16522
rect 18144 16458 18196 16464
rect 18248 16250 18276 17138
rect 19352 16658 19380 17750
rect 19904 17678 19932 18226
rect 19892 17672 19944 17678
rect 19892 17614 19944 17620
rect 19478 17436 19786 17456
rect 19478 17434 19484 17436
rect 19540 17434 19564 17436
rect 19620 17434 19644 17436
rect 19700 17434 19724 17436
rect 19780 17434 19786 17436
rect 19540 17382 19542 17434
rect 19722 17382 19724 17434
rect 19478 17380 19484 17382
rect 19540 17380 19564 17382
rect 19620 17380 19644 17382
rect 19700 17380 19724 17382
rect 19780 17380 19786 17382
rect 19478 17360 19786 17380
rect 19904 17338 19932 17614
rect 19892 17332 19944 17338
rect 19892 17274 19944 17280
rect 19340 16652 19392 16658
rect 19340 16594 19392 16600
rect 18236 16244 18288 16250
rect 18236 16186 18288 16192
rect 19352 16114 19380 16594
rect 19904 16590 19932 17274
rect 19892 16584 19944 16590
rect 19892 16526 19944 16532
rect 19478 16348 19786 16368
rect 19478 16346 19484 16348
rect 19540 16346 19564 16348
rect 19620 16346 19644 16348
rect 19700 16346 19724 16348
rect 19780 16346 19786 16348
rect 19540 16294 19542 16346
rect 19722 16294 19724 16346
rect 19478 16292 19484 16294
rect 19540 16292 19564 16294
rect 19620 16292 19644 16294
rect 19700 16292 19724 16294
rect 19780 16292 19786 16294
rect 19478 16272 19786 16292
rect 19340 16108 19392 16114
rect 19340 16050 19392 16056
rect 17960 16040 18012 16046
rect 17960 15982 18012 15988
rect 17776 15496 17828 15502
rect 17776 15438 17828 15444
rect 19478 15260 19786 15280
rect 19478 15258 19484 15260
rect 19540 15258 19564 15260
rect 19620 15258 19644 15260
rect 19700 15258 19724 15260
rect 19780 15258 19786 15260
rect 19540 15206 19542 15258
rect 19722 15206 19724 15258
rect 19478 15204 19484 15206
rect 19540 15204 19564 15206
rect 19620 15204 19644 15206
rect 19700 15204 19724 15206
rect 19780 15204 19786 15206
rect 19478 15184 19786 15204
rect 19478 14172 19786 14192
rect 19478 14170 19484 14172
rect 19540 14170 19564 14172
rect 19620 14170 19644 14172
rect 19700 14170 19724 14172
rect 19780 14170 19786 14172
rect 19540 14118 19542 14170
rect 19722 14118 19724 14170
rect 19478 14116 19484 14118
rect 19540 14116 19564 14118
rect 19620 14116 19644 14118
rect 19700 14116 19724 14118
rect 19780 14116 19786 14118
rect 19478 14096 19786 14116
rect 19478 13084 19786 13104
rect 19478 13082 19484 13084
rect 19540 13082 19564 13084
rect 19620 13082 19644 13084
rect 19700 13082 19724 13084
rect 19780 13082 19786 13084
rect 19540 13030 19542 13082
rect 19722 13030 19724 13082
rect 19478 13028 19484 13030
rect 19540 13028 19564 13030
rect 19620 13028 19644 13030
rect 19700 13028 19724 13030
rect 19780 13028 19786 13030
rect 19478 13008 19786 13028
rect 19478 11996 19786 12016
rect 19478 11994 19484 11996
rect 19540 11994 19564 11996
rect 19620 11994 19644 11996
rect 19700 11994 19724 11996
rect 19780 11994 19786 11996
rect 19540 11942 19542 11994
rect 19722 11942 19724 11994
rect 19478 11940 19484 11942
rect 19540 11940 19564 11942
rect 19620 11940 19644 11942
rect 19700 11940 19724 11942
rect 19780 11940 19786 11942
rect 19478 11920 19786 11940
rect 19478 10908 19786 10928
rect 19478 10906 19484 10908
rect 19540 10906 19564 10908
rect 19620 10906 19644 10908
rect 19700 10906 19724 10908
rect 19780 10906 19786 10908
rect 19540 10854 19542 10906
rect 19722 10854 19724 10906
rect 19478 10852 19484 10854
rect 19540 10852 19564 10854
rect 19620 10852 19644 10854
rect 19700 10852 19724 10854
rect 19780 10852 19786 10854
rect 19478 10832 19786 10852
rect 19478 9820 19786 9840
rect 19478 9818 19484 9820
rect 19540 9818 19564 9820
rect 19620 9818 19644 9820
rect 19700 9818 19724 9820
rect 19780 9818 19786 9820
rect 19540 9766 19542 9818
rect 19722 9766 19724 9818
rect 19478 9764 19484 9766
rect 19540 9764 19564 9766
rect 19620 9764 19644 9766
rect 19700 9764 19724 9766
rect 19780 9764 19786 9766
rect 19478 9744 19786 9764
rect 19478 8732 19786 8752
rect 19478 8730 19484 8732
rect 19540 8730 19564 8732
rect 19620 8730 19644 8732
rect 19700 8730 19724 8732
rect 19780 8730 19786 8732
rect 19540 8678 19542 8730
rect 19722 8678 19724 8730
rect 19478 8676 19484 8678
rect 19540 8676 19564 8678
rect 19620 8676 19644 8678
rect 19700 8676 19724 8678
rect 19780 8676 19786 8678
rect 19478 8656 19786 8676
rect 19478 7644 19786 7664
rect 19478 7642 19484 7644
rect 19540 7642 19564 7644
rect 19620 7642 19644 7644
rect 19700 7642 19724 7644
rect 19780 7642 19786 7644
rect 19540 7590 19542 7642
rect 19722 7590 19724 7642
rect 19478 7588 19484 7590
rect 19540 7588 19564 7590
rect 19620 7588 19644 7590
rect 19700 7588 19724 7590
rect 19780 7588 19786 7590
rect 19478 7568 19786 7588
rect 19478 6556 19786 6576
rect 19478 6554 19484 6556
rect 19540 6554 19564 6556
rect 19620 6554 19644 6556
rect 19700 6554 19724 6556
rect 19780 6554 19786 6556
rect 19540 6502 19542 6554
rect 19722 6502 19724 6554
rect 19478 6500 19484 6502
rect 19540 6500 19564 6502
rect 19620 6500 19644 6502
rect 19700 6500 19724 6502
rect 19780 6500 19786 6502
rect 19478 6480 19786 6500
rect 19478 5468 19786 5488
rect 19478 5466 19484 5468
rect 19540 5466 19564 5468
rect 19620 5466 19644 5468
rect 19700 5466 19724 5468
rect 19780 5466 19786 5468
rect 19540 5414 19542 5466
rect 19722 5414 19724 5466
rect 19478 5412 19484 5414
rect 19540 5412 19564 5414
rect 19620 5412 19644 5414
rect 19700 5412 19724 5414
rect 19780 5412 19786 5414
rect 19478 5392 19786 5412
rect 17132 5092 17184 5098
rect 17132 5034 17184 5040
rect 17592 5092 17644 5098
rect 17592 5034 17644 5040
rect 17144 4690 17172 5034
rect 17132 4684 17184 4690
rect 17132 4626 17184 4632
rect 19478 4380 19786 4400
rect 19478 4378 19484 4380
rect 19540 4378 19564 4380
rect 19620 4378 19644 4380
rect 19700 4378 19724 4380
rect 19780 4378 19786 4380
rect 19540 4326 19542 4378
rect 19722 4326 19724 4378
rect 19478 4324 19484 4326
rect 19540 4324 19564 4326
rect 19620 4324 19644 4326
rect 19700 4324 19724 4326
rect 19780 4324 19786 4326
rect 19478 4304 19786 4324
rect 17684 4072 17736 4078
rect 17684 4014 17736 4020
rect 18052 4072 18104 4078
rect 18052 4014 18104 4020
rect 17408 4004 17460 4010
rect 17408 3946 17460 3952
rect 17420 3738 17448 3946
rect 17408 3732 17460 3738
rect 17408 3674 17460 3680
rect 16672 3664 16724 3670
rect 16672 3606 16724 3612
rect 17696 3126 17724 4014
rect 17960 4004 18012 4010
rect 17960 3946 18012 3952
rect 17684 3120 17736 3126
rect 17684 3062 17736 3068
rect 17972 2650 18000 3946
rect 16304 2644 16356 2650
rect 16304 2586 16356 2592
rect 17960 2644 18012 2650
rect 17960 2586 18012 2592
rect 16764 2372 16816 2378
rect 16764 2314 16816 2320
rect 16776 800 16804 2314
rect 18064 800 18092 4014
rect 19996 3670 20024 26982
rect 20076 26784 20128 26790
rect 20076 26726 20128 26732
rect 20088 26081 20116 26726
rect 20180 26586 20208 30126
rect 20272 30054 20300 30602
rect 20260 30048 20312 30054
rect 20260 29990 20312 29996
rect 20364 29866 20392 31622
rect 20272 29838 20392 29866
rect 20272 27946 20300 29838
rect 20352 29640 20404 29646
rect 20352 29582 20404 29588
rect 20260 27940 20312 27946
rect 20260 27882 20312 27888
rect 20272 26625 20300 27882
rect 20258 26616 20314 26625
rect 20168 26580 20220 26586
rect 20258 26551 20314 26560
rect 20168 26522 20220 26528
rect 20166 26480 20222 26489
rect 20166 26415 20222 26424
rect 20180 26382 20208 26415
rect 20168 26376 20220 26382
rect 20168 26318 20220 26324
rect 20074 26072 20130 26081
rect 20074 26007 20130 26016
rect 20074 25664 20130 25673
rect 20074 25599 20130 25608
rect 20088 23662 20116 25599
rect 20258 24848 20314 24857
rect 20258 24783 20314 24792
rect 20272 24342 20300 24783
rect 20260 24336 20312 24342
rect 20260 24278 20312 24284
rect 20260 23724 20312 23730
rect 20180 23684 20260 23712
rect 20076 23656 20128 23662
rect 20076 23598 20128 23604
rect 20076 23044 20128 23050
rect 20076 22986 20128 22992
rect 20088 22710 20116 22986
rect 20076 22704 20128 22710
rect 20076 22646 20128 22652
rect 20180 22506 20208 23684
rect 20260 23666 20312 23672
rect 20260 22636 20312 22642
rect 20260 22578 20312 22584
rect 20168 22500 20220 22506
rect 20168 22442 20220 22448
rect 20074 22128 20130 22137
rect 20074 22063 20076 22072
rect 20128 22063 20130 22072
rect 20076 22034 20128 22040
rect 20168 22024 20220 22030
rect 20168 21966 20220 21972
rect 20076 21956 20128 21962
rect 20076 21898 20128 21904
rect 20088 21486 20116 21898
rect 20076 21480 20128 21486
rect 20076 21422 20128 21428
rect 20180 21146 20208 21966
rect 20272 21622 20300 22578
rect 20364 21962 20392 29582
rect 20456 28121 20484 31844
rect 20824 31822 20852 31878
rect 20812 31816 20864 31822
rect 20534 31784 20590 31793
rect 20812 31758 20864 31764
rect 20534 31719 20590 31728
rect 20442 28112 20498 28121
rect 20442 28047 20498 28056
rect 20442 24848 20498 24857
rect 20442 24783 20498 24792
rect 20456 23730 20484 24783
rect 20444 23724 20496 23730
rect 20444 23666 20496 23672
rect 20444 22432 20496 22438
rect 20444 22374 20496 22380
rect 20456 22098 20484 22374
rect 20444 22092 20496 22098
rect 20444 22034 20496 22040
rect 20352 21956 20404 21962
rect 20352 21898 20404 21904
rect 20260 21616 20312 21622
rect 20260 21558 20312 21564
rect 20444 21616 20496 21622
rect 20444 21558 20496 21564
rect 20168 21140 20220 21146
rect 20168 21082 20220 21088
rect 20272 20942 20300 21558
rect 20352 21344 20404 21350
rect 20352 21286 20404 21292
rect 20260 20936 20312 20942
rect 20260 20878 20312 20884
rect 20272 20806 20300 20878
rect 20364 20874 20392 21286
rect 20352 20868 20404 20874
rect 20352 20810 20404 20816
rect 20076 20800 20128 20806
rect 20076 20742 20128 20748
rect 20260 20800 20312 20806
rect 20260 20742 20312 20748
rect 20088 19310 20116 20742
rect 20168 20256 20220 20262
rect 20168 20198 20220 20204
rect 20180 19854 20208 20198
rect 20168 19848 20220 19854
rect 20168 19790 20220 19796
rect 20272 19378 20300 20742
rect 20456 20262 20484 21558
rect 20548 20466 20576 31719
rect 20812 31680 20864 31686
rect 20812 31622 20864 31628
rect 20628 31136 20680 31142
rect 20628 31078 20680 31084
rect 20640 30190 20668 31078
rect 20720 30252 20772 30258
rect 20720 30194 20772 30200
rect 20628 30184 20680 30190
rect 20628 30126 20680 30132
rect 20732 29850 20760 30194
rect 20720 29844 20772 29850
rect 20720 29786 20772 29792
rect 20824 28914 20852 31622
rect 20916 30258 20944 32943
rect 21008 31754 21036 33374
rect 21088 33040 21140 33046
rect 21088 32982 21140 32988
rect 21100 32842 21128 32982
rect 21088 32836 21140 32842
rect 21088 32778 21140 32784
rect 21192 31754 21220 33510
rect 21284 33402 21312 34156
rect 21362 34096 21418 34105
rect 21362 34031 21418 34040
rect 21376 33561 21404 34031
rect 21362 33552 21418 33561
rect 21362 33487 21418 33496
rect 21284 33374 21404 33402
rect 21272 32904 21324 32910
rect 21272 32846 21324 32852
rect 21284 32434 21312 32846
rect 21272 32428 21324 32434
rect 21272 32370 21324 32376
rect 20996 31748 21048 31754
rect 21192 31726 21312 31754
rect 20996 31690 21048 31696
rect 21008 30394 21036 31690
rect 21088 31204 21140 31210
rect 21088 31146 21140 31152
rect 20996 30388 21048 30394
rect 20996 30330 21048 30336
rect 21100 30297 21128 31146
rect 21086 30288 21142 30297
rect 20904 30252 20956 30258
rect 21086 30223 21142 30232
rect 20904 30194 20956 30200
rect 21180 30184 21232 30190
rect 21180 30126 21232 30132
rect 20994 30016 21050 30025
rect 20994 29951 21050 29960
rect 20904 29844 20956 29850
rect 20904 29786 20956 29792
rect 20640 28886 20852 28914
rect 20640 28558 20668 28886
rect 20810 28792 20866 28801
rect 20810 28727 20866 28736
rect 20628 28552 20680 28558
rect 20628 28494 20680 28500
rect 20720 28552 20772 28558
rect 20720 28494 20772 28500
rect 20732 28257 20760 28494
rect 20824 28490 20852 28727
rect 20812 28484 20864 28490
rect 20812 28426 20864 28432
rect 20718 28248 20774 28257
rect 20718 28183 20774 28192
rect 20812 28008 20864 28014
rect 20718 27976 20774 27985
rect 20628 27940 20680 27946
rect 20812 27950 20864 27956
rect 20916 27962 20944 29786
rect 21008 28937 21036 29951
rect 21192 29850 21220 30126
rect 21180 29844 21232 29850
rect 21180 29786 21232 29792
rect 21180 28960 21232 28966
rect 20994 28928 21050 28937
rect 21180 28902 21232 28908
rect 20994 28863 21050 28872
rect 21192 28082 21220 28902
rect 21180 28076 21232 28082
rect 21180 28018 21232 28024
rect 20718 27911 20774 27920
rect 20628 27882 20680 27888
rect 20640 26926 20668 27882
rect 20732 27878 20760 27911
rect 20720 27872 20772 27878
rect 20720 27814 20772 27820
rect 20824 27402 20852 27950
rect 20916 27934 21036 27962
rect 20720 27396 20772 27402
rect 20720 27338 20772 27344
rect 20812 27396 20864 27402
rect 20812 27338 20864 27344
rect 20628 26920 20680 26926
rect 20628 26862 20680 26868
rect 20640 25294 20668 26862
rect 20628 25288 20680 25294
rect 20628 25230 20680 25236
rect 20628 24812 20680 24818
rect 20628 24754 20680 24760
rect 20640 24313 20668 24754
rect 20626 24304 20682 24313
rect 20626 24239 20682 24248
rect 20732 23322 20760 27338
rect 20812 26784 20864 26790
rect 20812 26726 20864 26732
rect 20824 26382 20852 26726
rect 20812 26376 20864 26382
rect 20812 26318 20864 26324
rect 20824 25906 20852 26318
rect 21008 26314 21036 27934
rect 21088 27396 21140 27402
rect 21088 27338 21140 27344
rect 20996 26308 21048 26314
rect 20996 26250 21048 26256
rect 20812 25900 20864 25906
rect 20812 25842 20864 25848
rect 20824 24818 20852 25842
rect 21008 25770 21036 26250
rect 21100 26246 21128 27338
rect 21192 26450 21220 28018
rect 21284 26790 21312 31726
rect 21376 31142 21404 33374
rect 21364 31136 21416 31142
rect 21364 31078 21416 31084
rect 21362 30424 21418 30433
rect 21362 30359 21418 30368
rect 21376 30122 21404 30359
rect 21364 30116 21416 30122
rect 21364 30058 21416 30064
rect 21364 28960 21416 28966
rect 21364 28902 21416 28908
rect 21376 28150 21404 28902
rect 21364 28144 21416 28150
rect 21364 28086 21416 28092
rect 21468 26976 21496 36722
rect 21560 36650 21588 38286
rect 21836 37874 21864 39743
rect 21824 37868 21876 37874
rect 21824 37810 21876 37816
rect 21640 37800 21692 37806
rect 21640 37742 21692 37748
rect 21548 36644 21600 36650
rect 21548 36586 21600 36592
rect 21546 36408 21602 36417
rect 21546 36343 21602 36352
rect 21560 36174 21588 36343
rect 21548 36168 21600 36174
rect 21548 36110 21600 36116
rect 21548 35760 21600 35766
rect 21546 35728 21548 35737
rect 21600 35728 21602 35737
rect 21546 35663 21602 35672
rect 21548 35488 21600 35494
rect 21548 35430 21600 35436
rect 21560 34610 21588 35430
rect 21548 34604 21600 34610
rect 21548 34546 21600 34552
rect 21548 34196 21600 34202
rect 21548 34138 21600 34144
rect 21560 30734 21588 34138
rect 21652 32502 21680 37742
rect 21928 37738 21956 41200
rect 22284 40452 22336 40458
rect 22284 40394 22336 40400
rect 22008 40384 22060 40390
rect 22008 40326 22060 40332
rect 22020 39506 22048 40326
rect 22192 39976 22244 39982
rect 22192 39918 22244 39924
rect 22204 39506 22232 39918
rect 22008 39500 22060 39506
rect 22008 39442 22060 39448
rect 22192 39500 22244 39506
rect 22192 39442 22244 39448
rect 22296 38962 22324 40394
rect 22284 38956 22336 38962
rect 22284 38898 22336 38904
rect 23216 38894 23244 41200
rect 23572 40860 23624 40866
rect 23572 40802 23624 40808
rect 23480 39840 23532 39846
rect 23480 39782 23532 39788
rect 23204 38888 23256 38894
rect 23204 38830 23256 38836
rect 22928 38412 22980 38418
rect 22928 38354 22980 38360
rect 22008 38276 22060 38282
rect 22008 38218 22060 38224
rect 22284 38276 22336 38282
rect 22284 38218 22336 38224
rect 22020 37806 22048 38218
rect 22008 37800 22060 37806
rect 22008 37742 22060 37748
rect 21732 37732 21784 37738
rect 21732 37674 21784 37680
rect 21916 37732 21968 37738
rect 21916 37674 21968 37680
rect 21744 32756 21772 37674
rect 22296 37233 22324 38218
rect 22940 38214 22968 38354
rect 22928 38208 22980 38214
rect 22928 38150 22980 38156
rect 23388 38004 23440 38010
rect 23388 37946 23440 37952
rect 22928 37664 22980 37670
rect 22928 37606 22980 37612
rect 22006 37224 22062 37233
rect 22006 37159 22008 37168
rect 22060 37159 22062 37168
rect 22282 37224 22338 37233
rect 22282 37159 22338 37168
rect 22560 37188 22612 37194
rect 22008 37130 22060 37136
rect 21914 36952 21970 36961
rect 21914 36887 21970 36896
rect 21928 36786 21956 36887
rect 22296 36802 22324 37159
rect 22560 37130 22612 37136
rect 22836 37188 22888 37194
rect 22836 37130 22888 37136
rect 22374 36952 22430 36961
rect 22572 36922 22600 37130
rect 22374 36887 22376 36896
rect 22428 36887 22430 36896
rect 22560 36916 22612 36922
rect 22376 36858 22428 36864
rect 22560 36858 22612 36864
rect 22652 36916 22704 36922
rect 22652 36858 22704 36864
rect 21916 36780 21968 36786
rect 22296 36774 22416 36802
rect 21916 36722 21968 36728
rect 21914 36680 21970 36689
rect 21824 36644 21876 36650
rect 21914 36615 21970 36624
rect 21824 36586 21876 36592
rect 21836 36310 21864 36586
rect 21824 36304 21876 36310
rect 21824 36246 21876 36252
rect 21928 36174 21956 36615
rect 22008 36304 22060 36310
rect 22008 36246 22060 36252
rect 21916 36168 21968 36174
rect 21916 36110 21968 36116
rect 21822 36000 21878 36009
rect 21822 35935 21878 35944
rect 21836 34898 21864 35935
rect 21928 35698 21956 36110
rect 21916 35692 21968 35698
rect 21916 35634 21968 35640
rect 21928 35329 21956 35634
rect 22020 35562 22048 36246
rect 22284 36168 22336 36174
rect 22284 36110 22336 36116
rect 22296 35873 22324 36110
rect 22282 35864 22338 35873
rect 22100 35828 22152 35834
rect 22282 35799 22338 35808
rect 22100 35770 22152 35776
rect 22008 35556 22060 35562
rect 22008 35498 22060 35504
rect 21914 35320 21970 35329
rect 21914 35255 21970 35264
rect 21928 35086 21956 35255
rect 21916 35080 21968 35086
rect 21916 35022 21968 35028
rect 22112 34898 22140 35770
rect 22296 35698 22324 35799
rect 22284 35692 22336 35698
rect 22284 35634 22336 35640
rect 22296 35136 22324 35634
rect 22388 35290 22416 36774
rect 22664 36174 22692 36858
rect 22848 36281 22876 37130
rect 22834 36272 22890 36281
rect 22940 36258 22968 37606
rect 23112 37120 23164 37126
rect 23112 37062 23164 37068
rect 23020 36780 23072 36786
rect 23020 36722 23072 36728
rect 23032 36378 23060 36722
rect 23124 36718 23152 37062
rect 23296 36848 23348 36854
rect 23296 36790 23348 36796
rect 23112 36712 23164 36718
rect 23112 36654 23164 36660
rect 23020 36372 23072 36378
rect 23020 36314 23072 36320
rect 22940 36230 23060 36258
rect 22834 36207 22890 36216
rect 22848 36174 22876 36207
rect 22652 36168 22704 36174
rect 22652 36110 22704 36116
rect 22836 36168 22888 36174
rect 22836 36110 22888 36116
rect 22560 36100 22612 36106
rect 22560 36042 22612 36048
rect 22572 35630 22600 36042
rect 22744 36032 22796 36038
rect 22744 35974 22796 35980
rect 22650 35728 22706 35737
rect 22756 35698 22784 35974
rect 22650 35663 22706 35672
rect 22744 35692 22796 35698
rect 22560 35624 22612 35630
rect 22560 35566 22612 35572
rect 22664 35578 22692 35663
rect 22744 35634 22796 35640
rect 22468 35556 22520 35562
rect 22664 35550 22784 35578
rect 22468 35498 22520 35504
rect 22376 35284 22428 35290
rect 22376 35226 22428 35232
rect 22296 35108 22416 35136
rect 22282 35048 22338 35057
rect 22388 35018 22416 35108
rect 22282 34983 22338 34992
rect 22376 35012 22428 35018
rect 21836 34870 21956 34898
rect 22112 34870 22232 34898
rect 21824 34604 21876 34610
rect 21824 34546 21876 34552
rect 21836 34066 21864 34546
rect 21928 34202 21956 34870
rect 22204 34649 22232 34870
rect 22190 34640 22246 34649
rect 22008 34604 22060 34610
rect 22190 34575 22246 34584
rect 22008 34546 22060 34552
rect 22020 34406 22048 34546
rect 22008 34400 22060 34406
rect 22008 34342 22060 34348
rect 21916 34196 21968 34202
rect 21916 34138 21968 34144
rect 21824 34060 21876 34066
rect 21824 34002 21876 34008
rect 22192 33992 22244 33998
rect 22192 33934 22244 33940
rect 22204 33522 22232 33934
rect 22008 33516 22060 33522
rect 22008 33458 22060 33464
rect 22192 33516 22244 33522
rect 22192 33458 22244 33464
rect 22020 33318 22048 33458
rect 21824 33312 21876 33318
rect 21824 33254 21876 33260
rect 22008 33312 22060 33318
rect 22008 33254 22060 33260
rect 21836 32910 21864 33254
rect 21824 32904 21876 32910
rect 21824 32846 21876 32852
rect 21916 32904 21968 32910
rect 21916 32846 21968 32852
rect 21744 32728 21864 32756
rect 21640 32496 21692 32502
rect 21692 32444 21772 32450
rect 21640 32438 21772 32444
rect 21652 32422 21772 32438
rect 21744 31754 21772 32422
rect 21652 31726 21772 31754
rect 21548 30728 21600 30734
rect 21548 30670 21600 30676
rect 21548 29776 21600 29782
rect 21546 29744 21548 29753
rect 21600 29744 21602 29753
rect 21546 29679 21602 29688
rect 21546 29336 21602 29345
rect 21546 29271 21548 29280
rect 21600 29271 21602 29280
rect 21548 29242 21600 29248
rect 21548 28688 21600 28694
rect 21548 28630 21600 28636
rect 21560 28082 21588 28630
rect 21548 28076 21600 28082
rect 21548 28018 21600 28024
rect 21376 26948 21496 26976
rect 21272 26784 21324 26790
rect 21272 26726 21324 26732
rect 21180 26444 21232 26450
rect 21180 26386 21232 26392
rect 21088 26240 21140 26246
rect 21088 26182 21140 26188
rect 21100 25945 21128 26182
rect 21086 25936 21142 25945
rect 21086 25871 21142 25880
rect 20996 25764 21048 25770
rect 20996 25706 21048 25712
rect 21100 25498 21128 25871
rect 21088 25492 21140 25498
rect 21088 25434 21140 25440
rect 21192 25378 21220 26386
rect 21008 25350 21220 25378
rect 20812 24812 20864 24818
rect 20812 24754 20864 24760
rect 20812 24676 20864 24682
rect 20812 24618 20864 24624
rect 20824 24313 20852 24618
rect 21008 24585 21036 25350
rect 21376 24818 21404 26948
rect 21652 26874 21680 31726
rect 21732 29708 21784 29714
rect 21732 29650 21784 29656
rect 21744 29617 21772 29650
rect 21730 29608 21786 29617
rect 21730 29543 21786 29552
rect 21732 29300 21784 29306
rect 21732 29242 21784 29248
rect 21744 29102 21772 29242
rect 21732 29096 21784 29102
rect 21732 29038 21784 29044
rect 21732 28688 21784 28694
rect 21836 28642 21864 32728
rect 21928 32434 21956 32846
rect 22098 32600 22154 32609
rect 22098 32535 22154 32544
rect 21916 32428 21968 32434
rect 21916 32370 21968 32376
rect 22112 32337 22140 32535
rect 22098 32328 22154 32337
rect 22098 32263 22154 32272
rect 21916 31748 21968 31754
rect 21916 31690 21968 31696
rect 21928 31210 21956 31690
rect 22296 31482 22324 34983
rect 22376 34954 22428 34960
rect 22480 34134 22508 35498
rect 22756 35494 22784 35550
rect 22652 35488 22704 35494
rect 22652 35430 22704 35436
rect 22744 35488 22796 35494
rect 22744 35430 22796 35436
rect 22560 35284 22612 35290
rect 22560 35226 22612 35232
rect 22572 34406 22600 35226
rect 22664 35086 22692 35430
rect 22756 35154 22784 35430
rect 22836 35284 22888 35290
rect 22836 35226 22888 35232
rect 22744 35148 22796 35154
rect 22744 35090 22796 35096
rect 22652 35080 22704 35086
rect 22652 35022 22704 35028
rect 22560 34400 22612 34406
rect 22560 34342 22612 34348
rect 22468 34128 22520 34134
rect 22468 34070 22520 34076
rect 22468 33516 22520 33522
rect 22468 33458 22520 33464
rect 22480 33153 22508 33458
rect 22560 33448 22612 33454
rect 22560 33390 22612 33396
rect 22466 33144 22522 33153
rect 22466 33079 22522 33088
rect 22572 32881 22600 33390
rect 22664 33318 22692 35022
rect 22848 34950 22876 35226
rect 22928 35080 22980 35086
rect 22926 35048 22928 35057
rect 22980 35048 22982 35057
rect 22926 34983 22982 34992
rect 22836 34944 22888 34950
rect 22836 34886 22888 34892
rect 22744 34740 22796 34746
rect 22744 34682 22796 34688
rect 22756 33998 22784 34682
rect 22848 34610 22876 34886
rect 22928 34672 22980 34678
rect 22928 34614 22980 34620
rect 22836 34604 22888 34610
rect 22836 34546 22888 34552
rect 22940 34490 22968 34614
rect 22848 34462 22968 34490
rect 22744 33992 22796 33998
rect 22744 33934 22796 33940
rect 22848 33454 22876 34462
rect 22928 33856 22980 33862
rect 22928 33798 22980 33804
rect 22836 33448 22888 33454
rect 22836 33390 22888 33396
rect 22652 33312 22704 33318
rect 22652 33254 22704 33260
rect 22664 33046 22692 33254
rect 22652 33040 22704 33046
rect 22652 32982 22704 32988
rect 22558 32872 22614 32881
rect 22558 32807 22614 32816
rect 22560 31816 22612 31822
rect 22560 31758 22612 31764
rect 22284 31476 22336 31482
rect 22284 31418 22336 31424
rect 21916 31204 21968 31210
rect 21916 31146 21968 31152
rect 22376 31136 22428 31142
rect 22376 31078 22428 31084
rect 22100 30252 22152 30258
rect 22020 30212 22100 30240
rect 21916 29708 21968 29714
rect 21916 29650 21968 29656
rect 21928 29073 21956 29650
rect 22020 29170 22048 30212
rect 22100 30194 22152 30200
rect 22100 29844 22152 29850
rect 22100 29786 22152 29792
rect 22112 29481 22140 29786
rect 22284 29776 22336 29782
rect 22190 29744 22246 29753
rect 22284 29718 22336 29724
rect 22190 29679 22246 29688
rect 22098 29472 22154 29481
rect 22098 29407 22154 29416
rect 22100 29232 22152 29238
rect 22100 29174 22152 29180
rect 22008 29164 22060 29170
rect 22008 29106 22060 29112
rect 22112 29073 22140 29174
rect 21914 29064 21970 29073
rect 21914 28999 21970 29008
rect 22098 29064 22154 29073
rect 22098 28999 22154 29008
rect 21916 28960 21968 28966
rect 21968 28908 22048 28914
rect 21916 28902 22048 28908
rect 21928 28886 22048 28902
rect 22020 28762 22048 28886
rect 22008 28756 22060 28762
rect 22008 28698 22060 28704
rect 21784 28636 21864 28642
rect 21732 28630 21864 28636
rect 21744 28614 21864 28630
rect 21732 28552 21784 28558
rect 21732 28494 21784 28500
rect 21836 28506 21864 28614
rect 22098 28520 22154 28529
rect 21744 27946 21772 28494
rect 21836 28478 22098 28506
rect 22098 28455 22154 28464
rect 22204 28422 22232 29679
rect 22296 29170 22324 29718
rect 22388 29646 22416 31078
rect 22466 30696 22522 30705
rect 22466 30631 22468 30640
rect 22520 30631 22522 30640
rect 22468 30602 22520 30608
rect 22376 29640 22428 29646
rect 22376 29582 22428 29588
rect 22284 29164 22336 29170
rect 22284 29106 22336 29112
rect 22284 28960 22336 28966
rect 22284 28902 22336 28908
rect 22192 28416 22244 28422
rect 22192 28358 22244 28364
rect 21914 28112 21970 28121
rect 21914 28047 21970 28056
rect 21732 27940 21784 27946
rect 21732 27882 21784 27888
rect 21824 27872 21876 27878
rect 21730 27840 21786 27849
rect 21824 27814 21876 27820
rect 21730 27775 21786 27784
rect 21744 27674 21772 27775
rect 21732 27668 21784 27674
rect 21732 27610 21784 27616
rect 21730 27568 21786 27577
rect 21730 27503 21786 27512
rect 21744 26994 21772 27503
rect 21836 26994 21864 27814
rect 21928 27538 21956 28047
rect 22296 27985 22324 28902
rect 22376 28144 22428 28150
rect 22376 28086 22428 28092
rect 22282 27976 22338 27985
rect 22282 27911 22338 27920
rect 22190 27840 22246 27849
rect 22190 27775 22246 27784
rect 22006 27704 22062 27713
rect 22006 27639 22008 27648
rect 22060 27639 22062 27648
rect 22008 27610 22060 27616
rect 22204 27554 22232 27775
rect 22296 27656 22324 27911
rect 22388 27878 22416 28086
rect 22376 27872 22428 27878
rect 22572 27849 22600 31758
rect 22848 31634 22876 33390
rect 22940 32434 22968 33798
rect 22928 32428 22980 32434
rect 22928 32370 22980 32376
rect 22928 31748 22980 31754
rect 22928 31690 22980 31696
rect 22756 31606 22876 31634
rect 22652 30932 22704 30938
rect 22652 30874 22704 30880
rect 22664 29170 22692 30874
rect 22652 29164 22704 29170
rect 22652 29106 22704 29112
rect 22376 27814 22428 27820
rect 22558 27840 22614 27849
rect 22558 27775 22614 27784
rect 22296 27628 22600 27656
rect 21916 27532 21968 27538
rect 22204 27526 22508 27554
rect 21916 27474 21968 27480
rect 22284 27464 22336 27470
rect 22284 27406 22336 27412
rect 22376 27464 22428 27470
rect 22376 27406 22428 27412
rect 22192 27328 22244 27334
rect 22192 27270 22244 27276
rect 22204 27062 22232 27270
rect 22192 27056 22244 27062
rect 22192 26998 22244 27004
rect 21732 26988 21784 26994
rect 21732 26930 21784 26936
rect 21824 26988 21876 26994
rect 21824 26930 21876 26936
rect 22100 26988 22152 26994
rect 22100 26930 22152 26936
rect 21468 26846 21680 26874
rect 21364 24812 21416 24818
rect 21192 24772 21364 24800
rect 21088 24676 21140 24682
rect 21088 24618 21140 24624
rect 20994 24576 21050 24585
rect 20994 24511 21050 24520
rect 20810 24304 20866 24313
rect 20810 24239 20866 24248
rect 21100 23730 21128 24618
rect 21088 23724 21140 23730
rect 21088 23666 21140 23672
rect 20628 23316 20680 23322
rect 20628 23258 20680 23264
rect 20720 23316 20772 23322
rect 20720 23258 20772 23264
rect 20640 23118 20668 23258
rect 20810 23216 20866 23225
rect 20810 23151 20866 23160
rect 20628 23112 20680 23118
rect 20628 23054 20680 23060
rect 20824 22438 20852 23151
rect 21100 23089 21128 23666
rect 21086 23080 21142 23089
rect 21086 23015 21142 23024
rect 20904 22976 20956 22982
rect 20904 22918 20956 22924
rect 20916 22574 20944 22918
rect 20994 22672 21050 22681
rect 20994 22607 20996 22616
rect 21048 22607 21050 22616
rect 20996 22578 21048 22584
rect 20904 22568 20956 22574
rect 20904 22510 20956 22516
rect 20812 22432 20864 22438
rect 20812 22374 20864 22380
rect 20720 21480 20772 21486
rect 20720 21422 20772 21428
rect 20628 21344 20680 21350
rect 20628 21286 20680 21292
rect 20536 20460 20588 20466
rect 20536 20402 20588 20408
rect 20640 20398 20668 21286
rect 20628 20392 20680 20398
rect 20628 20334 20680 20340
rect 20444 20256 20496 20262
rect 20444 20198 20496 20204
rect 20260 19372 20312 19378
rect 20260 19314 20312 19320
rect 20076 19304 20128 19310
rect 20076 19246 20128 19252
rect 20168 18692 20220 18698
rect 20168 18634 20220 18640
rect 20076 18284 20128 18290
rect 20076 18226 20128 18232
rect 20088 16250 20116 18226
rect 20076 16244 20128 16250
rect 20076 16186 20128 16192
rect 20180 16114 20208 18634
rect 20456 18630 20484 20198
rect 20640 19718 20668 20334
rect 20628 19712 20680 19718
rect 20628 19654 20680 19660
rect 20732 19334 20760 21422
rect 20824 21350 20852 22374
rect 20916 22012 20944 22510
rect 21008 22166 21036 22578
rect 20996 22160 21048 22166
rect 20996 22102 21048 22108
rect 20996 22024 21048 22030
rect 20916 21984 20996 22012
rect 20996 21966 21048 21972
rect 21100 21486 21128 23015
rect 21088 21480 21140 21486
rect 21088 21422 21140 21428
rect 20812 21344 20864 21350
rect 20812 21286 20864 21292
rect 20904 20868 20956 20874
rect 20904 20810 20956 20816
rect 20812 19508 20864 19514
rect 20812 19450 20864 19456
rect 20548 19306 20760 19334
rect 20260 18624 20312 18630
rect 20444 18624 20496 18630
rect 20260 18566 20312 18572
rect 20364 18584 20444 18612
rect 20272 17814 20300 18566
rect 20260 17808 20312 17814
rect 20260 17750 20312 17756
rect 20364 16114 20392 18584
rect 20444 18566 20496 18572
rect 20444 17196 20496 17202
rect 20444 17138 20496 17144
rect 20456 16794 20484 17138
rect 20444 16788 20496 16794
rect 20444 16730 20496 16736
rect 20548 16182 20576 19306
rect 20720 18964 20772 18970
rect 20720 18906 20772 18912
rect 20628 18760 20680 18766
rect 20628 18702 20680 18708
rect 20640 18426 20668 18702
rect 20628 18420 20680 18426
rect 20628 18362 20680 18368
rect 20732 18034 20760 18906
rect 20640 18006 20760 18034
rect 20536 16176 20588 16182
rect 20536 16118 20588 16124
rect 20168 16108 20220 16114
rect 20168 16050 20220 16056
rect 20352 16108 20404 16114
rect 20352 16050 20404 16056
rect 20640 13870 20668 18006
rect 20720 17876 20772 17882
rect 20720 17818 20772 17824
rect 20732 16658 20760 17818
rect 20720 16652 20772 16658
rect 20720 16594 20772 16600
rect 20824 16114 20852 19450
rect 20916 16250 20944 20810
rect 21088 20460 21140 20466
rect 21088 20402 21140 20408
rect 20996 19780 21048 19786
rect 20996 19722 21048 19728
rect 21008 19310 21036 19722
rect 20996 19304 21048 19310
rect 20996 19246 21048 19252
rect 20996 18760 21048 18766
rect 20996 18702 21048 18708
rect 21008 17882 21036 18702
rect 20996 17876 21048 17882
rect 20996 17818 21048 17824
rect 20996 17672 21048 17678
rect 20996 17614 21048 17620
rect 21008 17270 21036 17614
rect 20996 17264 21048 17270
rect 20996 17206 21048 17212
rect 20904 16244 20956 16250
rect 20904 16186 20956 16192
rect 20812 16108 20864 16114
rect 20812 16050 20864 16056
rect 20628 13864 20680 13870
rect 20628 13806 20680 13812
rect 21100 12434 21128 20402
rect 21192 18970 21220 24772
rect 21364 24754 21416 24760
rect 21364 23112 21416 23118
rect 21364 23054 21416 23060
rect 21376 22098 21404 23054
rect 21364 22092 21416 22098
rect 21364 22034 21416 22040
rect 21376 22001 21404 22034
rect 21362 21992 21418 22001
rect 21362 21927 21418 21936
rect 21364 21888 21416 21894
rect 21364 21830 21416 21836
rect 21376 21690 21404 21830
rect 21364 21684 21416 21690
rect 21364 21626 21416 21632
rect 21272 21616 21324 21622
rect 21272 21558 21324 21564
rect 21284 20942 21312 21558
rect 21364 21344 21416 21350
rect 21364 21286 21416 21292
rect 21272 20936 21324 20942
rect 21272 20878 21324 20884
rect 21284 19922 21312 20878
rect 21272 19916 21324 19922
rect 21272 19858 21324 19864
rect 21180 18964 21232 18970
rect 21180 18906 21232 18912
rect 21180 18828 21232 18834
rect 21180 18770 21232 18776
rect 21192 16726 21220 18770
rect 21180 16720 21232 16726
rect 21180 16662 21232 16668
rect 21376 16114 21404 21286
rect 21468 18086 21496 26846
rect 21548 26784 21600 26790
rect 21640 26784 21692 26790
rect 21548 26726 21600 26732
rect 21638 26752 21640 26761
rect 21692 26752 21694 26761
rect 21560 20262 21588 26726
rect 21638 26687 21694 26696
rect 21836 25974 21864 26930
rect 22008 26852 22060 26858
rect 22008 26794 22060 26800
rect 21824 25968 21876 25974
rect 21824 25910 21876 25916
rect 22020 25906 22048 26794
rect 22112 25906 22140 26930
rect 22192 26784 22244 26790
rect 22192 26726 22244 26732
rect 22204 26042 22232 26726
rect 22296 26586 22324 27406
rect 22388 27130 22416 27406
rect 22376 27124 22428 27130
rect 22376 27066 22428 27072
rect 22376 26988 22428 26994
rect 22376 26930 22428 26936
rect 22284 26580 22336 26586
rect 22284 26522 22336 26528
rect 22192 26036 22244 26042
rect 22192 25978 22244 25984
rect 22008 25900 22060 25906
rect 22008 25842 22060 25848
rect 22100 25900 22152 25906
rect 22100 25842 22152 25848
rect 21640 25832 21692 25838
rect 21640 25774 21692 25780
rect 21652 25498 21680 25774
rect 21640 25492 21692 25498
rect 21640 25434 21692 25440
rect 21638 24984 21694 24993
rect 21638 24919 21694 24928
rect 21652 24750 21680 24919
rect 21640 24744 21692 24750
rect 21640 24686 21692 24692
rect 21824 24132 21876 24138
rect 21824 24074 21876 24080
rect 21640 24064 21692 24070
rect 21640 24006 21692 24012
rect 21652 23866 21680 24006
rect 21836 23866 21864 24074
rect 21640 23860 21692 23866
rect 21640 23802 21692 23808
rect 21824 23860 21876 23866
rect 21824 23802 21876 23808
rect 21914 23760 21970 23769
rect 21732 23724 21784 23730
rect 22020 23730 22048 25842
rect 22112 25294 22140 25842
rect 22204 25838 22232 25978
rect 22192 25832 22244 25838
rect 22192 25774 22244 25780
rect 22296 25430 22324 26522
rect 22388 26246 22416 26930
rect 22376 26240 22428 26246
rect 22376 26182 22428 26188
rect 22388 25906 22416 26182
rect 22376 25900 22428 25906
rect 22376 25842 22428 25848
rect 22284 25424 22336 25430
rect 22284 25366 22336 25372
rect 22388 25294 22416 25842
rect 22480 25809 22508 27526
rect 22572 27334 22600 27628
rect 22652 27396 22704 27402
rect 22652 27338 22704 27344
rect 22560 27328 22612 27334
rect 22560 27270 22612 27276
rect 22560 26988 22612 26994
rect 22560 26930 22612 26936
rect 22466 25800 22522 25809
rect 22466 25735 22522 25744
rect 22468 25696 22520 25702
rect 22468 25638 22520 25644
rect 22100 25288 22152 25294
rect 22100 25230 22152 25236
rect 22376 25288 22428 25294
rect 22376 25230 22428 25236
rect 22112 24954 22140 25230
rect 22480 25106 22508 25638
rect 22572 25294 22600 26930
rect 22664 25838 22692 27338
rect 22756 26382 22784 31606
rect 22940 31414 22968 31690
rect 22928 31408 22980 31414
rect 22928 31350 22980 31356
rect 22836 31136 22888 31142
rect 22836 31078 22888 31084
rect 22848 29714 22876 31078
rect 22928 30728 22980 30734
rect 22928 30670 22980 30676
rect 22940 30394 22968 30670
rect 22928 30388 22980 30394
rect 22928 30330 22980 30336
rect 22940 30258 22968 30330
rect 22928 30252 22980 30258
rect 22928 30194 22980 30200
rect 22836 29708 22888 29714
rect 22836 29650 22888 29656
rect 22928 29164 22980 29170
rect 22928 29106 22980 29112
rect 22836 29096 22888 29102
rect 22836 29038 22888 29044
rect 22848 28966 22876 29038
rect 22940 28966 22968 29106
rect 22836 28960 22888 28966
rect 22836 28902 22888 28908
rect 22928 28960 22980 28966
rect 22928 28902 22980 28908
rect 22834 28520 22890 28529
rect 22834 28455 22890 28464
rect 22928 28484 22980 28490
rect 22744 26376 22796 26382
rect 22744 26318 22796 26324
rect 22848 26194 22876 28455
rect 22928 28426 22980 28432
rect 22756 26166 22876 26194
rect 22652 25832 22704 25838
rect 22652 25774 22704 25780
rect 22560 25288 22612 25294
rect 22560 25230 22612 25236
rect 22388 25078 22508 25106
rect 22100 24948 22152 24954
rect 22100 24890 22152 24896
rect 22284 24948 22336 24954
rect 22284 24890 22336 24896
rect 22192 24676 22244 24682
rect 22192 24618 22244 24624
rect 22204 24177 22232 24618
rect 22296 24410 22324 24890
rect 22388 24818 22416 25078
rect 22376 24812 22428 24818
rect 22376 24754 22428 24760
rect 22284 24404 22336 24410
rect 22284 24346 22336 24352
rect 22284 24268 22336 24274
rect 22284 24210 22336 24216
rect 22190 24168 22246 24177
rect 22190 24103 22246 24112
rect 22296 24070 22324 24210
rect 22284 24064 22336 24070
rect 22284 24006 22336 24012
rect 22100 23860 22152 23866
rect 22100 23802 22152 23808
rect 21914 23695 21970 23704
rect 22008 23724 22060 23730
rect 21732 23666 21784 23672
rect 21638 23352 21694 23361
rect 21638 23287 21694 23296
rect 21652 22778 21680 23287
rect 21640 22772 21692 22778
rect 21640 22714 21692 22720
rect 21744 22658 21772 23666
rect 21824 23044 21876 23050
rect 21824 22986 21876 22992
rect 21836 22778 21864 22986
rect 21824 22772 21876 22778
rect 21824 22714 21876 22720
rect 21652 22630 21772 22658
rect 21548 20256 21600 20262
rect 21548 20198 21600 20204
rect 21652 20058 21680 22630
rect 21928 22080 21956 23695
rect 22008 23666 22060 23672
rect 22112 23118 22140 23802
rect 22284 23724 22336 23730
rect 22204 23684 22284 23712
rect 22204 23254 22232 23684
rect 22284 23666 22336 23672
rect 22388 23633 22416 24754
rect 22572 24410 22600 25230
rect 22652 25152 22704 25158
rect 22652 25094 22704 25100
rect 22664 24818 22692 25094
rect 22652 24812 22704 24818
rect 22652 24754 22704 24760
rect 22560 24404 22612 24410
rect 22560 24346 22612 24352
rect 22652 24200 22704 24206
rect 22652 24142 22704 24148
rect 22756 24154 22784 26166
rect 22836 25832 22888 25838
rect 22836 25774 22888 25780
rect 22848 24818 22876 25774
rect 22940 25770 22968 28426
rect 23032 26874 23060 36230
rect 23204 36168 23256 36174
rect 23204 36110 23256 36116
rect 23110 35592 23166 35601
rect 23110 35527 23166 35536
rect 23124 34542 23152 35527
rect 23112 34536 23164 34542
rect 23112 34478 23164 34484
rect 23112 34400 23164 34406
rect 23216 34377 23244 36110
rect 23112 34342 23164 34348
rect 23202 34368 23258 34377
rect 23124 33862 23152 34342
rect 23202 34303 23258 34312
rect 23308 34134 23336 36790
rect 23400 36718 23428 37946
rect 23492 37330 23520 39782
rect 23480 37324 23532 37330
rect 23480 37266 23532 37272
rect 23480 36780 23532 36786
rect 23480 36722 23532 36728
rect 23388 36712 23440 36718
rect 23388 36654 23440 36660
rect 23386 36272 23442 36281
rect 23386 36207 23388 36216
rect 23440 36207 23442 36216
rect 23388 36178 23440 36184
rect 23388 35556 23440 35562
rect 23388 35498 23440 35504
rect 23400 34950 23428 35498
rect 23492 35494 23520 36722
rect 23584 36378 23612 40802
rect 23664 40316 23716 40322
rect 23664 40258 23716 40264
rect 23676 38962 23704 40258
rect 23860 39506 23888 41200
rect 23940 40588 23992 40594
rect 23940 40530 23992 40536
rect 23848 39500 23900 39506
rect 23848 39442 23900 39448
rect 23664 38956 23716 38962
rect 23664 38898 23716 38904
rect 23664 38548 23716 38554
rect 23664 38490 23716 38496
rect 23676 38350 23704 38490
rect 23848 38412 23900 38418
rect 23848 38354 23900 38360
rect 23664 38344 23716 38350
rect 23860 38321 23888 38354
rect 23664 38286 23716 38292
rect 23846 38312 23902 38321
rect 23756 38276 23808 38282
rect 23846 38247 23902 38256
rect 23756 38218 23808 38224
rect 23664 37120 23716 37126
rect 23662 37088 23664 37097
rect 23716 37088 23718 37097
rect 23662 37023 23718 37032
rect 23664 36712 23716 36718
rect 23664 36654 23716 36660
rect 23572 36372 23624 36378
rect 23572 36314 23624 36320
rect 23572 35624 23624 35630
rect 23572 35566 23624 35572
rect 23480 35488 23532 35494
rect 23480 35430 23532 35436
rect 23388 34944 23440 34950
rect 23388 34886 23440 34892
rect 23584 34728 23612 35566
rect 23676 34746 23704 36654
rect 23768 36242 23796 38218
rect 23848 38208 23900 38214
rect 23848 38150 23900 38156
rect 23860 37806 23888 38150
rect 23848 37800 23900 37806
rect 23848 37742 23900 37748
rect 23848 37324 23900 37330
rect 23848 37266 23900 37272
rect 23756 36236 23808 36242
rect 23756 36178 23808 36184
rect 23756 36032 23808 36038
rect 23756 35974 23808 35980
rect 23768 35698 23796 35974
rect 23860 35834 23888 37266
rect 23848 35828 23900 35834
rect 23848 35770 23900 35776
rect 23756 35692 23808 35698
rect 23756 35634 23808 35640
rect 23756 35488 23808 35494
rect 23756 35430 23808 35436
rect 23848 35488 23900 35494
rect 23848 35430 23900 35436
rect 23492 34700 23612 34728
rect 23664 34740 23716 34746
rect 23386 34232 23442 34241
rect 23386 34167 23442 34176
rect 23296 34128 23348 34134
rect 23296 34070 23348 34076
rect 23112 33856 23164 33862
rect 23112 33798 23164 33804
rect 23308 33590 23336 34070
rect 23400 34066 23428 34167
rect 23388 34060 23440 34066
rect 23388 34002 23440 34008
rect 23296 33584 23348 33590
rect 23296 33526 23348 33532
rect 23400 33130 23428 34002
rect 23492 33289 23520 34700
rect 23664 34682 23716 34688
rect 23572 34604 23624 34610
rect 23572 34546 23624 34552
rect 23584 33504 23612 34546
rect 23662 34368 23718 34377
rect 23662 34303 23718 34312
rect 23676 34202 23704 34303
rect 23664 34196 23716 34202
rect 23664 34138 23716 34144
rect 23768 34134 23796 35430
rect 23756 34128 23808 34134
rect 23756 34070 23808 34076
rect 23860 33522 23888 35430
rect 23952 34066 23980 40530
rect 26884 40520 26936 40526
rect 26884 40462 26936 40468
rect 26332 40248 26384 40254
rect 26332 40190 26384 40196
rect 24768 40180 24820 40186
rect 24768 40122 24820 40128
rect 24110 39740 24418 39760
rect 24110 39738 24116 39740
rect 24172 39738 24196 39740
rect 24252 39738 24276 39740
rect 24332 39738 24356 39740
rect 24412 39738 24418 39740
rect 24172 39686 24174 39738
rect 24354 39686 24356 39738
rect 24110 39684 24116 39686
rect 24172 39684 24196 39686
rect 24252 39684 24276 39686
rect 24332 39684 24356 39686
rect 24412 39684 24418 39686
rect 24110 39664 24418 39684
rect 24780 39506 24808 40122
rect 24768 39500 24820 39506
rect 24768 39442 24820 39448
rect 26056 39500 26108 39506
rect 26056 39442 26108 39448
rect 24584 39432 24636 39438
rect 24582 39400 24584 39409
rect 24636 39400 24638 39409
rect 24582 39335 24638 39344
rect 24030 39264 24086 39273
rect 24030 39199 24086 39208
rect 24044 35086 24072 39199
rect 24490 39128 24546 39137
rect 24490 39063 24546 39072
rect 24110 38652 24418 38672
rect 24110 38650 24116 38652
rect 24172 38650 24196 38652
rect 24252 38650 24276 38652
rect 24332 38650 24356 38652
rect 24412 38650 24418 38652
rect 24172 38598 24174 38650
rect 24354 38598 24356 38650
rect 24110 38596 24116 38598
rect 24172 38596 24196 38598
rect 24252 38596 24276 38598
rect 24332 38596 24356 38598
rect 24412 38596 24418 38598
rect 24110 38576 24418 38596
rect 24504 37754 24532 39063
rect 25964 38888 26016 38894
rect 25964 38830 26016 38836
rect 24582 38448 24638 38457
rect 24582 38383 24638 38392
rect 24596 37874 24624 38383
rect 24860 38344 24912 38350
rect 24860 38286 24912 38292
rect 25044 38344 25096 38350
rect 25044 38286 25096 38292
rect 25596 38344 25648 38350
rect 25872 38344 25924 38350
rect 25596 38286 25648 38292
rect 25870 38312 25872 38321
rect 25924 38312 25926 38321
rect 24676 38208 24728 38214
rect 24676 38150 24728 38156
rect 24768 38208 24820 38214
rect 24768 38150 24820 38156
rect 24584 37868 24636 37874
rect 24584 37810 24636 37816
rect 24504 37726 24624 37754
rect 24110 37564 24418 37584
rect 24110 37562 24116 37564
rect 24172 37562 24196 37564
rect 24252 37562 24276 37564
rect 24332 37562 24356 37564
rect 24412 37562 24418 37564
rect 24172 37510 24174 37562
rect 24354 37510 24356 37562
rect 24110 37508 24116 37510
rect 24172 37508 24196 37510
rect 24252 37508 24276 37510
rect 24332 37508 24356 37510
rect 24412 37508 24418 37510
rect 24110 37488 24418 37508
rect 24492 37256 24544 37262
rect 24492 37198 24544 37204
rect 24122 36952 24178 36961
rect 24122 36887 24124 36896
rect 24176 36887 24178 36896
rect 24124 36858 24176 36864
rect 24124 36780 24176 36786
rect 24124 36722 24176 36728
rect 24136 36689 24164 36722
rect 24122 36680 24178 36689
rect 24122 36615 24178 36624
rect 24110 36476 24418 36496
rect 24110 36474 24116 36476
rect 24172 36474 24196 36476
rect 24252 36474 24276 36476
rect 24332 36474 24356 36476
rect 24412 36474 24418 36476
rect 24172 36422 24174 36474
rect 24354 36422 24356 36474
rect 24110 36420 24116 36422
rect 24172 36420 24196 36422
rect 24252 36420 24276 36422
rect 24332 36420 24356 36422
rect 24412 36420 24418 36422
rect 24110 36400 24418 36420
rect 24504 35698 24532 37198
rect 24596 36786 24624 37726
rect 24688 37262 24716 38150
rect 24676 37256 24728 37262
rect 24676 37198 24728 37204
rect 24584 36780 24636 36786
rect 24584 36722 24636 36728
rect 24780 36582 24808 38150
rect 24768 36576 24820 36582
rect 24768 36518 24820 36524
rect 24676 36372 24728 36378
rect 24676 36314 24728 36320
rect 24584 35760 24636 35766
rect 24584 35702 24636 35708
rect 24492 35692 24544 35698
rect 24492 35634 24544 35640
rect 24492 35556 24544 35562
rect 24492 35498 24544 35504
rect 24110 35388 24418 35408
rect 24110 35386 24116 35388
rect 24172 35386 24196 35388
rect 24252 35386 24276 35388
rect 24332 35386 24356 35388
rect 24412 35386 24418 35388
rect 24172 35334 24174 35386
rect 24354 35334 24356 35386
rect 24110 35332 24116 35334
rect 24172 35332 24196 35334
rect 24252 35332 24276 35334
rect 24332 35332 24356 35334
rect 24412 35332 24418 35334
rect 24110 35312 24418 35332
rect 24398 35184 24454 35193
rect 24308 35148 24360 35154
rect 24504 35154 24532 35498
rect 24398 35119 24454 35128
rect 24492 35148 24544 35154
rect 24308 35090 24360 35096
rect 24032 35080 24084 35086
rect 24032 35022 24084 35028
rect 24320 34542 24348 35090
rect 24412 34592 24440 35119
rect 24492 35090 24544 35096
rect 24492 34604 24544 34610
rect 24412 34564 24492 34592
rect 24492 34546 24544 34552
rect 24308 34536 24360 34542
rect 24044 34474 24256 34490
rect 24308 34478 24360 34484
rect 24596 34490 24624 35702
rect 24688 34649 24716 36314
rect 24780 35562 24808 36518
rect 24872 36378 24900 38286
rect 24952 38276 25004 38282
rect 24952 38218 25004 38224
rect 24964 36854 24992 38218
rect 25056 38010 25084 38286
rect 25044 38004 25096 38010
rect 25044 37946 25096 37952
rect 25136 38004 25188 38010
rect 25136 37946 25188 37952
rect 25044 37800 25096 37806
rect 25044 37742 25096 37748
rect 24952 36848 25004 36854
rect 24952 36790 25004 36796
rect 24860 36372 24912 36378
rect 24860 36314 24912 36320
rect 24768 35556 24820 35562
rect 24768 35498 24820 35504
rect 24952 34944 25004 34950
rect 24766 34912 24822 34921
rect 24952 34886 25004 34892
rect 24766 34847 24822 34856
rect 24674 34640 24730 34649
rect 24780 34610 24808 34847
rect 24964 34746 24992 34886
rect 24952 34740 25004 34746
rect 24952 34682 25004 34688
rect 24950 34640 25006 34649
rect 24674 34575 24730 34584
rect 24768 34604 24820 34610
rect 24950 34575 25006 34584
rect 24768 34546 24820 34552
rect 24860 34536 24912 34542
rect 24044 34468 24268 34474
rect 24044 34462 24216 34468
rect 23940 34060 23992 34066
rect 23940 34002 23992 34008
rect 23644 33516 23696 33522
rect 23584 33476 23644 33504
rect 23644 33458 23696 33464
rect 23848 33516 23900 33522
rect 23848 33458 23900 33464
rect 23756 33312 23808 33318
rect 23478 33280 23534 33289
rect 23756 33254 23808 33260
rect 23478 33215 23534 33224
rect 23400 33102 23520 33130
rect 23492 32910 23520 33102
rect 23480 32904 23532 32910
rect 23110 32872 23166 32881
rect 23480 32846 23532 32852
rect 23110 32807 23166 32816
rect 23124 32026 23152 32807
rect 23492 32298 23520 32846
rect 23768 32434 23796 33254
rect 23940 33108 23992 33114
rect 23940 33050 23992 33056
rect 23952 33017 23980 33050
rect 23938 33008 23994 33017
rect 23938 32943 23994 32952
rect 23756 32428 23808 32434
rect 23756 32370 23808 32376
rect 23480 32292 23532 32298
rect 23480 32234 23532 32240
rect 23112 32020 23164 32026
rect 23112 31962 23164 31968
rect 23480 32020 23532 32026
rect 23480 31962 23532 31968
rect 23124 31822 23152 31962
rect 23112 31816 23164 31822
rect 23388 31816 23440 31822
rect 23112 31758 23164 31764
rect 23386 31784 23388 31793
rect 23440 31784 23442 31793
rect 23492 31754 23520 31962
rect 24044 31754 24072 34462
rect 24596 34462 24808 34490
rect 24860 34478 24912 34484
rect 24216 34410 24268 34416
rect 24492 34400 24544 34406
rect 24492 34342 24544 34348
rect 24110 34300 24418 34320
rect 24110 34298 24116 34300
rect 24172 34298 24196 34300
rect 24252 34298 24276 34300
rect 24332 34298 24356 34300
rect 24412 34298 24418 34300
rect 24172 34246 24174 34298
rect 24354 34246 24356 34298
rect 24110 34244 24116 34246
rect 24172 34244 24196 34246
rect 24252 34244 24276 34246
rect 24332 34244 24356 34246
rect 24412 34244 24418 34246
rect 24110 34224 24418 34244
rect 24124 34060 24176 34066
rect 24124 34002 24176 34008
rect 24136 33454 24164 34002
rect 24504 33930 24532 34342
rect 24492 33924 24544 33930
rect 24492 33866 24544 33872
rect 24780 33674 24808 34462
rect 24872 34406 24900 34478
rect 24860 34400 24912 34406
rect 24860 34342 24912 34348
rect 24780 33646 24900 33674
rect 24768 33584 24820 33590
rect 24768 33526 24820 33532
rect 24124 33448 24176 33454
rect 24124 33390 24176 33396
rect 24110 33212 24418 33232
rect 24110 33210 24116 33212
rect 24172 33210 24196 33212
rect 24252 33210 24276 33212
rect 24332 33210 24356 33212
rect 24412 33210 24418 33212
rect 24172 33158 24174 33210
rect 24354 33158 24356 33210
rect 24110 33156 24116 33158
rect 24172 33156 24196 33158
rect 24252 33156 24276 33158
rect 24332 33156 24356 33158
rect 24412 33156 24418 33158
rect 24110 33136 24418 33156
rect 24676 32972 24728 32978
rect 24676 32914 24728 32920
rect 24584 32768 24636 32774
rect 24584 32710 24636 32716
rect 24110 32124 24418 32144
rect 24110 32122 24116 32124
rect 24172 32122 24196 32124
rect 24252 32122 24276 32124
rect 24332 32122 24356 32124
rect 24412 32122 24418 32124
rect 24172 32070 24174 32122
rect 24354 32070 24356 32122
rect 24110 32068 24116 32070
rect 24172 32068 24196 32070
rect 24252 32068 24276 32070
rect 24332 32068 24356 32070
rect 24412 32068 24418 32070
rect 24110 32048 24418 32068
rect 24596 31822 24624 32710
rect 24688 32434 24716 32914
rect 24676 32428 24728 32434
rect 24676 32370 24728 32376
rect 24676 32292 24728 32298
rect 24676 32234 24728 32240
rect 24492 31816 24544 31822
rect 24492 31758 24544 31764
rect 24584 31816 24636 31822
rect 24584 31758 24636 31764
rect 23386 31719 23442 31728
rect 23480 31748 23532 31754
rect 23480 31690 23532 31696
rect 23952 31726 24072 31754
rect 23204 31408 23256 31414
rect 23204 31350 23256 31356
rect 23112 31340 23164 31346
rect 23112 31282 23164 31288
rect 23124 30666 23152 31282
rect 23216 30938 23244 31350
rect 23388 31340 23440 31346
rect 23388 31282 23440 31288
rect 23204 30932 23256 30938
rect 23204 30874 23256 30880
rect 23294 30832 23350 30841
rect 23294 30767 23350 30776
rect 23308 30734 23336 30767
rect 23204 30728 23256 30734
rect 23204 30670 23256 30676
rect 23296 30728 23348 30734
rect 23296 30670 23348 30676
rect 23112 30660 23164 30666
rect 23112 30602 23164 30608
rect 23216 29170 23244 30670
rect 23294 29744 23350 29753
rect 23294 29679 23350 29688
rect 23308 29170 23336 29679
rect 23400 29578 23428 31282
rect 23492 31142 23520 31690
rect 23848 31680 23900 31686
rect 23848 31622 23900 31628
rect 23756 31476 23808 31482
rect 23756 31418 23808 31424
rect 23480 31136 23532 31142
rect 23480 31078 23532 31084
rect 23480 30592 23532 30598
rect 23480 30534 23532 30540
rect 23492 29646 23520 30534
rect 23572 30320 23624 30326
rect 23572 30262 23624 30268
rect 23480 29640 23532 29646
rect 23480 29582 23532 29588
rect 23388 29572 23440 29578
rect 23388 29514 23440 29520
rect 23480 29232 23532 29238
rect 23480 29174 23532 29180
rect 23204 29164 23256 29170
rect 23204 29106 23256 29112
rect 23296 29164 23348 29170
rect 23296 29106 23348 29112
rect 23110 29064 23166 29073
rect 23110 28999 23166 29008
rect 23124 28626 23152 28999
rect 23216 28762 23244 29106
rect 23388 29096 23440 29102
rect 23388 29038 23440 29044
rect 23296 28960 23348 28966
rect 23400 28937 23428 29038
rect 23296 28902 23348 28908
rect 23386 28928 23442 28937
rect 23204 28756 23256 28762
rect 23204 28698 23256 28704
rect 23112 28620 23164 28626
rect 23112 28562 23164 28568
rect 23308 27674 23336 28902
rect 23386 28863 23442 28872
rect 23492 28257 23520 29174
rect 23584 29170 23612 30262
rect 23768 30122 23796 31418
rect 23860 31414 23888 31622
rect 23848 31408 23900 31414
rect 23848 31350 23900 31356
rect 23952 31210 23980 31726
rect 24504 31346 24532 31758
rect 24688 31362 24716 32234
rect 24032 31340 24084 31346
rect 24032 31282 24084 31288
rect 24492 31340 24544 31346
rect 24492 31282 24544 31288
rect 24596 31334 24716 31362
rect 23940 31204 23992 31210
rect 23940 31146 23992 31152
rect 23848 30864 23900 30870
rect 23848 30806 23900 30812
rect 23860 30190 23888 30806
rect 23848 30184 23900 30190
rect 23848 30126 23900 30132
rect 23756 30116 23808 30122
rect 23756 30058 23808 30064
rect 23768 29889 23796 30058
rect 23754 29880 23810 29889
rect 23754 29815 23810 29824
rect 23952 29646 23980 31146
rect 24044 29850 24072 31282
rect 24110 31036 24418 31056
rect 24110 31034 24116 31036
rect 24172 31034 24196 31036
rect 24252 31034 24276 31036
rect 24332 31034 24356 31036
rect 24412 31034 24418 31036
rect 24172 30982 24174 31034
rect 24354 30982 24356 31034
rect 24110 30980 24116 30982
rect 24172 30980 24196 30982
rect 24252 30980 24276 30982
rect 24332 30980 24356 30982
rect 24412 30980 24418 30982
rect 24110 30960 24418 30980
rect 24110 29948 24418 29968
rect 24110 29946 24116 29948
rect 24172 29946 24196 29948
rect 24252 29946 24276 29948
rect 24332 29946 24356 29948
rect 24412 29946 24418 29948
rect 24172 29894 24174 29946
rect 24354 29894 24356 29946
rect 24110 29892 24116 29894
rect 24172 29892 24196 29894
rect 24252 29892 24276 29894
rect 24332 29892 24356 29894
rect 24412 29892 24418 29894
rect 24110 29872 24418 29892
rect 24032 29844 24084 29850
rect 24032 29786 24084 29792
rect 24400 29708 24452 29714
rect 24504 29696 24532 31282
rect 24452 29668 24532 29696
rect 24400 29650 24452 29656
rect 23940 29640 23992 29646
rect 23940 29582 23992 29588
rect 23754 29472 23810 29481
rect 23754 29407 23810 29416
rect 23662 29336 23718 29345
rect 23662 29271 23718 29280
rect 23572 29164 23624 29170
rect 23572 29106 23624 29112
rect 23676 28490 23704 29271
rect 23768 28490 23796 29407
rect 23664 28484 23716 28490
rect 23664 28426 23716 28432
rect 23756 28484 23808 28490
rect 23756 28426 23808 28432
rect 23478 28248 23534 28257
rect 23478 28183 23534 28192
rect 23848 28076 23900 28082
rect 23848 28018 23900 28024
rect 23480 28008 23532 28014
rect 23480 27950 23532 27956
rect 23204 27668 23256 27674
rect 23204 27610 23256 27616
rect 23296 27668 23348 27674
rect 23296 27610 23348 27616
rect 23112 27600 23164 27606
rect 23112 27542 23164 27548
rect 23216 27554 23244 27610
rect 23492 27554 23520 27950
rect 23756 27872 23808 27878
rect 23756 27814 23808 27820
rect 23768 27674 23796 27814
rect 23756 27668 23808 27674
rect 23756 27610 23808 27616
rect 23124 27305 23152 27542
rect 23216 27526 23520 27554
rect 23572 27464 23624 27470
rect 23572 27406 23624 27412
rect 23110 27296 23166 27305
rect 23110 27231 23166 27240
rect 23584 26926 23612 27406
rect 23860 27146 23888 28018
rect 23952 27946 23980 29582
rect 24030 29200 24086 29209
rect 24412 29170 24440 29650
rect 24596 29345 24624 31334
rect 24676 31272 24728 31278
rect 24676 31214 24728 31220
rect 24688 30734 24716 31214
rect 24676 30728 24728 30734
rect 24676 30670 24728 30676
rect 24582 29336 24638 29345
rect 24582 29271 24638 29280
rect 24030 29135 24086 29144
rect 24400 29164 24452 29170
rect 23940 27940 23992 27946
rect 23940 27882 23992 27888
rect 23952 27402 23980 27882
rect 23940 27396 23992 27402
rect 23940 27338 23992 27344
rect 23768 27118 23888 27146
rect 23572 26920 23624 26926
rect 23032 26846 23152 26874
rect 23572 26862 23624 26868
rect 22928 25764 22980 25770
rect 22928 25706 22980 25712
rect 22926 25664 22982 25673
rect 22926 25599 22982 25608
rect 22836 24812 22888 24818
rect 22836 24754 22888 24760
rect 22848 24274 22876 24754
rect 22836 24268 22888 24274
rect 22836 24210 22888 24216
rect 22468 24132 22520 24138
rect 22468 24074 22520 24080
rect 22374 23624 22430 23633
rect 22374 23559 22430 23568
rect 22284 23520 22336 23526
rect 22480 23474 22508 24074
rect 22664 23905 22692 24142
rect 22756 24126 22876 24154
rect 22650 23896 22706 23905
rect 22650 23831 22706 23840
rect 22560 23724 22612 23730
rect 22560 23666 22612 23672
rect 22284 23462 22336 23468
rect 22192 23248 22244 23254
rect 22192 23190 22244 23196
rect 22296 23118 22324 23462
rect 22388 23446 22508 23474
rect 22100 23112 22152 23118
rect 22100 23054 22152 23060
rect 22284 23112 22336 23118
rect 22284 23054 22336 23060
rect 21836 22052 21956 22080
rect 21732 22024 21784 22030
rect 21732 21966 21784 21972
rect 21744 21622 21772 21966
rect 21732 21616 21784 21622
rect 21732 21558 21784 21564
rect 21836 21536 21864 22052
rect 22008 21684 22060 21690
rect 22008 21626 22060 21632
rect 21916 21548 21968 21554
rect 21836 21508 21916 21536
rect 21836 20505 21864 21508
rect 21916 21490 21968 21496
rect 22020 21146 22048 21626
rect 22388 21554 22416 23446
rect 22572 23361 22600 23666
rect 22652 23656 22704 23662
rect 22652 23598 22704 23604
rect 22664 23497 22692 23598
rect 22650 23488 22706 23497
rect 22650 23423 22706 23432
rect 22558 23352 22614 23361
rect 22558 23287 22614 23296
rect 22468 23248 22520 23254
rect 22468 23190 22520 23196
rect 22376 21548 22428 21554
rect 22376 21490 22428 21496
rect 22388 21418 22416 21490
rect 22192 21412 22244 21418
rect 22192 21354 22244 21360
rect 22376 21412 22428 21418
rect 22376 21354 22428 21360
rect 22008 21140 22060 21146
rect 22008 21082 22060 21088
rect 22204 20913 22232 21354
rect 22374 21176 22430 21185
rect 22374 21111 22430 21120
rect 22388 20942 22416 21111
rect 22376 20936 22428 20942
rect 22190 20904 22246 20913
rect 22376 20878 22428 20884
rect 22190 20839 22246 20848
rect 21822 20496 21878 20505
rect 21822 20431 21878 20440
rect 22008 20324 22060 20330
rect 22008 20266 22060 20272
rect 21640 20052 21692 20058
rect 21640 19994 21692 20000
rect 22020 19854 22048 20266
rect 22008 19848 22060 19854
rect 22008 19790 22060 19796
rect 21548 19780 21600 19786
rect 21548 19722 21600 19728
rect 21456 18080 21508 18086
rect 21456 18022 21508 18028
rect 21364 16108 21416 16114
rect 21364 16050 21416 16056
rect 21468 12434 21496 18022
rect 21560 16794 21588 19722
rect 22192 19372 22244 19378
rect 22192 19314 22244 19320
rect 22100 19304 22152 19310
rect 22100 19246 22152 19252
rect 21732 19168 21784 19174
rect 21732 19110 21784 19116
rect 21744 18766 21772 19110
rect 22112 18970 22140 19246
rect 22100 18964 22152 18970
rect 22100 18906 22152 18912
rect 22100 18828 22152 18834
rect 22100 18770 22152 18776
rect 21732 18760 21784 18766
rect 21732 18702 21784 18708
rect 21824 18624 21876 18630
rect 21824 18566 21876 18572
rect 21836 18290 21864 18566
rect 21824 18284 21876 18290
rect 21824 18226 21876 18232
rect 21824 18080 21876 18086
rect 21824 18022 21876 18028
rect 21836 17678 21864 18022
rect 21824 17672 21876 17678
rect 21824 17614 21876 17620
rect 21640 16992 21692 16998
rect 21640 16934 21692 16940
rect 21548 16788 21600 16794
rect 21548 16730 21600 16736
rect 21652 16590 21680 16934
rect 22112 16794 22140 18770
rect 22204 18766 22232 19314
rect 22192 18760 22244 18766
rect 22192 18702 22244 18708
rect 22204 18290 22232 18702
rect 22284 18692 22336 18698
rect 22284 18634 22336 18640
rect 22192 18284 22244 18290
rect 22192 18226 22244 18232
rect 22204 18086 22232 18226
rect 22296 18222 22324 18634
rect 22284 18216 22336 18222
rect 22284 18158 22336 18164
rect 22296 18086 22324 18158
rect 22192 18080 22244 18086
rect 22192 18022 22244 18028
rect 22284 18080 22336 18086
rect 22284 18022 22336 18028
rect 22100 16788 22152 16794
rect 22100 16730 22152 16736
rect 22008 16720 22060 16726
rect 22006 16688 22008 16697
rect 22060 16688 22062 16697
rect 22204 16658 22232 18022
rect 22296 17542 22324 18022
rect 22284 17536 22336 17542
rect 22284 17478 22336 17484
rect 22006 16623 22062 16632
rect 22192 16652 22244 16658
rect 22192 16594 22244 16600
rect 21640 16584 21692 16590
rect 21640 16526 21692 16532
rect 22296 16454 22324 17478
rect 22284 16448 22336 16454
rect 22284 16390 22336 16396
rect 22388 16114 22416 20878
rect 22480 18970 22508 23190
rect 22664 22710 22692 23423
rect 22744 23180 22796 23186
rect 22744 23122 22796 23128
rect 22652 22704 22704 22710
rect 22652 22646 22704 22652
rect 22652 21888 22704 21894
rect 22652 21830 22704 21836
rect 22664 21486 22692 21830
rect 22652 21480 22704 21486
rect 22652 21422 22704 21428
rect 22652 21140 22704 21146
rect 22652 21082 22704 21088
rect 22560 20936 22612 20942
rect 22560 20878 22612 20884
rect 22572 19718 22600 20878
rect 22664 20369 22692 21082
rect 22756 21049 22784 23122
rect 22848 22166 22876 24126
rect 22940 23254 22968 25599
rect 23018 24712 23074 24721
rect 23018 24647 23074 24656
rect 23032 24206 23060 24647
rect 23020 24200 23072 24206
rect 23020 24142 23072 24148
rect 22928 23248 22980 23254
rect 22928 23190 22980 23196
rect 22928 23044 22980 23050
rect 22928 22986 22980 22992
rect 22836 22160 22888 22166
rect 22836 22102 22888 22108
rect 22940 21593 22968 22986
rect 23032 22642 23060 24142
rect 23020 22636 23072 22642
rect 23020 22578 23072 22584
rect 23020 22432 23072 22438
rect 23020 22374 23072 22380
rect 22926 21584 22982 21593
rect 22836 21548 22888 21554
rect 23032 21554 23060 22374
rect 22926 21519 22982 21528
rect 23020 21548 23072 21554
rect 22836 21490 22888 21496
rect 23020 21490 23072 21496
rect 22848 21434 22876 21490
rect 22848 21406 23060 21434
rect 22742 21040 22798 21049
rect 22742 20975 22798 20984
rect 22744 20800 22796 20806
rect 22744 20742 22796 20748
rect 22756 20466 22784 20742
rect 22836 20528 22888 20534
rect 22836 20470 22888 20476
rect 22744 20460 22796 20466
rect 22744 20402 22796 20408
rect 22650 20360 22706 20369
rect 22650 20295 22706 20304
rect 22848 20058 22876 20470
rect 22928 20460 22980 20466
rect 22928 20402 22980 20408
rect 22836 20052 22888 20058
rect 22836 19994 22888 20000
rect 22560 19712 22612 19718
rect 22560 19654 22612 19660
rect 22572 19242 22600 19654
rect 22560 19236 22612 19242
rect 22560 19178 22612 19184
rect 22468 18964 22520 18970
rect 22468 18906 22520 18912
rect 22468 18624 22520 18630
rect 22468 18566 22520 18572
rect 22480 17202 22508 18566
rect 22468 17196 22520 17202
rect 22468 17138 22520 17144
rect 22572 16182 22600 19178
rect 22836 18760 22888 18766
rect 22836 18702 22888 18708
rect 22848 18426 22876 18702
rect 22836 18420 22888 18426
rect 22836 18362 22888 18368
rect 22744 18352 22796 18358
rect 22744 18294 22796 18300
rect 22756 17338 22784 18294
rect 22744 17332 22796 17338
rect 22744 17274 22796 17280
rect 22756 16522 22784 17274
rect 22848 16658 22876 18362
rect 22836 16652 22888 16658
rect 22836 16594 22888 16600
rect 22744 16516 22796 16522
rect 22744 16458 22796 16464
rect 22560 16176 22612 16182
rect 22560 16118 22612 16124
rect 22756 16114 22784 16458
rect 22940 16250 22968 20402
rect 23032 16454 23060 21406
rect 23020 16448 23072 16454
rect 23020 16390 23072 16396
rect 22928 16244 22980 16250
rect 22928 16186 22980 16192
rect 22376 16108 22428 16114
rect 22376 16050 22428 16056
rect 22744 16108 22796 16114
rect 22744 16050 22796 16056
rect 23124 12434 23152 26846
rect 23572 26784 23624 26790
rect 23624 26744 23704 26772
rect 23572 26726 23624 26732
rect 23296 26512 23348 26518
rect 23296 26454 23348 26460
rect 23204 24608 23256 24614
rect 23204 24550 23256 24556
rect 23216 23662 23244 24550
rect 23308 24138 23336 26454
rect 23388 26444 23440 26450
rect 23388 26386 23440 26392
rect 23572 26444 23624 26450
rect 23572 26386 23624 26392
rect 23400 25498 23428 26386
rect 23584 26353 23612 26386
rect 23676 26382 23704 26744
rect 23664 26376 23716 26382
rect 23570 26344 23626 26353
rect 23664 26318 23716 26324
rect 23570 26279 23626 26288
rect 23478 26072 23534 26081
rect 23478 26007 23534 26016
rect 23492 25702 23520 26007
rect 23572 25900 23624 25906
rect 23572 25842 23624 25848
rect 23480 25696 23532 25702
rect 23480 25638 23532 25644
rect 23388 25492 23440 25498
rect 23388 25434 23440 25440
rect 23492 25294 23520 25638
rect 23480 25288 23532 25294
rect 23480 25230 23532 25236
rect 23480 25152 23532 25158
rect 23480 25094 23532 25100
rect 23388 24268 23440 24274
rect 23388 24210 23440 24216
rect 23296 24132 23348 24138
rect 23296 24074 23348 24080
rect 23204 23656 23256 23662
rect 23204 23598 23256 23604
rect 23400 23610 23428 24210
rect 23492 24041 23520 25094
rect 23478 24032 23534 24041
rect 23478 23967 23534 23976
rect 23492 23730 23520 23967
rect 23480 23724 23532 23730
rect 23480 23666 23532 23672
rect 23400 23582 23520 23610
rect 23388 23520 23440 23526
rect 23388 23462 23440 23468
rect 23296 23112 23348 23118
rect 23296 23054 23348 23060
rect 23204 22636 23256 22642
rect 23204 22578 23256 22584
rect 23216 22250 23244 22578
rect 23308 22438 23336 23054
rect 23400 22642 23428 23462
rect 23388 22636 23440 22642
rect 23388 22578 23440 22584
rect 23296 22432 23348 22438
rect 23296 22374 23348 22380
rect 23216 22222 23428 22250
rect 23296 22160 23348 22166
rect 23296 22102 23348 22108
rect 23308 20482 23336 22102
rect 23216 20454 23336 20482
rect 23216 18902 23244 20454
rect 23296 20392 23348 20398
rect 23296 20334 23348 20340
rect 23308 19854 23336 20334
rect 23296 19848 23348 19854
rect 23296 19790 23348 19796
rect 23308 19446 23336 19790
rect 23296 19440 23348 19446
rect 23296 19382 23348 19388
rect 23400 19378 23428 22222
rect 23492 21146 23520 23582
rect 23584 23118 23612 25842
rect 23676 25838 23704 26318
rect 23664 25832 23716 25838
rect 23664 25774 23716 25780
rect 23662 25392 23718 25401
rect 23662 25327 23718 25336
rect 23676 25226 23704 25327
rect 23664 25220 23716 25226
rect 23664 25162 23716 25168
rect 23664 24744 23716 24750
rect 23662 24712 23664 24721
rect 23716 24712 23718 24721
rect 23662 24647 23718 24656
rect 23664 24064 23716 24070
rect 23664 24006 23716 24012
rect 23676 23186 23704 24006
rect 23768 23338 23796 27118
rect 23848 26988 23900 26994
rect 23848 26930 23900 26936
rect 23860 26586 23888 26930
rect 24044 26874 24072 29135
rect 24400 29106 24452 29112
rect 24584 29164 24636 29170
rect 24584 29106 24636 29112
rect 24412 28948 24440 29106
rect 24412 28920 24532 28948
rect 24110 28860 24418 28880
rect 24110 28858 24116 28860
rect 24172 28858 24196 28860
rect 24252 28858 24276 28860
rect 24332 28858 24356 28860
rect 24412 28858 24418 28860
rect 24172 28806 24174 28858
rect 24354 28806 24356 28858
rect 24110 28804 24116 28806
rect 24172 28804 24196 28806
rect 24252 28804 24276 28806
rect 24332 28804 24356 28806
rect 24412 28804 24418 28806
rect 24110 28784 24418 28804
rect 24504 28558 24532 28920
rect 24492 28552 24544 28558
rect 24492 28494 24544 28500
rect 24124 28484 24176 28490
rect 24124 28426 24176 28432
rect 24136 27946 24164 28426
rect 24492 28076 24544 28082
rect 24492 28018 24544 28024
rect 24124 27940 24176 27946
rect 24124 27882 24176 27888
rect 24110 27772 24418 27792
rect 24110 27770 24116 27772
rect 24172 27770 24196 27772
rect 24252 27770 24276 27772
rect 24332 27770 24356 27772
rect 24412 27770 24418 27772
rect 24172 27718 24174 27770
rect 24354 27718 24356 27770
rect 24110 27716 24116 27718
rect 24172 27716 24196 27718
rect 24252 27716 24276 27718
rect 24332 27716 24356 27718
rect 24412 27716 24418 27718
rect 24110 27696 24418 27716
rect 24504 27577 24532 28018
rect 24490 27568 24546 27577
rect 24124 27532 24176 27538
rect 24490 27503 24546 27512
rect 24124 27474 24176 27480
rect 24136 26994 24164 27474
rect 24596 27130 24624 29106
rect 24688 27334 24716 30670
rect 24676 27328 24728 27334
rect 24676 27270 24728 27276
rect 24584 27124 24636 27130
rect 24584 27066 24636 27072
rect 24780 27033 24808 33526
rect 24872 32298 24900 33646
rect 24964 33454 24992 34575
rect 25056 33998 25084 37742
rect 25148 36038 25176 37946
rect 25608 37806 25636 38286
rect 25780 38276 25832 38282
rect 25870 38247 25926 38256
rect 25780 38218 25832 38224
rect 25596 37800 25648 37806
rect 25596 37742 25648 37748
rect 25608 37466 25636 37742
rect 25688 37664 25740 37670
rect 25688 37606 25740 37612
rect 25412 37460 25464 37466
rect 25412 37402 25464 37408
rect 25596 37460 25648 37466
rect 25596 37402 25648 37408
rect 25318 37088 25374 37097
rect 25318 37023 25374 37032
rect 25228 36236 25280 36242
rect 25228 36178 25280 36184
rect 25136 36032 25188 36038
rect 25136 35974 25188 35980
rect 25240 35834 25268 36178
rect 25228 35828 25280 35834
rect 25228 35770 25280 35776
rect 25332 35494 25360 37023
rect 25320 35488 25372 35494
rect 25320 35430 25372 35436
rect 25424 35086 25452 37402
rect 25596 36168 25648 36174
rect 25596 36110 25648 36116
rect 25504 36100 25556 36106
rect 25504 36042 25556 36048
rect 25516 35290 25544 36042
rect 25608 35601 25636 36110
rect 25594 35592 25650 35601
rect 25594 35527 25650 35536
rect 25504 35284 25556 35290
rect 25504 35226 25556 35232
rect 25504 35148 25556 35154
rect 25504 35090 25556 35096
rect 25412 35080 25464 35086
rect 25412 35022 25464 35028
rect 25516 34746 25544 35090
rect 25594 34776 25650 34785
rect 25504 34740 25556 34746
rect 25594 34711 25650 34720
rect 25504 34682 25556 34688
rect 25516 34542 25544 34682
rect 25608 34610 25636 34711
rect 25596 34604 25648 34610
rect 25596 34546 25648 34552
rect 25504 34536 25556 34542
rect 25504 34478 25556 34484
rect 25136 34400 25188 34406
rect 25136 34342 25188 34348
rect 25044 33992 25096 33998
rect 25044 33934 25096 33940
rect 24952 33448 25004 33454
rect 24952 33390 25004 33396
rect 25044 32972 25096 32978
rect 25044 32914 25096 32920
rect 24952 32768 25004 32774
rect 24952 32710 25004 32716
rect 24860 32292 24912 32298
rect 24860 32234 24912 32240
rect 24964 32230 24992 32710
rect 25056 32609 25084 32914
rect 25042 32600 25098 32609
rect 25042 32535 25098 32544
rect 25148 32298 25176 34342
rect 25228 33856 25280 33862
rect 25228 33798 25280 33804
rect 25240 32366 25268 33798
rect 25320 33448 25372 33454
rect 25320 33390 25372 33396
rect 25332 32910 25360 33390
rect 25412 32972 25464 32978
rect 25412 32914 25464 32920
rect 25320 32904 25372 32910
rect 25320 32846 25372 32852
rect 25320 32428 25372 32434
rect 25320 32370 25372 32376
rect 25228 32360 25280 32366
rect 25228 32302 25280 32308
rect 25136 32292 25188 32298
rect 25136 32234 25188 32240
rect 24952 32224 25004 32230
rect 24952 32166 25004 32172
rect 25148 31793 25176 32234
rect 25134 31784 25190 31793
rect 25134 31719 25190 31728
rect 25332 31686 25360 32370
rect 24860 31680 24912 31686
rect 24860 31622 24912 31628
rect 25320 31680 25372 31686
rect 25320 31622 25372 31628
rect 24872 31482 24900 31622
rect 24860 31476 24912 31482
rect 24860 31418 24912 31424
rect 24872 30666 24900 31418
rect 25424 31414 25452 32914
rect 25504 32904 25556 32910
rect 25608 32892 25636 34546
rect 25700 34066 25728 37606
rect 25792 35290 25820 38218
rect 25872 36304 25924 36310
rect 25870 36272 25872 36281
rect 25924 36272 25926 36281
rect 25870 36207 25926 36216
rect 25780 35284 25832 35290
rect 25780 35226 25832 35232
rect 25870 34776 25926 34785
rect 25870 34711 25926 34720
rect 25688 34060 25740 34066
rect 25688 34002 25740 34008
rect 25780 32972 25832 32978
rect 25780 32914 25832 32920
rect 25608 32864 25728 32892
rect 25792 32881 25820 32914
rect 25504 32846 25556 32852
rect 25516 31482 25544 32846
rect 25596 32360 25648 32366
rect 25596 32302 25648 32308
rect 25504 31476 25556 31482
rect 25504 31418 25556 31424
rect 24952 31408 25004 31414
rect 24952 31350 25004 31356
rect 25412 31408 25464 31414
rect 25412 31350 25464 31356
rect 24860 30660 24912 30666
rect 24860 30602 24912 30608
rect 24872 28540 24900 30602
rect 24964 30326 24992 31350
rect 25608 31346 25636 32302
rect 25320 31340 25372 31346
rect 25320 31282 25372 31288
rect 25596 31340 25648 31346
rect 25596 31282 25648 31288
rect 25228 31136 25280 31142
rect 25228 31078 25280 31084
rect 25044 30932 25096 30938
rect 25044 30874 25096 30880
rect 24952 30320 25004 30326
rect 24952 30262 25004 30268
rect 25056 30274 25084 30874
rect 25136 30728 25188 30734
rect 25136 30670 25188 30676
rect 25148 30394 25176 30670
rect 25136 30388 25188 30394
rect 25136 30330 25188 30336
rect 25056 30246 25176 30274
rect 25240 30258 25268 31078
rect 24950 30016 25006 30025
rect 24950 29951 25006 29960
rect 24964 29306 24992 29951
rect 25044 29640 25096 29646
rect 25148 29617 25176 30246
rect 25228 30252 25280 30258
rect 25228 30194 25280 30200
rect 25332 30054 25360 31282
rect 25700 30870 25728 32864
rect 25778 32872 25834 32881
rect 25778 32807 25834 32816
rect 25780 31136 25832 31142
rect 25780 31078 25832 31084
rect 25688 30864 25740 30870
rect 25688 30806 25740 30812
rect 25504 30660 25556 30666
rect 25504 30602 25556 30608
rect 25516 30326 25544 30602
rect 25504 30320 25556 30326
rect 25504 30262 25556 30268
rect 25412 30252 25464 30258
rect 25412 30194 25464 30200
rect 25320 30048 25372 30054
rect 25320 29990 25372 29996
rect 25044 29582 25096 29588
rect 25134 29608 25190 29617
rect 24952 29300 25004 29306
rect 24952 29242 25004 29248
rect 24952 28552 25004 28558
rect 24872 28512 24952 28540
rect 24952 28494 25004 28500
rect 25056 28150 25084 29582
rect 25134 29543 25190 29552
rect 25044 28144 25096 28150
rect 24950 28112 25006 28121
rect 25044 28086 25096 28092
rect 24950 28047 25006 28056
rect 24860 27328 24912 27334
rect 24860 27270 24912 27276
rect 24766 27024 24822 27033
rect 24124 26988 24176 26994
rect 24766 26959 24822 26968
rect 24124 26930 24176 26936
rect 24584 26920 24636 26926
rect 24044 26846 24532 26874
rect 24584 26862 24636 26868
rect 24110 26684 24418 26704
rect 24110 26682 24116 26684
rect 24172 26682 24196 26684
rect 24252 26682 24276 26684
rect 24332 26682 24356 26684
rect 24412 26682 24418 26684
rect 24172 26630 24174 26682
rect 24354 26630 24356 26682
rect 24110 26628 24116 26630
rect 24172 26628 24196 26630
rect 24252 26628 24276 26630
rect 24332 26628 24356 26630
rect 24412 26628 24418 26630
rect 24110 26608 24418 26628
rect 23848 26580 23900 26586
rect 23848 26522 23900 26528
rect 24504 26058 24532 26846
rect 24596 26314 24624 26862
rect 24768 26852 24820 26858
rect 24768 26794 24820 26800
rect 24780 26586 24808 26794
rect 24768 26580 24820 26586
rect 24768 26522 24820 26528
rect 24872 26314 24900 27270
rect 24964 26586 24992 28047
rect 25044 28008 25096 28014
rect 25044 27950 25096 27956
rect 25056 27470 25084 27950
rect 25044 27464 25096 27470
rect 25044 27406 25096 27412
rect 24952 26580 25004 26586
rect 24952 26522 25004 26528
rect 24584 26308 24636 26314
rect 24584 26250 24636 26256
rect 24860 26308 24912 26314
rect 24860 26250 24912 26256
rect 24504 26030 24808 26058
rect 24492 25900 24544 25906
rect 24492 25842 24544 25848
rect 24676 25900 24728 25906
rect 24676 25842 24728 25848
rect 24032 25832 24084 25838
rect 24032 25774 24084 25780
rect 23848 25696 23900 25702
rect 23848 25638 23900 25644
rect 23860 24274 23888 25638
rect 24044 25276 24072 25774
rect 24110 25596 24418 25616
rect 24110 25594 24116 25596
rect 24172 25594 24196 25596
rect 24252 25594 24276 25596
rect 24332 25594 24356 25596
rect 24412 25594 24418 25596
rect 24172 25542 24174 25594
rect 24354 25542 24356 25594
rect 24110 25540 24116 25542
rect 24172 25540 24196 25542
rect 24252 25540 24276 25542
rect 24332 25540 24356 25542
rect 24412 25540 24418 25542
rect 24110 25520 24418 25540
rect 24044 25248 24164 25276
rect 23940 24812 23992 24818
rect 23940 24754 23992 24760
rect 23848 24268 23900 24274
rect 23848 24210 23900 24216
rect 23768 23310 23888 23338
rect 23664 23180 23716 23186
rect 23664 23122 23716 23128
rect 23860 23118 23888 23310
rect 23572 23112 23624 23118
rect 23756 23112 23808 23118
rect 23572 23054 23624 23060
rect 23662 23080 23718 23089
rect 23584 22488 23612 23054
rect 23756 23054 23808 23060
rect 23848 23112 23900 23118
rect 23848 23054 23900 23060
rect 23662 23015 23718 23024
rect 23676 22681 23704 23015
rect 23768 22817 23796 23054
rect 23952 22982 23980 24754
rect 24136 24750 24164 25248
rect 24124 24744 24176 24750
rect 24124 24686 24176 24692
rect 24136 24596 24164 24686
rect 24044 24568 24164 24596
rect 23940 22976 23992 22982
rect 23940 22918 23992 22924
rect 23754 22808 23810 22817
rect 24044 22794 24072 24568
rect 24110 24508 24418 24528
rect 24110 24506 24116 24508
rect 24172 24506 24196 24508
rect 24252 24506 24276 24508
rect 24332 24506 24356 24508
rect 24412 24506 24418 24508
rect 24172 24454 24174 24506
rect 24354 24454 24356 24506
rect 24110 24452 24116 24454
rect 24172 24452 24196 24454
rect 24252 24452 24276 24454
rect 24332 24452 24356 24454
rect 24412 24452 24418 24454
rect 24110 24432 24418 24452
rect 24504 24070 24532 25842
rect 24584 25696 24636 25702
rect 24584 25638 24636 25644
rect 24492 24064 24544 24070
rect 24306 24032 24362 24041
rect 24492 24006 24544 24012
rect 24306 23967 24362 23976
rect 24320 23866 24348 23967
rect 24596 23866 24624 25638
rect 24688 25498 24716 25842
rect 24676 25492 24728 25498
rect 24676 25434 24728 25440
rect 24780 25378 24808 26030
rect 24688 25350 24808 25378
rect 24688 24614 24716 25350
rect 24872 25276 24900 26250
rect 25056 25838 25084 27406
rect 25148 26858 25176 29543
rect 25424 29034 25452 30194
rect 25412 29028 25464 29034
rect 25412 28970 25464 28976
rect 25516 27606 25544 30262
rect 25700 30258 25728 30806
rect 25688 30252 25740 30258
rect 25688 30194 25740 30200
rect 25792 29850 25820 31078
rect 25780 29844 25832 29850
rect 25780 29786 25832 29792
rect 25596 29776 25648 29782
rect 25594 29744 25596 29753
rect 25648 29744 25650 29753
rect 25884 29714 25912 34711
rect 25976 33658 26004 38830
rect 26068 38185 26096 39442
rect 26148 38888 26200 38894
rect 26146 38856 26148 38865
rect 26200 38856 26202 38865
rect 26146 38791 26202 38800
rect 26238 38720 26294 38729
rect 26238 38655 26294 38664
rect 26054 38176 26110 38185
rect 26054 38111 26110 38120
rect 26252 37262 26280 38655
rect 26344 38418 26372 40190
rect 26606 39944 26662 39953
rect 26606 39879 26662 39888
rect 26332 38412 26384 38418
rect 26332 38354 26384 38360
rect 26424 37732 26476 37738
rect 26424 37674 26476 37680
rect 26240 37256 26292 37262
rect 26240 37198 26292 37204
rect 26436 36922 26464 37674
rect 26514 37360 26570 37369
rect 26514 37295 26516 37304
rect 26568 37295 26570 37304
rect 26516 37266 26568 37272
rect 26424 36916 26476 36922
rect 26424 36858 26476 36864
rect 26330 36816 26386 36825
rect 26330 36751 26386 36760
rect 26344 36174 26372 36751
rect 26332 36168 26384 36174
rect 26332 36110 26384 36116
rect 26436 35562 26464 36858
rect 26424 35556 26476 35562
rect 26424 35498 26476 35504
rect 26620 35154 26648 39879
rect 26792 39364 26844 39370
rect 26792 39306 26844 39312
rect 26804 37874 26832 39306
rect 26792 37868 26844 37874
rect 26792 37810 26844 37816
rect 26608 35148 26660 35154
rect 26608 35090 26660 35096
rect 26804 34746 26832 37810
rect 26896 36718 26924 40462
rect 26976 39024 27028 39030
rect 26976 38966 27028 38972
rect 26988 38554 27016 38966
rect 26976 38548 27028 38554
rect 26976 38490 27028 38496
rect 26988 36922 27016 38490
rect 27080 37942 27108 41200
rect 27620 39364 27672 39370
rect 27620 39306 27672 39312
rect 27160 39024 27212 39030
rect 27160 38966 27212 38972
rect 27068 37936 27120 37942
rect 27068 37878 27120 37884
rect 26976 36916 27028 36922
rect 26976 36858 27028 36864
rect 27172 36786 27200 38966
rect 27436 38820 27488 38826
rect 27436 38762 27488 38768
rect 27344 38752 27396 38758
rect 27344 38694 27396 38700
rect 27160 36780 27212 36786
rect 27160 36722 27212 36728
rect 26884 36712 26936 36718
rect 26884 36654 26936 36660
rect 27068 36712 27120 36718
rect 27068 36654 27120 36660
rect 26974 36000 27030 36009
rect 26974 35935 27030 35944
rect 26988 35698 27016 35935
rect 26976 35692 27028 35698
rect 26976 35634 27028 35640
rect 26988 35290 27016 35634
rect 26976 35284 27028 35290
rect 26976 35226 27028 35232
rect 26792 34740 26844 34746
rect 26792 34682 26844 34688
rect 26240 34468 26292 34474
rect 26240 34410 26292 34416
rect 26252 34134 26280 34410
rect 26330 34232 26386 34241
rect 26330 34167 26386 34176
rect 26240 34128 26292 34134
rect 26146 34096 26202 34105
rect 26240 34070 26292 34076
rect 26344 34066 26372 34167
rect 26146 34031 26202 34040
rect 26332 34060 26384 34066
rect 25964 33652 26016 33658
rect 25964 33594 26016 33600
rect 26160 33454 26188 34031
rect 26332 34002 26384 34008
rect 26514 33960 26570 33969
rect 26514 33895 26516 33904
rect 26568 33895 26570 33904
rect 26516 33866 26568 33872
rect 26976 33516 27028 33522
rect 26976 33458 27028 33464
rect 26148 33448 26200 33454
rect 26148 33390 26200 33396
rect 26330 33416 26386 33425
rect 26330 33351 26386 33360
rect 26344 32978 26372 33351
rect 26332 32972 26384 32978
rect 26332 32914 26384 32920
rect 26146 32464 26202 32473
rect 26146 32399 26202 32408
rect 25964 32224 26016 32230
rect 25964 32166 26016 32172
rect 26056 32224 26108 32230
rect 26056 32166 26108 32172
rect 25976 32026 26004 32166
rect 25964 32020 26016 32026
rect 25964 31962 26016 31968
rect 26068 30433 26096 32166
rect 26160 31346 26188 32399
rect 26988 32337 27016 33458
rect 26974 32328 27030 32337
rect 26896 32286 26974 32314
rect 26330 31920 26386 31929
rect 26330 31855 26332 31864
rect 26384 31855 26386 31864
rect 26332 31826 26384 31832
rect 26424 31476 26476 31482
rect 26424 31418 26476 31424
rect 26436 31385 26464 31418
rect 26422 31376 26478 31385
rect 26148 31340 26200 31346
rect 26422 31311 26478 31320
rect 26148 31282 26200 31288
rect 26332 30728 26384 30734
rect 26332 30670 26384 30676
rect 26344 30433 26372 30670
rect 26054 30424 26110 30433
rect 26054 30359 26110 30368
rect 26330 30424 26386 30433
rect 26330 30359 26386 30368
rect 26896 30326 26924 32286
rect 26974 32263 27030 32272
rect 27080 30870 27108 36654
rect 27172 34474 27200 36722
rect 27252 36032 27304 36038
rect 27252 35974 27304 35980
rect 27264 35698 27292 35974
rect 27356 35766 27384 38694
rect 27448 36786 27476 38762
rect 27528 38752 27580 38758
rect 27528 38694 27580 38700
rect 27436 36780 27488 36786
rect 27436 36722 27488 36728
rect 27448 36378 27476 36722
rect 27436 36372 27488 36378
rect 27436 36314 27488 36320
rect 27344 35760 27396 35766
rect 27344 35702 27396 35708
rect 27252 35692 27304 35698
rect 27252 35634 27304 35640
rect 27436 35624 27488 35630
rect 27540 35612 27568 38694
rect 27632 36802 27660 39306
rect 27724 38418 27752 41200
rect 28170 40896 28226 40905
rect 28170 40831 28226 40840
rect 27988 38956 28040 38962
rect 27988 38898 28040 38904
rect 27712 38412 27764 38418
rect 27712 38354 27764 38360
rect 28000 37942 28028 38898
rect 27988 37936 28040 37942
rect 27988 37878 28040 37884
rect 28080 37664 28132 37670
rect 28080 37606 28132 37612
rect 28092 37126 28120 37606
rect 28184 37262 28212 40831
rect 28262 39536 28318 39545
rect 28262 39471 28318 39480
rect 28172 37256 28224 37262
rect 28172 37198 28224 37204
rect 28080 37120 28132 37126
rect 28080 37062 28132 37068
rect 28170 36816 28226 36825
rect 27632 36774 27752 36802
rect 27620 36644 27672 36650
rect 27620 36586 27672 36592
rect 27488 35584 27568 35612
rect 27436 35566 27488 35572
rect 27344 35488 27396 35494
rect 27344 35430 27396 35436
rect 27356 34474 27384 35430
rect 27160 34468 27212 34474
rect 27160 34410 27212 34416
rect 27344 34468 27396 34474
rect 27344 34410 27396 34416
rect 27252 33312 27304 33318
rect 27252 33254 27304 33260
rect 27160 32428 27212 32434
rect 27160 32370 27212 32376
rect 27172 31482 27200 32370
rect 27264 32366 27292 33254
rect 27448 33114 27476 35566
rect 27632 33590 27660 36586
rect 27620 33584 27672 33590
rect 27620 33526 27672 33532
rect 27724 33454 27752 36774
rect 28170 36751 28226 36760
rect 27896 36576 27948 36582
rect 27896 36518 27948 36524
rect 27804 35284 27856 35290
rect 27804 35226 27856 35232
rect 27712 33448 27764 33454
rect 27712 33390 27764 33396
rect 27712 33312 27764 33318
rect 27712 33254 27764 33260
rect 27436 33108 27488 33114
rect 27436 33050 27488 33056
rect 27344 32496 27396 32502
rect 27344 32438 27396 32444
rect 27252 32360 27304 32366
rect 27252 32302 27304 32308
rect 27356 31482 27384 32438
rect 27528 32224 27580 32230
rect 27528 32166 27580 32172
rect 27160 31476 27212 31482
rect 27160 31418 27212 31424
rect 27344 31476 27396 31482
rect 27344 31418 27396 31424
rect 27068 30864 27120 30870
rect 27068 30806 27120 30812
rect 26976 30592 27028 30598
rect 26976 30534 27028 30540
rect 26884 30320 26936 30326
rect 26804 30280 26884 30308
rect 25976 30190 26004 30221
rect 25964 30184 26016 30190
rect 25962 30152 25964 30161
rect 26016 30152 26018 30161
rect 25962 30087 26018 30096
rect 25976 29850 26004 30087
rect 25964 29844 26016 29850
rect 25964 29786 26016 29792
rect 25594 29679 25650 29688
rect 25872 29708 25924 29714
rect 25872 29650 25924 29656
rect 26332 29640 26384 29646
rect 26332 29582 26384 29588
rect 26344 29238 26372 29582
rect 26606 29336 26662 29345
rect 26804 29306 26832 30280
rect 26884 30262 26936 30268
rect 26988 30258 27016 30534
rect 27080 30258 27108 30806
rect 27540 30802 27568 32166
rect 27620 31340 27672 31346
rect 27620 31282 27672 31288
rect 27528 30796 27580 30802
rect 27528 30738 27580 30744
rect 27252 30660 27304 30666
rect 27252 30602 27304 30608
rect 27264 30258 27292 30602
rect 26976 30252 27028 30258
rect 26976 30194 27028 30200
rect 27068 30252 27120 30258
rect 27068 30194 27120 30200
rect 27252 30252 27304 30258
rect 27252 30194 27304 30200
rect 26884 30184 26936 30190
rect 26884 30126 26936 30132
rect 26606 29271 26662 29280
rect 26792 29300 26844 29306
rect 26332 29232 26384 29238
rect 26332 29174 26384 29180
rect 26056 29164 26108 29170
rect 26056 29106 26108 29112
rect 26068 29034 26096 29106
rect 25872 29028 25924 29034
rect 25872 28970 25924 28976
rect 26056 29028 26108 29034
rect 26056 28970 26108 28976
rect 25688 28552 25740 28558
rect 25688 28494 25740 28500
rect 25700 28422 25728 28494
rect 25596 28416 25648 28422
rect 25596 28358 25648 28364
rect 25688 28416 25740 28422
rect 25688 28358 25740 28364
rect 25608 28082 25636 28358
rect 25596 28076 25648 28082
rect 25596 28018 25648 28024
rect 25504 27600 25556 27606
rect 25504 27542 25556 27548
rect 25412 27396 25464 27402
rect 25412 27338 25464 27344
rect 25136 26852 25188 26858
rect 25136 26794 25188 26800
rect 25424 26432 25452 27338
rect 25594 27296 25650 27305
rect 25594 27231 25650 27240
rect 25424 26404 25544 26432
rect 25410 26344 25466 26353
rect 25410 26279 25466 26288
rect 25044 25832 25096 25838
rect 25044 25774 25096 25780
rect 24780 25248 24900 25276
rect 24676 24608 24728 24614
rect 24676 24550 24728 24556
rect 24674 23896 24730 23905
rect 24308 23860 24360 23866
rect 24308 23802 24360 23808
rect 24584 23860 24636 23866
rect 24674 23831 24676 23840
rect 24584 23802 24636 23808
rect 24728 23831 24730 23840
rect 24676 23802 24728 23808
rect 24320 23730 24348 23802
rect 24780 23746 24808 25248
rect 24860 25152 24912 25158
rect 24860 25094 24912 25100
rect 24872 24041 24900 25094
rect 24952 24200 25004 24206
rect 24950 24168 24952 24177
rect 25004 24168 25006 24177
rect 24950 24103 25006 24112
rect 24858 24032 24914 24041
rect 24858 23967 24914 23976
rect 24308 23724 24360 23730
rect 24308 23666 24360 23672
rect 24504 23718 24808 23746
rect 25056 23730 25084 25774
rect 25228 25696 25280 25702
rect 25228 25638 25280 25644
rect 25240 25294 25268 25638
rect 25228 25288 25280 25294
rect 25228 25230 25280 25236
rect 25320 25288 25372 25294
rect 25320 25230 25372 25236
rect 25228 24880 25280 24886
rect 25228 24822 25280 24828
rect 25240 24410 25268 24822
rect 25228 24404 25280 24410
rect 25228 24346 25280 24352
rect 25226 24304 25282 24313
rect 25226 24239 25282 24248
rect 24860 23724 24912 23730
rect 24110 23420 24418 23440
rect 24110 23418 24116 23420
rect 24172 23418 24196 23420
rect 24252 23418 24276 23420
rect 24332 23418 24356 23420
rect 24412 23418 24418 23420
rect 24172 23366 24174 23418
rect 24354 23366 24356 23418
rect 24110 23364 24116 23366
rect 24172 23364 24196 23366
rect 24252 23364 24276 23366
rect 24332 23364 24356 23366
rect 24412 23364 24418 23366
rect 24110 23344 24418 23364
rect 24124 23112 24176 23118
rect 24124 23054 24176 23060
rect 24400 23112 24452 23118
rect 24504 23100 24532 23718
rect 24860 23666 24912 23672
rect 25044 23724 25096 23730
rect 25044 23666 25096 23672
rect 24584 23520 24636 23526
rect 24584 23462 24636 23468
rect 24452 23072 24532 23100
rect 24400 23054 24452 23060
rect 24136 22982 24164 23054
rect 24124 22976 24176 22982
rect 24124 22918 24176 22924
rect 23754 22743 23810 22752
rect 23860 22766 24072 22794
rect 24492 22772 24544 22778
rect 23662 22672 23718 22681
rect 23662 22607 23664 22616
rect 23716 22607 23718 22616
rect 23664 22578 23716 22584
rect 23676 22547 23704 22578
rect 23664 22500 23716 22506
rect 23584 22460 23664 22488
rect 23584 21962 23612 22460
rect 23664 22442 23716 22448
rect 23662 22128 23718 22137
rect 23662 22063 23718 22072
rect 23676 22030 23704 22063
rect 23664 22024 23716 22030
rect 23664 21966 23716 21972
rect 23572 21956 23624 21962
rect 23572 21898 23624 21904
rect 23664 21684 23716 21690
rect 23664 21626 23716 21632
rect 23676 21146 23704 21626
rect 23756 21344 23808 21350
rect 23756 21286 23808 21292
rect 23480 21140 23532 21146
rect 23480 21082 23532 21088
rect 23664 21140 23716 21146
rect 23664 21082 23716 21088
rect 23480 21004 23532 21010
rect 23480 20946 23532 20952
rect 23664 20974 23716 20980
rect 23492 19514 23520 20946
rect 23572 20936 23624 20942
rect 23664 20916 23716 20922
rect 23572 20878 23624 20884
rect 23584 20058 23612 20878
rect 23676 20602 23704 20916
rect 23664 20596 23716 20602
rect 23664 20538 23716 20544
rect 23572 20052 23624 20058
rect 23572 19994 23624 20000
rect 23664 19984 23716 19990
rect 23664 19926 23716 19932
rect 23480 19508 23532 19514
rect 23480 19450 23532 19456
rect 23676 19378 23704 19926
rect 23768 19854 23796 21286
rect 23860 20398 23888 22766
rect 24492 22714 24544 22720
rect 24110 22332 24418 22352
rect 24110 22330 24116 22332
rect 24172 22330 24196 22332
rect 24252 22330 24276 22332
rect 24332 22330 24356 22332
rect 24412 22330 24418 22332
rect 24172 22278 24174 22330
rect 24354 22278 24356 22330
rect 24110 22276 24116 22278
rect 24172 22276 24196 22278
rect 24252 22276 24276 22278
rect 24332 22276 24356 22278
rect 24412 22276 24418 22278
rect 24110 22256 24418 22276
rect 24504 22234 24532 22714
rect 24032 22228 24084 22234
rect 24032 22170 24084 22176
rect 24492 22228 24544 22234
rect 24492 22170 24544 22176
rect 24044 21690 24072 22170
rect 24032 21684 24084 21690
rect 24032 21626 24084 21632
rect 24504 21536 24532 22170
rect 24596 21962 24624 23462
rect 24768 23112 24820 23118
rect 24674 23080 24730 23089
rect 24768 23054 24820 23060
rect 24674 23015 24676 23024
rect 24728 23015 24730 23024
rect 24676 22986 24728 22992
rect 24780 22642 24808 23054
rect 24872 22982 24900 23666
rect 25044 23588 25096 23594
rect 25044 23530 25096 23536
rect 25056 23186 25084 23530
rect 25044 23180 25096 23186
rect 25044 23122 25096 23128
rect 25240 23050 25268 24239
rect 25228 23044 25280 23050
rect 25228 22986 25280 22992
rect 24860 22976 24912 22982
rect 24860 22918 24912 22924
rect 25136 22704 25188 22710
rect 24950 22672 25006 22681
rect 24768 22636 24820 22642
rect 25188 22664 25268 22692
rect 25332 22681 25360 25230
rect 25424 22692 25452 26279
rect 25516 26246 25544 26404
rect 25608 26382 25636 27231
rect 25700 26790 25728 28358
rect 25884 26994 25912 28970
rect 26068 27878 26096 28970
rect 26332 28552 26384 28558
rect 26332 28494 26384 28500
rect 26056 27872 26108 27878
rect 26056 27814 26108 27820
rect 26344 27713 26372 28494
rect 26516 28484 26568 28490
rect 26516 28426 26568 28432
rect 26528 28218 26556 28426
rect 26516 28212 26568 28218
rect 26516 28154 26568 28160
rect 26330 27704 26386 27713
rect 26330 27639 26386 27648
rect 25964 27600 26016 27606
rect 25964 27542 26016 27548
rect 25872 26988 25924 26994
rect 25872 26930 25924 26936
rect 25688 26784 25740 26790
rect 25688 26726 25740 26732
rect 25780 26580 25832 26586
rect 25780 26522 25832 26528
rect 25596 26376 25648 26382
rect 25596 26318 25648 26324
rect 25504 26240 25556 26246
rect 25504 26182 25556 26188
rect 25792 25906 25820 26522
rect 25976 26382 26004 27542
rect 26332 27464 26384 27470
rect 26054 27432 26110 27441
rect 26332 27406 26384 27412
rect 26054 27367 26110 27376
rect 26068 26382 26096 27367
rect 26344 26897 26372 27406
rect 26330 26888 26386 26897
rect 26330 26823 26386 26832
rect 25964 26376 26016 26382
rect 25964 26318 26016 26324
rect 26056 26376 26108 26382
rect 26056 26318 26108 26324
rect 25780 25900 25832 25906
rect 25780 25842 25832 25848
rect 25976 25820 26004 26318
rect 26422 25936 26478 25945
rect 26422 25871 26478 25880
rect 26056 25832 26108 25838
rect 25976 25792 26056 25820
rect 26056 25774 26108 25780
rect 26436 25770 26464 25871
rect 26424 25764 26476 25770
rect 26424 25706 26476 25712
rect 26332 25288 26384 25294
rect 26330 25256 26332 25265
rect 26384 25256 26386 25265
rect 25504 25220 25556 25226
rect 26330 25191 26386 25200
rect 25504 25162 25556 25168
rect 25516 24750 25544 25162
rect 26056 24880 26108 24886
rect 26056 24822 26108 24828
rect 26146 24848 26202 24857
rect 25504 24744 25556 24750
rect 25504 24686 25556 24692
rect 25596 24608 25648 24614
rect 25596 24550 25648 24556
rect 25608 23730 25636 24550
rect 25780 24064 25832 24070
rect 25780 24006 25832 24012
rect 25792 23798 25820 24006
rect 25780 23792 25832 23798
rect 25780 23734 25832 23740
rect 25596 23724 25648 23730
rect 25596 23666 25648 23672
rect 25688 23316 25740 23322
rect 25688 23258 25740 23264
rect 25700 23225 25728 23258
rect 25686 23216 25742 23225
rect 26068 23186 26096 24822
rect 26146 24783 26148 24792
rect 26200 24783 26202 24792
rect 26148 24754 26200 24760
rect 26332 24200 26384 24206
rect 26332 24142 26384 24148
rect 26344 23497 26372 24142
rect 26330 23488 26386 23497
rect 26330 23423 26386 23432
rect 25686 23151 25742 23160
rect 26056 23180 26108 23186
rect 26056 23122 26108 23128
rect 25136 22646 25188 22652
rect 24950 22607 25006 22616
rect 24768 22578 24820 22584
rect 24674 22536 24730 22545
rect 24674 22471 24676 22480
rect 24728 22471 24730 22480
rect 24676 22442 24728 22448
rect 24676 22024 24728 22030
rect 24780 21978 24808 22578
rect 24964 22030 24992 22607
rect 25044 22568 25096 22574
rect 25044 22510 25096 22516
rect 24952 22024 25004 22030
rect 24728 21972 24900 21978
rect 24676 21966 24900 21972
rect 24952 21966 25004 21972
rect 24584 21956 24636 21962
rect 24688 21950 24900 21966
rect 24584 21898 24636 21904
rect 24676 21888 24728 21894
rect 24676 21830 24728 21836
rect 24504 21508 24624 21536
rect 24110 21244 24418 21264
rect 24110 21242 24116 21244
rect 24172 21242 24196 21244
rect 24252 21242 24276 21244
rect 24332 21242 24356 21244
rect 24412 21242 24418 21244
rect 24172 21190 24174 21242
rect 24354 21190 24356 21242
rect 24110 21188 24116 21190
rect 24172 21188 24196 21190
rect 24252 21188 24276 21190
rect 24332 21188 24356 21190
rect 24412 21188 24418 21190
rect 24110 21168 24418 21188
rect 24596 21185 24624 21508
rect 24582 21176 24638 21185
rect 24582 21111 24638 21120
rect 24584 20868 24636 20874
rect 24584 20810 24636 20816
rect 23940 20460 23992 20466
rect 23940 20402 23992 20408
rect 23848 20392 23900 20398
rect 23848 20334 23900 20340
rect 23756 19848 23808 19854
rect 23756 19790 23808 19796
rect 23388 19372 23440 19378
rect 23388 19314 23440 19320
rect 23572 19372 23624 19378
rect 23572 19314 23624 19320
rect 23664 19372 23716 19378
rect 23664 19314 23716 19320
rect 23584 18970 23612 19314
rect 23388 18964 23440 18970
rect 23388 18906 23440 18912
rect 23572 18964 23624 18970
rect 23572 18906 23624 18912
rect 23204 18896 23256 18902
rect 23204 18838 23256 18844
rect 23296 18692 23348 18698
rect 23296 18634 23348 18640
rect 23308 17338 23336 18634
rect 23400 18086 23428 18906
rect 23388 18080 23440 18086
rect 23388 18022 23440 18028
rect 23572 17672 23624 17678
rect 23572 17614 23624 17620
rect 23296 17332 23348 17338
rect 23296 17274 23348 17280
rect 23308 16794 23336 17274
rect 23388 16992 23440 16998
rect 23388 16934 23440 16940
rect 23296 16788 23348 16794
rect 23296 16730 23348 16736
rect 23202 16688 23258 16697
rect 23202 16623 23258 16632
rect 23296 16652 23348 16658
rect 23216 16182 23244 16623
rect 23296 16594 23348 16600
rect 23204 16176 23256 16182
rect 23204 16118 23256 16124
rect 23308 15978 23336 16594
rect 23400 16590 23428 16934
rect 23388 16584 23440 16590
rect 23388 16526 23440 16532
rect 23400 16114 23428 16526
rect 23388 16108 23440 16114
rect 23388 16050 23440 16056
rect 23296 15972 23348 15978
rect 23296 15914 23348 15920
rect 23400 15026 23428 16050
rect 23480 15904 23532 15910
rect 23480 15846 23532 15852
rect 23492 15570 23520 15846
rect 23480 15564 23532 15570
rect 23480 15506 23532 15512
rect 23584 15366 23612 17614
rect 23676 16114 23704 19314
rect 23768 18766 23796 19790
rect 23860 19446 23888 20334
rect 23848 19440 23900 19446
rect 23848 19382 23900 19388
rect 23952 19378 23980 20402
rect 24032 20256 24084 20262
rect 24032 20198 24084 20204
rect 24492 20256 24544 20262
rect 24492 20198 24544 20204
rect 23940 19372 23992 19378
rect 23940 19314 23992 19320
rect 23848 19236 23900 19242
rect 23848 19178 23900 19184
rect 23756 18760 23808 18766
rect 23756 18702 23808 18708
rect 23756 17672 23808 17678
rect 23756 17614 23808 17620
rect 23768 17542 23796 17614
rect 23756 17536 23808 17542
rect 23756 17478 23808 17484
rect 23756 17196 23808 17202
rect 23756 17138 23808 17144
rect 23664 16108 23716 16114
rect 23664 16050 23716 16056
rect 23768 15722 23796 17138
rect 23676 15706 23796 15722
rect 23664 15700 23796 15706
rect 23716 15694 23796 15700
rect 23664 15642 23716 15648
rect 23860 15434 23888 19178
rect 23848 15428 23900 15434
rect 23848 15370 23900 15376
rect 23572 15360 23624 15366
rect 23572 15302 23624 15308
rect 23952 15162 23980 19314
rect 23940 15156 23992 15162
rect 23940 15098 23992 15104
rect 23388 15020 23440 15026
rect 23388 14962 23440 14968
rect 24044 12434 24072 20198
rect 24110 20156 24418 20176
rect 24110 20154 24116 20156
rect 24172 20154 24196 20156
rect 24252 20154 24276 20156
rect 24332 20154 24356 20156
rect 24412 20154 24418 20156
rect 24172 20102 24174 20154
rect 24354 20102 24356 20154
rect 24110 20100 24116 20102
rect 24172 20100 24196 20102
rect 24252 20100 24276 20102
rect 24332 20100 24356 20102
rect 24412 20100 24418 20102
rect 24110 20080 24418 20100
rect 24306 19952 24362 19961
rect 24306 19887 24362 19896
rect 24320 19242 24348 19887
rect 24308 19236 24360 19242
rect 24308 19178 24360 19184
rect 24110 19068 24418 19088
rect 24110 19066 24116 19068
rect 24172 19066 24196 19068
rect 24252 19066 24276 19068
rect 24332 19066 24356 19068
rect 24412 19066 24418 19068
rect 24172 19014 24174 19066
rect 24354 19014 24356 19066
rect 24110 19012 24116 19014
rect 24172 19012 24196 19014
rect 24252 19012 24276 19014
rect 24332 19012 24356 19014
rect 24412 19012 24418 19014
rect 24110 18992 24418 19012
rect 24308 18624 24360 18630
rect 24308 18566 24360 18572
rect 24320 18290 24348 18566
rect 24504 18426 24532 20198
rect 24492 18420 24544 18426
rect 24492 18362 24544 18368
rect 24596 18290 24624 20810
rect 24688 19854 24716 21830
rect 24768 21684 24820 21690
rect 24768 21626 24820 21632
rect 24780 21486 24808 21626
rect 24768 21480 24820 21486
rect 24768 21422 24820 21428
rect 24872 21350 24900 21950
rect 25056 21622 25084 22510
rect 25044 21616 25096 21622
rect 25044 21558 25096 21564
rect 24860 21344 24912 21350
rect 24860 21286 24912 21292
rect 24858 21176 24914 21185
rect 24858 21111 24914 21120
rect 24676 19848 24728 19854
rect 24676 19790 24728 19796
rect 24872 19334 24900 21111
rect 24952 20256 25004 20262
rect 24952 20198 25004 20204
rect 24688 19306 24900 19334
rect 24308 18284 24360 18290
rect 24308 18226 24360 18232
rect 24584 18284 24636 18290
rect 24584 18226 24636 18232
rect 24110 17980 24418 18000
rect 24110 17978 24116 17980
rect 24172 17978 24196 17980
rect 24252 17978 24276 17980
rect 24332 17978 24356 17980
rect 24412 17978 24418 17980
rect 24172 17926 24174 17978
rect 24354 17926 24356 17978
rect 24110 17924 24116 17926
rect 24172 17924 24196 17926
rect 24252 17924 24276 17926
rect 24332 17924 24356 17926
rect 24412 17924 24418 17926
rect 24110 17904 24418 17924
rect 24306 17776 24362 17785
rect 24306 17711 24308 17720
rect 24360 17711 24362 17720
rect 24400 17740 24452 17746
rect 24308 17682 24360 17688
rect 24400 17682 24452 17688
rect 24412 17626 24440 17682
rect 24412 17598 24532 17626
rect 24504 17270 24532 17598
rect 24492 17264 24544 17270
rect 24492 17206 24544 17212
rect 24110 16892 24418 16912
rect 24110 16890 24116 16892
rect 24172 16890 24196 16892
rect 24252 16890 24276 16892
rect 24332 16890 24356 16892
rect 24412 16890 24418 16892
rect 24172 16838 24174 16890
rect 24354 16838 24356 16890
rect 24110 16836 24116 16838
rect 24172 16836 24196 16838
rect 24252 16836 24276 16838
rect 24332 16836 24356 16838
rect 24412 16836 24418 16838
rect 24110 16816 24418 16836
rect 24504 16658 24532 17206
rect 24492 16652 24544 16658
rect 24492 16594 24544 16600
rect 24110 15804 24418 15824
rect 24110 15802 24116 15804
rect 24172 15802 24196 15804
rect 24252 15802 24276 15804
rect 24332 15802 24356 15804
rect 24412 15802 24418 15804
rect 24172 15750 24174 15802
rect 24354 15750 24356 15802
rect 24110 15748 24116 15750
rect 24172 15748 24196 15750
rect 24252 15748 24276 15750
rect 24332 15748 24356 15750
rect 24412 15748 24418 15750
rect 24110 15728 24418 15748
rect 24504 15638 24532 16594
rect 24688 16250 24716 19306
rect 24860 19168 24912 19174
rect 24860 19110 24912 19116
rect 24872 18358 24900 19110
rect 24964 18698 24992 20198
rect 25056 19786 25084 21558
rect 25240 21486 25268 22664
rect 25318 22672 25374 22681
rect 25424 22664 25544 22692
rect 25318 22607 25374 22616
rect 25412 22024 25464 22030
rect 25412 21966 25464 21972
rect 25228 21480 25280 21486
rect 25228 21422 25280 21428
rect 25240 21010 25268 21422
rect 25228 21004 25280 21010
rect 25228 20946 25280 20952
rect 25136 20936 25188 20942
rect 25136 20878 25188 20884
rect 25148 20534 25176 20878
rect 25136 20528 25188 20534
rect 25136 20470 25188 20476
rect 25044 19780 25096 19786
rect 25044 19722 25096 19728
rect 25056 19378 25084 19722
rect 25044 19372 25096 19378
rect 25044 19314 25096 19320
rect 24952 18692 25004 18698
rect 24952 18634 25004 18640
rect 24860 18352 24912 18358
rect 24860 18294 24912 18300
rect 24768 18284 24820 18290
rect 24768 18226 24820 18232
rect 24780 17882 24808 18226
rect 24768 17876 24820 17882
rect 24768 17818 24820 17824
rect 24768 17604 24820 17610
rect 24768 17546 24820 17552
rect 24676 16244 24728 16250
rect 24676 16186 24728 16192
rect 24584 16040 24636 16046
rect 24584 15982 24636 15988
rect 24492 15632 24544 15638
rect 24492 15574 24544 15580
rect 24110 14716 24418 14736
rect 24110 14714 24116 14716
rect 24172 14714 24196 14716
rect 24252 14714 24276 14716
rect 24332 14714 24356 14716
rect 24412 14714 24418 14716
rect 24172 14662 24174 14714
rect 24354 14662 24356 14714
rect 24110 14660 24116 14662
rect 24172 14660 24196 14662
rect 24252 14660 24276 14662
rect 24332 14660 24356 14662
rect 24412 14660 24418 14662
rect 24110 14640 24418 14660
rect 24110 13628 24418 13648
rect 24110 13626 24116 13628
rect 24172 13626 24196 13628
rect 24252 13626 24276 13628
rect 24332 13626 24356 13628
rect 24412 13626 24418 13628
rect 24172 13574 24174 13626
rect 24354 13574 24356 13626
rect 24110 13572 24116 13574
rect 24172 13572 24196 13574
rect 24252 13572 24276 13574
rect 24332 13572 24356 13574
rect 24412 13572 24418 13574
rect 24110 13552 24418 13572
rect 24596 13530 24624 15982
rect 24780 15026 24808 17546
rect 24860 16448 24912 16454
rect 24860 16390 24912 16396
rect 24872 16046 24900 16390
rect 24860 16040 24912 16046
rect 24860 15982 24912 15988
rect 24860 15360 24912 15366
rect 24860 15302 24912 15308
rect 24768 15020 24820 15026
rect 24768 14962 24820 14968
rect 24872 14414 24900 15302
rect 24964 14618 24992 18634
rect 25056 18290 25084 19314
rect 25148 18698 25176 20470
rect 25320 20460 25372 20466
rect 25320 20402 25372 20408
rect 25228 20392 25280 20398
rect 25228 20334 25280 20340
rect 25240 18873 25268 20334
rect 25332 19174 25360 20402
rect 25320 19168 25372 19174
rect 25320 19110 25372 19116
rect 25226 18864 25282 18873
rect 25226 18799 25282 18808
rect 25136 18692 25188 18698
rect 25136 18634 25188 18640
rect 25044 18284 25096 18290
rect 25044 18226 25096 18232
rect 25042 18184 25098 18193
rect 25042 18119 25098 18128
rect 25056 15162 25084 18119
rect 25148 18068 25176 18634
rect 25240 18193 25268 18799
rect 25226 18184 25282 18193
rect 25226 18119 25282 18128
rect 25148 18040 25268 18068
rect 25136 16448 25188 16454
rect 25136 16390 25188 16396
rect 25148 15434 25176 16390
rect 25136 15428 25188 15434
rect 25136 15370 25188 15376
rect 25044 15156 25096 15162
rect 25044 15098 25096 15104
rect 25148 15026 25176 15370
rect 25240 15094 25268 18040
rect 25320 17876 25372 17882
rect 25320 17818 25372 17824
rect 25228 15088 25280 15094
rect 25228 15030 25280 15036
rect 25136 15020 25188 15026
rect 25136 14962 25188 14968
rect 25044 14952 25096 14958
rect 25044 14894 25096 14900
rect 24952 14612 25004 14618
rect 24952 14554 25004 14560
rect 24860 14408 24912 14414
rect 24860 14350 24912 14356
rect 25056 13870 25084 14894
rect 25332 14550 25360 17818
rect 25320 14544 25372 14550
rect 25320 14486 25372 14492
rect 25424 13938 25452 21966
rect 25516 21962 25544 22664
rect 25688 22636 25740 22642
rect 25688 22578 25740 22584
rect 25700 22438 25728 22578
rect 25688 22432 25740 22438
rect 25688 22374 25740 22380
rect 25596 22092 25648 22098
rect 25596 22034 25648 22040
rect 25504 21956 25556 21962
rect 25504 21898 25556 21904
rect 25608 20602 25636 22034
rect 25700 21146 25728 22374
rect 26056 22228 26108 22234
rect 26056 22170 26108 22176
rect 25964 21888 26016 21894
rect 25964 21830 26016 21836
rect 25688 21140 25740 21146
rect 25688 21082 25740 21088
rect 25596 20596 25648 20602
rect 25596 20538 25648 20544
rect 25688 20392 25740 20398
rect 25688 20334 25740 20340
rect 25502 18864 25558 18873
rect 25502 18799 25504 18808
rect 25556 18799 25558 18808
rect 25504 18770 25556 18776
rect 25700 18170 25728 20334
rect 25780 20324 25832 20330
rect 25780 20266 25832 20272
rect 25792 19718 25820 20266
rect 25872 20256 25924 20262
rect 25872 20198 25924 20204
rect 25780 19712 25832 19718
rect 25780 19654 25832 19660
rect 25792 19446 25820 19654
rect 25780 19440 25832 19446
rect 25780 19382 25832 19388
rect 25700 18142 25820 18170
rect 25688 17672 25740 17678
rect 25688 17614 25740 17620
rect 25596 17536 25648 17542
rect 25596 17478 25648 17484
rect 25608 17270 25636 17478
rect 25504 17264 25556 17270
rect 25504 17206 25556 17212
rect 25596 17264 25648 17270
rect 25596 17206 25648 17212
rect 25516 16454 25544 17206
rect 25608 16522 25636 17206
rect 25700 16998 25728 17614
rect 25688 16992 25740 16998
rect 25688 16934 25740 16940
rect 25596 16516 25648 16522
rect 25596 16458 25648 16464
rect 25504 16448 25556 16454
rect 25504 16390 25556 16396
rect 25608 15502 25636 16458
rect 25596 15496 25648 15502
rect 25596 15438 25648 15444
rect 25700 15434 25728 16934
rect 25688 15428 25740 15434
rect 25688 15370 25740 15376
rect 25792 14074 25820 18142
rect 25884 14618 25912 20198
rect 25872 14612 25924 14618
rect 25872 14554 25924 14560
rect 25780 14068 25832 14074
rect 25780 14010 25832 14016
rect 25412 13932 25464 13938
rect 25412 13874 25464 13880
rect 25044 13864 25096 13870
rect 25044 13806 25096 13812
rect 24584 13524 24636 13530
rect 24584 13466 24636 13472
rect 24110 12540 24418 12560
rect 24110 12538 24116 12540
rect 24172 12538 24196 12540
rect 24252 12538 24276 12540
rect 24332 12538 24356 12540
rect 24412 12538 24418 12540
rect 24172 12486 24174 12538
rect 24354 12486 24356 12538
rect 24110 12484 24116 12486
rect 24172 12484 24196 12486
rect 24252 12484 24276 12486
rect 24332 12484 24356 12486
rect 24412 12484 24418 12486
rect 24110 12464 24418 12484
rect 25056 12434 25084 13806
rect 25976 13258 26004 21830
rect 26068 20806 26096 22170
rect 26146 21856 26202 21865
rect 26146 21791 26202 21800
rect 26160 21486 26188 21791
rect 26148 21480 26200 21486
rect 26148 21422 26200 21428
rect 26240 21480 26292 21486
rect 26240 21422 26292 21428
rect 26252 20942 26280 21422
rect 26240 20936 26292 20942
rect 26240 20878 26292 20884
rect 26056 20800 26108 20806
rect 26056 20742 26108 20748
rect 26068 19514 26096 20742
rect 26436 20534 26464 25706
rect 26516 25220 26568 25226
rect 26516 25162 26568 25168
rect 26528 24993 26556 25162
rect 26514 24984 26570 24993
rect 26514 24919 26570 24928
rect 26620 24818 26648 29271
rect 26792 29242 26844 29248
rect 26896 29170 26924 30126
rect 26884 29164 26936 29170
rect 26936 29124 27016 29152
rect 26884 29106 26936 29112
rect 26988 28014 27016 29124
rect 26976 28008 27028 28014
rect 26976 27950 27028 27956
rect 27080 27878 27108 30194
rect 27252 30048 27304 30054
rect 27252 29990 27304 29996
rect 27264 29170 27292 29990
rect 27252 29164 27304 29170
rect 27252 29106 27304 29112
rect 27632 28966 27660 31282
rect 27620 28960 27672 28966
rect 27620 28902 27672 28908
rect 27620 28756 27672 28762
rect 27620 28698 27672 28704
rect 27436 28144 27488 28150
rect 27436 28086 27488 28092
rect 27068 27872 27120 27878
rect 27068 27814 27120 27820
rect 27080 25974 27108 27814
rect 27344 27124 27396 27130
rect 27344 27066 27396 27072
rect 27356 26042 27384 27066
rect 27448 26994 27476 28086
rect 27632 28082 27660 28698
rect 27620 28076 27672 28082
rect 27620 28018 27672 28024
rect 27436 26988 27488 26994
rect 27436 26930 27488 26936
rect 27448 26489 27476 26930
rect 27434 26480 27490 26489
rect 27434 26415 27490 26424
rect 27632 26042 27660 28018
rect 27344 26036 27396 26042
rect 27344 25978 27396 25984
rect 27620 26036 27672 26042
rect 27620 25978 27672 25984
rect 27068 25968 27120 25974
rect 27068 25910 27120 25916
rect 26608 24812 26660 24818
rect 26608 24754 26660 24760
rect 26976 24812 27028 24818
rect 26976 24754 27028 24760
rect 26516 24676 26568 24682
rect 26516 24618 26568 24624
rect 26424 20528 26476 20534
rect 26424 20470 26476 20476
rect 26436 20398 26464 20470
rect 26424 20392 26476 20398
rect 26424 20334 26476 20340
rect 26528 19922 26556 24618
rect 26988 23866 27016 24754
rect 27160 24608 27212 24614
rect 27160 24550 27212 24556
rect 27252 24608 27304 24614
rect 27252 24550 27304 24556
rect 26608 23860 26660 23866
rect 26608 23802 26660 23808
rect 26976 23860 27028 23866
rect 26976 23802 27028 23808
rect 26620 20534 26648 23802
rect 27172 23730 27200 24550
rect 27160 23724 27212 23730
rect 27160 23666 27212 23672
rect 27264 23662 27292 24550
rect 27252 23656 27304 23662
rect 27252 23598 27304 23604
rect 27160 23180 27212 23186
rect 27160 23122 27212 23128
rect 27068 22976 27120 22982
rect 27068 22918 27120 22924
rect 26974 22808 27030 22817
rect 26974 22743 27030 22752
rect 26988 21690 27016 22743
rect 27080 22574 27108 22918
rect 27068 22568 27120 22574
rect 27068 22510 27120 22516
rect 26976 21684 27028 21690
rect 26976 21626 27028 21632
rect 27068 21412 27120 21418
rect 27068 21354 27120 21360
rect 26792 20868 26844 20874
rect 26792 20810 26844 20816
rect 26608 20528 26660 20534
rect 26608 20470 26660 20476
rect 26516 19916 26568 19922
rect 26516 19858 26568 19864
rect 26056 19508 26108 19514
rect 26056 19450 26108 19456
rect 26620 19174 26648 20470
rect 26424 19168 26476 19174
rect 26424 19110 26476 19116
rect 26608 19168 26660 19174
rect 26608 19110 26660 19116
rect 26332 18760 26384 18766
rect 26332 18702 26384 18708
rect 26240 18692 26292 18698
rect 26240 18634 26292 18640
rect 26056 18284 26108 18290
rect 26056 18226 26108 18232
rect 26068 13530 26096 18226
rect 26148 17060 26200 17066
rect 26148 17002 26200 17008
rect 26160 16590 26188 17002
rect 26148 16584 26200 16590
rect 26148 16526 26200 16532
rect 26148 16040 26200 16046
rect 26148 15982 26200 15988
rect 26160 15745 26188 15982
rect 26146 15736 26202 15745
rect 26146 15671 26202 15680
rect 26252 15162 26280 18634
rect 26344 17882 26372 18702
rect 26436 18222 26464 19110
rect 26424 18216 26476 18222
rect 26424 18158 26476 18164
rect 26332 17876 26384 17882
rect 26332 17818 26384 17824
rect 26332 16584 26384 16590
rect 26332 16526 26384 16532
rect 26344 15638 26372 16526
rect 26332 15632 26384 15638
rect 26332 15574 26384 15580
rect 26332 15496 26384 15502
rect 26332 15438 26384 15444
rect 26240 15156 26292 15162
rect 26240 15098 26292 15104
rect 26056 13524 26108 13530
rect 26056 13466 26108 13472
rect 25964 13252 26016 13258
rect 25964 13194 26016 13200
rect 26344 12850 26372 15438
rect 26436 14550 26464 18158
rect 26700 16992 26752 16998
rect 26700 16934 26752 16940
rect 26516 15428 26568 15434
rect 26516 15370 26568 15376
rect 26528 15162 26556 15370
rect 26516 15156 26568 15162
rect 26516 15098 26568 15104
rect 26424 14544 26476 14550
rect 26424 14486 26476 14492
rect 26712 13326 26740 16934
rect 26700 13320 26752 13326
rect 26700 13262 26752 13268
rect 26332 12844 26384 12850
rect 26332 12786 26384 12792
rect 26804 12782 26832 20810
rect 26884 19372 26936 19378
rect 26884 19314 26936 19320
rect 26896 18426 26924 19314
rect 26884 18420 26936 18426
rect 26884 18362 26936 18368
rect 27080 18086 27108 21354
rect 26976 18080 27028 18086
rect 26976 18022 27028 18028
rect 27068 18080 27120 18086
rect 27068 18022 27120 18028
rect 26988 17134 27016 18022
rect 27068 17604 27120 17610
rect 27068 17546 27120 17552
rect 26976 17128 27028 17134
rect 26976 17070 27028 17076
rect 26884 16516 26936 16522
rect 26884 16458 26936 16464
rect 26896 14074 26924 16458
rect 26884 14068 26936 14074
rect 26884 14010 26936 14016
rect 26988 13938 27016 17070
rect 27080 15162 27108 17546
rect 27068 15156 27120 15162
rect 27068 15098 27120 15104
rect 26976 13932 27028 13938
rect 26976 13874 27028 13880
rect 27172 13530 27200 23122
rect 27724 22642 27752 33254
rect 27816 27062 27844 35226
rect 27908 27130 27936 36518
rect 28184 36242 28212 36751
rect 28172 36236 28224 36242
rect 28172 36178 28224 36184
rect 28170 35456 28226 35465
rect 28170 35391 28226 35400
rect 27988 35216 28040 35222
rect 27988 35158 28040 35164
rect 28000 32434 28028 35158
rect 28184 35154 28212 35391
rect 28172 35148 28224 35154
rect 28172 35090 28224 35096
rect 28276 34762 28304 39471
rect 28368 36854 28396 41200
rect 28906 39536 28962 39545
rect 28906 39471 28962 39480
rect 28356 36848 28408 36854
rect 28356 36790 28408 36796
rect 28356 36712 28408 36718
rect 28356 36654 28408 36660
rect 28184 34734 28304 34762
rect 28080 34604 28132 34610
rect 28080 34546 28132 34552
rect 27988 32428 28040 32434
rect 27988 32370 28040 32376
rect 27896 27124 27948 27130
rect 27896 27066 27948 27072
rect 27804 27056 27856 27062
rect 27804 26998 27856 27004
rect 28000 23730 28028 32370
rect 28092 31482 28120 34546
rect 28184 33522 28212 34734
rect 28264 34604 28316 34610
rect 28264 34546 28316 34552
rect 28172 33516 28224 33522
rect 28172 33458 28224 33464
rect 28170 33416 28226 33425
rect 28170 33351 28226 33360
rect 28184 32978 28212 33351
rect 28172 32972 28224 32978
rect 28172 32914 28224 32920
rect 28170 32736 28226 32745
rect 28170 32671 28226 32680
rect 28184 31890 28212 32671
rect 28172 31884 28224 31890
rect 28172 31826 28224 31832
rect 28080 31476 28132 31482
rect 28080 31418 28132 31424
rect 28092 30938 28120 31418
rect 28276 31346 28304 34546
rect 28368 33046 28396 36654
rect 28448 34536 28500 34542
rect 28448 34478 28500 34484
rect 28356 33040 28408 33046
rect 28356 32982 28408 32988
rect 28264 31340 28316 31346
rect 28264 31282 28316 31288
rect 28080 30932 28132 30938
rect 28080 30874 28132 30880
rect 28276 29782 28304 31282
rect 28264 29776 28316 29782
rect 28264 29718 28316 29724
rect 28170 29336 28226 29345
rect 28170 29271 28226 29280
rect 28184 28626 28212 29271
rect 28172 28620 28224 28626
rect 28172 28562 28224 28568
rect 28078 28384 28134 28393
rect 28078 28319 28134 28328
rect 28092 28218 28120 28319
rect 28080 28212 28132 28218
rect 28132 28172 28304 28200
rect 28080 28154 28132 28160
rect 28172 27396 28224 27402
rect 28172 27338 28224 27344
rect 28184 27305 28212 27338
rect 28170 27296 28226 27305
rect 28170 27231 28226 27240
rect 28170 26616 28226 26625
rect 28170 26551 28226 26560
rect 28184 26450 28212 26551
rect 28172 26444 28224 26450
rect 28172 26386 28224 26392
rect 28170 25936 28226 25945
rect 28170 25871 28226 25880
rect 28184 25362 28212 25871
rect 28172 25356 28224 25362
rect 28172 25298 28224 25304
rect 28170 24576 28226 24585
rect 28170 24511 28226 24520
rect 28184 24274 28212 24511
rect 28172 24268 28224 24274
rect 28172 24210 28224 24216
rect 28080 24132 28132 24138
rect 28080 24074 28132 24080
rect 28092 23866 28120 24074
rect 28080 23860 28132 23866
rect 28080 23802 28132 23808
rect 27988 23724 28040 23730
rect 27988 23666 28040 23672
rect 27712 22636 27764 22642
rect 27712 22578 27764 22584
rect 28170 22536 28226 22545
rect 28170 22471 28226 22480
rect 27252 22432 27304 22438
rect 27252 22374 27304 22380
rect 27436 22432 27488 22438
rect 27436 22374 27488 22380
rect 27528 22432 27580 22438
rect 27528 22374 27580 22380
rect 27264 21486 27292 22374
rect 27344 21616 27396 21622
rect 27344 21558 27396 21564
rect 27252 21480 27304 21486
rect 27252 21422 27304 21428
rect 27252 21344 27304 21350
rect 27252 21286 27304 21292
rect 27264 19174 27292 21286
rect 27356 19378 27384 21558
rect 27448 21078 27476 22374
rect 27436 21072 27488 21078
rect 27436 21014 27488 21020
rect 27540 21010 27568 22374
rect 28184 22098 28212 22471
rect 28172 22092 28224 22098
rect 28172 22034 28224 22040
rect 27712 21888 27764 21894
rect 27712 21830 27764 21836
rect 27620 21344 27672 21350
rect 27620 21286 27672 21292
rect 27528 21004 27580 21010
rect 27528 20946 27580 20952
rect 27436 19780 27488 19786
rect 27436 19722 27488 19728
rect 27344 19372 27396 19378
rect 27344 19314 27396 19320
rect 27252 19168 27304 19174
rect 27252 19110 27304 19116
rect 27264 18902 27292 19110
rect 27252 18896 27304 18902
rect 27252 18838 27304 18844
rect 27344 18080 27396 18086
rect 27344 18022 27396 18028
rect 27356 16998 27384 18022
rect 27344 16992 27396 16998
rect 27344 16934 27396 16940
rect 27344 16176 27396 16182
rect 27344 16118 27396 16124
rect 27252 15020 27304 15026
rect 27252 14962 27304 14968
rect 27264 13938 27292 14962
rect 27252 13932 27304 13938
rect 27252 13874 27304 13880
rect 27160 13524 27212 13530
rect 27160 13466 27212 13472
rect 26792 12776 26844 12782
rect 26792 12718 26844 12724
rect 27264 12434 27292 13874
rect 27356 13530 27384 16118
rect 27344 13524 27396 13530
rect 27344 13466 27396 13472
rect 27448 12850 27476 19722
rect 27632 18290 27660 21286
rect 27724 20602 27752 21830
rect 27896 21548 27948 21554
rect 27896 21490 27948 21496
rect 27712 20596 27764 20602
rect 27712 20538 27764 20544
rect 27908 19961 27936 21490
rect 28170 21176 28226 21185
rect 28170 21111 28226 21120
rect 28184 21010 28212 21111
rect 28172 21004 28224 21010
rect 28172 20946 28224 20952
rect 27894 19952 27950 19961
rect 27894 19887 27950 19896
rect 28172 19848 28224 19854
rect 28170 19816 28172 19825
rect 28224 19816 28226 19825
rect 28170 19751 28226 19760
rect 28170 19136 28226 19145
rect 28170 19071 28226 19080
rect 27712 18964 27764 18970
rect 27712 18906 27764 18912
rect 27620 18284 27672 18290
rect 27620 18226 27672 18232
rect 27620 18148 27672 18154
rect 27620 18090 27672 18096
rect 27528 17128 27580 17134
rect 27528 17070 27580 17076
rect 27540 15706 27568 17070
rect 27528 15700 27580 15706
rect 27528 15642 27580 15648
rect 27632 13394 27660 18090
rect 27620 13388 27672 13394
rect 27620 13330 27672 13336
rect 27436 12844 27488 12850
rect 27436 12786 27488 12792
rect 20732 12406 21128 12434
rect 21376 12406 21496 12434
rect 23032 12406 23152 12434
rect 23768 12406 24072 12434
rect 24872 12406 25084 12434
rect 27172 12406 27292 12434
rect 19984 3664 20036 3670
rect 19984 3606 20036 3612
rect 19996 3534 20024 3606
rect 20732 3602 20760 12406
rect 21376 8430 21404 12406
rect 21364 8424 21416 8430
rect 21364 8366 21416 8372
rect 22192 3936 22244 3942
rect 22192 3878 22244 3884
rect 20720 3596 20772 3602
rect 20720 3538 20772 3544
rect 18880 3528 18932 3534
rect 18880 3470 18932 3476
rect 19984 3528 20036 3534
rect 19984 3470 20036 3476
rect 20168 3528 20220 3534
rect 20168 3470 20220 3476
rect 21916 3528 21968 3534
rect 21916 3470 21968 3476
rect 18236 3460 18288 3466
rect 18236 3402 18288 3408
rect 18248 3058 18276 3402
rect 18892 3058 18920 3470
rect 20076 3392 20128 3398
rect 20076 3334 20128 3340
rect 19478 3292 19786 3312
rect 19478 3290 19484 3292
rect 19540 3290 19564 3292
rect 19620 3290 19644 3292
rect 19700 3290 19724 3292
rect 19780 3290 19786 3292
rect 19540 3238 19542 3290
rect 19722 3238 19724 3290
rect 19478 3236 19484 3238
rect 19540 3236 19564 3238
rect 19620 3236 19644 3238
rect 19700 3236 19724 3238
rect 19780 3236 19786 3238
rect 19478 3216 19786 3236
rect 18236 3052 18288 3058
rect 18236 2994 18288 3000
rect 18880 3052 18932 3058
rect 18880 2994 18932 3000
rect 19340 2984 19392 2990
rect 19340 2926 19392 2932
rect 18696 2576 18748 2582
rect 18696 2518 18748 2524
rect 18708 800 18736 2518
rect 19352 800 19380 2926
rect 20088 2514 20116 3334
rect 20076 2508 20128 2514
rect 20076 2450 20128 2456
rect 20180 2378 20208 3470
rect 21928 3058 21956 3470
rect 22100 3392 22152 3398
rect 22100 3334 22152 3340
rect 22112 3126 22140 3334
rect 22100 3120 22152 3126
rect 22100 3062 22152 3068
rect 21916 3052 21968 3058
rect 21916 2994 21968 3000
rect 22204 2514 22232 3878
rect 23032 3534 23060 12406
rect 23768 11762 23796 12406
rect 23756 11756 23808 11762
rect 23756 11698 23808 11704
rect 24110 11452 24418 11472
rect 24110 11450 24116 11452
rect 24172 11450 24196 11452
rect 24252 11450 24276 11452
rect 24332 11450 24356 11452
rect 24412 11450 24418 11452
rect 24172 11398 24174 11450
rect 24354 11398 24356 11450
rect 24110 11396 24116 11398
rect 24172 11396 24196 11398
rect 24252 11396 24276 11398
rect 24332 11396 24356 11398
rect 24412 11396 24418 11398
rect 24110 11376 24418 11396
rect 24110 10364 24418 10384
rect 24110 10362 24116 10364
rect 24172 10362 24196 10364
rect 24252 10362 24276 10364
rect 24332 10362 24356 10364
rect 24412 10362 24418 10364
rect 24172 10310 24174 10362
rect 24354 10310 24356 10362
rect 24110 10308 24116 10310
rect 24172 10308 24196 10310
rect 24252 10308 24276 10310
rect 24332 10308 24356 10310
rect 24412 10308 24418 10310
rect 24110 10288 24418 10308
rect 24872 9654 24900 12406
rect 26332 12232 26384 12238
rect 26332 12174 26384 12180
rect 26344 11218 26372 12174
rect 26516 11552 26568 11558
rect 26516 11494 26568 11500
rect 26528 11218 26556 11494
rect 26332 11212 26384 11218
rect 26332 11154 26384 11160
rect 26516 11212 26568 11218
rect 26516 11154 26568 11160
rect 26332 10056 26384 10062
rect 26332 9998 26384 10004
rect 24860 9648 24912 9654
rect 24860 9590 24912 9596
rect 26344 9586 26372 9998
rect 26332 9580 26384 9586
rect 26332 9522 26384 9528
rect 24110 9276 24418 9296
rect 24110 9274 24116 9276
rect 24172 9274 24196 9276
rect 24252 9274 24276 9276
rect 24332 9274 24356 9276
rect 24412 9274 24418 9276
rect 24172 9222 24174 9274
rect 24354 9222 24356 9274
rect 24110 9220 24116 9222
rect 24172 9220 24196 9222
rect 24252 9220 24276 9222
rect 24332 9220 24356 9222
rect 24412 9220 24418 9222
rect 24110 9200 24418 9220
rect 24110 8188 24418 8208
rect 24110 8186 24116 8188
rect 24172 8186 24196 8188
rect 24252 8186 24276 8188
rect 24332 8186 24356 8188
rect 24412 8186 24418 8188
rect 24172 8134 24174 8186
rect 24354 8134 24356 8186
rect 24110 8132 24116 8134
rect 24172 8132 24196 8134
rect 24252 8132 24276 8134
rect 24332 8132 24356 8134
rect 24412 8132 24418 8134
rect 24110 8112 24418 8132
rect 24110 7100 24418 7120
rect 24110 7098 24116 7100
rect 24172 7098 24196 7100
rect 24252 7098 24276 7100
rect 24332 7098 24356 7100
rect 24412 7098 24418 7100
rect 24172 7046 24174 7098
rect 24354 7046 24356 7098
rect 24110 7044 24116 7046
rect 24172 7044 24196 7046
rect 24252 7044 24276 7046
rect 24332 7044 24356 7046
rect 24412 7044 24418 7046
rect 24110 7024 24418 7044
rect 27172 6914 27200 12406
rect 27344 10464 27396 10470
rect 27344 10406 27396 10412
rect 27356 9110 27384 10406
rect 27436 9988 27488 9994
rect 27436 9930 27488 9936
rect 27344 9104 27396 9110
rect 27344 9046 27396 9052
rect 27252 8288 27304 8294
rect 27252 8230 27304 8236
rect 27264 7954 27292 8230
rect 27252 7948 27304 7954
rect 27252 7890 27304 7896
rect 27252 7200 27304 7206
rect 27252 7142 27304 7148
rect 27080 6886 27200 6914
rect 24584 6248 24636 6254
rect 24584 6190 24636 6196
rect 24952 6248 25004 6254
rect 24952 6190 25004 6196
rect 26056 6248 26108 6254
rect 26056 6190 26108 6196
rect 24110 6012 24418 6032
rect 24110 6010 24116 6012
rect 24172 6010 24196 6012
rect 24252 6010 24276 6012
rect 24332 6010 24356 6012
rect 24412 6010 24418 6012
rect 24172 5958 24174 6010
rect 24354 5958 24356 6010
rect 24110 5956 24116 5958
rect 24172 5956 24196 5958
rect 24252 5956 24276 5958
rect 24332 5956 24356 5958
rect 24412 5956 24418 5958
rect 24110 5936 24418 5956
rect 24596 5914 24624 6190
rect 24584 5908 24636 5914
rect 24584 5850 24636 5856
rect 24860 5704 24912 5710
rect 24860 5646 24912 5652
rect 24872 5166 24900 5646
rect 24964 5370 24992 6190
rect 24952 5364 25004 5370
rect 24952 5306 25004 5312
rect 24860 5160 24912 5166
rect 24860 5102 24912 5108
rect 24110 4924 24418 4944
rect 24110 4922 24116 4924
rect 24172 4922 24196 4924
rect 24252 4922 24276 4924
rect 24332 4922 24356 4924
rect 24412 4922 24418 4924
rect 24172 4870 24174 4922
rect 24354 4870 24356 4922
rect 24110 4868 24116 4870
rect 24172 4868 24196 4870
rect 24252 4868 24276 4870
rect 24332 4868 24356 4870
rect 24412 4868 24418 4870
rect 24110 4848 24418 4868
rect 26068 4865 26096 6190
rect 26516 6112 26568 6118
rect 26516 6054 26568 6060
rect 26528 5778 26556 6054
rect 26516 5772 26568 5778
rect 26516 5714 26568 5720
rect 26148 5160 26200 5166
rect 26148 5102 26200 5108
rect 26054 4856 26110 4865
rect 26054 4791 26110 4800
rect 23848 4616 23900 4622
rect 23848 4558 23900 4564
rect 23480 4072 23532 4078
rect 23480 4014 23532 4020
rect 23112 4004 23164 4010
rect 23112 3946 23164 3952
rect 23124 3738 23152 3946
rect 23492 3738 23520 4014
rect 23112 3732 23164 3738
rect 23112 3674 23164 3680
rect 23480 3732 23532 3738
rect 23480 3674 23532 3680
rect 23020 3528 23072 3534
rect 23020 3470 23072 3476
rect 23756 3392 23808 3398
rect 23756 3334 23808 3340
rect 22560 2984 22612 2990
rect 22560 2926 22612 2932
rect 22192 2508 22244 2514
rect 22192 2450 22244 2456
rect 20168 2372 20220 2378
rect 20168 2314 20220 2320
rect 19478 2204 19786 2224
rect 19478 2202 19484 2204
rect 19540 2202 19564 2204
rect 19620 2202 19644 2204
rect 19700 2202 19724 2204
rect 19780 2202 19786 2204
rect 19540 2150 19542 2202
rect 19722 2150 19724 2202
rect 19478 2148 19484 2150
rect 19540 2148 19564 2150
rect 19620 2148 19644 2150
rect 19700 2148 19724 2150
rect 19780 2148 19786 2150
rect 19478 2128 19786 2148
rect 22572 800 22600 2926
rect 23768 2378 23796 3334
rect 23860 2514 23888 4558
rect 24860 4548 24912 4554
rect 24860 4490 24912 4496
rect 24872 4146 24900 4490
rect 24952 4480 25004 4486
rect 24952 4422 25004 4428
rect 24860 4140 24912 4146
rect 24860 4082 24912 4088
rect 24110 3836 24418 3856
rect 24110 3834 24116 3836
rect 24172 3834 24196 3836
rect 24252 3834 24276 3836
rect 24332 3834 24356 3836
rect 24412 3834 24418 3836
rect 24172 3782 24174 3834
rect 24354 3782 24356 3834
rect 24110 3780 24116 3782
rect 24172 3780 24196 3782
rect 24252 3780 24276 3782
rect 24332 3780 24356 3782
rect 24412 3780 24418 3782
rect 24110 3760 24418 3780
rect 24872 3670 24900 4082
rect 24860 3664 24912 3670
rect 24860 3606 24912 3612
rect 24964 3534 24992 4422
rect 26160 4185 26188 5102
rect 26146 4176 26202 4185
rect 26146 4111 26202 4120
rect 25136 3936 25188 3942
rect 25136 3878 25188 3884
rect 25148 3602 25176 3878
rect 25136 3596 25188 3602
rect 25136 3538 25188 3544
rect 26148 3596 26200 3602
rect 26148 3538 26200 3544
rect 24952 3528 25004 3534
rect 24952 3470 25004 3476
rect 26056 3052 26108 3058
rect 26056 2994 26108 3000
rect 24584 2984 24636 2990
rect 25504 2984 25556 2990
rect 24636 2944 24716 2972
rect 24584 2926 24636 2932
rect 24688 2938 24716 2944
rect 24688 2922 24808 2938
rect 25240 2932 25504 2938
rect 25240 2926 25556 2932
rect 25240 2922 25544 2926
rect 24688 2916 24820 2922
rect 24688 2910 24768 2916
rect 24768 2858 24820 2864
rect 25228 2916 25544 2922
rect 25280 2910 25544 2916
rect 25228 2858 25280 2864
rect 25044 2848 25096 2854
rect 25044 2790 25096 2796
rect 24110 2748 24418 2768
rect 24110 2746 24116 2748
rect 24172 2746 24196 2748
rect 24252 2746 24276 2748
rect 24332 2746 24356 2748
rect 24412 2746 24418 2748
rect 24172 2694 24174 2746
rect 24354 2694 24356 2746
rect 24110 2692 24116 2694
rect 24172 2692 24196 2694
rect 24252 2692 24276 2694
rect 24332 2692 24356 2694
rect 24412 2692 24418 2694
rect 24110 2672 24418 2692
rect 23848 2508 23900 2514
rect 23848 2450 23900 2456
rect 25056 2378 25084 2790
rect 23756 2372 23808 2378
rect 23756 2314 23808 2320
rect 25044 2372 25096 2378
rect 25044 2314 25096 2320
rect 26068 2145 26096 2994
rect 26160 2825 26188 3538
rect 26516 2984 26568 2990
rect 26516 2926 26568 2932
rect 26146 2816 26202 2825
rect 26146 2751 26202 2760
rect 26528 2650 26556 2926
rect 26516 2644 26568 2650
rect 26516 2586 26568 2592
rect 27080 2582 27108 6886
rect 27264 6866 27292 7142
rect 27252 6860 27304 6866
rect 27252 6802 27304 6808
rect 27160 5228 27212 5234
rect 27160 5170 27212 5176
rect 27172 4146 27200 5170
rect 27160 4140 27212 4146
rect 27160 4082 27212 4088
rect 27448 3505 27476 9930
rect 27724 9586 27752 18906
rect 28184 18834 28212 19071
rect 28172 18828 28224 18834
rect 28172 18770 28224 18776
rect 28170 18456 28226 18465
rect 28170 18391 28226 18400
rect 27804 18352 27856 18358
rect 27804 18294 27856 18300
rect 27816 14958 27844 18294
rect 27988 18080 28040 18086
rect 27988 18022 28040 18028
rect 28000 17202 28028 18022
rect 28184 17746 28212 18391
rect 28276 18222 28304 28172
rect 28460 23254 28488 34478
rect 28920 34066 28948 39471
rect 28908 34060 28960 34066
rect 28908 34002 28960 34008
rect 28722 32056 28778 32065
rect 28722 31991 28778 32000
rect 28736 30802 28764 31991
rect 28724 30796 28776 30802
rect 28724 30738 28776 30744
rect 28632 29028 28684 29034
rect 28632 28970 28684 28976
rect 28540 24812 28592 24818
rect 28540 24754 28592 24760
rect 28448 23248 28500 23254
rect 28448 23190 28500 23196
rect 28356 22636 28408 22642
rect 28356 22578 28408 22584
rect 28264 18216 28316 18222
rect 28264 18158 28316 18164
rect 28172 17740 28224 17746
rect 28172 17682 28224 17688
rect 27988 17196 28040 17202
rect 27988 17138 28040 17144
rect 28172 16516 28224 16522
rect 28172 16458 28224 16464
rect 28184 16425 28212 16458
rect 28170 16416 28226 16425
rect 28170 16351 28226 16360
rect 27988 16108 28040 16114
rect 27988 16050 28040 16056
rect 27804 14952 27856 14958
rect 27804 14894 27856 14900
rect 28000 14822 28028 16050
rect 28276 15978 28304 18158
rect 28264 15972 28316 15978
rect 28264 15914 28316 15920
rect 28172 15428 28224 15434
rect 28172 15370 28224 15376
rect 28184 15065 28212 15370
rect 28170 15056 28226 15065
rect 28170 14991 28226 15000
rect 27988 14816 28040 14822
rect 27988 14758 28040 14764
rect 28080 14476 28132 14482
rect 28080 14418 28132 14424
rect 27804 14340 27856 14346
rect 27804 14282 27856 14288
rect 27816 14074 27844 14282
rect 27804 14068 27856 14074
rect 27804 14010 27856 14016
rect 27804 13864 27856 13870
rect 27804 13806 27856 13812
rect 27816 13326 27844 13806
rect 27804 13320 27856 13326
rect 27804 13262 27856 13268
rect 28092 12442 28120 14418
rect 28170 14376 28226 14385
rect 28170 14311 28172 14320
rect 28224 14311 28226 14320
rect 28172 14282 28224 14288
rect 28080 12436 28132 12442
rect 28080 12378 28132 12384
rect 27988 11756 28040 11762
rect 27988 11698 28040 11704
rect 28000 11665 28028 11698
rect 27986 11656 28042 11665
rect 27986 11591 28042 11600
rect 28172 11076 28224 11082
rect 28172 11018 28224 11024
rect 28184 10985 28212 11018
rect 28170 10976 28226 10985
rect 28170 10911 28226 10920
rect 27896 10464 27948 10470
rect 27896 10406 27948 10412
rect 27908 10130 27936 10406
rect 27896 10124 27948 10130
rect 27896 10066 27948 10072
rect 28170 9616 28226 9625
rect 27712 9580 27764 9586
rect 28170 9551 28226 9560
rect 27712 9522 27764 9528
rect 27804 9376 27856 9382
rect 27804 9318 27856 9324
rect 27816 9042 27844 9318
rect 28184 9042 28212 9551
rect 27804 9036 27856 9042
rect 27804 8978 27856 8984
rect 28172 9036 28224 9042
rect 28172 8978 28224 8984
rect 27988 8424 28040 8430
rect 27988 8366 28040 8372
rect 27620 8356 27672 8362
rect 27620 8298 27672 8304
rect 27632 5846 27660 8298
rect 27804 7812 27856 7818
rect 27804 7754 27856 7760
rect 27816 7546 27844 7754
rect 27804 7540 27856 7546
rect 27804 7482 27856 7488
rect 27712 7404 27764 7410
rect 27712 7346 27764 7352
rect 27620 5840 27672 5846
rect 27620 5782 27672 5788
rect 27724 5098 27752 7346
rect 27896 6724 27948 6730
rect 27896 6666 27948 6672
rect 27908 6458 27936 6666
rect 27896 6452 27948 6458
rect 27896 6394 27948 6400
rect 27804 6180 27856 6186
rect 27804 6122 27856 6128
rect 27712 5092 27764 5098
rect 27712 5034 27764 5040
rect 27712 4548 27764 4554
rect 27712 4490 27764 4496
rect 27434 3496 27490 3505
rect 27434 3431 27490 3440
rect 27724 3194 27752 4490
rect 27712 3188 27764 3194
rect 27712 3130 27764 3136
rect 27816 3058 27844 6122
rect 28000 5234 28028 8366
rect 28172 7812 28224 7818
rect 28172 7754 28224 7760
rect 28184 7585 28212 7754
rect 28170 7576 28226 7585
rect 28170 7511 28226 7520
rect 28368 6914 28396 22578
rect 28552 15094 28580 24754
rect 28644 23769 28672 28970
rect 28722 25256 28778 25265
rect 28722 25191 28778 25200
rect 28630 23760 28686 23769
rect 28630 23695 28686 23704
rect 28736 23186 28764 25191
rect 28724 23180 28776 23186
rect 28724 23122 28776 23128
rect 28540 15088 28592 15094
rect 28540 15030 28592 15036
rect 28170 6896 28226 6905
rect 28170 6831 28172 6840
rect 28224 6831 28226 6840
rect 28276 6886 28396 6914
rect 28172 6802 28224 6808
rect 28170 6216 28226 6225
rect 28170 6151 28226 6160
rect 28184 5778 28212 6151
rect 28172 5772 28224 5778
rect 28172 5714 28224 5720
rect 27988 5228 28040 5234
rect 27988 5170 28040 5176
rect 28000 3534 28028 5170
rect 28276 4146 28304 6886
rect 28356 4548 28408 4554
rect 28356 4490 28408 4496
rect 28264 4140 28316 4146
rect 28264 4082 28316 4088
rect 27988 3528 28040 3534
rect 27988 3470 28040 3476
rect 27804 3052 27856 3058
rect 27804 2994 27856 3000
rect 27068 2576 27120 2582
rect 27068 2518 27120 2524
rect 28000 2446 28028 3470
rect 27988 2440 28040 2446
rect 27988 2382 28040 2388
rect 26148 2372 26200 2378
rect 26148 2314 26200 2320
rect 26054 2136 26110 2145
rect 26054 2071 26110 2080
rect -10 0 102 800
rect 634 0 746 800
rect 1278 0 1390 800
rect 1922 0 2034 800
rect 2566 0 2678 800
rect 3210 0 3322 800
rect 3854 0 3966 800
rect 4498 0 4610 800
rect 5142 0 5254 800
rect 5786 0 5898 800
rect 6430 0 6542 800
rect 7074 0 7186 800
rect 7718 0 7830 800
rect 8362 0 8474 800
rect 9006 0 9118 800
rect 9650 0 9762 800
rect 10294 0 10406 800
rect 10938 0 11050 800
rect 11582 0 11694 800
rect 12226 0 12338 800
rect 12870 0 12982 800
rect 13514 0 13626 800
rect 14158 0 14270 800
rect 14802 0 14914 800
rect 15446 0 15558 800
rect 16090 0 16202 800
rect 16734 0 16846 800
rect 17378 0 17490 800
rect 18022 0 18134 800
rect 18666 0 18778 800
rect 19310 0 19422 800
rect 19954 0 20066 800
rect 20598 0 20710 800
rect 21242 0 21354 800
rect 21886 0 21998 800
rect 22530 0 22642 800
rect 23818 0 23930 800
rect 24462 0 24574 800
rect 25106 0 25218 800
rect 25750 0 25862 800
rect 26160 105 26188 2314
rect 28368 800 28396 4490
rect 29000 4004 29052 4010
rect 29000 3946 29052 3952
rect 29012 800 29040 3946
rect 29644 2848 29696 2854
rect 29644 2790 29696 2796
rect 29656 800 29684 2790
rect 26146 96 26202 105
rect 26146 31 26202 40
rect 26394 0 26506 800
rect 27038 0 27150 800
rect 27682 0 27794 800
rect 28326 0 28438 800
rect 28970 0 29082 800
rect 29614 0 29726 800
<< via2 >>
rect 1766 39480 1822 39536
rect 1398 33360 1454 33416
rect 2778 40160 2834 40216
rect 2870 39344 2926 39400
rect 2778 38120 2834 38176
rect 1858 37440 1914 37496
rect 1858 17076 1860 17096
rect 1860 17076 1912 17096
rect 1912 17076 1914 17096
rect 1858 17040 1914 17076
rect 1858 14320 1914 14376
rect 1858 10920 1914 10976
rect 1858 5480 1914 5536
rect 2778 34720 2834 34776
rect 2778 34060 2834 34096
rect 2778 34040 2780 34060
rect 2780 34040 2832 34060
rect 2832 34040 2834 34060
rect 2870 32680 2926 32736
rect 2778 31320 2834 31376
rect 2778 29280 2834 29336
rect 2778 23180 2834 23216
rect 2778 23160 2780 23180
rect 2780 23160 2832 23180
rect 2832 23160 2834 23180
rect 2778 17740 2834 17776
rect 2778 17720 2780 17740
rect 2780 17720 2832 17740
rect 2832 17720 2834 17740
rect 2778 15680 2834 15736
rect 2778 12960 2834 13016
rect 2778 12300 2834 12336
rect 2778 12280 2780 12300
rect 2780 12280 2832 12300
rect 2832 12280 2834 12300
rect 4066 36080 4122 36136
rect 7102 39888 7158 39944
rect 5588 39738 5644 39740
rect 5668 39738 5724 39740
rect 5748 39738 5804 39740
rect 5828 39738 5884 39740
rect 5588 39686 5634 39738
rect 5634 39686 5644 39738
rect 5668 39686 5698 39738
rect 5698 39686 5710 39738
rect 5710 39686 5724 39738
rect 5748 39686 5762 39738
rect 5762 39686 5774 39738
rect 5774 39686 5804 39738
rect 5828 39686 5838 39738
rect 5838 39686 5884 39738
rect 5588 39684 5644 39686
rect 5668 39684 5724 39686
rect 5748 39684 5804 39686
rect 5828 39684 5884 39686
rect 3882 29960 3938 30016
rect 2870 10240 2926 10296
rect 2778 8200 2834 8256
rect 2778 7520 2834 7576
rect 2870 6860 2926 6896
rect 2870 6840 2872 6860
rect 2872 6840 2924 6860
rect 2924 6840 2926 6860
rect 2778 4800 2834 4856
rect 5588 38650 5644 38652
rect 5668 38650 5724 38652
rect 5748 38650 5804 38652
rect 5828 38650 5884 38652
rect 5588 38598 5634 38650
rect 5634 38598 5644 38650
rect 5668 38598 5698 38650
rect 5698 38598 5710 38650
rect 5710 38598 5724 38650
rect 5748 38598 5762 38650
rect 5762 38598 5774 38650
rect 5774 38598 5804 38650
rect 5828 38598 5838 38650
rect 5838 38598 5884 38650
rect 5588 38596 5644 38598
rect 5668 38596 5724 38598
rect 5748 38596 5804 38598
rect 5828 38596 5884 38598
rect 5588 37562 5644 37564
rect 5668 37562 5724 37564
rect 5748 37562 5804 37564
rect 5828 37562 5884 37564
rect 5588 37510 5634 37562
rect 5634 37510 5644 37562
rect 5668 37510 5698 37562
rect 5698 37510 5710 37562
rect 5710 37510 5724 37562
rect 5748 37510 5762 37562
rect 5762 37510 5774 37562
rect 5774 37510 5804 37562
rect 5828 37510 5838 37562
rect 5838 37510 5884 37562
rect 5588 37508 5644 37510
rect 5668 37508 5724 37510
rect 5748 37508 5804 37510
rect 5828 37508 5884 37510
rect 5588 36474 5644 36476
rect 5668 36474 5724 36476
rect 5748 36474 5804 36476
rect 5828 36474 5884 36476
rect 5588 36422 5634 36474
rect 5634 36422 5644 36474
rect 5668 36422 5698 36474
rect 5698 36422 5710 36474
rect 5710 36422 5724 36474
rect 5748 36422 5762 36474
rect 5762 36422 5774 36474
rect 5774 36422 5804 36474
rect 5828 36422 5838 36474
rect 5838 36422 5884 36474
rect 5588 36420 5644 36422
rect 5668 36420 5724 36422
rect 5748 36420 5804 36422
rect 5828 36420 5884 36422
rect 6274 36352 6330 36408
rect 5588 35386 5644 35388
rect 5668 35386 5724 35388
rect 5748 35386 5804 35388
rect 5828 35386 5884 35388
rect 5588 35334 5634 35386
rect 5634 35334 5644 35386
rect 5668 35334 5698 35386
rect 5698 35334 5710 35386
rect 5710 35334 5724 35386
rect 5748 35334 5762 35386
rect 5762 35334 5774 35386
rect 5774 35334 5804 35386
rect 5828 35334 5838 35386
rect 5838 35334 5884 35386
rect 5588 35332 5644 35334
rect 5668 35332 5724 35334
rect 5748 35332 5804 35334
rect 5828 35332 5884 35334
rect 5998 35400 6054 35456
rect 5588 34298 5644 34300
rect 5668 34298 5724 34300
rect 5748 34298 5804 34300
rect 5828 34298 5884 34300
rect 5588 34246 5634 34298
rect 5634 34246 5644 34298
rect 5668 34246 5698 34298
rect 5698 34246 5710 34298
rect 5710 34246 5724 34298
rect 5748 34246 5762 34298
rect 5762 34246 5774 34298
rect 5774 34246 5804 34298
rect 5828 34246 5838 34298
rect 5838 34246 5884 34298
rect 5588 34244 5644 34246
rect 5668 34244 5724 34246
rect 5748 34244 5804 34246
rect 5828 34244 5884 34246
rect 5588 33210 5644 33212
rect 5668 33210 5724 33212
rect 5748 33210 5804 33212
rect 5828 33210 5884 33212
rect 5588 33158 5634 33210
rect 5634 33158 5644 33210
rect 5668 33158 5698 33210
rect 5698 33158 5710 33210
rect 5710 33158 5724 33210
rect 5748 33158 5762 33210
rect 5762 33158 5774 33210
rect 5774 33158 5804 33210
rect 5828 33158 5838 33210
rect 5838 33158 5884 33210
rect 5588 33156 5644 33158
rect 5668 33156 5724 33158
rect 5748 33156 5804 33158
rect 5828 33156 5884 33158
rect 5588 32122 5644 32124
rect 5668 32122 5724 32124
rect 5748 32122 5804 32124
rect 5828 32122 5884 32124
rect 5588 32070 5634 32122
rect 5634 32070 5644 32122
rect 5668 32070 5698 32122
rect 5698 32070 5710 32122
rect 5710 32070 5724 32122
rect 5748 32070 5762 32122
rect 5762 32070 5774 32122
rect 5774 32070 5804 32122
rect 5828 32070 5838 32122
rect 5838 32070 5884 32122
rect 5588 32068 5644 32070
rect 5668 32068 5724 32070
rect 5748 32068 5804 32070
rect 5828 32068 5884 32070
rect 5588 31034 5644 31036
rect 5668 31034 5724 31036
rect 5748 31034 5804 31036
rect 5828 31034 5884 31036
rect 5588 30982 5634 31034
rect 5634 30982 5644 31034
rect 5668 30982 5698 31034
rect 5698 30982 5710 31034
rect 5710 30982 5724 31034
rect 5748 30982 5762 31034
rect 5762 30982 5774 31034
rect 5774 30982 5804 31034
rect 5828 30982 5838 31034
rect 5838 30982 5884 31034
rect 5588 30980 5644 30982
rect 5668 30980 5724 30982
rect 5748 30980 5804 30982
rect 5828 30980 5884 30982
rect 5588 29946 5644 29948
rect 5668 29946 5724 29948
rect 5748 29946 5804 29948
rect 5828 29946 5884 29948
rect 5588 29894 5634 29946
rect 5634 29894 5644 29946
rect 5668 29894 5698 29946
rect 5698 29894 5710 29946
rect 5710 29894 5724 29946
rect 5748 29894 5762 29946
rect 5762 29894 5774 29946
rect 5774 29894 5804 29946
rect 5828 29894 5838 29946
rect 5838 29894 5884 29946
rect 5588 29892 5644 29894
rect 5668 29892 5724 29894
rect 5748 29892 5804 29894
rect 5828 29892 5884 29894
rect 5588 28858 5644 28860
rect 5668 28858 5724 28860
rect 5748 28858 5804 28860
rect 5828 28858 5884 28860
rect 5588 28806 5634 28858
rect 5634 28806 5644 28858
rect 5668 28806 5698 28858
rect 5698 28806 5710 28858
rect 5710 28806 5724 28858
rect 5748 28806 5762 28858
rect 5762 28806 5774 28858
rect 5774 28806 5804 28858
rect 5828 28806 5838 28858
rect 5838 28806 5884 28858
rect 5588 28804 5644 28806
rect 5668 28804 5724 28806
rect 5748 28804 5804 28806
rect 5828 28804 5884 28806
rect 5588 27770 5644 27772
rect 5668 27770 5724 27772
rect 5748 27770 5804 27772
rect 5828 27770 5884 27772
rect 5588 27718 5634 27770
rect 5634 27718 5644 27770
rect 5668 27718 5698 27770
rect 5698 27718 5710 27770
rect 5710 27718 5724 27770
rect 5748 27718 5762 27770
rect 5762 27718 5774 27770
rect 5774 27718 5804 27770
rect 5828 27718 5838 27770
rect 5838 27718 5884 27770
rect 5588 27716 5644 27718
rect 5668 27716 5724 27718
rect 5748 27716 5804 27718
rect 5828 27716 5884 27718
rect 5588 26682 5644 26684
rect 5668 26682 5724 26684
rect 5748 26682 5804 26684
rect 5828 26682 5884 26684
rect 5588 26630 5634 26682
rect 5634 26630 5644 26682
rect 5668 26630 5698 26682
rect 5698 26630 5710 26682
rect 5710 26630 5724 26682
rect 5748 26630 5762 26682
rect 5762 26630 5774 26682
rect 5774 26630 5804 26682
rect 5828 26630 5838 26682
rect 5838 26630 5884 26682
rect 5588 26628 5644 26630
rect 5668 26628 5724 26630
rect 5748 26628 5804 26630
rect 5828 26628 5884 26630
rect 5588 25594 5644 25596
rect 5668 25594 5724 25596
rect 5748 25594 5804 25596
rect 5828 25594 5884 25596
rect 5588 25542 5634 25594
rect 5634 25542 5644 25594
rect 5668 25542 5698 25594
rect 5698 25542 5710 25594
rect 5710 25542 5724 25594
rect 5748 25542 5762 25594
rect 5762 25542 5774 25594
rect 5774 25542 5804 25594
rect 5828 25542 5838 25594
rect 5838 25542 5884 25594
rect 5588 25540 5644 25542
rect 5668 25540 5724 25542
rect 5748 25540 5804 25542
rect 5828 25540 5884 25542
rect 5588 24506 5644 24508
rect 5668 24506 5724 24508
rect 5748 24506 5804 24508
rect 5828 24506 5884 24508
rect 5588 24454 5634 24506
rect 5634 24454 5644 24506
rect 5668 24454 5698 24506
rect 5698 24454 5710 24506
rect 5710 24454 5724 24506
rect 5748 24454 5762 24506
rect 5762 24454 5774 24506
rect 5774 24454 5804 24506
rect 5828 24454 5838 24506
rect 5838 24454 5884 24506
rect 5588 24452 5644 24454
rect 5668 24452 5724 24454
rect 5748 24452 5804 24454
rect 5828 24452 5884 24454
rect 5588 23418 5644 23420
rect 5668 23418 5724 23420
rect 5748 23418 5804 23420
rect 5828 23418 5884 23420
rect 5588 23366 5634 23418
rect 5634 23366 5644 23418
rect 5668 23366 5698 23418
rect 5698 23366 5710 23418
rect 5710 23366 5724 23418
rect 5748 23366 5762 23418
rect 5762 23366 5774 23418
rect 5774 23366 5804 23418
rect 5828 23366 5838 23418
rect 5838 23366 5884 23418
rect 5588 23364 5644 23366
rect 5668 23364 5724 23366
rect 5748 23364 5804 23366
rect 5828 23364 5884 23366
rect 5588 22330 5644 22332
rect 5668 22330 5724 22332
rect 5748 22330 5804 22332
rect 5828 22330 5884 22332
rect 5588 22278 5634 22330
rect 5634 22278 5644 22330
rect 5668 22278 5698 22330
rect 5698 22278 5710 22330
rect 5710 22278 5724 22330
rect 5748 22278 5762 22330
rect 5762 22278 5774 22330
rect 5774 22278 5804 22330
rect 5828 22278 5838 22330
rect 5838 22278 5884 22330
rect 5588 22276 5644 22278
rect 5668 22276 5724 22278
rect 5748 22276 5804 22278
rect 5828 22276 5884 22278
rect 5588 21242 5644 21244
rect 5668 21242 5724 21244
rect 5748 21242 5804 21244
rect 5828 21242 5884 21244
rect 5588 21190 5634 21242
rect 5634 21190 5644 21242
rect 5668 21190 5698 21242
rect 5698 21190 5710 21242
rect 5710 21190 5724 21242
rect 5748 21190 5762 21242
rect 5762 21190 5774 21242
rect 5774 21190 5804 21242
rect 5828 21190 5838 21242
rect 5838 21190 5884 21242
rect 5588 21188 5644 21190
rect 5668 21188 5724 21190
rect 5748 21188 5804 21190
rect 5828 21188 5884 21190
rect 5588 20154 5644 20156
rect 5668 20154 5724 20156
rect 5748 20154 5804 20156
rect 5828 20154 5884 20156
rect 5588 20102 5634 20154
rect 5634 20102 5644 20154
rect 5668 20102 5698 20154
rect 5698 20102 5710 20154
rect 5710 20102 5724 20154
rect 5748 20102 5762 20154
rect 5762 20102 5774 20154
rect 5774 20102 5804 20154
rect 5828 20102 5838 20154
rect 5838 20102 5884 20154
rect 5588 20100 5644 20102
rect 5668 20100 5724 20102
rect 5748 20100 5804 20102
rect 5828 20100 5884 20102
rect 5588 19066 5644 19068
rect 5668 19066 5724 19068
rect 5748 19066 5804 19068
rect 5828 19066 5884 19068
rect 5588 19014 5634 19066
rect 5634 19014 5644 19066
rect 5668 19014 5698 19066
rect 5698 19014 5710 19066
rect 5710 19014 5724 19066
rect 5748 19014 5762 19066
rect 5762 19014 5774 19066
rect 5774 19014 5804 19066
rect 5828 19014 5838 19066
rect 5838 19014 5884 19066
rect 5588 19012 5644 19014
rect 5668 19012 5724 19014
rect 5748 19012 5804 19014
rect 5828 19012 5884 19014
rect 5588 17978 5644 17980
rect 5668 17978 5724 17980
rect 5748 17978 5804 17980
rect 5828 17978 5884 17980
rect 5588 17926 5634 17978
rect 5634 17926 5644 17978
rect 5668 17926 5698 17978
rect 5698 17926 5710 17978
rect 5710 17926 5724 17978
rect 5748 17926 5762 17978
rect 5762 17926 5774 17978
rect 5774 17926 5804 17978
rect 5828 17926 5838 17978
rect 5838 17926 5884 17978
rect 5588 17924 5644 17926
rect 5668 17924 5724 17926
rect 5748 17924 5804 17926
rect 5828 17924 5884 17926
rect 7286 39752 7342 39808
rect 7378 38256 7434 38312
rect 7286 36624 7342 36680
rect 7102 34584 7158 34640
rect 7562 35692 7618 35728
rect 7562 35672 7564 35692
rect 7564 35672 7616 35692
rect 7616 35672 7618 35692
rect 7562 34584 7618 34640
rect 7562 34040 7618 34096
rect 8666 40432 8722 40488
rect 7838 39344 7894 39400
rect 7746 38428 7748 38448
rect 7748 38428 7800 38448
rect 7800 38428 7802 38448
rect 7746 38392 7802 38428
rect 8298 38936 8354 38992
rect 8022 38820 8078 38856
rect 8022 38800 8024 38820
rect 8024 38800 8076 38820
rect 8076 38800 8078 38820
rect 8206 37984 8262 38040
rect 8666 37712 8722 37768
rect 8022 37440 8078 37496
rect 7562 33224 7618 33280
rect 7562 17720 7618 17776
rect 5588 16890 5644 16892
rect 5668 16890 5724 16892
rect 5748 16890 5804 16892
rect 5828 16890 5884 16892
rect 5588 16838 5634 16890
rect 5634 16838 5644 16890
rect 5668 16838 5698 16890
rect 5698 16838 5710 16890
rect 5710 16838 5724 16890
rect 5748 16838 5762 16890
rect 5762 16838 5774 16890
rect 5774 16838 5804 16890
rect 5828 16838 5838 16890
rect 5838 16838 5884 16890
rect 5588 16836 5644 16838
rect 5668 16836 5724 16838
rect 5748 16836 5804 16838
rect 5828 16836 5884 16838
rect 8206 37168 8262 37224
rect 8206 35692 8262 35728
rect 8206 35672 8208 35692
rect 8208 35672 8260 35692
rect 8260 35672 8262 35692
rect 8114 33496 8170 33552
rect 8390 35128 8446 35184
rect 8390 34856 8446 34912
rect 8482 34176 8538 34232
rect 8482 33940 8484 33960
rect 8484 33940 8536 33960
rect 8536 33940 8538 33960
rect 8482 33904 8538 33940
rect 8114 31204 8170 31240
rect 8114 31184 8116 31204
rect 8116 31184 8168 31204
rect 8168 31184 8170 31204
rect 8206 30504 8262 30560
rect 8758 37304 8814 37360
rect 8850 36488 8906 36544
rect 8758 34312 8814 34368
rect 8942 36252 8944 36272
rect 8944 36252 8996 36272
rect 8996 36252 8998 36272
rect 8942 36216 8998 36252
rect 9494 38292 9496 38312
rect 9496 38292 9548 38312
rect 9548 38292 9550 38312
rect 9494 38256 9550 38292
rect 9678 38256 9734 38312
rect 9218 37848 9274 37904
rect 9494 37576 9550 37632
rect 9402 36216 9458 36272
rect 9310 36080 9366 36136
rect 9126 35944 9182 36000
rect 9034 35808 9090 35864
rect 9586 36896 9642 36952
rect 9586 36760 9642 36816
rect 10220 39194 10276 39196
rect 10300 39194 10356 39196
rect 10380 39194 10436 39196
rect 10460 39194 10516 39196
rect 10220 39142 10266 39194
rect 10266 39142 10276 39194
rect 10300 39142 10330 39194
rect 10330 39142 10342 39194
rect 10342 39142 10356 39194
rect 10380 39142 10394 39194
rect 10394 39142 10406 39194
rect 10406 39142 10436 39194
rect 10460 39142 10470 39194
rect 10470 39142 10516 39194
rect 10220 39140 10276 39142
rect 10300 39140 10356 39142
rect 10380 39140 10436 39142
rect 10460 39140 10516 39142
rect 10690 38664 10746 38720
rect 9954 37984 10010 38040
rect 10220 38106 10276 38108
rect 10300 38106 10356 38108
rect 10380 38106 10436 38108
rect 10460 38106 10516 38108
rect 10220 38054 10266 38106
rect 10266 38054 10276 38106
rect 10300 38054 10330 38106
rect 10330 38054 10342 38106
rect 10342 38054 10356 38106
rect 10380 38054 10394 38106
rect 10394 38054 10406 38106
rect 10406 38054 10436 38106
rect 10460 38054 10470 38106
rect 10470 38054 10516 38106
rect 10220 38052 10276 38054
rect 10300 38052 10356 38054
rect 10380 38052 10436 38054
rect 10460 38052 10516 38054
rect 10874 39072 10930 39128
rect 11426 40296 11482 40352
rect 10782 38120 10838 38176
rect 10874 37984 10930 38040
rect 9862 37032 9918 37088
rect 9770 36216 9826 36272
rect 10690 37032 10746 37088
rect 10220 37018 10276 37020
rect 10300 37018 10356 37020
rect 10380 37018 10436 37020
rect 10460 37018 10516 37020
rect 10220 36966 10266 37018
rect 10266 36966 10276 37018
rect 10300 36966 10330 37018
rect 10330 36966 10342 37018
rect 10342 36966 10356 37018
rect 10380 36966 10394 37018
rect 10394 36966 10406 37018
rect 10406 36966 10436 37018
rect 10460 36966 10470 37018
rect 10470 36966 10516 37018
rect 10220 36964 10276 36966
rect 10300 36964 10356 36966
rect 10380 36964 10436 36966
rect 10460 36964 10516 36966
rect 10046 36896 10102 36952
rect 10046 35980 10048 36000
rect 10048 35980 10100 36000
rect 10100 35980 10102 36000
rect 10046 35944 10102 35980
rect 10322 36216 10378 36272
rect 9218 35284 9274 35320
rect 9218 35264 9220 35284
rect 9220 35264 9272 35284
rect 9272 35264 9274 35284
rect 9862 35808 9918 35864
rect 10598 35944 10654 36000
rect 10220 35930 10276 35932
rect 10300 35930 10356 35932
rect 10380 35930 10436 35932
rect 10460 35930 10516 35932
rect 10220 35878 10266 35930
rect 10266 35878 10276 35930
rect 10300 35878 10330 35930
rect 10330 35878 10342 35930
rect 10342 35878 10356 35930
rect 10380 35878 10394 35930
rect 10394 35878 10406 35930
rect 10406 35878 10436 35930
rect 10460 35878 10470 35930
rect 10470 35878 10516 35930
rect 10220 35876 10276 35878
rect 10300 35876 10356 35878
rect 10380 35876 10436 35878
rect 10460 35876 10516 35878
rect 9494 35536 9550 35592
rect 9494 35264 9550 35320
rect 11058 35944 11114 36000
rect 10874 35808 10930 35864
rect 8942 33632 8998 33688
rect 8666 32292 8722 32328
rect 8666 32272 8668 32292
rect 8668 32272 8720 32292
rect 8720 32272 8722 32292
rect 8574 30776 8630 30832
rect 8574 29824 8630 29880
rect 8666 29688 8722 29744
rect 8390 29588 8392 29608
rect 8392 29588 8444 29608
rect 8444 29588 8446 29608
rect 8390 29552 8446 29588
rect 8942 31456 8998 31512
rect 9126 32172 9128 32192
rect 9128 32172 9180 32192
rect 9180 32172 9182 32192
rect 9126 32136 9182 32172
rect 9126 32000 9182 32056
rect 8298 28056 8354 28112
rect 9126 30640 9182 30696
rect 9586 35128 9642 35184
rect 9862 34992 9918 35048
rect 9954 34856 10010 34912
rect 10046 34720 10102 34776
rect 9310 34448 9366 34504
rect 10598 34856 10654 34912
rect 10874 34856 10930 34912
rect 10220 34842 10276 34844
rect 10300 34842 10356 34844
rect 10380 34842 10436 34844
rect 10460 34842 10516 34844
rect 10220 34790 10266 34842
rect 10266 34790 10276 34842
rect 10300 34790 10330 34842
rect 10330 34790 10342 34842
rect 10342 34790 10356 34842
rect 10380 34790 10394 34842
rect 10394 34790 10406 34842
rect 10406 34790 10436 34842
rect 10460 34790 10470 34842
rect 10470 34790 10516 34842
rect 10220 34788 10276 34790
rect 10300 34788 10356 34790
rect 10380 34788 10436 34790
rect 10460 34788 10516 34790
rect 12162 40160 12218 40216
rect 12162 39616 12218 39672
rect 12530 40160 12586 40216
rect 12530 39888 12586 39944
rect 12346 39616 12402 39672
rect 11978 37984 12034 38040
rect 12530 37984 12586 38040
rect 12070 37712 12126 37768
rect 12990 38548 13046 38584
rect 12990 38528 12992 38548
rect 12992 38528 13044 38548
rect 13044 38528 13046 38548
rect 12990 37984 13046 38040
rect 11518 37032 11574 37088
rect 12254 37032 12310 37088
rect 11610 35944 11666 36000
rect 12070 36624 12126 36680
rect 12438 37032 12494 37088
rect 12070 36488 12126 36544
rect 11886 35944 11942 36000
rect 11242 34584 11298 34640
rect 9678 33904 9734 33960
rect 10414 33940 10416 33960
rect 10416 33940 10468 33960
rect 10468 33940 10470 33960
rect 9770 33768 9826 33824
rect 9402 33088 9458 33144
rect 9770 32952 9826 33008
rect 10414 33904 10470 33940
rect 11058 34176 11114 34232
rect 10874 34040 10930 34096
rect 10598 33768 10654 33824
rect 10966 33768 11022 33824
rect 10220 33754 10276 33756
rect 10300 33754 10356 33756
rect 10380 33754 10436 33756
rect 10460 33754 10516 33756
rect 10220 33702 10266 33754
rect 10266 33702 10276 33754
rect 10300 33702 10330 33754
rect 10330 33702 10342 33754
rect 10342 33702 10356 33754
rect 10380 33702 10394 33754
rect 10394 33702 10406 33754
rect 10406 33702 10436 33754
rect 10460 33702 10470 33754
rect 10470 33702 10516 33754
rect 10220 33700 10276 33702
rect 10300 33700 10356 33702
rect 10380 33700 10436 33702
rect 10460 33700 10516 33702
rect 10046 33632 10102 33688
rect 10598 33632 10654 33688
rect 10046 33360 10102 33416
rect 10414 33496 10470 33552
rect 9678 32816 9734 32872
rect 9770 32408 9826 32464
rect 9402 31592 9458 31648
rect 10322 33224 10378 33280
rect 11426 33496 11482 33552
rect 11058 33224 11114 33280
rect 10874 33088 10930 33144
rect 10220 32666 10276 32668
rect 10300 32666 10356 32668
rect 10380 32666 10436 32668
rect 10460 32666 10516 32668
rect 10220 32614 10266 32666
rect 10266 32614 10276 32666
rect 10300 32614 10330 32666
rect 10330 32614 10342 32666
rect 10342 32614 10356 32666
rect 10380 32614 10394 32666
rect 10394 32614 10406 32666
rect 10406 32614 10436 32666
rect 10460 32614 10470 32666
rect 10470 32614 10516 32666
rect 10220 32612 10276 32614
rect 10300 32612 10356 32614
rect 10380 32612 10436 32614
rect 10460 32612 10516 32614
rect 11702 34076 11704 34096
rect 11704 34076 11756 34096
rect 11756 34076 11758 34096
rect 11702 34040 11758 34076
rect 11058 32816 11114 32872
rect 9954 31864 10010 31920
rect 11242 32680 11298 32736
rect 12254 36080 12310 36136
rect 12714 36352 12770 36408
rect 12162 35808 12218 35864
rect 12162 35264 12218 35320
rect 11978 34448 12034 34504
rect 12254 34448 12310 34504
rect 12254 33904 12310 33960
rect 11794 32680 11850 32736
rect 9862 31456 9918 31512
rect 9954 31320 10010 31376
rect 9402 30912 9458 30968
rect 10046 30504 10102 30560
rect 9862 30368 9918 30424
rect 9494 30232 9550 30288
rect 9310 29960 9366 30016
rect 9402 29144 9458 29200
rect 9126 29008 9182 29064
rect 9126 28908 9128 28928
rect 9128 28908 9180 28928
rect 9180 28908 9182 28928
rect 9126 28872 9182 28908
rect 9034 28464 9090 28520
rect 8942 27512 8998 27568
rect 9770 29280 9826 29336
rect 9586 27648 9642 27704
rect 9494 27412 9496 27432
rect 9496 27412 9548 27432
rect 9548 27412 9550 27432
rect 9494 27376 9550 27412
rect 9678 26852 9734 26888
rect 9678 26832 9680 26852
rect 9680 26832 9732 26852
rect 9732 26832 9734 26852
rect 9954 30096 10010 30152
rect 10220 31578 10276 31580
rect 10300 31578 10356 31580
rect 10380 31578 10436 31580
rect 10460 31578 10516 31580
rect 10220 31526 10266 31578
rect 10266 31526 10276 31578
rect 10300 31526 10330 31578
rect 10330 31526 10342 31578
rect 10342 31526 10356 31578
rect 10380 31526 10394 31578
rect 10394 31526 10406 31578
rect 10406 31526 10436 31578
rect 10460 31526 10470 31578
rect 10470 31526 10516 31578
rect 10220 31524 10276 31526
rect 10300 31524 10356 31526
rect 10380 31524 10436 31526
rect 10460 31524 10516 31526
rect 10782 31748 10838 31784
rect 10782 31728 10784 31748
rect 10784 31728 10836 31748
rect 10836 31728 10838 31748
rect 10874 31048 10930 31104
rect 10782 30640 10838 30696
rect 10220 30490 10276 30492
rect 10300 30490 10356 30492
rect 10380 30490 10436 30492
rect 10460 30490 10516 30492
rect 10220 30438 10266 30490
rect 10266 30438 10276 30490
rect 10300 30438 10330 30490
rect 10330 30438 10342 30490
rect 10342 30438 10356 30490
rect 10380 30438 10394 30490
rect 10394 30438 10406 30490
rect 10406 30438 10436 30490
rect 10460 30438 10470 30490
rect 10470 30438 10516 30490
rect 10220 30436 10276 30438
rect 10300 30436 10356 30438
rect 10380 30436 10436 30438
rect 10460 30436 10516 30438
rect 10220 29402 10276 29404
rect 10300 29402 10356 29404
rect 10380 29402 10436 29404
rect 10460 29402 10516 29404
rect 10220 29350 10266 29402
rect 10266 29350 10276 29402
rect 10300 29350 10330 29402
rect 10330 29350 10342 29402
rect 10342 29350 10356 29402
rect 10380 29350 10394 29402
rect 10394 29350 10406 29402
rect 10406 29350 10436 29402
rect 10460 29350 10470 29402
rect 10470 29350 10516 29402
rect 10220 29348 10276 29350
rect 10300 29348 10356 29350
rect 10380 29348 10436 29350
rect 10460 29348 10516 29350
rect 10598 29280 10654 29336
rect 10874 29416 10930 29472
rect 9954 28736 10010 28792
rect 10046 28600 10102 28656
rect 10046 27920 10102 27976
rect 10506 28736 10562 28792
rect 10220 28314 10276 28316
rect 10300 28314 10356 28316
rect 10380 28314 10436 28316
rect 10460 28314 10516 28316
rect 10220 28262 10266 28314
rect 10266 28262 10276 28314
rect 10300 28262 10330 28314
rect 10330 28262 10342 28314
rect 10342 28262 10356 28314
rect 10380 28262 10394 28314
rect 10394 28262 10406 28314
rect 10406 28262 10436 28314
rect 10460 28262 10470 28314
rect 10470 28262 10516 28314
rect 10220 28260 10276 28262
rect 10300 28260 10356 28262
rect 10380 28260 10436 28262
rect 10460 28260 10516 28262
rect 10598 27920 10654 27976
rect 10138 27784 10194 27840
rect 9034 26288 9090 26344
rect 7838 24792 7894 24848
rect 7746 16496 7802 16552
rect 9586 16088 9642 16144
rect 5588 15802 5644 15804
rect 5668 15802 5724 15804
rect 5748 15802 5804 15804
rect 5828 15802 5884 15804
rect 5588 15750 5634 15802
rect 5634 15750 5644 15802
rect 5668 15750 5698 15802
rect 5698 15750 5710 15802
rect 5710 15750 5724 15802
rect 5748 15750 5762 15802
rect 5762 15750 5774 15802
rect 5774 15750 5804 15802
rect 5828 15750 5838 15802
rect 5838 15750 5884 15802
rect 5588 15748 5644 15750
rect 5668 15748 5724 15750
rect 5748 15748 5804 15750
rect 5828 15748 5884 15750
rect 5588 14714 5644 14716
rect 5668 14714 5724 14716
rect 5748 14714 5804 14716
rect 5828 14714 5884 14716
rect 5588 14662 5634 14714
rect 5634 14662 5644 14714
rect 5668 14662 5698 14714
rect 5698 14662 5710 14714
rect 5710 14662 5724 14714
rect 5748 14662 5762 14714
rect 5762 14662 5774 14714
rect 5774 14662 5804 14714
rect 5828 14662 5838 14714
rect 5838 14662 5884 14714
rect 5588 14660 5644 14662
rect 5668 14660 5724 14662
rect 5748 14660 5804 14662
rect 5828 14660 5884 14662
rect 5588 13626 5644 13628
rect 5668 13626 5724 13628
rect 5748 13626 5804 13628
rect 5828 13626 5884 13628
rect 5588 13574 5634 13626
rect 5634 13574 5644 13626
rect 5668 13574 5698 13626
rect 5698 13574 5710 13626
rect 5710 13574 5724 13626
rect 5748 13574 5762 13626
rect 5762 13574 5774 13626
rect 5774 13574 5804 13626
rect 5828 13574 5838 13626
rect 5838 13574 5884 13626
rect 5588 13572 5644 13574
rect 5668 13572 5724 13574
rect 5748 13572 5804 13574
rect 5828 13572 5884 13574
rect 5588 12538 5644 12540
rect 5668 12538 5724 12540
rect 5748 12538 5804 12540
rect 5828 12538 5884 12540
rect 5588 12486 5634 12538
rect 5634 12486 5644 12538
rect 5668 12486 5698 12538
rect 5698 12486 5710 12538
rect 5710 12486 5724 12538
rect 5748 12486 5762 12538
rect 5762 12486 5774 12538
rect 5774 12486 5804 12538
rect 5828 12486 5838 12538
rect 5838 12486 5884 12538
rect 5588 12484 5644 12486
rect 5668 12484 5724 12486
rect 5748 12484 5804 12486
rect 5828 12484 5884 12486
rect 5588 11450 5644 11452
rect 5668 11450 5724 11452
rect 5748 11450 5804 11452
rect 5828 11450 5884 11452
rect 5588 11398 5634 11450
rect 5634 11398 5644 11450
rect 5668 11398 5698 11450
rect 5698 11398 5710 11450
rect 5710 11398 5724 11450
rect 5748 11398 5762 11450
rect 5762 11398 5774 11450
rect 5774 11398 5804 11450
rect 5828 11398 5838 11450
rect 5838 11398 5884 11450
rect 5588 11396 5644 11398
rect 5668 11396 5724 11398
rect 5748 11396 5804 11398
rect 5828 11396 5884 11398
rect 5588 10362 5644 10364
rect 5668 10362 5724 10364
rect 5748 10362 5804 10364
rect 5828 10362 5884 10364
rect 5588 10310 5634 10362
rect 5634 10310 5644 10362
rect 5668 10310 5698 10362
rect 5698 10310 5710 10362
rect 5710 10310 5724 10362
rect 5748 10310 5762 10362
rect 5762 10310 5774 10362
rect 5774 10310 5804 10362
rect 5828 10310 5838 10362
rect 5838 10310 5884 10362
rect 5588 10308 5644 10310
rect 5668 10308 5724 10310
rect 5748 10308 5804 10310
rect 5828 10308 5884 10310
rect 5588 9274 5644 9276
rect 5668 9274 5724 9276
rect 5748 9274 5804 9276
rect 5828 9274 5884 9276
rect 5588 9222 5634 9274
rect 5634 9222 5644 9274
rect 5668 9222 5698 9274
rect 5698 9222 5710 9274
rect 5710 9222 5724 9274
rect 5748 9222 5762 9274
rect 5762 9222 5774 9274
rect 5774 9222 5804 9274
rect 5828 9222 5838 9274
rect 5838 9222 5884 9274
rect 5588 9220 5644 9222
rect 5668 9220 5724 9222
rect 5748 9220 5804 9222
rect 5828 9220 5884 9222
rect 5588 8186 5644 8188
rect 5668 8186 5724 8188
rect 5748 8186 5804 8188
rect 5828 8186 5884 8188
rect 5588 8134 5634 8186
rect 5634 8134 5644 8186
rect 5668 8134 5698 8186
rect 5698 8134 5710 8186
rect 5710 8134 5724 8186
rect 5748 8134 5762 8186
rect 5762 8134 5774 8186
rect 5774 8134 5804 8186
rect 5828 8134 5838 8186
rect 5838 8134 5884 8186
rect 5588 8132 5644 8134
rect 5668 8132 5724 8134
rect 5748 8132 5804 8134
rect 5828 8132 5884 8134
rect 5588 7098 5644 7100
rect 5668 7098 5724 7100
rect 5748 7098 5804 7100
rect 5828 7098 5884 7100
rect 5588 7046 5634 7098
rect 5634 7046 5644 7098
rect 5668 7046 5698 7098
rect 5698 7046 5710 7098
rect 5710 7046 5724 7098
rect 5748 7046 5762 7098
rect 5762 7046 5774 7098
rect 5774 7046 5804 7098
rect 5828 7046 5838 7098
rect 5838 7046 5884 7098
rect 5588 7044 5644 7046
rect 5668 7044 5724 7046
rect 5748 7044 5804 7046
rect 5828 7044 5884 7046
rect 4066 4120 4122 4176
rect 2962 3440 3018 3496
rect 2778 2760 2834 2816
rect 3238 2080 3294 2136
rect 3054 1400 3110 1456
rect 5588 6010 5644 6012
rect 5668 6010 5724 6012
rect 5748 6010 5804 6012
rect 5828 6010 5884 6012
rect 5588 5958 5634 6010
rect 5634 5958 5644 6010
rect 5668 5958 5698 6010
rect 5698 5958 5710 6010
rect 5710 5958 5724 6010
rect 5748 5958 5762 6010
rect 5762 5958 5774 6010
rect 5774 5958 5804 6010
rect 5828 5958 5838 6010
rect 5838 5958 5884 6010
rect 5588 5956 5644 5958
rect 5668 5956 5724 5958
rect 5748 5956 5804 5958
rect 5828 5956 5884 5958
rect 5588 4922 5644 4924
rect 5668 4922 5724 4924
rect 5748 4922 5804 4924
rect 5828 4922 5884 4924
rect 5588 4870 5634 4922
rect 5634 4870 5644 4922
rect 5668 4870 5698 4922
rect 5698 4870 5710 4922
rect 5710 4870 5724 4922
rect 5748 4870 5762 4922
rect 5762 4870 5774 4922
rect 5774 4870 5804 4922
rect 5828 4870 5838 4922
rect 5838 4870 5884 4922
rect 5588 4868 5644 4870
rect 5668 4868 5724 4870
rect 5748 4868 5804 4870
rect 5828 4868 5884 4870
rect 5588 3834 5644 3836
rect 5668 3834 5724 3836
rect 5748 3834 5804 3836
rect 5828 3834 5884 3836
rect 5588 3782 5634 3834
rect 5634 3782 5644 3834
rect 5668 3782 5698 3834
rect 5698 3782 5710 3834
rect 5710 3782 5724 3834
rect 5748 3782 5762 3834
rect 5762 3782 5774 3834
rect 5774 3782 5804 3834
rect 5828 3782 5838 3834
rect 5838 3782 5884 3834
rect 5588 3780 5644 3782
rect 5668 3780 5724 3782
rect 5748 3780 5804 3782
rect 5828 3780 5884 3782
rect 5588 2746 5644 2748
rect 5668 2746 5724 2748
rect 5748 2746 5804 2748
rect 5828 2746 5884 2748
rect 5588 2694 5634 2746
rect 5634 2694 5644 2746
rect 5668 2694 5698 2746
rect 5698 2694 5710 2746
rect 5710 2694 5724 2746
rect 5748 2694 5762 2746
rect 5762 2694 5774 2746
rect 5774 2694 5804 2746
rect 5828 2694 5838 2746
rect 5838 2694 5884 2746
rect 5588 2692 5644 2694
rect 5668 2692 5724 2694
rect 5748 2692 5804 2694
rect 5828 2692 5884 2694
rect 10220 27226 10276 27228
rect 10300 27226 10356 27228
rect 10380 27226 10436 27228
rect 10460 27226 10516 27228
rect 10220 27174 10266 27226
rect 10266 27174 10276 27226
rect 10300 27174 10330 27226
rect 10330 27174 10342 27226
rect 10342 27174 10356 27226
rect 10380 27174 10394 27226
rect 10394 27174 10406 27226
rect 10406 27174 10436 27226
rect 10460 27174 10470 27226
rect 10470 27174 10516 27226
rect 10220 27172 10276 27174
rect 10300 27172 10356 27174
rect 10380 27172 10436 27174
rect 10460 27172 10516 27174
rect 10230 26560 10286 26616
rect 10220 26138 10276 26140
rect 10300 26138 10356 26140
rect 10380 26138 10436 26140
rect 10460 26138 10516 26140
rect 10220 26086 10266 26138
rect 10266 26086 10276 26138
rect 10300 26086 10330 26138
rect 10330 26086 10342 26138
rect 10342 26086 10356 26138
rect 10380 26086 10394 26138
rect 10394 26086 10406 26138
rect 10406 26086 10436 26138
rect 10460 26086 10470 26138
rect 10470 26086 10516 26138
rect 10220 26084 10276 26086
rect 10300 26084 10356 26086
rect 10380 26084 10436 26086
rect 10460 26084 10516 26086
rect 10782 28192 10838 28248
rect 10874 27920 10930 27976
rect 10782 26988 10838 27024
rect 10782 26968 10784 26988
rect 10784 26968 10836 26988
rect 10836 26968 10838 26988
rect 10690 26016 10746 26072
rect 10782 25608 10838 25664
rect 10598 25336 10654 25392
rect 10782 25236 10784 25256
rect 10784 25236 10836 25256
rect 10836 25236 10838 25256
rect 10220 25050 10276 25052
rect 10300 25050 10356 25052
rect 10380 25050 10436 25052
rect 10460 25050 10516 25052
rect 10220 24998 10266 25050
rect 10266 24998 10276 25050
rect 10300 24998 10330 25050
rect 10330 24998 10342 25050
rect 10342 24998 10356 25050
rect 10380 24998 10394 25050
rect 10394 24998 10406 25050
rect 10406 24998 10436 25050
rect 10460 24998 10470 25050
rect 10470 24998 10516 25050
rect 10220 24996 10276 24998
rect 10300 24996 10356 24998
rect 10380 24996 10436 24998
rect 10460 24996 10516 24998
rect 10782 25200 10838 25236
rect 12254 32680 12310 32736
rect 11426 31728 11482 31784
rect 11426 30912 11482 30968
rect 11702 31048 11758 31104
rect 11702 30368 11758 30424
rect 11058 28736 11114 28792
rect 11518 29688 11574 29744
rect 11978 31728 12034 31784
rect 12898 37032 12954 37088
rect 13082 37068 13084 37088
rect 13084 37068 13136 37088
rect 13136 37068 13138 37088
rect 13082 37032 13138 37068
rect 12990 36488 13046 36544
rect 12898 35944 12954 36000
rect 12806 35436 12808 35456
rect 12808 35436 12860 35456
rect 12860 35436 12862 35456
rect 12806 35400 12862 35436
rect 13726 37440 13782 37496
rect 13542 37032 13598 37088
rect 13542 36488 13598 36544
rect 13082 35536 13138 35592
rect 13266 35556 13322 35592
rect 13266 35536 13268 35556
rect 13268 35536 13320 35556
rect 13320 35536 13322 35556
rect 13266 35400 13322 35456
rect 13266 34992 13322 35048
rect 15382 40432 15438 40488
rect 15290 40024 15346 40080
rect 14646 39752 14702 39808
rect 14554 39616 14610 39672
rect 14370 39072 14426 39128
rect 15290 39752 15346 39808
rect 14852 39738 14908 39740
rect 14932 39738 14988 39740
rect 15012 39738 15068 39740
rect 15092 39738 15148 39740
rect 14852 39686 14898 39738
rect 14898 39686 14908 39738
rect 14932 39686 14962 39738
rect 14962 39686 14974 39738
rect 14974 39686 14988 39738
rect 15012 39686 15026 39738
rect 15026 39686 15038 39738
rect 15038 39686 15068 39738
rect 15092 39686 15102 39738
rect 15102 39686 15148 39738
rect 14852 39684 14908 39686
rect 14932 39684 14988 39686
rect 15012 39684 15068 39686
rect 15092 39684 15148 39686
rect 14646 39072 14702 39128
rect 14646 38664 14702 38720
rect 15290 38664 15346 38720
rect 14852 38650 14908 38652
rect 14932 38650 14988 38652
rect 15012 38650 15068 38652
rect 15092 38650 15148 38652
rect 14852 38598 14898 38650
rect 14898 38598 14908 38650
rect 14932 38598 14962 38650
rect 14962 38598 14974 38650
rect 14974 38598 14988 38650
rect 15012 38598 15026 38650
rect 15026 38598 15038 38650
rect 15038 38598 15068 38650
rect 15092 38598 15102 38650
rect 15102 38598 15148 38650
rect 14852 38596 14908 38598
rect 14932 38596 14988 38598
rect 15012 38596 15068 38598
rect 15092 38596 15148 38598
rect 14186 38528 14242 38584
rect 15290 38528 15346 38584
rect 14002 36252 14004 36272
rect 14004 36252 14056 36272
rect 14056 36252 14058 36272
rect 14002 36216 14058 36252
rect 15198 37712 15254 37768
rect 15382 37712 15438 37768
rect 14852 37562 14908 37564
rect 14932 37562 14988 37564
rect 15012 37562 15068 37564
rect 15092 37562 15148 37564
rect 14852 37510 14898 37562
rect 14898 37510 14908 37562
rect 14932 37510 14962 37562
rect 14962 37510 14974 37562
rect 14974 37510 14988 37562
rect 15012 37510 15026 37562
rect 15026 37510 15038 37562
rect 15038 37510 15068 37562
rect 15092 37510 15102 37562
rect 15102 37510 15148 37562
rect 14852 37508 14908 37510
rect 14932 37508 14988 37510
rect 15012 37508 15068 37510
rect 15092 37508 15148 37510
rect 15474 37440 15530 37496
rect 14370 36624 14426 36680
rect 14462 36488 14518 36544
rect 14852 36474 14908 36476
rect 14932 36474 14988 36476
rect 15012 36474 15068 36476
rect 15092 36474 15148 36476
rect 14852 36422 14898 36474
rect 14898 36422 14908 36474
rect 14932 36422 14962 36474
rect 14962 36422 14974 36474
rect 14974 36422 14988 36474
rect 15012 36422 15026 36474
rect 15026 36422 15038 36474
rect 15038 36422 15068 36474
rect 15092 36422 15102 36474
rect 15102 36422 15148 36474
rect 14852 36420 14908 36422
rect 14932 36420 14988 36422
rect 15012 36420 15068 36422
rect 15092 36420 15148 36422
rect 14646 36352 14702 36408
rect 15382 36372 15438 36408
rect 15382 36352 15384 36372
rect 15384 36352 15436 36372
rect 15436 36352 15438 36372
rect 13726 34992 13782 35048
rect 13910 35400 13966 35456
rect 13910 35028 13912 35048
rect 13912 35028 13964 35048
rect 13964 35028 13966 35048
rect 13910 34992 13966 35028
rect 12990 33632 13046 33688
rect 12990 33224 13046 33280
rect 13266 33224 13322 33280
rect 12714 32952 12770 33008
rect 14002 34312 14058 34368
rect 13910 34176 13966 34232
rect 13818 33496 13874 33552
rect 14094 34176 14150 34232
rect 14554 35536 14610 35592
rect 14738 35536 14794 35592
rect 14646 35264 14702 35320
rect 14852 35386 14908 35388
rect 14932 35386 14988 35388
rect 15012 35386 15068 35388
rect 15092 35386 15148 35388
rect 14852 35334 14898 35386
rect 14898 35334 14908 35386
rect 14932 35334 14962 35386
rect 14962 35334 14974 35386
rect 14974 35334 14988 35386
rect 15012 35334 15026 35386
rect 15026 35334 15038 35386
rect 15038 35334 15068 35386
rect 15092 35334 15102 35386
rect 15102 35334 15148 35386
rect 14852 35332 14908 35334
rect 14932 35332 14988 35334
rect 15012 35332 15068 35334
rect 15092 35332 15148 35334
rect 15290 35436 15292 35456
rect 15292 35436 15344 35456
rect 15344 35436 15346 35456
rect 15290 35400 15346 35436
rect 15290 35264 15346 35320
rect 19062 40296 19118 40352
rect 17038 39616 17094 39672
rect 17038 39344 17094 39400
rect 17314 39244 17316 39264
rect 17316 39244 17368 39264
rect 17368 39244 17370 39264
rect 17314 39208 17370 39244
rect 16118 37304 16174 37360
rect 15934 36216 15990 36272
rect 16210 36660 16212 36680
rect 16212 36660 16264 36680
rect 16264 36660 16266 36680
rect 16210 36624 16266 36660
rect 16486 35400 16542 35456
rect 15106 34584 15162 34640
rect 14852 34298 14908 34300
rect 14932 34298 14988 34300
rect 15012 34298 15068 34300
rect 15092 34298 15148 34300
rect 14852 34246 14898 34298
rect 14898 34246 14908 34298
rect 14932 34246 14962 34298
rect 14962 34246 14974 34298
rect 14974 34246 14988 34298
rect 15012 34246 15026 34298
rect 15026 34246 15038 34298
rect 15038 34246 15068 34298
rect 15092 34246 15102 34298
rect 15102 34246 15148 34298
rect 14852 34244 14908 34246
rect 14932 34244 14988 34246
rect 15012 34244 15068 34246
rect 15092 34244 15148 34246
rect 14646 34176 14702 34232
rect 15382 34312 15438 34368
rect 15198 34040 15254 34096
rect 14554 33904 14610 33960
rect 13910 33360 13966 33416
rect 12530 32136 12586 32192
rect 13542 32836 13598 32872
rect 13542 32816 13544 32836
rect 13544 32816 13596 32836
rect 13596 32816 13598 32836
rect 13726 32816 13782 32872
rect 13358 32564 13414 32600
rect 13358 32544 13360 32564
rect 13360 32544 13412 32564
rect 13412 32544 13414 32564
rect 13450 31864 13506 31920
rect 11886 31048 11942 31104
rect 11886 30504 11942 30560
rect 12714 30932 12770 30968
rect 12714 30912 12716 30932
rect 12716 30912 12768 30932
rect 12768 30912 12770 30932
rect 12898 30912 12954 30968
rect 12346 30540 12348 30560
rect 12348 30540 12400 30560
rect 12400 30540 12402 30560
rect 12346 30504 12402 30540
rect 12070 30096 12126 30152
rect 12438 30096 12494 30152
rect 12714 30640 12770 30696
rect 12714 30116 12770 30152
rect 12714 30096 12716 30116
rect 12716 30096 12768 30116
rect 12768 30096 12770 30116
rect 14002 32172 14004 32192
rect 14004 32172 14056 32192
rect 14056 32172 14058 32192
rect 14002 32136 14058 32172
rect 15106 33396 15108 33416
rect 15108 33396 15160 33416
rect 15160 33396 15162 33416
rect 15106 33360 15162 33396
rect 14646 33224 14702 33280
rect 14462 33088 14518 33144
rect 14852 33210 14908 33212
rect 14932 33210 14988 33212
rect 15012 33210 15068 33212
rect 15092 33210 15148 33212
rect 14852 33158 14898 33210
rect 14898 33158 14908 33210
rect 14932 33158 14962 33210
rect 14962 33158 14974 33210
rect 14974 33158 14988 33210
rect 15012 33158 15026 33210
rect 15026 33158 15038 33210
rect 15038 33158 15068 33210
rect 15092 33158 15102 33210
rect 15102 33158 15148 33210
rect 14852 33156 14908 33158
rect 14932 33156 14988 33158
rect 15012 33156 15068 33158
rect 15092 33156 15148 33158
rect 14278 32136 14334 32192
rect 13818 31864 13874 31920
rect 14278 31864 14334 31920
rect 13818 31592 13874 31648
rect 13726 31356 13728 31376
rect 13728 31356 13780 31376
rect 13780 31356 13782 31376
rect 13726 31320 13782 31356
rect 14002 31592 14058 31648
rect 13082 30640 13138 30696
rect 13174 30368 13230 30424
rect 13358 30368 13414 30424
rect 11978 29552 12034 29608
rect 11794 29416 11850 29472
rect 12254 29572 12310 29608
rect 12622 29688 12678 29744
rect 12254 29552 12256 29572
rect 12256 29552 12308 29572
rect 12308 29552 12310 29572
rect 12438 29416 12494 29472
rect 11610 29044 11612 29064
rect 11612 29044 11664 29064
rect 11664 29044 11666 29064
rect 11610 29008 11666 29044
rect 11978 29008 12034 29064
rect 11058 28464 11114 28520
rect 11334 28056 11390 28112
rect 10966 27240 11022 27296
rect 10220 23962 10276 23964
rect 10300 23962 10356 23964
rect 10380 23962 10436 23964
rect 10460 23962 10516 23964
rect 10220 23910 10266 23962
rect 10266 23910 10276 23962
rect 10300 23910 10330 23962
rect 10330 23910 10342 23962
rect 10342 23910 10356 23962
rect 10380 23910 10394 23962
rect 10394 23910 10406 23962
rect 10406 23910 10436 23962
rect 10460 23910 10470 23962
rect 10470 23910 10516 23962
rect 10220 23908 10276 23910
rect 10300 23908 10356 23910
rect 10380 23908 10436 23910
rect 10460 23908 10516 23910
rect 10322 23296 10378 23352
rect 10230 23160 10286 23216
rect 10220 22874 10276 22876
rect 10300 22874 10356 22876
rect 10380 22874 10436 22876
rect 10460 22874 10516 22876
rect 10220 22822 10266 22874
rect 10266 22822 10276 22874
rect 10300 22822 10330 22874
rect 10330 22822 10342 22874
rect 10342 22822 10356 22874
rect 10380 22822 10394 22874
rect 10394 22822 10406 22874
rect 10406 22822 10436 22874
rect 10460 22822 10470 22874
rect 10470 22822 10516 22874
rect 10220 22820 10276 22822
rect 10300 22820 10356 22822
rect 10380 22820 10436 22822
rect 10460 22820 10516 22822
rect 10220 21786 10276 21788
rect 10300 21786 10356 21788
rect 10380 21786 10436 21788
rect 10460 21786 10516 21788
rect 10220 21734 10266 21786
rect 10266 21734 10276 21786
rect 10300 21734 10330 21786
rect 10330 21734 10342 21786
rect 10342 21734 10356 21786
rect 10380 21734 10394 21786
rect 10394 21734 10406 21786
rect 10406 21734 10436 21786
rect 10460 21734 10470 21786
rect 10470 21734 10516 21786
rect 10220 21732 10276 21734
rect 10300 21732 10356 21734
rect 10380 21732 10436 21734
rect 10460 21732 10516 21734
rect 10220 20698 10276 20700
rect 10300 20698 10356 20700
rect 10380 20698 10436 20700
rect 10460 20698 10516 20700
rect 10220 20646 10266 20698
rect 10266 20646 10276 20698
rect 10300 20646 10330 20698
rect 10330 20646 10342 20698
rect 10342 20646 10356 20698
rect 10380 20646 10394 20698
rect 10394 20646 10406 20698
rect 10406 20646 10436 20698
rect 10460 20646 10470 20698
rect 10470 20646 10516 20698
rect 10220 20644 10276 20646
rect 10300 20644 10356 20646
rect 10380 20644 10436 20646
rect 10460 20644 10516 20646
rect 10220 19610 10276 19612
rect 10300 19610 10356 19612
rect 10380 19610 10436 19612
rect 10460 19610 10516 19612
rect 10220 19558 10266 19610
rect 10266 19558 10276 19610
rect 10300 19558 10330 19610
rect 10330 19558 10342 19610
rect 10342 19558 10356 19610
rect 10380 19558 10394 19610
rect 10394 19558 10406 19610
rect 10406 19558 10436 19610
rect 10460 19558 10470 19610
rect 10470 19558 10516 19610
rect 10220 19556 10276 19558
rect 10300 19556 10356 19558
rect 10380 19556 10436 19558
rect 10460 19556 10516 19558
rect 10220 18522 10276 18524
rect 10300 18522 10356 18524
rect 10380 18522 10436 18524
rect 10460 18522 10516 18524
rect 10220 18470 10266 18522
rect 10266 18470 10276 18522
rect 10300 18470 10330 18522
rect 10330 18470 10342 18522
rect 10342 18470 10356 18522
rect 10380 18470 10394 18522
rect 10394 18470 10406 18522
rect 10406 18470 10436 18522
rect 10460 18470 10470 18522
rect 10470 18470 10516 18522
rect 10220 18468 10276 18470
rect 10300 18468 10356 18470
rect 10380 18468 10436 18470
rect 10460 18468 10516 18470
rect 11334 26424 11390 26480
rect 11610 27920 11666 27976
rect 11794 28056 11850 28112
rect 12622 29144 12678 29200
rect 12438 28872 12494 28928
rect 12438 28636 12440 28656
rect 12440 28636 12492 28656
rect 12492 28636 12494 28656
rect 12438 28600 12494 28636
rect 11886 27940 11942 27976
rect 11886 27920 11888 27940
rect 11888 27920 11940 27940
rect 11940 27920 11942 27940
rect 11702 27104 11758 27160
rect 11794 26696 11850 26752
rect 12438 28056 12494 28112
rect 12622 28600 12678 28656
rect 12622 28464 12678 28520
rect 12622 28056 12678 28112
rect 12530 27920 12586 27976
rect 12990 29824 13046 29880
rect 13266 29824 13322 29880
rect 12990 29552 13046 29608
rect 12898 28500 12900 28520
rect 12900 28500 12952 28520
rect 12952 28500 12954 28520
rect 12898 28464 12954 28500
rect 13082 29008 13138 29064
rect 13450 29824 13506 29880
rect 13450 29552 13506 29608
rect 14186 30504 14242 30560
rect 12254 27240 12310 27296
rect 12438 27276 12440 27296
rect 12440 27276 12492 27296
rect 12492 27276 12494 27296
rect 12438 27240 12494 27276
rect 11058 25880 11114 25936
rect 11150 25744 11206 25800
rect 11058 25492 11114 25528
rect 11058 25472 11060 25492
rect 11060 25472 11112 25492
rect 11112 25472 11114 25492
rect 11058 24928 11114 24984
rect 12622 26424 12678 26480
rect 12070 26152 12126 26208
rect 12070 24656 12126 24712
rect 11518 24520 11574 24576
rect 10690 23976 10746 24032
rect 10782 23840 10838 23896
rect 11426 23704 11482 23760
rect 13266 27376 13322 27432
rect 12990 27240 13046 27296
rect 12806 25880 12862 25936
rect 12530 25472 12586 25528
rect 14094 29960 14150 30016
rect 13450 27240 13506 27296
rect 13634 27240 13690 27296
rect 12438 23724 12494 23760
rect 12438 23704 12440 23724
rect 12440 23704 12492 23724
rect 12492 23704 12494 23724
rect 11334 22752 11390 22808
rect 11978 22636 12034 22672
rect 11978 22616 11980 22636
rect 11980 22616 12032 22636
rect 12032 22616 12034 22636
rect 12162 23060 12164 23080
rect 12164 23060 12216 23080
rect 12216 23060 12218 23080
rect 12162 23024 12218 23060
rect 11242 21664 11298 21720
rect 12070 20848 12126 20904
rect 10874 20440 10930 20496
rect 12254 22072 12310 22128
rect 12162 20304 12218 20360
rect 12438 19352 12494 19408
rect 10598 17584 10654 17640
rect 10220 17434 10276 17436
rect 10300 17434 10356 17436
rect 10380 17434 10436 17436
rect 10460 17434 10516 17436
rect 10220 17382 10266 17434
rect 10266 17382 10276 17434
rect 10300 17382 10330 17434
rect 10330 17382 10342 17434
rect 10342 17382 10356 17434
rect 10380 17382 10394 17434
rect 10394 17382 10406 17434
rect 10406 17382 10436 17434
rect 10460 17382 10470 17434
rect 10470 17382 10516 17434
rect 10220 17380 10276 17382
rect 10300 17380 10356 17382
rect 10380 17380 10436 17382
rect 10460 17380 10516 17382
rect 10220 16346 10276 16348
rect 10300 16346 10356 16348
rect 10380 16346 10436 16348
rect 10460 16346 10516 16348
rect 10220 16294 10266 16346
rect 10266 16294 10276 16346
rect 10300 16294 10330 16346
rect 10330 16294 10342 16346
rect 10342 16294 10356 16346
rect 10380 16294 10394 16346
rect 10394 16294 10406 16346
rect 10406 16294 10436 16346
rect 10460 16294 10470 16346
rect 10470 16294 10516 16346
rect 10220 16292 10276 16294
rect 10300 16292 10356 16294
rect 10380 16292 10436 16294
rect 10460 16292 10516 16294
rect 10220 15258 10276 15260
rect 10300 15258 10356 15260
rect 10380 15258 10436 15260
rect 10460 15258 10516 15260
rect 10220 15206 10266 15258
rect 10266 15206 10276 15258
rect 10300 15206 10330 15258
rect 10330 15206 10342 15258
rect 10342 15206 10356 15258
rect 10380 15206 10394 15258
rect 10394 15206 10406 15258
rect 10406 15206 10436 15258
rect 10460 15206 10470 15258
rect 10470 15206 10516 15258
rect 10220 15204 10276 15206
rect 10300 15204 10356 15206
rect 10380 15204 10436 15206
rect 10460 15204 10516 15206
rect 10220 14170 10276 14172
rect 10300 14170 10356 14172
rect 10380 14170 10436 14172
rect 10460 14170 10516 14172
rect 10220 14118 10266 14170
rect 10266 14118 10276 14170
rect 10300 14118 10330 14170
rect 10330 14118 10342 14170
rect 10342 14118 10356 14170
rect 10380 14118 10394 14170
rect 10394 14118 10406 14170
rect 10406 14118 10436 14170
rect 10460 14118 10470 14170
rect 10470 14118 10516 14170
rect 10220 14116 10276 14118
rect 10300 14116 10356 14118
rect 10380 14116 10436 14118
rect 10460 14116 10516 14118
rect 10220 13082 10276 13084
rect 10300 13082 10356 13084
rect 10380 13082 10436 13084
rect 10460 13082 10516 13084
rect 10220 13030 10266 13082
rect 10266 13030 10276 13082
rect 10300 13030 10330 13082
rect 10330 13030 10342 13082
rect 10342 13030 10356 13082
rect 10380 13030 10394 13082
rect 10394 13030 10406 13082
rect 10406 13030 10436 13082
rect 10460 13030 10470 13082
rect 10470 13030 10516 13082
rect 10220 13028 10276 13030
rect 10300 13028 10356 13030
rect 10380 13028 10436 13030
rect 10460 13028 10516 13030
rect 10220 11994 10276 11996
rect 10300 11994 10356 11996
rect 10380 11994 10436 11996
rect 10460 11994 10516 11996
rect 10220 11942 10266 11994
rect 10266 11942 10276 11994
rect 10300 11942 10330 11994
rect 10330 11942 10342 11994
rect 10342 11942 10356 11994
rect 10380 11942 10394 11994
rect 10394 11942 10406 11994
rect 10406 11942 10436 11994
rect 10460 11942 10470 11994
rect 10470 11942 10516 11994
rect 10220 11940 10276 11942
rect 10300 11940 10356 11942
rect 10380 11940 10436 11942
rect 10460 11940 10516 11942
rect 10220 10906 10276 10908
rect 10300 10906 10356 10908
rect 10380 10906 10436 10908
rect 10460 10906 10516 10908
rect 10220 10854 10266 10906
rect 10266 10854 10276 10906
rect 10300 10854 10330 10906
rect 10330 10854 10342 10906
rect 10342 10854 10356 10906
rect 10380 10854 10394 10906
rect 10394 10854 10406 10906
rect 10406 10854 10436 10906
rect 10460 10854 10470 10906
rect 10470 10854 10516 10906
rect 10220 10852 10276 10854
rect 10300 10852 10356 10854
rect 10380 10852 10436 10854
rect 10460 10852 10516 10854
rect 10220 9818 10276 9820
rect 10300 9818 10356 9820
rect 10380 9818 10436 9820
rect 10460 9818 10516 9820
rect 10220 9766 10266 9818
rect 10266 9766 10276 9818
rect 10300 9766 10330 9818
rect 10330 9766 10342 9818
rect 10342 9766 10356 9818
rect 10380 9766 10394 9818
rect 10394 9766 10406 9818
rect 10406 9766 10436 9818
rect 10460 9766 10470 9818
rect 10470 9766 10516 9818
rect 10220 9764 10276 9766
rect 10300 9764 10356 9766
rect 10380 9764 10436 9766
rect 10460 9764 10516 9766
rect 10220 8730 10276 8732
rect 10300 8730 10356 8732
rect 10380 8730 10436 8732
rect 10460 8730 10516 8732
rect 10220 8678 10266 8730
rect 10266 8678 10276 8730
rect 10300 8678 10330 8730
rect 10330 8678 10342 8730
rect 10342 8678 10356 8730
rect 10380 8678 10394 8730
rect 10394 8678 10406 8730
rect 10406 8678 10436 8730
rect 10460 8678 10470 8730
rect 10470 8678 10516 8730
rect 10220 8676 10276 8678
rect 10300 8676 10356 8678
rect 10380 8676 10436 8678
rect 10460 8676 10516 8678
rect 10220 7642 10276 7644
rect 10300 7642 10356 7644
rect 10380 7642 10436 7644
rect 10460 7642 10516 7644
rect 10220 7590 10266 7642
rect 10266 7590 10276 7642
rect 10300 7590 10330 7642
rect 10330 7590 10342 7642
rect 10342 7590 10356 7642
rect 10380 7590 10394 7642
rect 10394 7590 10406 7642
rect 10406 7590 10436 7642
rect 10460 7590 10470 7642
rect 10470 7590 10516 7642
rect 10220 7588 10276 7590
rect 10300 7588 10356 7590
rect 10380 7588 10436 7590
rect 10460 7588 10516 7590
rect 12622 25064 12678 25120
rect 12990 24948 13046 24984
rect 12990 24928 12992 24948
rect 12992 24928 13044 24948
rect 13044 24928 13046 24948
rect 13174 24928 13230 24984
rect 12622 23024 12678 23080
rect 12622 21392 12678 21448
rect 13082 24384 13138 24440
rect 12898 24248 12954 24304
rect 13266 24112 13322 24168
rect 14186 28736 14242 28792
rect 16118 34720 16174 34776
rect 15566 33360 15622 33416
rect 14646 32136 14702 32192
rect 14852 32122 14908 32124
rect 14932 32122 14988 32124
rect 15012 32122 15068 32124
rect 15092 32122 15148 32124
rect 14852 32070 14898 32122
rect 14898 32070 14908 32122
rect 14932 32070 14962 32122
rect 14962 32070 14974 32122
rect 14974 32070 14988 32122
rect 15012 32070 15026 32122
rect 15026 32070 15038 32122
rect 15038 32070 15068 32122
rect 15092 32070 15102 32122
rect 15102 32070 15148 32122
rect 14852 32068 14908 32070
rect 14932 32068 14988 32070
rect 15012 32068 15068 32070
rect 15092 32068 15148 32070
rect 15290 32000 15346 32056
rect 14830 31748 14886 31784
rect 14830 31728 14832 31748
rect 14832 31728 14884 31748
rect 14884 31728 14886 31748
rect 15198 31728 15254 31784
rect 15106 31320 15162 31376
rect 15198 31184 15254 31240
rect 14462 30912 14518 30968
rect 14646 31048 14702 31104
rect 14852 31034 14908 31036
rect 14932 31034 14988 31036
rect 15012 31034 15068 31036
rect 15092 31034 15148 31036
rect 14852 30982 14898 31034
rect 14898 30982 14908 31034
rect 14932 30982 14962 31034
rect 14962 30982 14974 31034
rect 14974 30982 14988 31034
rect 15012 30982 15026 31034
rect 15026 30982 15038 31034
rect 15038 30982 15068 31034
rect 15092 30982 15102 31034
rect 15102 30982 15148 31034
rect 14852 30980 14908 30982
rect 14932 30980 14988 30982
rect 15012 30980 15068 30982
rect 15092 30980 15148 30982
rect 15474 30912 15530 30968
rect 14462 30504 14518 30560
rect 14370 29824 14426 29880
rect 14462 29552 14518 29608
rect 14186 27784 14242 27840
rect 13818 25900 13874 25936
rect 13818 25880 13820 25900
rect 13820 25880 13872 25900
rect 13872 25880 13874 25900
rect 14002 24828 14004 24848
rect 14004 24828 14056 24848
rect 14056 24828 14058 24848
rect 14002 24792 14058 24828
rect 14186 24656 14242 24712
rect 14462 27648 14518 27704
rect 14852 29946 14908 29948
rect 14932 29946 14988 29948
rect 15012 29946 15068 29948
rect 15092 29946 15148 29948
rect 14852 29894 14898 29946
rect 14898 29894 14908 29946
rect 14932 29894 14962 29946
rect 14962 29894 14974 29946
rect 14974 29894 14988 29946
rect 15012 29894 15026 29946
rect 15026 29894 15038 29946
rect 15038 29894 15068 29946
rect 15092 29894 15102 29946
rect 15102 29894 15148 29946
rect 14852 29892 14908 29894
rect 14932 29892 14988 29894
rect 15012 29892 15068 29894
rect 15092 29892 15148 29894
rect 15290 29824 15346 29880
rect 15198 29144 15254 29200
rect 15290 28872 15346 28928
rect 14852 28858 14908 28860
rect 14932 28858 14988 28860
rect 15012 28858 15068 28860
rect 15092 28858 15148 28860
rect 14852 28806 14898 28858
rect 14898 28806 14908 28858
rect 14932 28806 14962 28858
rect 14962 28806 14974 28858
rect 14974 28806 14988 28858
rect 15012 28806 15026 28858
rect 15026 28806 15038 28858
rect 15038 28806 15068 28858
rect 15092 28806 15102 28858
rect 15102 28806 15148 28858
rect 14852 28804 14908 28806
rect 14932 28804 14988 28806
rect 15012 28804 15068 28806
rect 15092 28804 15148 28806
rect 15290 28736 15346 28792
rect 14852 27770 14908 27772
rect 14932 27770 14988 27772
rect 15012 27770 15068 27772
rect 15092 27770 15148 27772
rect 14852 27718 14898 27770
rect 14898 27718 14908 27770
rect 14932 27718 14962 27770
rect 14962 27718 14974 27770
rect 14974 27718 14988 27770
rect 15012 27718 15026 27770
rect 15026 27718 15038 27770
rect 15038 27718 15068 27770
rect 15092 27718 15102 27770
rect 15102 27718 15148 27770
rect 14852 27716 14908 27718
rect 14932 27716 14988 27718
rect 15012 27716 15068 27718
rect 15092 27716 15148 27718
rect 14554 25744 14610 25800
rect 14852 26682 14908 26684
rect 14932 26682 14988 26684
rect 15012 26682 15068 26684
rect 15092 26682 15148 26684
rect 14852 26630 14898 26682
rect 14898 26630 14908 26682
rect 14932 26630 14962 26682
rect 14962 26630 14974 26682
rect 14974 26630 14988 26682
rect 15012 26630 15026 26682
rect 15026 26630 15038 26682
rect 15038 26630 15068 26682
rect 15092 26630 15102 26682
rect 15102 26630 15148 26682
rect 14852 26628 14908 26630
rect 14932 26628 14988 26630
rect 15012 26628 15068 26630
rect 15092 26628 15148 26630
rect 15842 29960 15898 30016
rect 15474 29144 15530 29200
rect 16302 31320 16358 31376
rect 16210 31184 16266 31240
rect 15934 29280 15990 29336
rect 15382 27940 15438 27976
rect 15382 27920 15384 27940
rect 15384 27920 15436 27940
rect 15436 27920 15438 27940
rect 15382 26288 15438 26344
rect 15658 26696 15714 26752
rect 15566 26288 15622 26344
rect 16210 27784 16266 27840
rect 15474 25744 15530 25800
rect 14646 25608 14702 25664
rect 14852 25594 14908 25596
rect 14932 25594 14988 25596
rect 15012 25594 15068 25596
rect 15092 25594 15148 25596
rect 14852 25542 14898 25594
rect 14898 25542 14908 25594
rect 14932 25542 14962 25594
rect 14962 25542 14974 25594
rect 14974 25542 14988 25594
rect 15012 25542 15026 25594
rect 15026 25542 15038 25594
rect 15038 25542 15068 25594
rect 15092 25542 15102 25594
rect 15102 25542 15148 25594
rect 14852 25540 14908 25542
rect 14932 25540 14988 25542
rect 15012 25540 15068 25542
rect 15092 25540 15148 25542
rect 15290 25608 15346 25664
rect 13910 23568 13966 23624
rect 13266 22480 13322 22536
rect 13358 21972 13360 21992
rect 13360 21972 13412 21992
rect 13412 21972 13414 21992
rect 13358 21936 13414 21972
rect 13726 22752 13782 22808
rect 12990 20712 13046 20768
rect 13266 20576 13322 20632
rect 13634 21800 13690 21856
rect 13634 20440 13690 20496
rect 14186 23160 14242 23216
rect 14186 22924 14188 22944
rect 14188 22924 14240 22944
rect 14240 22924 14242 22944
rect 14186 22888 14242 22924
rect 14186 21936 14242 21992
rect 13910 20984 13966 21040
rect 14186 18300 14188 18320
rect 14188 18300 14240 18320
rect 14240 18300 14242 18320
rect 14186 18264 14242 18300
rect 10220 6554 10276 6556
rect 10300 6554 10356 6556
rect 10380 6554 10436 6556
rect 10460 6554 10516 6556
rect 10220 6502 10266 6554
rect 10266 6502 10276 6554
rect 10300 6502 10330 6554
rect 10330 6502 10342 6554
rect 10342 6502 10356 6554
rect 10380 6502 10394 6554
rect 10394 6502 10406 6554
rect 10406 6502 10436 6554
rect 10460 6502 10470 6554
rect 10470 6502 10516 6554
rect 10220 6500 10276 6502
rect 10300 6500 10356 6502
rect 10380 6500 10436 6502
rect 10460 6500 10516 6502
rect 10220 5466 10276 5468
rect 10300 5466 10356 5468
rect 10380 5466 10436 5468
rect 10460 5466 10516 5468
rect 10220 5414 10266 5466
rect 10266 5414 10276 5466
rect 10300 5414 10330 5466
rect 10330 5414 10342 5466
rect 10342 5414 10356 5466
rect 10380 5414 10394 5466
rect 10394 5414 10406 5466
rect 10406 5414 10436 5466
rect 10460 5414 10470 5466
rect 10470 5414 10516 5466
rect 10220 5412 10276 5414
rect 10300 5412 10356 5414
rect 10380 5412 10436 5414
rect 10460 5412 10516 5414
rect 10220 4378 10276 4380
rect 10300 4378 10356 4380
rect 10380 4378 10436 4380
rect 10460 4378 10516 4380
rect 10220 4326 10266 4378
rect 10266 4326 10276 4378
rect 10300 4326 10330 4378
rect 10330 4326 10342 4378
rect 10342 4326 10356 4378
rect 10380 4326 10394 4378
rect 10394 4326 10406 4378
rect 10406 4326 10436 4378
rect 10460 4326 10470 4378
rect 10470 4326 10516 4378
rect 10220 4324 10276 4326
rect 10300 4324 10356 4326
rect 10380 4324 10436 4326
rect 10460 4324 10516 4326
rect 10220 3290 10276 3292
rect 10300 3290 10356 3292
rect 10380 3290 10436 3292
rect 10460 3290 10516 3292
rect 10220 3238 10266 3290
rect 10266 3238 10276 3290
rect 10300 3238 10330 3290
rect 10330 3238 10342 3290
rect 10342 3238 10356 3290
rect 10380 3238 10394 3290
rect 10394 3238 10406 3290
rect 10406 3238 10436 3290
rect 10460 3238 10470 3290
rect 10470 3238 10516 3290
rect 10220 3236 10276 3238
rect 10300 3236 10356 3238
rect 10380 3236 10436 3238
rect 10460 3236 10516 3238
rect 10220 2202 10276 2204
rect 10300 2202 10356 2204
rect 10380 2202 10436 2204
rect 10460 2202 10516 2204
rect 10220 2150 10266 2202
rect 10266 2150 10276 2202
rect 10300 2150 10330 2202
rect 10330 2150 10342 2202
rect 10342 2150 10356 2202
rect 10380 2150 10394 2202
rect 10394 2150 10406 2202
rect 10406 2150 10436 2202
rect 10460 2150 10470 2202
rect 10470 2150 10516 2202
rect 10220 2148 10276 2150
rect 10300 2148 10356 2150
rect 10380 2148 10436 2150
rect 10460 2148 10516 2150
rect 14370 24112 14426 24168
rect 15566 25336 15622 25392
rect 14738 24656 14794 24712
rect 14646 24520 14702 24576
rect 14646 24384 14702 24440
rect 16026 25608 16082 25664
rect 15750 25200 15806 25256
rect 15382 24520 15438 24576
rect 14852 24506 14908 24508
rect 14932 24506 14988 24508
rect 15012 24506 15068 24508
rect 15092 24506 15148 24508
rect 14852 24454 14898 24506
rect 14898 24454 14908 24506
rect 14932 24454 14962 24506
rect 14962 24454 14974 24506
rect 14974 24454 14988 24506
rect 15012 24454 15026 24506
rect 15026 24454 15038 24506
rect 15038 24454 15068 24506
rect 15092 24454 15102 24506
rect 15102 24454 15148 24506
rect 14852 24452 14908 24454
rect 14932 24452 14988 24454
rect 15012 24452 15068 24454
rect 15092 24452 15148 24454
rect 15290 24384 15346 24440
rect 14738 23724 14794 23760
rect 14738 23704 14740 23724
rect 14740 23704 14792 23724
rect 14792 23704 14794 23724
rect 16118 24828 16120 24848
rect 16120 24828 16172 24848
rect 16172 24828 16174 24848
rect 16118 24792 16174 24828
rect 15842 24520 15898 24576
rect 16026 24520 16082 24576
rect 15934 24384 15990 24440
rect 16118 24384 16174 24440
rect 15014 23840 15070 23896
rect 15198 23840 15254 23896
rect 14922 23704 14978 23760
rect 15842 23840 15898 23896
rect 14462 23160 14518 23216
rect 14852 23418 14908 23420
rect 14932 23418 14988 23420
rect 15012 23418 15068 23420
rect 15092 23418 15148 23420
rect 14852 23366 14898 23418
rect 14898 23366 14908 23418
rect 14932 23366 14962 23418
rect 14962 23366 14974 23418
rect 14974 23366 14988 23418
rect 15012 23366 15026 23418
rect 15026 23366 15038 23418
rect 15038 23366 15068 23418
rect 15092 23366 15102 23418
rect 15102 23366 15148 23418
rect 14852 23364 14908 23366
rect 14932 23364 14988 23366
rect 15012 23364 15068 23366
rect 15092 23364 15148 23366
rect 14646 23296 14702 23352
rect 15278 23296 15334 23352
rect 14852 22330 14908 22332
rect 14932 22330 14988 22332
rect 15012 22330 15068 22332
rect 15092 22330 15148 22332
rect 14852 22278 14898 22330
rect 14898 22278 14908 22330
rect 14932 22278 14962 22330
rect 14962 22278 14974 22330
rect 14974 22278 14988 22330
rect 15012 22278 15026 22330
rect 15026 22278 15038 22330
rect 15038 22278 15068 22330
rect 15092 22278 15102 22330
rect 15102 22278 15148 22330
rect 14852 22276 14908 22278
rect 14932 22276 14988 22278
rect 15012 22276 15068 22278
rect 15092 22276 15148 22278
rect 15750 22636 15806 22672
rect 15750 22616 15752 22636
rect 15752 22616 15804 22636
rect 15804 22616 15806 22636
rect 15290 22344 15346 22400
rect 14370 21528 14426 21584
rect 14738 21664 14794 21720
rect 15474 22208 15530 22264
rect 14922 21664 14978 21720
rect 15474 21936 15530 21992
rect 14852 21242 14908 21244
rect 14932 21242 14988 21244
rect 15012 21242 15068 21244
rect 15092 21242 15148 21244
rect 14852 21190 14898 21242
rect 14898 21190 14908 21242
rect 14932 21190 14962 21242
rect 14962 21190 14974 21242
rect 14974 21190 14988 21242
rect 15012 21190 15026 21242
rect 15026 21190 15038 21242
rect 15038 21190 15068 21242
rect 15092 21190 15102 21242
rect 15102 21190 15148 21242
rect 14852 21188 14908 21190
rect 14932 21188 14988 21190
rect 15012 21188 15068 21190
rect 15092 21188 15148 21190
rect 14830 20848 14886 20904
rect 15382 20984 15438 21040
rect 14852 20154 14908 20156
rect 14932 20154 14988 20156
rect 15012 20154 15068 20156
rect 15092 20154 15148 20156
rect 14852 20102 14898 20154
rect 14898 20102 14908 20154
rect 14932 20102 14962 20154
rect 14962 20102 14974 20154
rect 14974 20102 14988 20154
rect 15012 20102 15026 20154
rect 15026 20102 15038 20154
rect 15038 20102 15068 20154
rect 15092 20102 15102 20154
rect 15102 20102 15148 20154
rect 14852 20100 14908 20102
rect 14932 20100 14988 20102
rect 15012 20100 15068 20102
rect 15092 20100 15148 20102
rect 15106 19896 15162 19952
rect 15106 19624 15162 19680
rect 14852 19066 14908 19068
rect 14932 19066 14988 19068
rect 15012 19066 15068 19068
rect 15092 19066 15148 19068
rect 14852 19014 14898 19066
rect 14898 19014 14908 19066
rect 14932 19014 14962 19066
rect 14962 19014 14974 19066
rect 14974 19014 14988 19066
rect 15012 19014 15026 19066
rect 15026 19014 15038 19066
rect 15038 19014 15068 19066
rect 15092 19014 15102 19066
rect 15102 19014 15148 19066
rect 14852 19012 14908 19014
rect 14932 19012 14988 19014
rect 15012 19012 15068 19014
rect 15092 19012 15148 19014
rect 14852 17978 14908 17980
rect 14932 17978 14988 17980
rect 15012 17978 15068 17980
rect 15092 17978 15148 17980
rect 14852 17926 14898 17978
rect 14898 17926 14908 17978
rect 14932 17926 14962 17978
rect 14962 17926 14974 17978
rect 14974 17926 14988 17978
rect 15012 17926 15026 17978
rect 15026 17926 15038 17978
rect 15038 17926 15068 17978
rect 15092 17926 15102 17978
rect 15102 17926 15148 17978
rect 14852 17924 14908 17926
rect 14932 17924 14988 17926
rect 15012 17924 15068 17926
rect 15092 17924 15148 17926
rect 16026 21936 16082 21992
rect 16118 21664 16174 21720
rect 15750 20984 15806 21040
rect 16026 21256 16082 21312
rect 16486 34720 16542 34776
rect 16762 35128 16818 35184
rect 16486 31864 16542 31920
rect 18418 39208 18474 39264
rect 17130 37984 17186 38040
rect 16946 37032 17002 37088
rect 16946 35944 17002 36000
rect 17866 37304 17922 37360
rect 17130 36352 17186 36408
rect 17038 35672 17094 35728
rect 17590 36216 17646 36272
rect 17774 36216 17830 36272
rect 17590 35944 17646 36000
rect 17498 35400 17554 35456
rect 17314 34856 17370 34912
rect 17590 35128 17646 35184
rect 17314 33224 17370 33280
rect 17314 32544 17370 32600
rect 16486 31340 16542 31376
rect 16486 31320 16488 31340
rect 16488 31320 16540 31340
rect 16540 31320 16542 31340
rect 16394 26288 16450 26344
rect 16578 26288 16634 26344
rect 16578 26036 16634 26072
rect 16578 26016 16580 26036
rect 16580 26016 16632 26036
rect 16632 26016 16634 26036
rect 14852 16890 14908 16892
rect 14932 16890 14988 16892
rect 15012 16890 15068 16892
rect 15092 16890 15148 16892
rect 14852 16838 14898 16890
rect 14898 16838 14908 16890
rect 14932 16838 14962 16890
rect 14962 16838 14974 16890
rect 14974 16838 14988 16890
rect 15012 16838 15026 16890
rect 15026 16838 15038 16890
rect 15038 16838 15068 16890
rect 15092 16838 15102 16890
rect 15102 16838 15148 16890
rect 14852 16836 14908 16838
rect 14932 16836 14988 16838
rect 15012 16836 15068 16838
rect 15092 16836 15148 16838
rect 14852 15802 14908 15804
rect 14932 15802 14988 15804
rect 15012 15802 15068 15804
rect 15092 15802 15148 15804
rect 14852 15750 14898 15802
rect 14898 15750 14908 15802
rect 14932 15750 14962 15802
rect 14962 15750 14974 15802
rect 14974 15750 14988 15802
rect 15012 15750 15026 15802
rect 15026 15750 15038 15802
rect 15038 15750 15068 15802
rect 15092 15750 15102 15802
rect 15102 15750 15148 15802
rect 14852 15748 14908 15750
rect 14932 15748 14988 15750
rect 15012 15748 15068 15750
rect 15092 15748 15148 15750
rect 14852 14714 14908 14716
rect 14932 14714 14988 14716
rect 15012 14714 15068 14716
rect 15092 14714 15148 14716
rect 14852 14662 14898 14714
rect 14898 14662 14908 14714
rect 14932 14662 14962 14714
rect 14962 14662 14974 14714
rect 14974 14662 14988 14714
rect 15012 14662 15026 14714
rect 15026 14662 15038 14714
rect 15038 14662 15068 14714
rect 15092 14662 15102 14714
rect 15102 14662 15148 14714
rect 14852 14660 14908 14662
rect 14932 14660 14988 14662
rect 15012 14660 15068 14662
rect 15092 14660 15148 14662
rect 14852 13626 14908 13628
rect 14932 13626 14988 13628
rect 15012 13626 15068 13628
rect 15092 13626 15148 13628
rect 14852 13574 14898 13626
rect 14898 13574 14908 13626
rect 14932 13574 14962 13626
rect 14962 13574 14974 13626
rect 14974 13574 14988 13626
rect 15012 13574 15026 13626
rect 15026 13574 15038 13626
rect 15038 13574 15068 13626
rect 15092 13574 15102 13626
rect 15102 13574 15148 13626
rect 14852 13572 14908 13574
rect 14932 13572 14988 13574
rect 15012 13572 15068 13574
rect 15092 13572 15148 13574
rect 14852 12538 14908 12540
rect 14932 12538 14988 12540
rect 15012 12538 15068 12540
rect 15092 12538 15148 12540
rect 14852 12486 14898 12538
rect 14898 12486 14908 12538
rect 14932 12486 14962 12538
rect 14962 12486 14974 12538
rect 14974 12486 14988 12538
rect 15012 12486 15026 12538
rect 15026 12486 15038 12538
rect 15038 12486 15068 12538
rect 15092 12486 15102 12538
rect 15102 12486 15148 12538
rect 14852 12484 14908 12486
rect 14932 12484 14988 12486
rect 15012 12484 15068 12486
rect 15092 12484 15148 12486
rect 17498 32444 17500 32464
rect 17500 32444 17552 32464
rect 17552 32444 17554 32464
rect 17498 32408 17554 32444
rect 17498 31592 17554 31648
rect 16946 30368 17002 30424
rect 16762 30232 16818 30288
rect 18234 35944 18290 36000
rect 18418 35944 18474 36000
rect 18878 36896 18934 36952
rect 18786 36624 18842 36680
rect 18234 35536 18290 35592
rect 17774 35128 17830 35184
rect 18050 34448 18106 34504
rect 20074 39616 20130 39672
rect 20074 39344 20130 39400
rect 19484 39194 19540 39196
rect 19564 39194 19620 39196
rect 19644 39194 19700 39196
rect 19724 39194 19780 39196
rect 19484 39142 19530 39194
rect 19530 39142 19540 39194
rect 19564 39142 19594 39194
rect 19594 39142 19606 39194
rect 19606 39142 19620 39194
rect 19644 39142 19658 39194
rect 19658 39142 19670 39194
rect 19670 39142 19700 39194
rect 19724 39142 19734 39194
rect 19734 39142 19780 39194
rect 19484 39140 19540 39142
rect 19564 39140 19620 39142
rect 19644 39140 19700 39142
rect 19724 39140 19780 39142
rect 19338 39072 19394 39128
rect 19062 38120 19118 38176
rect 19062 37440 19118 37496
rect 19484 38106 19540 38108
rect 19564 38106 19620 38108
rect 19644 38106 19700 38108
rect 19724 38106 19780 38108
rect 19484 38054 19530 38106
rect 19530 38054 19540 38106
rect 19564 38054 19594 38106
rect 19594 38054 19606 38106
rect 19606 38054 19620 38106
rect 19644 38054 19658 38106
rect 19658 38054 19670 38106
rect 19670 38054 19700 38106
rect 19724 38054 19734 38106
rect 19734 38054 19780 38106
rect 19484 38052 19540 38054
rect 19564 38052 19620 38054
rect 19644 38052 19700 38054
rect 19724 38052 19780 38054
rect 19982 38664 20038 38720
rect 19614 37732 19670 37768
rect 19614 37712 19616 37732
rect 19616 37712 19668 37732
rect 19668 37712 19670 37732
rect 19614 37188 19670 37224
rect 19614 37168 19616 37188
rect 19616 37168 19668 37188
rect 19668 37168 19670 37188
rect 19484 37018 19540 37020
rect 19564 37018 19620 37020
rect 19644 37018 19700 37020
rect 19724 37018 19780 37020
rect 19484 36966 19530 37018
rect 19530 36966 19540 37018
rect 19564 36966 19594 37018
rect 19594 36966 19606 37018
rect 19606 36966 19620 37018
rect 19644 36966 19658 37018
rect 19658 36966 19670 37018
rect 19670 36966 19700 37018
rect 19724 36966 19734 37018
rect 19734 36966 19780 37018
rect 19484 36964 19540 36966
rect 19564 36964 19620 36966
rect 19644 36964 19700 36966
rect 19724 36964 19780 36966
rect 19338 36896 19394 36952
rect 19062 36624 19118 36680
rect 19246 36644 19302 36680
rect 19246 36624 19248 36644
rect 19248 36624 19300 36644
rect 19300 36624 19302 36644
rect 19154 36080 19210 36136
rect 19338 35944 19394 36000
rect 19890 35944 19946 36000
rect 19484 35930 19540 35932
rect 19564 35930 19620 35932
rect 19644 35930 19700 35932
rect 19724 35930 19780 35932
rect 19484 35878 19530 35930
rect 19530 35878 19540 35930
rect 19564 35878 19594 35930
rect 19594 35878 19606 35930
rect 19606 35878 19620 35930
rect 19644 35878 19658 35930
rect 19658 35878 19670 35930
rect 19670 35878 19700 35930
rect 19724 35878 19734 35930
rect 19734 35878 19780 35930
rect 19484 35876 19540 35878
rect 19564 35876 19620 35878
rect 19644 35876 19700 35878
rect 19724 35876 19780 35878
rect 19338 35808 19394 35864
rect 18418 34856 18474 34912
rect 18786 34720 18842 34776
rect 17866 34176 17922 34232
rect 18234 34448 18290 34504
rect 18050 33108 18106 33144
rect 18050 33088 18052 33108
rect 18052 33088 18104 33108
rect 18104 33088 18106 33108
rect 16946 29824 17002 29880
rect 16854 29280 16910 29336
rect 17130 30096 17186 30152
rect 16762 28600 16818 28656
rect 16946 28600 17002 28656
rect 16854 28056 16910 28112
rect 17130 28192 17186 28248
rect 16854 27648 16910 27704
rect 16946 26560 17002 26616
rect 17774 30912 17830 30968
rect 19522 35400 19578 35456
rect 19484 34842 19540 34844
rect 19564 34842 19620 34844
rect 19644 34842 19700 34844
rect 19724 34842 19780 34844
rect 19484 34790 19530 34842
rect 19530 34790 19540 34842
rect 19564 34790 19594 34842
rect 19594 34790 19606 34842
rect 19606 34790 19620 34842
rect 19644 34790 19658 34842
rect 19658 34790 19670 34842
rect 19670 34790 19700 34842
rect 19724 34790 19734 34842
rect 19734 34790 19780 34842
rect 19484 34788 19540 34790
rect 19564 34788 19620 34790
rect 19644 34788 19700 34790
rect 19724 34788 19780 34790
rect 19062 34312 19118 34368
rect 18418 32952 18474 33008
rect 18694 33632 18750 33688
rect 18694 32952 18750 33008
rect 17774 29960 17830 30016
rect 17498 29688 17554 29744
rect 17590 28872 17646 28928
rect 17406 28328 17462 28384
rect 17314 27512 17370 27568
rect 17406 27240 17462 27296
rect 17222 25608 17278 25664
rect 16946 25064 17002 25120
rect 17130 24948 17186 24984
rect 17130 24928 17132 24948
rect 17132 24928 17184 24948
rect 17184 24928 17186 24948
rect 17958 29688 18014 29744
rect 18050 29008 18106 29064
rect 18418 30096 18474 30152
rect 18418 29280 18474 29336
rect 18418 28464 18474 28520
rect 18142 27512 18198 27568
rect 17958 27276 17960 27296
rect 17960 27276 18012 27296
rect 18012 27276 18014 27296
rect 17958 27240 18014 27276
rect 16762 22888 16818 22944
rect 16486 22208 16542 22264
rect 16578 21800 16634 21856
rect 16578 21664 16634 21720
rect 16578 21120 16634 21176
rect 16762 21664 16818 21720
rect 14852 11450 14908 11452
rect 14932 11450 14988 11452
rect 15012 11450 15068 11452
rect 15092 11450 15148 11452
rect 14852 11398 14898 11450
rect 14898 11398 14908 11450
rect 14932 11398 14962 11450
rect 14962 11398 14974 11450
rect 14974 11398 14988 11450
rect 15012 11398 15026 11450
rect 15026 11398 15038 11450
rect 15038 11398 15068 11450
rect 15092 11398 15102 11450
rect 15102 11398 15148 11450
rect 14852 11396 14908 11398
rect 14932 11396 14988 11398
rect 15012 11396 15068 11398
rect 15092 11396 15148 11398
rect 14852 10362 14908 10364
rect 14932 10362 14988 10364
rect 15012 10362 15068 10364
rect 15092 10362 15148 10364
rect 14852 10310 14898 10362
rect 14898 10310 14908 10362
rect 14932 10310 14962 10362
rect 14962 10310 14974 10362
rect 14974 10310 14988 10362
rect 15012 10310 15026 10362
rect 15026 10310 15038 10362
rect 15038 10310 15068 10362
rect 15092 10310 15102 10362
rect 15102 10310 15148 10362
rect 14852 10308 14908 10310
rect 14932 10308 14988 10310
rect 15012 10308 15068 10310
rect 15092 10308 15148 10310
rect 14852 9274 14908 9276
rect 14932 9274 14988 9276
rect 15012 9274 15068 9276
rect 15092 9274 15148 9276
rect 14852 9222 14898 9274
rect 14898 9222 14908 9274
rect 14932 9222 14962 9274
rect 14962 9222 14974 9274
rect 14974 9222 14988 9274
rect 15012 9222 15026 9274
rect 15026 9222 15038 9274
rect 15038 9222 15068 9274
rect 15092 9222 15102 9274
rect 15102 9222 15148 9274
rect 14852 9220 14908 9222
rect 14932 9220 14988 9222
rect 15012 9220 15068 9222
rect 15092 9220 15148 9222
rect 14852 8186 14908 8188
rect 14932 8186 14988 8188
rect 15012 8186 15068 8188
rect 15092 8186 15148 8188
rect 14852 8134 14898 8186
rect 14898 8134 14908 8186
rect 14932 8134 14962 8186
rect 14962 8134 14974 8186
rect 14974 8134 14988 8186
rect 15012 8134 15026 8186
rect 15026 8134 15038 8186
rect 15038 8134 15068 8186
rect 15092 8134 15102 8186
rect 15102 8134 15148 8186
rect 14852 8132 14908 8134
rect 14932 8132 14988 8134
rect 15012 8132 15068 8134
rect 15092 8132 15148 8134
rect 14852 7098 14908 7100
rect 14932 7098 14988 7100
rect 15012 7098 15068 7100
rect 15092 7098 15148 7100
rect 14852 7046 14898 7098
rect 14898 7046 14908 7098
rect 14932 7046 14962 7098
rect 14962 7046 14974 7098
rect 14974 7046 14988 7098
rect 15012 7046 15026 7098
rect 15026 7046 15038 7098
rect 15038 7046 15068 7098
rect 15092 7046 15102 7098
rect 15102 7046 15148 7098
rect 14852 7044 14908 7046
rect 14932 7044 14988 7046
rect 15012 7044 15068 7046
rect 15092 7044 15148 7046
rect 14852 6010 14908 6012
rect 14932 6010 14988 6012
rect 15012 6010 15068 6012
rect 15092 6010 15148 6012
rect 14852 5958 14898 6010
rect 14898 5958 14908 6010
rect 14932 5958 14962 6010
rect 14962 5958 14974 6010
rect 14974 5958 14988 6010
rect 15012 5958 15026 6010
rect 15026 5958 15038 6010
rect 15038 5958 15068 6010
rect 15092 5958 15102 6010
rect 15102 5958 15148 6010
rect 14852 5956 14908 5958
rect 14932 5956 14988 5958
rect 15012 5956 15068 5958
rect 15092 5956 15148 5958
rect 14852 4922 14908 4924
rect 14932 4922 14988 4924
rect 15012 4922 15068 4924
rect 15092 4922 15148 4924
rect 14852 4870 14898 4922
rect 14898 4870 14908 4922
rect 14932 4870 14962 4922
rect 14962 4870 14974 4922
rect 14974 4870 14988 4922
rect 15012 4870 15026 4922
rect 15026 4870 15038 4922
rect 15038 4870 15068 4922
rect 15092 4870 15102 4922
rect 15102 4870 15148 4922
rect 14852 4868 14908 4870
rect 14932 4868 14988 4870
rect 15012 4868 15068 4870
rect 15092 4868 15148 4870
rect 14852 3834 14908 3836
rect 14932 3834 14988 3836
rect 15012 3834 15068 3836
rect 15092 3834 15148 3836
rect 14852 3782 14898 3834
rect 14898 3782 14908 3834
rect 14932 3782 14962 3834
rect 14962 3782 14974 3834
rect 14974 3782 14988 3834
rect 15012 3782 15026 3834
rect 15026 3782 15038 3834
rect 15038 3782 15068 3834
rect 15092 3782 15102 3834
rect 15102 3782 15148 3834
rect 14852 3780 14908 3782
rect 14932 3780 14988 3782
rect 15012 3780 15068 3782
rect 15092 3780 15148 3782
rect 14852 2746 14908 2748
rect 14932 2746 14988 2748
rect 15012 2746 15068 2748
rect 15092 2746 15148 2748
rect 14852 2694 14898 2746
rect 14898 2694 14908 2746
rect 14932 2694 14962 2746
rect 14962 2694 14974 2746
rect 14974 2694 14988 2746
rect 15012 2694 15026 2746
rect 15026 2694 15038 2746
rect 15038 2694 15068 2746
rect 15092 2694 15102 2746
rect 15102 2694 15148 2746
rect 14852 2692 14908 2694
rect 14932 2692 14988 2694
rect 15012 2692 15068 2694
rect 15092 2692 15148 2694
rect 16946 23296 17002 23352
rect 16946 23160 17002 23216
rect 16854 19896 16910 19952
rect 16854 19352 16910 19408
rect 17038 19624 17094 19680
rect 17498 22208 17554 22264
rect 18142 26732 18144 26752
rect 18144 26732 18196 26752
rect 18196 26732 18198 26752
rect 17958 26152 18014 26208
rect 18142 26696 18198 26732
rect 18418 27240 18474 27296
rect 19338 34312 19394 34368
rect 19338 33768 19394 33824
rect 19484 33754 19540 33756
rect 19564 33754 19620 33756
rect 19644 33754 19700 33756
rect 19724 33754 19780 33756
rect 19484 33702 19530 33754
rect 19530 33702 19540 33754
rect 19564 33702 19594 33754
rect 19594 33702 19606 33754
rect 19606 33702 19620 33754
rect 19644 33702 19658 33754
rect 19658 33702 19670 33754
rect 19670 33702 19700 33754
rect 19724 33702 19734 33754
rect 19734 33702 19780 33754
rect 19484 33700 19540 33702
rect 19564 33700 19620 33702
rect 19644 33700 19700 33702
rect 19724 33700 19780 33702
rect 20166 35944 20222 36000
rect 20350 35808 20406 35864
rect 20534 37304 20590 37360
rect 20534 35128 20590 35184
rect 20166 34856 20222 34912
rect 19338 32716 19340 32736
rect 19340 32716 19392 32736
rect 19392 32716 19394 32736
rect 19338 32680 19394 32716
rect 19484 32666 19540 32668
rect 19564 32666 19620 32668
rect 19644 32666 19700 32668
rect 19724 32666 19780 32668
rect 19484 32614 19530 32666
rect 19530 32614 19540 32666
rect 19564 32614 19594 32666
rect 19594 32614 19606 32666
rect 19606 32614 19620 32666
rect 19644 32614 19658 32666
rect 19658 32614 19670 32666
rect 19670 32614 19700 32666
rect 19724 32614 19734 32666
rect 19734 32614 19780 32666
rect 19484 32612 19540 32614
rect 19564 32612 19620 32614
rect 19644 32612 19700 32614
rect 19724 32612 19780 32614
rect 19338 32408 19394 32464
rect 19522 32136 19578 32192
rect 19246 32000 19302 32056
rect 19154 31184 19210 31240
rect 19062 30640 19118 30696
rect 18878 30504 18934 30560
rect 18602 27648 18658 27704
rect 18418 26580 18474 26616
rect 18418 26560 18420 26580
rect 18420 26560 18472 26580
rect 18472 26560 18474 26580
rect 18142 24792 18198 24848
rect 18878 27376 18934 27432
rect 18878 26424 18934 26480
rect 17682 22888 17738 22944
rect 17774 22752 17830 22808
rect 18234 23976 18290 24032
rect 18418 23976 18474 24032
rect 18142 23160 18198 23216
rect 18326 23296 18382 23352
rect 18326 23160 18382 23216
rect 17958 22616 18014 22672
rect 18050 22344 18106 22400
rect 19484 31578 19540 31580
rect 19564 31578 19620 31580
rect 19644 31578 19700 31580
rect 19724 31578 19780 31580
rect 19484 31526 19530 31578
rect 19530 31526 19540 31578
rect 19564 31526 19594 31578
rect 19594 31526 19606 31578
rect 19606 31526 19620 31578
rect 19644 31526 19658 31578
rect 19658 31526 19670 31578
rect 19670 31526 19700 31578
rect 19724 31526 19734 31578
rect 19734 31526 19780 31578
rect 19484 31524 19540 31526
rect 19564 31524 19620 31526
rect 19644 31524 19700 31526
rect 19724 31524 19780 31526
rect 19614 30676 19616 30696
rect 19616 30676 19668 30696
rect 19668 30676 19670 30696
rect 19614 30640 19670 30676
rect 20534 34720 20590 34776
rect 20350 32000 20406 32056
rect 20902 37848 20958 37904
rect 20810 36660 20812 36680
rect 20812 36660 20864 36680
rect 20864 36660 20866 36680
rect 20810 36624 20866 36660
rect 20810 36524 20812 36544
rect 20812 36524 20864 36544
rect 20864 36524 20866 36544
rect 20810 36488 20866 36524
rect 20902 36216 20958 36272
rect 20810 35672 20866 35728
rect 21178 38528 21234 38584
rect 20994 35672 21050 35728
rect 21086 35400 21142 35456
rect 20902 35128 20958 35184
rect 20810 34856 20866 34912
rect 20810 34584 20866 34640
rect 20902 34312 20958 34368
rect 21822 39752 21878 39808
rect 21270 35944 21326 36000
rect 21270 34892 21272 34912
rect 21272 34892 21324 34912
rect 21324 34892 21326 34912
rect 21270 34856 21326 34892
rect 21178 34312 21234 34368
rect 21178 34040 21234 34096
rect 20902 32952 20958 33008
rect 19484 30490 19540 30492
rect 19564 30490 19620 30492
rect 19644 30490 19700 30492
rect 19724 30490 19780 30492
rect 19484 30438 19530 30490
rect 19530 30438 19540 30490
rect 19564 30438 19594 30490
rect 19594 30438 19606 30490
rect 19606 30438 19620 30490
rect 19644 30438 19658 30490
rect 19658 30438 19670 30490
rect 19670 30438 19700 30490
rect 19724 30438 19734 30490
rect 19734 30438 19780 30490
rect 19484 30436 19540 30438
rect 19564 30436 19620 30438
rect 19644 30436 19700 30438
rect 19724 30436 19780 30438
rect 19430 30096 19486 30152
rect 19246 29688 19302 29744
rect 19338 29552 19394 29608
rect 19062 29416 19118 29472
rect 19484 29402 19540 29404
rect 19564 29402 19620 29404
rect 19644 29402 19700 29404
rect 19724 29402 19780 29404
rect 19484 29350 19530 29402
rect 19530 29350 19540 29402
rect 19564 29350 19594 29402
rect 19594 29350 19606 29402
rect 19606 29350 19620 29402
rect 19644 29350 19658 29402
rect 19658 29350 19670 29402
rect 19670 29350 19700 29402
rect 19724 29350 19734 29402
rect 19734 29350 19780 29402
rect 19484 29348 19540 29350
rect 19564 29348 19620 29350
rect 19644 29348 19700 29350
rect 19724 29348 19780 29350
rect 19982 30096 20038 30152
rect 19338 28736 19394 28792
rect 19890 28736 19946 28792
rect 19798 28600 19854 28656
rect 19062 28464 19118 28520
rect 19062 26696 19118 26752
rect 19706 28464 19762 28520
rect 19246 27784 19302 27840
rect 19484 28314 19540 28316
rect 19564 28314 19620 28316
rect 19644 28314 19700 28316
rect 19724 28314 19780 28316
rect 19484 28262 19530 28314
rect 19530 28262 19540 28314
rect 19564 28262 19594 28314
rect 19594 28262 19606 28314
rect 19606 28262 19620 28314
rect 19644 28262 19658 28314
rect 19658 28262 19670 28314
rect 19670 28262 19700 28314
rect 19724 28262 19734 28314
rect 19734 28262 19780 28314
rect 19484 28260 19540 28262
rect 19564 28260 19620 28262
rect 19644 28260 19700 28262
rect 19724 28260 19780 28262
rect 19484 27226 19540 27228
rect 19564 27226 19620 27228
rect 19644 27226 19700 27228
rect 19724 27226 19780 27228
rect 19484 27174 19530 27226
rect 19530 27174 19540 27226
rect 19564 27174 19594 27226
rect 19594 27174 19606 27226
rect 19606 27174 19620 27226
rect 19644 27174 19658 27226
rect 19658 27174 19670 27226
rect 19670 27174 19700 27226
rect 19724 27174 19734 27226
rect 19734 27174 19780 27226
rect 19484 27172 19540 27174
rect 19564 27172 19620 27174
rect 19644 27172 19700 27174
rect 19724 27172 19780 27174
rect 18602 23160 18658 23216
rect 18510 22636 18566 22672
rect 18510 22616 18512 22636
rect 18512 22616 18564 22636
rect 18564 22616 18566 22636
rect 18326 21972 18328 21992
rect 18328 21972 18380 21992
rect 18380 21972 18382 21992
rect 17774 20848 17830 20904
rect 18326 21936 18382 21972
rect 18510 21664 18566 21720
rect 18786 23976 18842 24032
rect 18786 23860 18842 23896
rect 19154 25744 19210 25800
rect 19154 25356 19210 25392
rect 19154 25336 19156 25356
rect 19156 25336 19208 25356
rect 19208 25336 19210 25356
rect 19706 26308 19762 26344
rect 19706 26288 19708 26308
rect 19708 26288 19760 26308
rect 19760 26288 19762 26308
rect 19484 26138 19540 26140
rect 19564 26138 19620 26140
rect 19644 26138 19700 26140
rect 19724 26138 19780 26140
rect 19484 26086 19530 26138
rect 19530 26086 19540 26138
rect 19564 26086 19594 26138
rect 19594 26086 19606 26138
rect 19606 26086 19620 26138
rect 19644 26086 19658 26138
rect 19658 26086 19670 26138
rect 19670 26086 19700 26138
rect 19724 26086 19734 26138
rect 19734 26086 19780 26138
rect 19484 26084 19540 26086
rect 19564 26084 19620 26086
rect 19644 26084 19700 26086
rect 19724 26084 19780 26086
rect 19890 25336 19946 25392
rect 18786 23840 18788 23860
rect 18788 23840 18840 23860
rect 18840 23840 18842 23860
rect 19062 22888 19118 22944
rect 19890 25100 19892 25120
rect 19892 25100 19944 25120
rect 19944 25100 19946 25120
rect 19890 25064 19946 25100
rect 19484 25050 19540 25052
rect 19564 25050 19620 25052
rect 19644 25050 19700 25052
rect 19724 25050 19780 25052
rect 19484 24998 19530 25050
rect 19530 24998 19540 25050
rect 19564 24998 19594 25050
rect 19594 24998 19606 25050
rect 19606 24998 19620 25050
rect 19644 24998 19658 25050
rect 19658 24998 19670 25050
rect 19670 24998 19700 25050
rect 19724 24998 19734 25050
rect 19734 24998 19780 25050
rect 19484 24996 19540 24998
rect 19564 24996 19620 24998
rect 19644 24996 19700 24998
rect 19724 24996 19780 24998
rect 19338 24384 19394 24440
rect 19484 23962 19540 23964
rect 19564 23962 19620 23964
rect 19644 23962 19700 23964
rect 19724 23962 19780 23964
rect 19484 23910 19530 23962
rect 19530 23910 19540 23962
rect 19564 23910 19594 23962
rect 19594 23910 19606 23962
rect 19606 23910 19620 23962
rect 19644 23910 19658 23962
rect 19658 23910 19670 23962
rect 19670 23910 19700 23962
rect 19724 23910 19734 23962
rect 19734 23910 19780 23962
rect 19484 23908 19540 23910
rect 19564 23908 19620 23910
rect 19644 23908 19700 23910
rect 19724 23908 19780 23910
rect 19706 23296 19762 23352
rect 19798 23180 19854 23216
rect 19798 23160 19800 23180
rect 19800 23160 19852 23180
rect 19852 23160 19854 23180
rect 19484 22874 19540 22876
rect 19564 22874 19620 22876
rect 19644 22874 19700 22876
rect 19724 22874 19780 22876
rect 19484 22822 19530 22874
rect 19530 22822 19540 22874
rect 19564 22822 19594 22874
rect 19594 22822 19606 22874
rect 19606 22822 19620 22874
rect 19644 22822 19658 22874
rect 19658 22822 19670 22874
rect 19670 22822 19700 22874
rect 19724 22822 19734 22874
rect 19734 22822 19780 22874
rect 19484 22820 19540 22822
rect 19564 22820 19620 22822
rect 19644 22820 19700 22822
rect 19724 22820 19780 22822
rect 19614 22480 19670 22536
rect 19798 22480 19854 22536
rect 19614 22092 19670 22128
rect 19614 22072 19616 22092
rect 19616 22072 19668 22092
rect 19668 22072 19670 22092
rect 19484 21786 19540 21788
rect 19564 21786 19620 21788
rect 19644 21786 19700 21788
rect 19724 21786 19780 21788
rect 19484 21734 19530 21786
rect 19530 21734 19540 21786
rect 19564 21734 19594 21786
rect 19594 21734 19606 21786
rect 19606 21734 19620 21786
rect 19644 21734 19658 21786
rect 19658 21734 19670 21786
rect 19670 21734 19700 21786
rect 19724 21734 19734 21786
rect 19734 21734 19780 21786
rect 19484 21732 19540 21734
rect 19564 21732 19620 21734
rect 19644 21732 19700 21734
rect 19724 21732 19780 21734
rect 19154 21256 19210 21312
rect 18510 20748 18512 20768
rect 18512 20748 18564 20768
rect 18564 20748 18566 20768
rect 18510 20712 18566 20748
rect 18878 20576 18934 20632
rect 19484 20698 19540 20700
rect 19564 20698 19620 20700
rect 19644 20698 19700 20700
rect 19724 20698 19780 20700
rect 19484 20646 19530 20698
rect 19530 20646 19540 20698
rect 19564 20646 19594 20698
rect 19594 20646 19606 20698
rect 19606 20646 19620 20698
rect 19644 20646 19658 20698
rect 19658 20646 19670 20698
rect 19670 20646 19700 20698
rect 19724 20646 19734 20698
rect 19734 20646 19780 20698
rect 19484 20644 19540 20646
rect 19564 20644 19620 20646
rect 19644 20644 19700 20646
rect 19724 20644 19780 20646
rect 18326 18264 18382 18320
rect 19484 19610 19540 19612
rect 19564 19610 19620 19612
rect 19644 19610 19700 19612
rect 19724 19610 19780 19612
rect 19484 19558 19530 19610
rect 19530 19558 19540 19610
rect 19564 19558 19594 19610
rect 19594 19558 19606 19610
rect 19606 19558 19620 19610
rect 19644 19558 19658 19610
rect 19658 19558 19670 19610
rect 19670 19558 19700 19610
rect 19724 19558 19734 19610
rect 19734 19558 19780 19610
rect 19484 19556 19540 19558
rect 19564 19556 19620 19558
rect 19644 19556 19700 19558
rect 19724 19556 19780 19558
rect 19484 18522 19540 18524
rect 19564 18522 19620 18524
rect 19644 18522 19700 18524
rect 19724 18522 19780 18524
rect 19484 18470 19530 18522
rect 19530 18470 19540 18522
rect 19564 18470 19594 18522
rect 19594 18470 19606 18522
rect 19606 18470 19620 18522
rect 19644 18470 19658 18522
rect 19658 18470 19670 18522
rect 19670 18470 19700 18522
rect 19724 18470 19734 18522
rect 19734 18470 19780 18522
rect 19484 18468 19540 18470
rect 19564 18468 19620 18470
rect 19644 18468 19700 18470
rect 19724 18468 19780 18470
rect 19484 17434 19540 17436
rect 19564 17434 19620 17436
rect 19644 17434 19700 17436
rect 19724 17434 19780 17436
rect 19484 17382 19530 17434
rect 19530 17382 19540 17434
rect 19564 17382 19594 17434
rect 19594 17382 19606 17434
rect 19606 17382 19620 17434
rect 19644 17382 19658 17434
rect 19658 17382 19670 17434
rect 19670 17382 19700 17434
rect 19724 17382 19734 17434
rect 19734 17382 19780 17434
rect 19484 17380 19540 17382
rect 19564 17380 19620 17382
rect 19644 17380 19700 17382
rect 19724 17380 19780 17382
rect 19484 16346 19540 16348
rect 19564 16346 19620 16348
rect 19644 16346 19700 16348
rect 19724 16346 19780 16348
rect 19484 16294 19530 16346
rect 19530 16294 19540 16346
rect 19564 16294 19594 16346
rect 19594 16294 19606 16346
rect 19606 16294 19620 16346
rect 19644 16294 19658 16346
rect 19658 16294 19670 16346
rect 19670 16294 19700 16346
rect 19724 16294 19734 16346
rect 19734 16294 19780 16346
rect 19484 16292 19540 16294
rect 19564 16292 19620 16294
rect 19644 16292 19700 16294
rect 19724 16292 19780 16294
rect 19484 15258 19540 15260
rect 19564 15258 19620 15260
rect 19644 15258 19700 15260
rect 19724 15258 19780 15260
rect 19484 15206 19530 15258
rect 19530 15206 19540 15258
rect 19564 15206 19594 15258
rect 19594 15206 19606 15258
rect 19606 15206 19620 15258
rect 19644 15206 19658 15258
rect 19658 15206 19670 15258
rect 19670 15206 19700 15258
rect 19724 15206 19734 15258
rect 19734 15206 19780 15258
rect 19484 15204 19540 15206
rect 19564 15204 19620 15206
rect 19644 15204 19700 15206
rect 19724 15204 19780 15206
rect 19484 14170 19540 14172
rect 19564 14170 19620 14172
rect 19644 14170 19700 14172
rect 19724 14170 19780 14172
rect 19484 14118 19530 14170
rect 19530 14118 19540 14170
rect 19564 14118 19594 14170
rect 19594 14118 19606 14170
rect 19606 14118 19620 14170
rect 19644 14118 19658 14170
rect 19658 14118 19670 14170
rect 19670 14118 19700 14170
rect 19724 14118 19734 14170
rect 19734 14118 19780 14170
rect 19484 14116 19540 14118
rect 19564 14116 19620 14118
rect 19644 14116 19700 14118
rect 19724 14116 19780 14118
rect 19484 13082 19540 13084
rect 19564 13082 19620 13084
rect 19644 13082 19700 13084
rect 19724 13082 19780 13084
rect 19484 13030 19530 13082
rect 19530 13030 19540 13082
rect 19564 13030 19594 13082
rect 19594 13030 19606 13082
rect 19606 13030 19620 13082
rect 19644 13030 19658 13082
rect 19658 13030 19670 13082
rect 19670 13030 19700 13082
rect 19724 13030 19734 13082
rect 19734 13030 19780 13082
rect 19484 13028 19540 13030
rect 19564 13028 19620 13030
rect 19644 13028 19700 13030
rect 19724 13028 19780 13030
rect 19484 11994 19540 11996
rect 19564 11994 19620 11996
rect 19644 11994 19700 11996
rect 19724 11994 19780 11996
rect 19484 11942 19530 11994
rect 19530 11942 19540 11994
rect 19564 11942 19594 11994
rect 19594 11942 19606 11994
rect 19606 11942 19620 11994
rect 19644 11942 19658 11994
rect 19658 11942 19670 11994
rect 19670 11942 19700 11994
rect 19724 11942 19734 11994
rect 19734 11942 19780 11994
rect 19484 11940 19540 11942
rect 19564 11940 19620 11942
rect 19644 11940 19700 11942
rect 19724 11940 19780 11942
rect 19484 10906 19540 10908
rect 19564 10906 19620 10908
rect 19644 10906 19700 10908
rect 19724 10906 19780 10908
rect 19484 10854 19530 10906
rect 19530 10854 19540 10906
rect 19564 10854 19594 10906
rect 19594 10854 19606 10906
rect 19606 10854 19620 10906
rect 19644 10854 19658 10906
rect 19658 10854 19670 10906
rect 19670 10854 19700 10906
rect 19724 10854 19734 10906
rect 19734 10854 19780 10906
rect 19484 10852 19540 10854
rect 19564 10852 19620 10854
rect 19644 10852 19700 10854
rect 19724 10852 19780 10854
rect 19484 9818 19540 9820
rect 19564 9818 19620 9820
rect 19644 9818 19700 9820
rect 19724 9818 19780 9820
rect 19484 9766 19530 9818
rect 19530 9766 19540 9818
rect 19564 9766 19594 9818
rect 19594 9766 19606 9818
rect 19606 9766 19620 9818
rect 19644 9766 19658 9818
rect 19658 9766 19670 9818
rect 19670 9766 19700 9818
rect 19724 9766 19734 9818
rect 19734 9766 19780 9818
rect 19484 9764 19540 9766
rect 19564 9764 19620 9766
rect 19644 9764 19700 9766
rect 19724 9764 19780 9766
rect 19484 8730 19540 8732
rect 19564 8730 19620 8732
rect 19644 8730 19700 8732
rect 19724 8730 19780 8732
rect 19484 8678 19530 8730
rect 19530 8678 19540 8730
rect 19564 8678 19594 8730
rect 19594 8678 19606 8730
rect 19606 8678 19620 8730
rect 19644 8678 19658 8730
rect 19658 8678 19670 8730
rect 19670 8678 19700 8730
rect 19724 8678 19734 8730
rect 19734 8678 19780 8730
rect 19484 8676 19540 8678
rect 19564 8676 19620 8678
rect 19644 8676 19700 8678
rect 19724 8676 19780 8678
rect 19484 7642 19540 7644
rect 19564 7642 19620 7644
rect 19644 7642 19700 7644
rect 19724 7642 19780 7644
rect 19484 7590 19530 7642
rect 19530 7590 19540 7642
rect 19564 7590 19594 7642
rect 19594 7590 19606 7642
rect 19606 7590 19620 7642
rect 19644 7590 19658 7642
rect 19658 7590 19670 7642
rect 19670 7590 19700 7642
rect 19724 7590 19734 7642
rect 19734 7590 19780 7642
rect 19484 7588 19540 7590
rect 19564 7588 19620 7590
rect 19644 7588 19700 7590
rect 19724 7588 19780 7590
rect 19484 6554 19540 6556
rect 19564 6554 19620 6556
rect 19644 6554 19700 6556
rect 19724 6554 19780 6556
rect 19484 6502 19530 6554
rect 19530 6502 19540 6554
rect 19564 6502 19594 6554
rect 19594 6502 19606 6554
rect 19606 6502 19620 6554
rect 19644 6502 19658 6554
rect 19658 6502 19670 6554
rect 19670 6502 19700 6554
rect 19724 6502 19734 6554
rect 19734 6502 19780 6554
rect 19484 6500 19540 6502
rect 19564 6500 19620 6502
rect 19644 6500 19700 6502
rect 19724 6500 19780 6502
rect 19484 5466 19540 5468
rect 19564 5466 19620 5468
rect 19644 5466 19700 5468
rect 19724 5466 19780 5468
rect 19484 5414 19530 5466
rect 19530 5414 19540 5466
rect 19564 5414 19594 5466
rect 19594 5414 19606 5466
rect 19606 5414 19620 5466
rect 19644 5414 19658 5466
rect 19658 5414 19670 5466
rect 19670 5414 19700 5466
rect 19724 5414 19734 5466
rect 19734 5414 19780 5466
rect 19484 5412 19540 5414
rect 19564 5412 19620 5414
rect 19644 5412 19700 5414
rect 19724 5412 19780 5414
rect 19484 4378 19540 4380
rect 19564 4378 19620 4380
rect 19644 4378 19700 4380
rect 19724 4378 19780 4380
rect 19484 4326 19530 4378
rect 19530 4326 19540 4378
rect 19564 4326 19594 4378
rect 19594 4326 19606 4378
rect 19606 4326 19620 4378
rect 19644 4326 19658 4378
rect 19658 4326 19670 4378
rect 19670 4326 19700 4378
rect 19724 4326 19734 4378
rect 19734 4326 19780 4378
rect 19484 4324 19540 4326
rect 19564 4324 19620 4326
rect 19644 4324 19700 4326
rect 19724 4324 19780 4326
rect 20258 26560 20314 26616
rect 20166 26424 20222 26480
rect 20074 26016 20130 26072
rect 20074 25608 20130 25664
rect 20258 24792 20314 24848
rect 20074 22092 20130 22128
rect 20074 22072 20076 22092
rect 20076 22072 20128 22092
rect 20128 22072 20130 22092
rect 20534 31728 20590 31784
rect 20442 28056 20498 28112
rect 20442 24792 20498 24848
rect 21362 34040 21418 34096
rect 21362 33496 21418 33552
rect 21086 30232 21142 30288
rect 20994 29960 21050 30016
rect 20810 28736 20866 28792
rect 20718 28192 20774 28248
rect 20718 27920 20774 27976
rect 20994 28872 21050 28928
rect 20626 24248 20682 24304
rect 21362 30368 21418 30424
rect 21546 36352 21602 36408
rect 21546 35708 21548 35728
rect 21548 35708 21600 35728
rect 21600 35708 21602 35728
rect 21546 35672 21602 35708
rect 22006 37188 22062 37224
rect 22006 37168 22008 37188
rect 22008 37168 22060 37188
rect 22060 37168 22062 37188
rect 22282 37168 22338 37224
rect 21914 36896 21970 36952
rect 22374 36916 22430 36952
rect 22374 36896 22376 36916
rect 22376 36896 22428 36916
rect 22428 36896 22430 36916
rect 21914 36624 21970 36680
rect 21822 35944 21878 36000
rect 22282 35808 22338 35864
rect 21914 35264 21970 35320
rect 22834 36216 22890 36272
rect 22650 35672 22706 35728
rect 22282 34992 22338 35048
rect 22190 34584 22246 34640
rect 21546 29724 21548 29744
rect 21548 29724 21600 29744
rect 21600 29724 21602 29744
rect 21546 29688 21602 29724
rect 21546 29300 21602 29336
rect 21546 29280 21548 29300
rect 21548 29280 21600 29300
rect 21600 29280 21602 29300
rect 21086 25880 21142 25936
rect 21730 29552 21786 29608
rect 22098 32544 22154 32600
rect 22098 32272 22154 32328
rect 22466 33088 22522 33144
rect 22926 35028 22928 35048
rect 22928 35028 22980 35048
rect 22980 35028 22982 35048
rect 22926 34992 22982 35028
rect 22558 32816 22614 32872
rect 22190 29688 22246 29744
rect 22098 29416 22154 29472
rect 21914 29008 21970 29064
rect 22098 29008 22154 29064
rect 22098 28464 22154 28520
rect 22466 30660 22522 30696
rect 22466 30640 22468 30660
rect 22468 30640 22520 30660
rect 22520 30640 22522 30660
rect 21914 28056 21970 28112
rect 21730 27784 21786 27840
rect 21730 27512 21786 27568
rect 22282 27920 22338 27976
rect 22190 27784 22246 27840
rect 22006 27668 22062 27704
rect 22006 27648 22008 27668
rect 22008 27648 22060 27668
rect 22060 27648 22062 27668
rect 22558 27784 22614 27840
rect 20994 24520 21050 24576
rect 20810 24248 20866 24304
rect 20810 23160 20866 23216
rect 21086 23024 21142 23080
rect 20994 22636 21050 22672
rect 20994 22616 20996 22636
rect 20996 22616 21048 22636
rect 21048 22616 21050 22636
rect 21362 21936 21418 21992
rect 21638 26732 21640 26752
rect 21640 26732 21692 26752
rect 21692 26732 21694 26752
rect 21638 26696 21694 26732
rect 21638 24928 21694 24984
rect 21914 23704 21970 23760
rect 22466 25744 22522 25800
rect 22834 28464 22890 28520
rect 22190 24112 22246 24168
rect 21638 23296 21694 23352
rect 23110 35536 23166 35592
rect 23202 34312 23258 34368
rect 23386 36236 23442 36272
rect 23386 36216 23388 36236
rect 23388 36216 23440 36236
rect 23440 36216 23442 36236
rect 23846 38256 23902 38312
rect 23662 37068 23664 37088
rect 23664 37068 23716 37088
rect 23716 37068 23718 37088
rect 23662 37032 23718 37068
rect 23386 34176 23442 34232
rect 23662 34312 23718 34368
rect 24116 39738 24172 39740
rect 24196 39738 24252 39740
rect 24276 39738 24332 39740
rect 24356 39738 24412 39740
rect 24116 39686 24162 39738
rect 24162 39686 24172 39738
rect 24196 39686 24226 39738
rect 24226 39686 24238 39738
rect 24238 39686 24252 39738
rect 24276 39686 24290 39738
rect 24290 39686 24302 39738
rect 24302 39686 24332 39738
rect 24356 39686 24366 39738
rect 24366 39686 24412 39738
rect 24116 39684 24172 39686
rect 24196 39684 24252 39686
rect 24276 39684 24332 39686
rect 24356 39684 24412 39686
rect 24582 39380 24584 39400
rect 24584 39380 24636 39400
rect 24636 39380 24638 39400
rect 24582 39344 24638 39380
rect 24030 39208 24086 39264
rect 24490 39072 24546 39128
rect 24116 38650 24172 38652
rect 24196 38650 24252 38652
rect 24276 38650 24332 38652
rect 24356 38650 24412 38652
rect 24116 38598 24162 38650
rect 24162 38598 24172 38650
rect 24196 38598 24226 38650
rect 24226 38598 24238 38650
rect 24238 38598 24252 38650
rect 24276 38598 24290 38650
rect 24290 38598 24302 38650
rect 24302 38598 24332 38650
rect 24356 38598 24366 38650
rect 24366 38598 24412 38650
rect 24116 38596 24172 38598
rect 24196 38596 24252 38598
rect 24276 38596 24332 38598
rect 24356 38596 24412 38598
rect 24582 38392 24638 38448
rect 25870 38292 25872 38312
rect 25872 38292 25924 38312
rect 25924 38292 25926 38312
rect 24116 37562 24172 37564
rect 24196 37562 24252 37564
rect 24276 37562 24332 37564
rect 24356 37562 24412 37564
rect 24116 37510 24162 37562
rect 24162 37510 24172 37562
rect 24196 37510 24226 37562
rect 24226 37510 24238 37562
rect 24238 37510 24252 37562
rect 24276 37510 24290 37562
rect 24290 37510 24302 37562
rect 24302 37510 24332 37562
rect 24356 37510 24366 37562
rect 24366 37510 24412 37562
rect 24116 37508 24172 37510
rect 24196 37508 24252 37510
rect 24276 37508 24332 37510
rect 24356 37508 24412 37510
rect 24122 36916 24178 36952
rect 24122 36896 24124 36916
rect 24124 36896 24176 36916
rect 24176 36896 24178 36916
rect 24122 36624 24178 36680
rect 24116 36474 24172 36476
rect 24196 36474 24252 36476
rect 24276 36474 24332 36476
rect 24356 36474 24412 36476
rect 24116 36422 24162 36474
rect 24162 36422 24172 36474
rect 24196 36422 24226 36474
rect 24226 36422 24238 36474
rect 24238 36422 24252 36474
rect 24276 36422 24290 36474
rect 24290 36422 24302 36474
rect 24302 36422 24332 36474
rect 24356 36422 24366 36474
rect 24366 36422 24412 36474
rect 24116 36420 24172 36422
rect 24196 36420 24252 36422
rect 24276 36420 24332 36422
rect 24356 36420 24412 36422
rect 24116 35386 24172 35388
rect 24196 35386 24252 35388
rect 24276 35386 24332 35388
rect 24356 35386 24412 35388
rect 24116 35334 24162 35386
rect 24162 35334 24172 35386
rect 24196 35334 24226 35386
rect 24226 35334 24238 35386
rect 24238 35334 24252 35386
rect 24276 35334 24290 35386
rect 24290 35334 24302 35386
rect 24302 35334 24332 35386
rect 24356 35334 24366 35386
rect 24366 35334 24412 35386
rect 24116 35332 24172 35334
rect 24196 35332 24252 35334
rect 24276 35332 24332 35334
rect 24356 35332 24412 35334
rect 24398 35128 24454 35184
rect 24766 34856 24822 34912
rect 24674 34584 24730 34640
rect 24950 34584 25006 34640
rect 23478 33224 23534 33280
rect 23110 32816 23166 32872
rect 23938 32952 23994 33008
rect 23386 31764 23388 31784
rect 23388 31764 23440 31784
rect 23440 31764 23442 31784
rect 23386 31728 23442 31764
rect 24116 34298 24172 34300
rect 24196 34298 24252 34300
rect 24276 34298 24332 34300
rect 24356 34298 24412 34300
rect 24116 34246 24162 34298
rect 24162 34246 24172 34298
rect 24196 34246 24226 34298
rect 24226 34246 24238 34298
rect 24238 34246 24252 34298
rect 24276 34246 24290 34298
rect 24290 34246 24302 34298
rect 24302 34246 24332 34298
rect 24356 34246 24366 34298
rect 24366 34246 24412 34298
rect 24116 34244 24172 34246
rect 24196 34244 24252 34246
rect 24276 34244 24332 34246
rect 24356 34244 24412 34246
rect 24116 33210 24172 33212
rect 24196 33210 24252 33212
rect 24276 33210 24332 33212
rect 24356 33210 24412 33212
rect 24116 33158 24162 33210
rect 24162 33158 24172 33210
rect 24196 33158 24226 33210
rect 24226 33158 24238 33210
rect 24238 33158 24252 33210
rect 24276 33158 24290 33210
rect 24290 33158 24302 33210
rect 24302 33158 24332 33210
rect 24356 33158 24366 33210
rect 24366 33158 24412 33210
rect 24116 33156 24172 33158
rect 24196 33156 24252 33158
rect 24276 33156 24332 33158
rect 24356 33156 24412 33158
rect 24116 32122 24172 32124
rect 24196 32122 24252 32124
rect 24276 32122 24332 32124
rect 24356 32122 24412 32124
rect 24116 32070 24162 32122
rect 24162 32070 24172 32122
rect 24196 32070 24226 32122
rect 24226 32070 24238 32122
rect 24238 32070 24252 32122
rect 24276 32070 24290 32122
rect 24290 32070 24302 32122
rect 24302 32070 24332 32122
rect 24356 32070 24366 32122
rect 24366 32070 24412 32122
rect 24116 32068 24172 32070
rect 24196 32068 24252 32070
rect 24276 32068 24332 32070
rect 24356 32068 24412 32070
rect 23294 30776 23350 30832
rect 23294 29688 23350 29744
rect 23110 29008 23166 29064
rect 23386 28872 23442 28928
rect 23754 29824 23810 29880
rect 24116 31034 24172 31036
rect 24196 31034 24252 31036
rect 24276 31034 24332 31036
rect 24356 31034 24412 31036
rect 24116 30982 24162 31034
rect 24162 30982 24172 31034
rect 24196 30982 24226 31034
rect 24226 30982 24238 31034
rect 24238 30982 24252 31034
rect 24276 30982 24290 31034
rect 24290 30982 24302 31034
rect 24302 30982 24332 31034
rect 24356 30982 24366 31034
rect 24366 30982 24412 31034
rect 24116 30980 24172 30982
rect 24196 30980 24252 30982
rect 24276 30980 24332 30982
rect 24356 30980 24412 30982
rect 24116 29946 24172 29948
rect 24196 29946 24252 29948
rect 24276 29946 24332 29948
rect 24356 29946 24412 29948
rect 24116 29894 24162 29946
rect 24162 29894 24172 29946
rect 24196 29894 24226 29946
rect 24226 29894 24238 29946
rect 24238 29894 24252 29946
rect 24276 29894 24290 29946
rect 24290 29894 24302 29946
rect 24302 29894 24332 29946
rect 24356 29894 24366 29946
rect 24366 29894 24412 29946
rect 24116 29892 24172 29894
rect 24196 29892 24252 29894
rect 24276 29892 24332 29894
rect 24356 29892 24412 29894
rect 23754 29416 23810 29472
rect 23662 29280 23718 29336
rect 23478 28192 23534 28248
rect 23110 27240 23166 27296
rect 24030 29144 24086 29200
rect 24582 29280 24638 29336
rect 22926 25608 22982 25664
rect 22374 23568 22430 23624
rect 22650 23840 22706 23896
rect 22650 23432 22706 23488
rect 22558 23296 22614 23352
rect 22374 21120 22430 21176
rect 22190 20848 22246 20904
rect 21822 20440 21878 20496
rect 22006 16668 22008 16688
rect 22008 16668 22060 16688
rect 22060 16668 22062 16688
rect 22006 16632 22062 16668
rect 23018 24656 23074 24712
rect 22926 21528 22982 21584
rect 22742 20984 22798 21040
rect 22650 20304 22706 20360
rect 23570 26288 23626 26344
rect 23478 26016 23534 26072
rect 23478 23976 23534 24032
rect 23662 25336 23718 25392
rect 23662 24692 23664 24712
rect 23664 24692 23716 24712
rect 23716 24692 23718 24712
rect 23662 24656 23718 24692
rect 24116 28858 24172 28860
rect 24196 28858 24252 28860
rect 24276 28858 24332 28860
rect 24356 28858 24412 28860
rect 24116 28806 24162 28858
rect 24162 28806 24172 28858
rect 24196 28806 24226 28858
rect 24226 28806 24238 28858
rect 24238 28806 24252 28858
rect 24276 28806 24290 28858
rect 24290 28806 24302 28858
rect 24302 28806 24332 28858
rect 24356 28806 24366 28858
rect 24366 28806 24412 28858
rect 24116 28804 24172 28806
rect 24196 28804 24252 28806
rect 24276 28804 24332 28806
rect 24356 28804 24412 28806
rect 24116 27770 24172 27772
rect 24196 27770 24252 27772
rect 24276 27770 24332 27772
rect 24356 27770 24412 27772
rect 24116 27718 24162 27770
rect 24162 27718 24172 27770
rect 24196 27718 24226 27770
rect 24226 27718 24238 27770
rect 24238 27718 24252 27770
rect 24276 27718 24290 27770
rect 24290 27718 24302 27770
rect 24302 27718 24332 27770
rect 24356 27718 24366 27770
rect 24366 27718 24412 27770
rect 24116 27716 24172 27718
rect 24196 27716 24252 27718
rect 24276 27716 24332 27718
rect 24356 27716 24412 27718
rect 24490 27512 24546 27568
rect 25870 38256 25926 38292
rect 25318 37032 25374 37088
rect 25594 35536 25650 35592
rect 25594 34720 25650 34776
rect 25042 32544 25098 32600
rect 25134 31728 25190 31784
rect 25870 36252 25872 36272
rect 25872 36252 25924 36272
rect 25924 36252 25926 36272
rect 25870 36216 25926 36252
rect 25870 34720 25926 34776
rect 24950 29960 25006 30016
rect 25778 32816 25834 32872
rect 25134 29552 25190 29608
rect 24950 28056 25006 28112
rect 24766 26968 24822 27024
rect 24116 26682 24172 26684
rect 24196 26682 24252 26684
rect 24276 26682 24332 26684
rect 24356 26682 24412 26684
rect 24116 26630 24162 26682
rect 24162 26630 24172 26682
rect 24196 26630 24226 26682
rect 24226 26630 24238 26682
rect 24238 26630 24252 26682
rect 24276 26630 24290 26682
rect 24290 26630 24302 26682
rect 24302 26630 24332 26682
rect 24356 26630 24366 26682
rect 24366 26630 24412 26682
rect 24116 26628 24172 26630
rect 24196 26628 24252 26630
rect 24276 26628 24332 26630
rect 24356 26628 24412 26630
rect 24116 25594 24172 25596
rect 24196 25594 24252 25596
rect 24276 25594 24332 25596
rect 24356 25594 24412 25596
rect 24116 25542 24162 25594
rect 24162 25542 24172 25594
rect 24196 25542 24226 25594
rect 24226 25542 24238 25594
rect 24238 25542 24252 25594
rect 24276 25542 24290 25594
rect 24290 25542 24302 25594
rect 24302 25542 24332 25594
rect 24356 25542 24366 25594
rect 24366 25542 24412 25594
rect 24116 25540 24172 25542
rect 24196 25540 24252 25542
rect 24276 25540 24332 25542
rect 24356 25540 24412 25542
rect 23662 23024 23718 23080
rect 23754 22752 23810 22808
rect 24116 24506 24172 24508
rect 24196 24506 24252 24508
rect 24276 24506 24332 24508
rect 24356 24506 24412 24508
rect 24116 24454 24162 24506
rect 24162 24454 24172 24506
rect 24196 24454 24226 24506
rect 24226 24454 24238 24506
rect 24238 24454 24252 24506
rect 24276 24454 24290 24506
rect 24290 24454 24302 24506
rect 24302 24454 24332 24506
rect 24356 24454 24366 24506
rect 24366 24454 24412 24506
rect 24116 24452 24172 24454
rect 24196 24452 24252 24454
rect 24276 24452 24332 24454
rect 24356 24452 24412 24454
rect 24306 23976 24362 24032
rect 25594 29724 25596 29744
rect 25596 29724 25648 29744
rect 25648 29724 25650 29744
rect 25594 29688 25650 29724
rect 26146 38836 26148 38856
rect 26148 38836 26200 38856
rect 26200 38836 26202 38856
rect 26146 38800 26202 38836
rect 26238 38664 26294 38720
rect 26054 38120 26110 38176
rect 26606 39888 26662 39944
rect 26514 37324 26570 37360
rect 26514 37304 26516 37324
rect 26516 37304 26568 37324
rect 26568 37304 26570 37324
rect 26330 36760 26386 36816
rect 26974 35944 27030 36000
rect 26330 34176 26386 34232
rect 26146 34040 26202 34096
rect 26514 33924 26570 33960
rect 26514 33904 26516 33924
rect 26516 33904 26568 33924
rect 26568 33904 26570 33924
rect 26330 33360 26386 33416
rect 26146 32408 26202 32464
rect 26330 31884 26386 31920
rect 26330 31864 26332 31884
rect 26332 31864 26384 31884
rect 26384 31864 26386 31884
rect 26422 31320 26478 31376
rect 26054 30368 26110 30424
rect 26330 30368 26386 30424
rect 26974 32272 27030 32328
rect 28170 40840 28226 40896
rect 28262 39480 28318 39536
rect 28170 36760 28226 36816
rect 25962 30132 25964 30152
rect 25964 30132 26016 30152
rect 26016 30132 26018 30152
rect 25962 30096 26018 30132
rect 26606 29280 26662 29336
rect 25594 27240 25650 27296
rect 25410 26288 25466 26344
rect 24674 23860 24730 23896
rect 24674 23840 24676 23860
rect 24676 23840 24728 23860
rect 24728 23840 24730 23860
rect 24950 24148 24952 24168
rect 24952 24148 25004 24168
rect 25004 24148 25006 24168
rect 24950 24112 25006 24148
rect 24858 23976 24914 24032
rect 25226 24248 25282 24304
rect 24116 23418 24172 23420
rect 24196 23418 24252 23420
rect 24276 23418 24332 23420
rect 24356 23418 24412 23420
rect 24116 23366 24162 23418
rect 24162 23366 24172 23418
rect 24196 23366 24226 23418
rect 24226 23366 24238 23418
rect 24238 23366 24252 23418
rect 24276 23366 24290 23418
rect 24290 23366 24302 23418
rect 24302 23366 24332 23418
rect 24356 23366 24366 23418
rect 24366 23366 24412 23418
rect 24116 23364 24172 23366
rect 24196 23364 24252 23366
rect 24276 23364 24332 23366
rect 24356 23364 24412 23366
rect 23662 22636 23718 22672
rect 23662 22616 23664 22636
rect 23664 22616 23716 22636
rect 23716 22616 23718 22636
rect 23662 22072 23718 22128
rect 24116 22330 24172 22332
rect 24196 22330 24252 22332
rect 24276 22330 24332 22332
rect 24356 22330 24412 22332
rect 24116 22278 24162 22330
rect 24162 22278 24172 22330
rect 24196 22278 24226 22330
rect 24226 22278 24238 22330
rect 24238 22278 24252 22330
rect 24276 22278 24290 22330
rect 24290 22278 24302 22330
rect 24302 22278 24332 22330
rect 24356 22278 24366 22330
rect 24366 22278 24412 22330
rect 24116 22276 24172 22278
rect 24196 22276 24252 22278
rect 24276 22276 24332 22278
rect 24356 22276 24412 22278
rect 24674 23044 24730 23080
rect 24674 23024 24676 23044
rect 24676 23024 24728 23044
rect 24728 23024 24730 23044
rect 24950 22616 25006 22672
rect 26330 27648 26386 27704
rect 26054 27376 26110 27432
rect 26330 26832 26386 26888
rect 26422 25880 26478 25936
rect 26330 25236 26332 25256
rect 26332 25236 26384 25256
rect 26384 25236 26386 25256
rect 26330 25200 26386 25236
rect 25686 23160 25742 23216
rect 26146 24812 26202 24848
rect 26146 24792 26148 24812
rect 26148 24792 26200 24812
rect 26200 24792 26202 24812
rect 26330 23432 26386 23488
rect 24674 22500 24730 22536
rect 24674 22480 24676 22500
rect 24676 22480 24728 22500
rect 24728 22480 24730 22500
rect 24116 21242 24172 21244
rect 24196 21242 24252 21244
rect 24276 21242 24332 21244
rect 24356 21242 24412 21244
rect 24116 21190 24162 21242
rect 24162 21190 24172 21242
rect 24196 21190 24226 21242
rect 24226 21190 24238 21242
rect 24238 21190 24252 21242
rect 24276 21190 24290 21242
rect 24290 21190 24302 21242
rect 24302 21190 24332 21242
rect 24356 21190 24366 21242
rect 24366 21190 24412 21242
rect 24116 21188 24172 21190
rect 24196 21188 24252 21190
rect 24276 21188 24332 21190
rect 24356 21188 24412 21190
rect 24582 21120 24638 21176
rect 23202 16632 23258 16688
rect 24116 20154 24172 20156
rect 24196 20154 24252 20156
rect 24276 20154 24332 20156
rect 24356 20154 24412 20156
rect 24116 20102 24162 20154
rect 24162 20102 24172 20154
rect 24196 20102 24226 20154
rect 24226 20102 24238 20154
rect 24238 20102 24252 20154
rect 24276 20102 24290 20154
rect 24290 20102 24302 20154
rect 24302 20102 24332 20154
rect 24356 20102 24366 20154
rect 24366 20102 24412 20154
rect 24116 20100 24172 20102
rect 24196 20100 24252 20102
rect 24276 20100 24332 20102
rect 24356 20100 24412 20102
rect 24306 19896 24362 19952
rect 24116 19066 24172 19068
rect 24196 19066 24252 19068
rect 24276 19066 24332 19068
rect 24356 19066 24412 19068
rect 24116 19014 24162 19066
rect 24162 19014 24172 19066
rect 24196 19014 24226 19066
rect 24226 19014 24238 19066
rect 24238 19014 24252 19066
rect 24276 19014 24290 19066
rect 24290 19014 24302 19066
rect 24302 19014 24332 19066
rect 24356 19014 24366 19066
rect 24366 19014 24412 19066
rect 24116 19012 24172 19014
rect 24196 19012 24252 19014
rect 24276 19012 24332 19014
rect 24356 19012 24412 19014
rect 24858 21120 24914 21176
rect 24116 17978 24172 17980
rect 24196 17978 24252 17980
rect 24276 17978 24332 17980
rect 24356 17978 24412 17980
rect 24116 17926 24162 17978
rect 24162 17926 24172 17978
rect 24196 17926 24226 17978
rect 24226 17926 24238 17978
rect 24238 17926 24252 17978
rect 24276 17926 24290 17978
rect 24290 17926 24302 17978
rect 24302 17926 24332 17978
rect 24356 17926 24366 17978
rect 24366 17926 24412 17978
rect 24116 17924 24172 17926
rect 24196 17924 24252 17926
rect 24276 17924 24332 17926
rect 24356 17924 24412 17926
rect 24306 17740 24362 17776
rect 24306 17720 24308 17740
rect 24308 17720 24360 17740
rect 24360 17720 24362 17740
rect 24116 16890 24172 16892
rect 24196 16890 24252 16892
rect 24276 16890 24332 16892
rect 24356 16890 24412 16892
rect 24116 16838 24162 16890
rect 24162 16838 24172 16890
rect 24196 16838 24226 16890
rect 24226 16838 24238 16890
rect 24238 16838 24252 16890
rect 24276 16838 24290 16890
rect 24290 16838 24302 16890
rect 24302 16838 24332 16890
rect 24356 16838 24366 16890
rect 24366 16838 24412 16890
rect 24116 16836 24172 16838
rect 24196 16836 24252 16838
rect 24276 16836 24332 16838
rect 24356 16836 24412 16838
rect 24116 15802 24172 15804
rect 24196 15802 24252 15804
rect 24276 15802 24332 15804
rect 24356 15802 24412 15804
rect 24116 15750 24162 15802
rect 24162 15750 24172 15802
rect 24196 15750 24226 15802
rect 24226 15750 24238 15802
rect 24238 15750 24252 15802
rect 24276 15750 24290 15802
rect 24290 15750 24302 15802
rect 24302 15750 24332 15802
rect 24356 15750 24366 15802
rect 24366 15750 24412 15802
rect 24116 15748 24172 15750
rect 24196 15748 24252 15750
rect 24276 15748 24332 15750
rect 24356 15748 24412 15750
rect 25318 22616 25374 22672
rect 24116 14714 24172 14716
rect 24196 14714 24252 14716
rect 24276 14714 24332 14716
rect 24356 14714 24412 14716
rect 24116 14662 24162 14714
rect 24162 14662 24172 14714
rect 24196 14662 24226 14714
rect 24226 14662 24238 14714
rect 24238 14662 24252 14714
rect 24276 14662 24290 14714
rect 24290 14662 24302 14714
rect 24302 14662 24332 14714
rect 24356 14662 24366 14714
rect 24366 14662 24412 14714
rect 24116 14660 24172 14662
rect 24196 14660 24252 14662
rect 24276 14660 24332 14662
rect 24356 14660 24412 14662
rect 24116 13626 24172 13628
rect 24196 13626 24252 13628
rect 24276 13626 24332 13628
rect 24356 13626 24412 13628
rect 24116 13574 24162 13626
rect 24162 13574 24172 13626
rect 24196 13574 24226 13626
rect 24226 13574 24238 13626
rect 24238 13574 24252 13626
rect 24276 13574 24290 13626
rect 24290 13574 24302 13626
rect 24302 13574 24332 13626
rect 24356 13574 24366 13626
rect 24366 13574 24412 13626
rect 24116 13572 24172 13574
rect 24196 13572 24252 13574
rect 24276 13572 24332 13574
rect 24356 13572 24412 13574
rect 25226 18808 25282 18864
rect 25042 18128 25098 18184
rect 25226 18128 25282 18184
rect 25502 18828 25558 18864
rect 25502 18808 25504 18828
rect 25504 18808 25556 18828
rect 25556 18808 25558 18828
rect 24116 12538 24172 12540
rect 24196 12538 24252 12540
rect 24276 12538 24332 12540
rect 24356 12538 24412 12540
rect 24116 12486 24162 12538
rect 24162 12486 24172 12538
rect 24196 12486 24226 12538
rect 24226 12486 24238 12538
rect 24238 12486 24252 12538
rect 24276 12486 24290 12538
rect 24290 12486 24302 12538
rect 24302 12486 24332 12538
rect 24356 12486 24366 12538
rect 24366 12486 24412 12538
rect 24116 12484 24172 12486
rect 24196 12484 24252 12486
rect 24276 12484 24332 12486
rect 24356 12484 24412 12486
rect 26146 21800 26202 21856
rect 26514 24928 26570 24984
rect 27434 26424 27490 26480
rect 26974 22752 27030 22808
rect 26146 15680 26202 15736
rect 28170 35400 28226 35456
rect 28906 39480 28962 39536
rect 28170 33360 28226 33416
rect 28170 32680 28226 32736
rect 28170 29280 28226 29336
rect 28078 28328 28134 28384
rect 28170 27240 28226 27296
rect 28170 26560 28226 26616
rect 28170 25880 28226 25936
rect 28170 24520 28226 24576
rect 28170 22480 28226 22536
rect 28170 21120 28226 21176
rect 27894 19896 27950 19952
rect 28170 19796 28172 19816
rect 28172 19796 28224 19816
rect 28224 19796 28226 19816
rect 28170 19760 28226 19796
rect 28170 19080 28226 19136
rect 19484 3290 19540 3292
rect 19564 3290 19620 3292
rect 19644 3290 19700 3292
rect 19724 3290 19780 3292
rect 19484 3238 19530 3290
rect 19530 3238 19540 3290
rect 19564 3238 19594 3290
rect 19594 3238 19606 3290
rect 19606 3238 19620 3290
rect 19644 3238 19658 3290
rect 19658 3238 19670 3290
rect 19670 3238 19700 3290
rect 19724 3238 19734 3290
rect 19734 3238 19780 3290
rect 19484 3236 19540 3238
rect 19564 3236 19620 3238
rect 19644 3236 19700 3238
rect 19724 3236 19780 3238
rect 24116 11450 24172 11452
rect 24196 11450 24252 11452
rect 24276 11450 24332 11452
rect 24356 11450 24412 11452
rect 24116 11398 24162 11450
rect 24162 11398 24172 11450
rect 24196 11398 24226 11450
rect 24226 11398 24238 11450
rect 24238 11398 24252 11450
rect 24276 11398 24290 11450
rect 24290 11398 24302 11450
rect 24302 11398 24332 11450
rect 24356 11398 24366 11450
rect 24366 11398 24412 11450
rect 24116 11396 24172 11398
rect 24196 11396 24252 11398
rect 24276 11396 24332 11398
rect 24356 11396 24412 11398
rect 24116 10362 24172 10364
rect 24196 10362 24252 10364
rect 24276 10362 24332 10364
rect 24356 10362 24412 10364
rect 24116 10310 24162 10362
rect 24162 10310 24172 10362
rect 24196 10310 24226 10362
rect 24226 10310 24238 10362
rect 24238 10310 24252 10362
rect 24276 10310 24290 10362
rect 24290 10310 24302 10362
rect 24302 10310 24332 10362
rect 24356 10310 24366 10362
rect 24366 10310 24412 10362
rect 24116 10308 24172 10310
rect 24196 10308 24252 10310
rect 24276 10308 24332 10310
rect 24356 10308 24412 10310
rect 24116 9274 24172 9276
rect 24196 9274 24252 9276
rect 24276 9274 24332 9276
rect 24356 9274 24412 9276
rect 24116 9222 24162 9274
rect 24162 9222 24172 9274
rect 24196 9222 24226 9274
rect 24226 9222 24238 9274
rect 24238 9222 24252 9274
rect 24276 9222 24290 9274
rect 24290 9222 24302 9274
rect 24302 9222 24332 9274
rect 24356 9222 24366 9274
rect 24366 9222 24412 9274
rect 24116 9220 24172 9222
rect 24196 9220 24252 9222
rect 24276 9220 24332 9222
rect 24356 9220 24412 9222
rect 24116 8186 24172 8188
rect 24196 8186 24252 8188
rect 24276 8186 24332 8188
rect 24356 8186 24412 8188
rect 24116 8134 24162 8186
rect 24162 8134 24172 8186
rect 24196 8134 24226 8186
rect 24226 8134 24238 8186
rect 24238 8134 24252 8186
rect 24276 8134 24290 8186
rect 24290 8134 24302 8186
rect 24302 8134 24332 8186
rect 24356 8134 24366 8186
rect 24366 8134 24412 8186
rect 24116 8132 24172 8134
rect 24196 8132 24252 8134
rect 24276 8132 24332 8134
rect 24356 8132 24412 8134
rect 24116 7098 24172 7100
rect 24196 7098 24252 7100
rect 24276 7098 24332 7100
rect 24356 7098 24412 7100
rect 24116 7046 24162 7098
rect 24162 7046 24172 7098
rect 24196 7046 24226 7098
rect 24226 7046 24238 7098
rect 24238 7046 24252 7098
rect 24276 7046 24290 7098
rect 24290 7046 24302 7098
rect 24302 7046 24332 7098
rect 24356 7046 24366 7098
rect 24366 7046 24412 7098
rect 24116 7044 24172 7046
rect 24196 7044 24252 7046
rect 24276 7044 24332 7046
rect 24356 7044 24412 7046
rect 24116 6010 24172 6012
rect 24196 6010 24252 6012
rect 24276 6010 24332 6012
rect 24356 6010 24412 6012
rect 24116 5958 24162 6010
rect 24162 5958 24172 6010
rect 24196 5958 24226 6010
rect 24226 5958 24238 6010
rect 24238 5958 24252 6010
rect 24276 5958 24290 6010
rect 24290 5958 24302 6010
rect 24302 5958 24332 6010
rect 24356 5958 24366 6010
rect 24366 5958 24412 6010
rect 24116 5956 24172 5958
rect 24196 5956 24252 5958
rect 24276 5956 24332 5958
rect 24356 5956 24412 5958
rect 24116 4922 24172 4924
rect 24196 4922 24252 4924
rect 24276 4922 24332 4924
rect 24356 4922 24412 4924
rect 24116 4870 24162 4922
rect 24162 4870 24172 4922
rect 24196 4870 24226 4922
rect 24226 4870 24238 4922
rect 24238 4870 24252 4922
rect 24276 4870 24290 4922
rect 24290 4870 24302 4922
rect 24302 4870 24332 4922
rect 24356 4870 24366 4922
rect 24366 4870 24412 4922
rect 24116 4868 24172 4870
rect 24196 4868 24252 4870
rect 24276 4868 24332 4870
rect 24356 4868 24412 4870
rect 26054 4800 26110 4856
rect 19484 2202 19540 2204
rect 19564 2202 19620 2204
rect 19644 2202 19700 2204
rect 19724 2202 19780 2204
rect 19484 2150 19530 2202
rect 19530 2150 19540 2202
rect 19564 2150 19594 2202
rect 19594 2150 19606 2202
rect 19606 2150 19620 2202
rect 19644 2150 19658 2202
rect 19658 2150 19670 2202
rect 19670 2150 19700 2202
rect 19724 2150 19734 2202
rect 19734 2150 19780 2202
rect 19484 2148 19540 2150
rect 19564 2148 19620 2150
rect 19644 2148 19700 2150
rect 19724 2148 19780 2150
rect 24116 3834 24172 3836
rect 24196 3834 24252 3836
rect 24276 3834 24332 3836
rect 24356 3834 24412 3836
rect 24116 3782 24162 3834
rect 24162 3782 24172 3834
rect 24196 3782 24226 3834
rect 24226 3782 24238 3834
rect 24238 3782 24252 3834
rect 24276 3782 24290 3834
rect 24290 3782 24302 3834
rect 24302 3782 24332 3834
rect 24356 3782 24366 3834
rect 24366 3782 24412 3834
rect 24116 3780 24172 3782
rect 24196 3780 24252 3782
rect 24276 3780 24332 3782
rect 24356 3780 24412 3782
rect 26146 4120 26202 4176
rect 24116 2746 24172 2748
rect 24196 2746 24252 2748
rect 24276 2746 24332 2748
rect 24356 2746 24412 2748
rect 24116 2694 24162 2746
rect 24162 2694 24172 2746
rect 24196 2694 24226 2746
rect 24226 2694 24238 2746
rect 24238 2694 24252 2746
rect 24276 2694 24290 2746
rect 24290 2694 24302 2746
rect 24302 2694 24332 2746
rect 24356 2694 24366 2746
rect 24366 2694 24412 2746
rect 24116 2692 24172 2694
rect 24196 2692 24252 2694
rect 24276 2692 24332 2694
rect 24356 2692 24412 2694
rect 26146 2760 26202 2816
rect 28170 18400 28226 18456
rect 28722 32000 28778 32056
rect 28170 16360 28226 16416
rect 28170 15000 28226 15056
rect 28170 14340 28226 14376
rect 28170 14320 28172 14340
rect 28172 14320 28224 14340
rect 28224 14320 28226 14340
rect 27986 11600 28042 11656
rect 28170 10920 28226 10976
rect 28170 9560 28226 9616
rect 27434 3440 27490 3496
rect 28170 7520 28226 7576
rect 28722 25200 28778 25256
rect 28630 23704 28686 23760
rect 28170 6860 28226 6896
rect 28170 6840 28172 6860
rect 28172 6840 28224 6860
rect 28224 6840 28226 6860
rect 28170 6160 28226 6216
rect 26054 2080 26110 2136
rect 26146 40 26202 96
<< metal3 >>
rect 0 41428 800 41668
rect 0 40748 800 40988
rect 28165 40898 28231 40901
rect 29200 40898 30000 40988
rect 28165 40896 30000 40898
rect 28165 40840 28170 40896
rect 28226 40840 30000 40896
rect 28165 40838 30000 40840
rect 28165 40835 28231 40838
rect 29200 40748 30000 40838
rect 8661 40490 8727 40493
rect 15377 40490 15443 40493
rect 8661 40488 15443 40490
rect 8661 40432 8666 40488
rect 8722 40432 15382 40488
rect 15438 40432 15443 40488
rect 8661 40430 15443 40432
rect 8661 40427 8727 40430
rect 15377 40427 15443 40430
rect 11421 40354 11487 40357
rect 19057 40354 19123 40357
rect 11421 40352 19123 40354
rect 0 40218 800 40308
rect 11421 40296 11426 40352
rect 11482 40296 19062 40352
rect 19118 40296 19123 40352
rect 11421 40294 19123 40296
rect 11421 40291 11487 40294
rect 19057 40291 19123 40294
rect 2773 40218 2839 40221
rect 0 40216 2839 40218
rect 0 40160 2778 40216
rect 2834 40160 2839 40216
rect 0 40158 2839 40160
rect 0 40068 800 40158
rect 2773 40155 2839 40158
rect 12157 40218 12223 40221
rect 12525 40218 12591 40221
rect 12157 40216 12591 40218
rect 12157 40160 12162 40216
rect 12218 40160 12530 40216
rect 12586 40160 12591 40216
rect 12157 40158 12591 40160
rect 12157 40155 12223 40158
rect 12525 40155 12591 40158
rect 15285 40082 15351 40085
rect 12390 40080 15351 40082
rect 12390 40024 15290 40080
rect 15346 40024 15351 40080
rect 29200 40068 30000 40308
rect 12390 40022 15351 40024
rect 7097 39946 7163 39949
rect 12390 39946 12450 40022
rect 15285 40019 15351 40022
rect 7097 39944 12450 39946
rect 7097 39888 7102 39944
rect 7158 39888 12450 39944
rect 7097 39886 12450 39888
rect 12525 39946 12591 39949
rect 26601 39946 26667 39949
rect 12525 39944 26667 39946
rect 12525 39888 12530 39944
rect 12586 39888 26606 39944
rect 26662 39888 26667 39944
rect 12525 39886 26667 39888
rect 7097 39883 7163 39886
rect 12525 39883 12591 39886
rect 26601 39883 26667 39886
rect 7281 39810 7347 39813
rect 14641 39810 14707 39813
rect 7281 39808 14707 39810
rect 7281 39752 7286 39808
rect 7342 39752 14646 39808
rect 14702 39752 14707 39808
rect 7281 39750 14707 39752
rect 7281 39747 7347 39750
rect 14641 39747 14707 39750
rect 15285 39810 15351 39813
rect 21817 39810 21883 39813
rect 15285 39808 21883 39810
rect 15285 39752 15290 39808
rect 15346 39752 21822 39808
rect 21878 39752 21883 39808
rect 15285 39750 21883 39752
rect 15285 39747 15351 39750
rect 21817 39747 21883 39750
rect 5576 39744 5896 39745
rect 5576 39680 5584 39744
rect 5648 39680 5664 39744
rect 5728 39680 5744 39744
rect 5808 39680 5824 39744
rect 5888 39680 5896 39744
rect 5576 39679 5896 39680
rect 14840 39744 15160 39745
rect 14840 39680 14848 39744
rect 14912 39680 14928 39744
rect 14992 39680 15008 39744
rect 15072 39680 15088 39744
rect 15152 39680 15160 39744
rect 14840 39679 15160 39680
rect 24104 39744 24424 39745
rect 24104 39680 24112 39744
rect 24176 39680 24192 39744
rect 24256 39680 24272 39744
rect 24336 39680 24352 39744
rect 24416 39680 24424 39744
rect 24104 39679 24424 39680
rect 0 39538 800 39628
rect 7598 39612 7604 39676
rect 7668 39674 7674 39676
rect 12157 39674 12223 39677
rect 7668 39672 12223 39674
rect 7668 39616 12162 39672
rect 12218 39616 12223 39672
rect 7668 39614 12223 39616
rect 7668 39612 7674 39614
rect 12157 39611 12223 39614
rect 12341 39674 12407 39677
rect 14549 39674 14615 39677
rect 12341 39672 14615 39674
rect 12341 39616 12346 39672
rect 12402 39616 14554 39672
rect 14610 39616 14615 39672
rect 12341 39614 14615 39616
rect 12341 39611 12407 39614
rect 14549 39611 14615 39614
rect 17033 39674 17099 39677
rect 20069 39674 20135 39677
rect 17033 39672 20135 39674
rect 17033 39616 17038 39672
rect 17094 39616 20074 39672
rect 20130 39616 20135 39672
rect 17033 39614 20135 39616
rect 17033 39611 17099 39614
rect 20069 39611 20135 39614
rect 1761 39538 1827 39541
rect 28257 39538 28323 39541
rect 0 39478 1594 39538
rect 0 39388 800 39478
rect 1534 39402 1594 39478
rect 1761 39536 28323 39538
rect 1761 39480 1766 39536
rect 1822 39480 28262 39536
rect 28318 39480 28323 39536
rect 1761 39478 28323 39480
rect 1761 39475 1827 39478
rect 28257 39475 28323 39478
rect 28901 39538 28967 39541
rect 29200 39538 30000 39628
rect 28901 39536 30000 39538
rect 28901 39480 28906 39536
rect 28962 39480 30000 39536
rect 28901 39478 30000 39480
rect 28901 39475 28967 39478
rect 2865 39402 2931 39405
rect 1534 39400 2931 39402
rect 1534 39344 2870 39400
rect 2926 39344 2931 39400
rect 1534 39342 2931 39344
rect 2865 39339 2931 39342
rect 7833 39402 7899 39405
rect 17033 39402 17099 39405
rect 20069 39402 20135 39405
rect 24577 39402 24643 39405
rect 7833 39400 17099 39402
rect 7833 39344 7838 39400
rect 7894 39344 17038 39400
rect 17094 39344 17099 39400
rect 7833 39342 17099 39344
rect 7833 39339 7899 39342
rect 17033 39339 17099 39342
rect 17174 39342 19994 39402
rect 11462 39204 11468 39268
rect 11532 39266 11538 39268
rect 17174 39266 17234 39342
rect 11532 39206 17234 39266
rect 17309 39266 17375 39269
rect 18413 39266 18479 39269
rect 17309 39264 18479 39266
rect 17309 39208 17314 39264
rect 17370 39208 18418 39264
rect 18474 39208 18479 39264
rect 17309 39206 18479 39208
rect 19934 39266 19994 39342
rect 20069 39400 24643 39402
rect 20069 39344 20074 39400
rect 20130 39344 24582 39400
rect 24638 39344 24643 39400
rect 29200 39388 30000 39478
rect 20069 39342 24643 39344
rect 20069 39339 20135 39342
rect 24577 39339 24643 39342
rect 24025 39266 24091 39269
rect 19934 39264 24091 39266
rect 19934 39208 24030 39264
rect 24086 39208 24091 39264
rect 19934 39206 24091 39208
rect 11532 39204 11538 39206
rect 17309 39203 17375 39206
rect 18413 39203 18479 39206
rect 24025 39203 24091 39206
rect 10208 39200 10528 39201
rect 10208 39136 10216 39200
rect 10280 39136 10296 39200
rect 10360 39136 10376 39200
rect 10440 39136 10456 39200
rect 10520 39136 10528 39200
rect 10208 39135 10528 39136
rect 19472 39200 19792 39201
rect 19472 39136 19480 39200
rect 19544 39136 19560 39200
rect 19624 39136 19640 39200
rect 19704 39136 19720 39200
rect 19784 39136 19792 39200
rect 19472 39135 19792 39136
rect 10869 39130 10935 39133
rect 14365 39130 14431 39133
rect 10869 39128 14431 39130
rect 10869 39072 10874 39128
rect 10930 39072 14370 39128
rect 14426 39072 14431 39128
rect 10869 39070 14431 39072
rect 10869 39067 10935 39070
rect 14365 39067 14431 39070
rect 14641 39130 14707 39133
rect 19333 39130 19399 39133
rect 24485 39130 24551 39133
rect 14641 39128 19399 39130
rect 14641 39072 14646 39128
rect 14702 39072 19338 39128
rect 19394 39072 19399 39128
rect 14641 39070 19399 39072
rect 14641 39067 14707 39070
rect 19333 39067 19399 39070
rect 19934 39128 24551 39130
rect 19934 39072 24490 39128
rect 24546 39072 24551 39128
rect 19934 39070 24551 39072
rect 8293 38994 8359 38997
rect 19934 38994 19994 39070
rect 24485 39067 24551 39070
rect 8293 38992 19994 38994
rect 0 38708 800 38948
rect 8293 38936 8298 38992
rect 8354 38936 19994 38992
rect 8293 38934 19994 38936
rect 8293 38931 8359 38934
rect 8017 38858 8083 38861
rect 26141 38858 26207 38861
rect 29200 38858 30000 38948
rect 8017 38856 24594 38858
rect 8017 38800 8022 38856
rect 8078 38800 24594 38856
rect 8017 38798 24594 38800
rect 8017 38795 8083 38798
rect 9990 38660 9996 38724
rect 10060 38722 10066 38724
rect 10685 38722 10751 38725
rect 14641 38722 14707 38725
rect 10060 38720 12220 38722
rect 10060 38664 10690 38720
rect 10746 38664 12220 38720
rect 10060 38662 12220 38664
rect 10060 38660 10066 38662
rect 10685 38659 10751 38662
rect 5576 38656 5896 38657
rect 5576 38592 5584 38656
rect 5648 38592 5664 38656
rect 5728 38592 5744 38656
rect 5808 38592 5824 38656
rect 5888 38592 5896 38656
rect 5576 38591 5896 38592
rect 9254 38524 9260 38588
rect 9324 38586 9330 38588
rect 12014 38586 12020 38588
rect 9324 38526 12020 38586
rect 9324 38524 9330 38526
rect 12014 38524 12020 38526
rect 12084 38524 12090 38588
rect 12160 38586 12220 38662
rect 12758 38720 14707 38722
rect 12758 38664 14646 38720
rect 14702 38664 14707 38720
rect 12758 38662 14707 38664
rect 12758 38586 12818 38662
rect 14641 38659 14707 38662
rect 15285 38722 15351 38725
rect 19977 38722 20043 38725
rect 15285 38720 20043 38722
rect 15285 38664 15290 38720
rect 15346 38664 19982 38720
rect 20038 38664 20043 38720
rect 15285 38662 20043 38664
rect 24534 38722 24594 38798
rect 26141 38856 30000 38858
rect 26141 38800 26146 38856
rect 26202 38800 30000 38856
rect 26141 38798 30000 38800
rect 26141 38795 26207 38798
rect 26233 38722 26299 38725
rect 24534 38720 26299 38722
rect 24534 38664 26238 38720
rect 26294 38664 26299 38720
rect 29200 38708 30000 38798
rect 24534 38662 26299 38664
rect 15285 38659 15351 38662
rect 19977 38659 20043 38662
rect 26233 38659 26299 38662
rect 14840 38656 15160 38657
rect 14840 38592 14848 38656
rect 14912 38592 14928 38656
rect 14992 38592 15008 38656
rect 15072 38592 15088 38656
rect 15152 38592 15160 38656
rect 14840 38591 15160 38592
rect 24104 38656 24424 38657
rect 24104 38592 24112 38656
rect 24176 38592 24192 38656
rect 24256 38592 24272 38656
rect 24336 38592 24352 38656
rect 24416 38592 24424 38656
rect 24104 38591 24424 38592
rect 12160 38526 12818 38586
rect 12985 38586 13051 38589
rect 14181 38586 14247 38589
rect 12985 38584 14247 38586
rect 12985 38528 12990 38584
rect 13046 38528 14186 38584
rect 14242 38528 14247 38584
rect 12985 38526 14247 38528
rect 12985 38523 13051 38526
rect 14181 38523 14247 38526
rect 15285 38586 15351 38589
rect 21173 38586 21239 38589
rect 15285 38584 21239 38586
rect 15285 38528 15290 38584
rect 15346 38528 21178 38584
rect 21234 38528 21239 38584
rect 15285 38526 21239 38528
rect 15285 38523 15351 38526
rect 21173 38523 21239 38526
rect 7741 38450 7807 38453
rect 24577 38450 24643 38453
rect 7741 38448 24643 38450
rect 7741 38392 7746 38448
rect 7802 38392 24582 38448
rect 24638 38392 24643 38448
rect 7741 38390 24643 38392
rect 7741 38387 7807 38390
rect 24577 38387 24643 38390
rect 7373 38314 7439 38317
rect 9489 38314 9555 38317
rect 7373 38312 9555 38314
rect 0 38178 800 38268
rect 7373 38256 7378 38312
rect 7434 38256 9494 38312
rect 9550 38256 9555 38312
rect 7373 38254 9555 38256
rect 7373 38251 7439 38254
rect 9489 38251 9555 38254
rect 9673 38314 9739 38317
rect 19926 38314 19932 38316
rect 9673 38312 19932 38314
rect 9673 38256 9678 38312
rect 9734 38256 19932 38312
rect 9673 38254 19932 38256
rect 9673 38251 9739 38254
rect 19926 38252 19932 38254
rect 19996 38252 20002 38316
rect 23841 38314 23907 38317
rect 25865 38314 25931 38317
rect 23841 38312 25931 38314
rect 23841 38256 23846 38312
rect 23902 38256 25870 38312
rect 25926 38256 25931 38312
rect 23841 38254 25931 38256
rect 23841 38251 23907 38254
rect 25865 38251 25931 38254
rect 2773 38178 2839 38181
rect 0 38176 2839 38178
rect 0 38120 2778 38176
rect 2834 38120 2839 38176
rect 0 38118 2839 38120
rect 0 38028 800 38118
rect 2773 38115 2839 38118
rect 10777 38178 10843 38181
rect 19057 38178 19123 38181
rect 10777 38176 19123 38178
rect 10777 38120 10782 38176
rect 10838 38120 19062 38176
rect 19118 38120 19123 38176
rect 10777 38118 19123 38120
rect 10777 38115 10843 38118
rect 19057 38115 19123 38118
rect 26049 38178 26115 38181
rect 29200 38178 30000 38268
rect 26049 38176 30000 38178
rect 26049 38120 26054 38176
rect 26110 38120 30000 38176
rect 26049 38118 30000 38120
rect 26049 38115 26115 38118
rect 10208 38112 10528 38113
rect 10208 38048 10216 38112
rect 10280 38048 10296 38112
rect 10360 38048 10376 38112
rect 10440 38048 10456 38112
rect 10520 38048 10528 38112
rect 10208 38047 10528 38048
rect 19472 38112 19792 38113
rect 19472 38048 19480 38112
rect 19544 38048 19560 38112
rect 19624 38048 19640 38112
rect 19704 38048 19720 38112
rect 19784 38048 19792 38112
rect 19472 38047 19792 38048
rect 8201 38042 8267 38045
rect 9949 38042 10015 38045
rect 8201 38040 10015 38042
rect 8201 37984 8206 38040
rect 8262 37984 9954 38040
rect 10010 37984 10015 38040
rect 8201 37982 10015 37984
rect 8201 37979 8267 37982
rect 9949 37979 10015 37982
rect 10726 37980 10732 38044
rect 10796 38042 10802 38044
rect 10869 38042 10935 38045
rect 11973 38042 12039 38045
rect 10796 38040 12039 38042
rect 10796 37984 10874 38040
rect 10930 37984 11978 38040
rect 12034 37984 12039 38040
rect 10796 37982 12039 37984
rect 10796 37980 10802 37982
rect 10869 37979 10935 37982
rect 11973 37979 12039 37982
rect 12525 38042 12591 38045
rect 12985 38042 13051 38045
rect 17125 38042 17191 38045
rect 12525 38040 13051 38042
rect 12525 37984 12530 38040
rect 12586 37984 12990 38040
rect 13046 37984 13051 38040
rect 12525 37982 13051 37984
rect 12525 37979 12591 37982
rect 12985 37979 13051 37982
rect 13172 38040 17191 38042
rect 13172 37984 17130 38040
rect 17186 37984 17191 38040
rect 29200 38028 30000 38118
rect 13172 37982 17191 37984
rect 9213 37906 9279 37909
rect 13172 37906 13232 37982
rect 17125 37979 17191 37982
rect 20897 37906 20963 37909
rect 9213 37904 13232 37906
rect 9213 37848 9218 37904
rect 9274 37848 13232 37904
rect 9213 37846 13232 37848
rect 13310 37904 20963 37906
rect 13310 37848 20902 37904
rect 20958 37848 20963 37904
rect 13310 37846 20963 37848
rect 9213 37843 9279 37846
rect 8661 37770 8727 37773
rect 12065 37770 12131 37773
rect 8661 37768 12131 37770
rect 8661 37712 8666 37768
rect 8722 37712 12070 37768
rect 12126 37712 12131 37768
rect 8661 37710 12131 37712
rect 8661 37707 8727 37710
rect 12065 37707 12131 37710
rect 12198 37708 12204 37772
rect 12268 37770 12274 37772
rect 13310 37770 13370 37846
rect 20897 37843 20963 37846
rect 15193 37770 15259 37773
rect 12268 37710 13370 37770
rect 14460 37768 15259 37770
rect 14460 37712 15198 37768
rect 15254 37712 15259 37768
rect 14460 37710 15259 37712
rect 12268 37708 12274 37710
rect 9489 37634 9555 37637
rect 14460 37634 14520 37710
rect 15193 37707 15259 37710
rect 15377 37770 15443 37773
rect 19609 37770 19675 37773
rect 15377 37768 19675 37770
rect 15377 37712 15382 37768
rect 15438 37712 19614 37768
rect 19670 37712 19675 37768
rect 15377 37710 19675 37712
rect 15377 37707 15443 37710
rect 19609 37707 19675 37710
rect 9489 37632 14520 37634
rect 0 37498 800 37588
rect 9489 37576 9494 37632
rect 9550 37576 14520 37632
rect 9489 37574 14520 37576
rect 9489 37571 9555 37574
rect 5576 37568 5896 37569
rect 5576 37504 5584 37568
rect 5648 37504 5664 37568
rect 5728 37504 5744 37568
rect 5808 37504 5824 37568
rect 5888 37504 5896 37568
rect 5576 37503 5896 37504
rect 14840 37568 15160 37569
rect 14840 37504 14848 37568
rect 14912 37504 14928 37568
rect 14992 37504 15008 37568
rect 15072 37504 15088 37568
rect 15152 37504 15160 37568
rect 14840 37503 15160 37504
rect 24104 37568 24424 37569
rect 24104 37504 24112 37568
rect 24176 37504 24192 37568
rect 24256 37504 24272 37568
rect 24336 37504 24352 37568
rect 24416 37504 24424 37568
rect 24104 37503 24424 37504
rect 1853 37498 1919 37501
rect 0 37496 1919 37498
rect 0 37440 1858 37496
rect 1914 37440 1919 37496
rect 0 37438 1919 37440
rect 0 37348 800 37438
rect 1853 37435 1919 37438
rect 8017 37498 8083 37501
rect 13721 37498 13787 37501
rect 8017 37496 13787 37498
rect 8017 37440 8022 37496
rect 8078 37440 13726 37496
rect 13782 37440 13787 37496
rect 8017 37438 13787 37440
rect 8017 37435 8083 37438
rect 13721 37435 13787 37438
rect 15469 37498 15535 37501
rect 19057 37498 19123 37501
rect 15469 37496 19123 37498
rect 15469 37440 15474 37496
rect 15530 37440 19062 37496
rect 19118 37440 19123 37496
rect 15469 37438 19123 37440
rect 15469 37435 15535 37438
rect 19057 37435 19123 37438
rect 8753 37362 8819 37365
rect 16113 37362 16179 37365
rect 8753 37360 16179 37362
rect 8753 37304 8758 37360
rect 8814 37304 16118 37360
rect 16174 37304 16179 37360
rect 8753 37302 16179 37304
rect 8753 37299 8819 37302
rect 16113 37299 16179 37302
rect 17861 37362 17927 37365
rect 19190 37362 19196 37364
rect 17861 37360 19196 37362
rect 17861 37304 17866 37360
rect 17922 37304 19196 37360
rect 17861 37302 19196 37304
rect 17861 37299 17927 37302
rect 19190 37300 19196 37302
rect 19260 37300 19266 37364
rect 20529 37362 20595 37365
rect 26509 37362 26575 37365
rect 20529 37360 26575 37362
rect 20529 37304 20534 37360
rect 20590 37304 26514 37360
rect 26570 37304 26575 37360
rect 29200 37348 30000 37588
rect 20529 37302 26575 37304
rect 20529 37299 20595 37302
rect 26509 37299 26575 37302
rect 8201 37226 8267 37229
rect 19609 37226 19675 37229
rect 20110 37226 20116 37228
rect 8201 37224 17234 37226
rect 8201 37168 8206 37224
rect 8262 37168 17234 37224
rect 8201 37166 17234 37168
rect 8201 37163 8267 37166
rect 9622 37028 9628 37092
rect 9692 37090 9698 37092
rect 9857 37090 9923 37093
rect 9692 37088 9923 37090
rect 9692 37032 9862 37088
rect 9918 37032 9923 37088
rect 9692 37030 9923 37032
rect 9692 37028 9698 37030
rect 9857 37027 9923 37030
rect 10685 37090 10751 37093
rect 11513 37090 11579 37093
rect 10685 37088 11579 37090
rect 10685 37032 10690 37088
rect 10746 37032 11518 37088
rect 11574 37032 11579 37088
rect 10685 37030 11579 37032
rect 10685 37027 10751 37030
rect 11513 37027 11579 37030
rect 11646 37028 11652 37092
rect 11716 37090 11722 37092
rect 12249 37090 12315 37093
rect 11716 37088 12315 37090
rect 11716 37032 12254 37088
rect 12310 37032 12315 37088
rect 11716 37030 12315 37032
rect 11716 37028 11722 37030
rect 12249 37027 12315 37030
rect 12433 37090 12499 37093
rect 12893 37090 12959 37093
rect 12433 37088 12959 37090
rect 12433 37032 12438 37088
rect 12494 37032 12898 37088
rect 12954 37032 12959 37088
rect 12433 37030 12959 37032
rect 12433 37027 12499 37030
rect 12893 37027 12959 37030
rect 13077 37090 13143 37093
rect 13537 37090 13603 37093
rect 13077 37088 13603 37090
rect 13077 37032 13082 37088
rect 13138 37032 13542 37088
rect 13598 37032 13603 37088
rect 13077 37030 13603 37032
rect 13077 37027 13143 37030
rect 13537 37027 13603 37030
rect 14038 37028 14044 37092
rect 14108 37090 14114 37092
rect 16941 37090 17007 37093
rect 14108 37088 17007 37090
rect 14108 37032 16946 37088
rect 17002 37032 17007 37088
rect 14108 37030 17007 37032
rect 14108 37028 14114 37030
rect 16941 37027 17007 37030
rect 10208 37024 10528 37025
rect 10208 36960 10216 37024
rect 10280 36960 10296 37024
rect 10360 36960 10376 37024
rect 10440 36960 10456 37024
rect 10520 36960 10528 37024
rect 10208 36959 10528 36960
rect 9581 36954 9647 36957
rect 10041 36954 10107 36957
rect 9581 36952 10107 36954
rect 0 36668 800 36908
rect 9581 36896 9586 36952
rect 9642 36896 10046 36952
rect 10102 36896 10107 36952
rect 9581 36894 10107 36896
rect 9581 36891 9647 36894
rect 10041 36891 10107 36894
rect 10596 36894 17096 36954
rect 9581 36818 9647 36821
rect 10596 36818 10656 36894
rect 9581 36816 10656 36818
rect 9581 36760 9586 36816
rect 9642 36760 10656 36816
rect 9581 36758 10656 36760
rect 9581 36755 9647 36758
rect 10910 36756 10916 36820
rect 10980 36818 10986 36820
rect 10980 36758 16498 36818
rect 10980 36756 10986 36758
rect 7281 36682 7347 36685
rect 12065 36682 12131 36685
rect 7281 36680 12131 36682
rect 7281 36624 7286 36680
rect 7342 36624 12070 36680
rect 12126 36624 12131 36680
rect 7281 36622 12131 36624
rect 7281 36619 7347 36622
rect 12065 36619 12131 36622
rect 12198 36620 12204 36684
rect 12268 36682 12274 36684
rect 14365 36682 14431 36685
rect 16205 36682 16271 36685
rect 12268 36680 16271 36682
rect 12268 36624 14370 36680
rect 14426 36624 16210 36680
rect 16266 36624 16271 36680
rect 12268 36622 16271 36624
rect 12268 36620 12274 36622
rect 14365 36619 14431 36622
rect 16205 36619 16271 36622
rect 8845 36546 8911 36549
rect 12065 36546 12131 36549
rect 12985 36546 13051 36549
rect 8845 36544 11898 36546
rect 8845 36488 8850 36544
rect 8906 36488 11898 36544
rect 8845 36486 11898 36488
rect 8845 36483 8911 36486
rect 5576 36480 5896 36481
rect 5576 36416 5584 36480
rect 5648 36416 5664 36480
rect 5728 36416 5744 36480
rect 5808 36416 5824 36480
rect 5888 36416 5896 36480
rect 5576 36415 5896 36416
rect 6269 36410 6335 36413
rect 11646 36410 11652 36412
rect 6269 36408 11652 36410
rect 6269 36352 6274 36408
rect 6330 36352 11652 36408
rect 6269 36350 11652 36352
rect 6269 36347 6335 36350
rect 11646 36348 11652 36350
rect 11716 36348 11722 36412
rect 11838 36410 11898 36486
rect 12065 36544 13051 36546
rect 12065 36488 12070 36544
rect 12126 36488 12990 36544
rect 13046 36488 13051 36544
rect 12065 36486 13051 36488
rect 12065 36483 12131 36486
rect 12985 36483 13051 36486
rect 13537 36546 13603 36549
rect 14457 36546 14523 36549
rect 13537 36544 14523 36546
rect 13537 36488 13542 36544
rect 13598 36488 14462 36544
rect 14518 36488 14523 36544
rect 13537 36486 14523 36488
rect 16438 36546 16498 36758
rect 17036 36682 17096 36894
rect 17174 36818 17234 37166
rect 19609 37224 20116 37226
rect 19609 37168 19614 37224
rect 19670 37168 20116 37224
rect 19609 37166 20116 37168
rect 19609 37163 19675 37166
rect 20110 37164 20116 37166
rect 20180 37164 20186 37228
rect 22001 37226 22067 37229
rect 22277 37226 22343 37229
rect 22001 37224 22343 37226
rect 22001 37168 22006 37224
rect 22062 37168 22282 37224
rect 22338 37168 22343 37224
rect 22001 37166 22343 37168
rect 22001 37163 22067 37166
rect 22277 37163 22343 37166
rect 23657 37090 23723 37093
rect 25313 37090 25379 37093
rect 23657 37088 25379 37090
rect 23657 37032 23662 37088
rect 23718 37032 25318 37088
rect 25374 37032 25379 37088
rect 23657 37030 25379 37032
rect 23657 37027 23723 37030
rect 25313 37027 25379 37030
rect 19472 37024 19792 37025
rect 19472 36960 19480 37024
rect 19544 36960 19560 37024
rect 19624 36960 19640 37024
rect 19704 36960 19720 37024
rect 19784 36960 19792 37024
rect 19472 36959 19792 36960
rect 18873 36954 18939 36957
rect 19333 36954 19399 36957
rect 18873 36952 19399 36954
rect 18873 36896 18878 36952
rect 18934 36896 19338 36952
rect 19394 36896 19399 36952
rect 18873 36894 19399 36896
rect 18873 36891 18939 36894
rect 19333 36891 19399 36894
rect 19926 36892 19932 36956
rect 19996 36954 20002 36956
rect 21909 36954 21975 36957
rect 19996 36952 21975 36954
rect 19996 36896 21914 36952
rect 21970 36896 21975 36952
rect 19996 36894 21975 36896
rect 19996 36892 20002 36894
rect 21909 36891 21975 36894
rect 22369 36954 22435 36957
rect 24117 36954 24183 36957
rect 22369 36952 24183 36954
rect 22369 36896 22374 36952
rect 22430 36896 24122 36952
rect 24178 36896 24183 36952
rect 22369 36894 24183 36896
rect 22369 36891 22435 36894
rect 24117 36891 24183 36894
rect 26325 36818 26391 36821
rect 17174 36816 26391 36818
rect 17174 36760 26330 36816
rect 26386 36760 26391 36816
rect 17174 36758 26391 36760
rect 26325 36755 26391 36758
rect 28165 36818 28231 36821
rect 29200 36818 30000 36908
rect 28165 36816 30000 36818
rect 28165 36760 28170 36816
rect 28226 36760 30000 36816
rect 28165 36758 30000 36760
rect 28165 36755 28231 36758
rect 18781 36682 18847 36685
rect 19057 36682 19123 36685
rect 17036 36680 19123 36682
rect 17036 36624 18786 36680
rect 18842 36624 19062 36680
rect 19118 36624 19123 36680
rect 17036 36622 19123 36624
rect 18781 36619 18847 36622
rect 19057 36619 19123 36622
rect 19241 36682 19307 36685
rect 20805 36682 20871 36685
rect 19241 36680 20871 36682
rect 19241 36624 19246 36680
rect 19302 36624 20810 36680
rect 20866 36624 20871 36680
rect 19241 36622 20871 36624
rect 19241 36619 19307 36622
rect 20805 36619 20871 36622
rect 21909 36682 21975 36685
rect 24117 36682 24183 36685
rect 21909 36680 24183 36682
rect 21909 36624 21914 36680
rect 21970 36624 24122 36680
rect 24178 36624 24183 36680
rect 29200 36668 30000 36758
rect 21909 36622 24183 36624
rect 21909 36619 21975 36622
rect 24117 36619 24183 36622
rect 20805 36546 20871 36549
rect 16438 36544 20871 36546
rect 16438 36488 20810 36544
rect 20866 36488 20871 36544
rect 16438 36486 20871 36488
rect 13537 36483 13603 36486
rect 14457 36483 14523 36486
rect 20805 36483 20871 36486
rect 14840 36480 15160 36481
rect 14840 36416 14848 36480
rect 14912 36416 14928 36480
rect 14992 36416 15008 36480
rect 15072 36416 15088 36480
rect 15152 36416 15160 36480
rect 14840 36415 15160 36416
rect 24104 36480 24424 36481
rect 24104 36416 24112 36480
rect 24176 36416 24192 36480
rect 24256 36416 24272 36480
rect 24336 36416 24352 36480
rect 24416 36416 24424 36480
rect 24104 36415 24424 36416
rect 12198 36410 12204 36412
rect 11838 36350 12204 36410
rect 12198 36348 12204 36350
rect 12268 36348 12274 36412
rect 12709 36410 12775 36413
rect 14641 36410 14707 36413
rect 12709 36408 14707 36410
rect 12709 36352 12714 36408
rect 12770 36352 14646 36408
rect 14702 36352 14707 36408
rect 12709 36350 14707 36352
rect 12709 36347 12775 36350
rect 14641 36347 14707 36350
rect 15377 36410 15443 36413
rect 17125 36410 17191 36413
rect 21541 36410 21607 36413
rect 15377 36408 17050 36410
rect 15377 36352 15382 36408
rect 15438 36352 17050 36408
rect 15377 36350 17050 36352
rect 15377 36347 15443 36350
rect 8937 36274 9003 36277
rect 9397 36274 9463 36277
rect 9765 36276 9831 36277
rect 9765 36274 9812 36276
rect 8937 36272 9463 36274
rect 0 36138 800 36228
rect 8937 36216 8942 36272
rect 8998 36216 9402 36272
rect 9458 36216 9463 36272
rect 8937 36214 9463 36216
rect 9720 36272 9812 36274
rect 9720 36216 9770 36272
rect 9720 36214 9812 36216
rect 8937 36211 9003 36214
rect 9397 36211 9463 36214
rect 9765 36212 9812 36214
rect 9876 36212 9882 36276
rect 10317 36274 10383 36277
rect 12014 36274 12020 36276
rect 10317 36272 12020 36274
rect 10317 36216 10322 36272
rect 10378 36216 12020 36272
rect 10317 36214 12020 36216
rect 9765 36211 9831 36212
rect 10317 36211 10383 36214
rect 12014 36212 12020 36214
rect 12084 36212 12090 36276
rect 13854 36274 13860 36276
rect 12252 36214 13860 36274
rect 12252 36141 12312 36214
rect 13854 36212 13860 36214
rect 13924 36212 13930 36276
rect 13997 36274 14063 36277
rect 15929 36274 15995 36277
rect 13997 36272 15995 36274
rect 13997 36216 14002 36272
rect 14058 36216 15934 36272
rect 15990 36216 15995 36272
rect 13997 36214 15995 36216
rect 16990 36274 17050 36350
rect 17125 36408 21282 36410
rect 17125 36352 17130 36408
rect 17186 36352 21282 36408
rect 17125 36350 21282 36352
rect 17125 36347 17191 36350
rect 17585 36274 17651 36277
rect 16990 36272 17651 36274
rect 16990 36216 17590 36272
rect 17646 36216 17651 36272
rect 16990 36214 17651 36216
rect 13997 36211 14063 36214
rect 15929 36211 15995 36214
rect 17585 36211 17651 36214
rect 17769 36274 17835 36277
rect 20897 36274 20963 36277
rect 17769 36272 20963 36274
rect 17769 36216 17774 36272
rect 17830 36216 20902 36272
rect 20958 36216 20963 36272
rect 17769 36214 20963 36216
rect 21222 36274 21282 36350
rect 21541 36408 23306 36410
rect 21541 36352 21546 36408
rect 21602 36352 23306 36408
rect 21541 36350 23306 36352
rect 21541 36347 21607 36350
rect 22829 36274 22895 36277
rect 21222 36272 22895 36274
rect 21222 36216 22834 36272
rect 22890 36216 22895 36272
rect 21222 36214 22895 36216
rect 17769 36211 17835 36214
rect 20897 36211 20963 36214
rect 22829 36211 22895 36214
rect 4061 36138 4127 36141
rect 0 36136 4127 36138
rect 0 36080 4066 36136
rect 4122 36080 4127 36136
rect 0 36078 4127 36080
rect 0 35988 800 36078
rect 4061 36075 4127 36078
rect 9305 36138 9371 36141
rect 11830 36138 11836 36140
rect 9305 36136 11836 36138
rect 9305 36080 9310 36136
rect 9366 36080 11836 36136
rect 9305 36078 11836 36080
rect 9305 36075 9371 36078
rect 11830 36076 11836 36078
rect 11900 36076 11906 36140
rect 12249 36136 12315 36141
rect 18638 36138 18644 36140
rect 12249 36080 12254 36136
rect 12310 36080 12315 36136
rect 12249 36075 12315 36080
rect 12758 36078 18644 36138
rect 9121 36002 9187 36005
rect 10041 36002 10107 36005
rect 9121 36000 10107 36002
rect 9121 35944 9126 36000
rect 9182 35944 10046 36000
rect 10102 35944 10107 36000
rect 9121 35942 10107 35944
rect 9121 35939 9187 35942
rect 10041 35939 10107 35942
rect 10593 36002 10659 36005
rect 11053 36002 11119 36005
rect 10593 36000 11119 36002
rect 10593 35944 10598 36000
rect 10654 35944 11058 36000
rect 11114 35944 11119 36000
rect 10593 35942 11119 35944
rect 10593 35939 10659 35942
rect 11053 35939 11119 35942
rect 11462 35940 11468 36004
rect 11532 36002 11538 36004
rect 11605 36002 11671 36005
rect 11532 36000 11671 36002
rect 11532 35944 11610 36000
rect 11666 35944 11671 36000
rect 11532 35942 11671 35944
rect 11532 35940 11538 35942
rect 11605 35939 11671 35942
rect 11881 36002 11947 36005
rect 12758 36002 12818 36078
rect 18638 36076 18644 36078
rect 18708 36076 18714 36140
rect 19149 36138 19215 36141
rect 23246 36138 23306 36350
rect 23381 36274 23447 36277
rect 25865 36274 25931 36277
rect 23381 36272 25931 36274
rect 23381 36216 23386 36272
rect 23442 36216 25870 36272
rect 25926 36216 25931 36272
rect 23381 36214 25931 36216
rect 23381 36211 23447 36214
rect 25865 36211 25931 36214
rect 29200 36138 30000 36228
rect 18784 36136 22018 36138
rect 18784 36080 19154 36136
rect 19210 36080 22018 36136
rect 18784 36078 22018 36080
rect 23246 36078 30000 36138
rect 11881 36000 12818 36002
rect 11881 35944 11886 36000
rect 11942 35944 12818 36000
rect 11881 35942 12818 35944
rect 12893 36002 12959 36005
rect 16941 36002 17007 36005
rect 12893 36000 17007 36002
rect 12893 35944 12898 36000
rect 12954 35944 16946 36000
rect 17002 35944 17007 36000
rect 12893 35942 17007 35944
rect 11881 35939 11947 35942
rect 12893 35939 12959 35942
rect 16941 35939 17007 35942
rect 17585 36002 17651 36005
rect 18229 36002 18295 36005
rect 17585 36000 18295 36002
rect 17585 35944 17590 36000
rect 17646 35944 18234 36000
rect 18290 35944 18295 36000
rect 17585 35942 18295 35944
rect 17585 35939 17651 35942
rect 18229 35939 18295 35942
rect 18413 36002 18479 36005
rect 18784 36002 18844 36078
rect 19149 36075 19215 36078
rect 18413 36000 18844 36002
rect 18413 35944 18418 36000
rect 18474 35944 18844 36000
rect 18413 35942 18844 35944
rect 18413 35939 18479 35942
rect 19190 35940 19196 36004
rect 19260 36002 19266 36004
rect 19333 36002 19399 36005
rect 19260 36000 19399 36002
rect 19260 35944 19338 36000
rect 19394 35944 19399 36000
rect 19260 35942 19399 35944
rect 19260 35940 19266 35942
rect 19333 35939 19399 35942
rect 19885 36002 19951 36005
rect 20161 36002 20227 36005
rect 19885 36000 20227 36002
rect 19885 35944 19890 36000
rect 19946 35944 20166 36000
rect 20222 35944 20227 36000
rect 19885 35942 20227 35944
rect 19885 35939 19951 35942
rect 20161 35939 20227 35942
rect 21265 36002 21331 36005
rect 21817 36002 21883 36005
rect 21265 36000 21883 36002
rect 21265 35944 21270 36000
rect 21326 35944 21822 36000
rect 21878 35944 21883 36000
rect 21265 35942 21883 35944
rect 21958 36002 22018 36078
rect 26969 36002 27035 36005
rect 21958 36000 27035 36002
rect 21958 35944 26974 36000
rect 27030 35944 27035 36000
rect 29200 35988 30000 36078
rect 21958 35942 27035 35944
rect 21265 35939 21331 35942
rect 21817 35939 21883 35942
rect 26969 35939 27035 35942
rect 10208 35936 10528 35937
rect 10208 35872 10216 35936
rect 10280 35872 10296 35936
rect 10360 35872 10376 35936
rect 10440 35872 10456 35936
rect 10520 35872 10528 35936
rect 10208 35871 10528 35872
rect 19472 35936 19792 35937
rect 19472 35872 19480 35936
rect 19544 35872 19560 35936
rect 19624 35872 19640 35936
rect 19704 35872 19720 35936
rect 19784 35872 19792 35936
rect 19472 35871 19792 35872
rect 9029 35866 9095 35869
rect 9857 35866 9923 35869
rect 9029 35864 9923 35866
rect 9029 35808 9034 35864
rect 9090 35808 9862 35864
rect 9918 35808 9923 35864
rect 9029 35806 9923 35808
rect 9029 35803 9095 35806
rect 9857 35803 9923 35806
rect 10869 35866 10935 35869
rect 12157 35866 12223 35869
rect 10869 35864 12223 35866
rect 10869 35808 10874 35864
rect 10930 35808 12162 35864
rect 12218 35808 12223 35864
rect 10869 35806 12223 35808
rect 10869 35803 10935 35806
rect 12157 35803 12223 35806
rect 12382 35804 12388 35868
rect 12452 35866 12458 35868
rect 19333 35866 19399 35869
rect 12452 35864 19399 35866
rect 12452 35808 19338 35864
rect 19394 35808 19399 35864
rect 12452 35806 19399 35808
rect 12452 35804 12458 35806
rect 19333 35803 19399 35806
rect 20345 35866 20411 35869
rect 22277 35866 22343 35869
rect 20345 35864 22343 35866
rect 20345 35808 20350 35864
rect 20406 35808 22282 35864
rect 22338 35808 22343 35864
rect 20345 35806 22343 35808
rect 20345 35803 20411 35806
rect 22277 35803 22343 35806
rect 7557 35732 7623 35733
rect 7557 35730 7604 35732
rect 7512 35728 7604 35730
rect 7512 35672 7562 35728
rect 7512 35670 7604 35672
rect 7557 35668 7604 35670
rect 7668 35668 7674 35732
rect 8201 35730 8267 35733
rect 17033 35730 17099 35733
rect 20805 35730 20871 35733
rect 20989 35732 21055 35733
rect 20989 35730 21036 35732
rect 8201 35728 17099 35730
rect 8201 35672 8206 35728
rect 8262 35672 17038 35728
rect 17094 35672 17099 35728
rect 8201 35670 17099 35672
rect 7557 35667 7623 35668
rect 8201 35667 8267 35670
rect 17033 35667 17099 35670
rect 17174 35728 20871 35730
rect 17174 35672 20810 35728
rect 20866 35672 20871 35728
rect 17174 35670 20871 35672
rect 20944 35728 21036 35730
rect 20944 35672 20994 35728
rect 20944 35670 21036 35672
rect 9489 35594 9555 35597
rect 13077 35594 13143 35597
rect 9489 35592 13143 35594
rect 0 35308 800 35548
rect 9489 35536 9494 35592
rect 9550 35536 13082 35592
rect 13138 35536 13143 35592
rect 9489 35534 13143 35536
rect 9489 35531 9555 35534
rect 13077 35531 13143 35534
rect 13261 35594 13327 35597
rect 14549 35594 14615 35597
rect 13261 35592 14615 35594
rect 13261 35536 13266 35592
rect 13322 35536 14554 35592
rect 14610 35536 14615 35592
rect 13261 35534 14615 35536
rect 13261 35531 13327 35534
rect 14549 35531 14615 35534
rect 14733 35594 14799 35597
rect 17174 35594 17234 35670
rect 20805 35667 20871 35670
rect 20989 35668 21036 35670
rect 21100 35668 21106 35732
rect 21541 35730 21607 35733
rect 22645 35730 22711 35733
rect 21541 35728 22711 35730
rect 21541 35672 21546 35728
rect 21602 35672 22650 35728
rect 22706 35672 22711 35728
rect 21541 35670 22711 35672
rect 20989 35667 21055 35668
rect 21541 35667 21607 35670
rect 22645 35667 22711 35670
rect 14733 35592 17234 35594
rect 14733 35536 14738 35592
rect 14794 35536 17234 35592
rect 14733 35534 17234 35536
rect 18229 35594 18295 35597
rect 23105 35594 23171 35597
rect 25589 35594 25655 35597
rect 18229 35592 25655 35594
rect 18229 35536 18234 35592
rect 18290 35536 23110 35592
rect 23166 35536 25594 35592
rect 25650 35536 25655 35592
rect 18229 35534 25655 35536
rect 14733 35531 14799 35534
rect 18229 35531 18295 35534
rect 23105 35531 23171 35534
rect 25589 35531 25655 35534
rect 5993 35458 6059 35461
rect 12801 35458 12867 35461
rect 5993 35456 12867 35458
rect 5993 35400 5998 35456
rect 6054 35400 12806 35456
rect 12862 35400 12867 35456
rect 5993 35398 12867 35400
rect 5993 35395 6059 35398
rect 12801 35395 12867 35398
rect 13261 35458 13327 35461
rect 13905 35458 13971 35461
rect 13261 35456 13971 35458
rect 13261 35400 13266 35456
rect 13322 35400 13910 35456
rect 13966 35400 13971 35456
rect 13261 35398 13971 35400
rect 13261 35395 13327 35398
rect 13905 35395 13971 35398
rect 15285 35458 15351 35461
rect 16481 35458 16547 35461
rect 15285 35456 16547 35458
rect 15285 35400 15290 35456
rect 15346 35400 16486 35456
rect 16542 35400 16547 35456
rect 15285 35398 16547 35400
rect 15285 35395 15351 35398
rect 16481 35395 16547 35398
rect 17493 35458 17559 35461
rect 19517 35458 19583 35461
rect 21081 35458 21147 35461
rect 17493 35456 21147 35458
rect 17493 35400 17498 35456
rect 17554 35400 19522 35456
rect 19578 35400 21086 35456
rect 21142 35400 21147 35456
rect 17493 35398 21147 35400
rect 17493 35395 17559 35398
rect 19517 35395 19583 35398
rect 21081 35395 21147 35398
rect 28165 35458 28231 35461
rect 29200 35458 30000 35548
rect 28165 35456 30000 35458
rect 28165 35400 28170 35456
rect 28226 35400 30000 35456
rect 28165 35398 30000 35400
rect 28165 35395 28231 35398
rect 5576 35392 5896 35393
rect 5576 35328 5584 35392
rect 5648 35328 5664 35392
rect 5728 35328 5744 35392
rect 5808 35328 5824 35392
rect 5888 35328 5896 35392
rect 5576 35327 5896 35328
rect 14840 35392 15160 35393
rect 14840 35328 14848 35392
rect 14912 35328 14928 35392
rect 14992 35328 15008 35392
rect 15072 35328 15088 35392
rect 15152 35328 15160 35392
rect 14840 35327 15160 35328
rect 24104 35392 24424 35393
rect 24104 35328 24112 35392
rect 24176 35328 24192 35392
rect 24256 35328 24272 35392
rect 24336 35328 24352 35392
rect 24416 35328 24424 35392
rect 24104 35327 24424 35328
rect 9213 35324 9279 35325
rect 9213 35322 9260 35324
rect 9168 35320 9260 35322
rect 9168 35264 9218 35320
rect 9168 35262 9260 35264
rect 9213 35260 9260 35262
rect 9324 35260 9330 35324
rect 9489 35322 9555 35325
rect 12014 35322 12020 35324
rect 9489 35320 12020 35322
rect 9489 35264 9494 35320
rect 9550 35264 12020 35320
rect 9489 35262 12020 35264
rect 9213 35259 9279 35260
rect 9489 35259 9555 35262
rect 12014 35260 12020 35262
rect 12084 35260 12090 35324
rect 12157 35322 12223 35325
rect 14641 35322 14707 35325
rect 12157 35320 14707 35322
rect 12157 35264 12162 35320
rect 12218 35264 14646 35320
rect 14702 35264 14707 35320
rect 12157 35262 14707 35264
rect 12157 35259 12223 35262
rect 14641 35259 14707 35262
rect 15285 35322 15351 35325
rect 21909 35322 21975 35325
rect 15285 35320 21975 35322
rect 15285 35264 15290 35320
rect 15346 35264 21914 35320
rect 21970 35264 21975 35320
rect 29200 35308 30000 35398
rect 15285 35262 21975 35264
rect 15285 35259 15351 35262
rect 21909 35259 21975 35262
rect 8385 35186 8451 35189
rect 9581 35186 9647 35189
rect 8385 35184 9647 35186
rect 8385 35128 8390 35184
rect 8446 35128 9586 35184
rect 9642 35128 9647 35184
rect 8385 35126 9647 35128
rect 8385 35123 8451 35126
rect 9581 35123 9647 35126
rect 9806 35124 9812 35188
rect 9876 35186 9882 35188
rect 16757 35186 16823 35189
rect 17585 35186 17651 35189
rect 17769 35186 17835 35189
rect 9876 35184 16823 35186
rect 9876 35128 16762 35184
rect 16818 35128 16823 35184
rect 9876 35126 16823 35128
rect 9876 35124 9882 35126
rect 16757 35123 16823 35126
rect 16990 35184 17835 35186
rect 16990 35128 17590 35184
rect 17646 35128 17774 35184
rect 17830 35128 17835 35184
rect 16990 35126 17835 35128
rect 9857 35050 9923 35053
rect 13261 35050 13327 35053
rect 9857 35048 13327 35050
rect 9857 34992 9862 35048
rect 9918 34992 13266 35048
rect 13322 34992 13327 35048
rect 9857 34990 13327 34992
rect 9857 34987 9923 34990
rect 13261 34987 13327 34990
rect 13486 34988 13492 35052
rect 13556 35050 13562 35052
rect 13721 35050 13787 35053
rect 13556 35048 13787 35050
rect 13556 34992 13726 35048
rect 13782 34992 13787 35048
rect 13556 34990 13787 34992
rect 13556 34988 13562 34990
rect 13721 34987 13787 34990
rect 13905 35050 13971 35053
rect 16990 35050 17050 35126
rect 17585 35123 17651 35126
rect 17769 35123 17835 35126
rect 18638 35124 18644 35188
rect 18708 35186 18714 35188
rect 20529 35186 20595 35189
rect 18708 35184 20595 35186
rect 18708 35128 20534 35184
rect 20590 35128 20595 35184
rect 18708 35126 20595 35128
rect 18708 35124 18714 35126
rect 20529 35123 20595 35126
rect 20897 35186 20963 35189
rect 24393 35186 24459 35189
rect 20897 35184 24459 35186
rect 20897 35128 20902 35184
rect 20958 35128 24398 35184
rect 24454 35128 24459 35184
rect 20897 35126 24459 35128
rect 20897 35123 20963 35126
rect 24393 35123 24459 35126
rect 22277 35050 22343 35053
rect 22921 35050 22987 35053
rect 13905 35048 17050 35050
rect 13905 34992 13910 35048
rect 13966 34992 17050 35048
rect 13905 34990 17050 34992
rect 17128 35048 22987 35050
rect 17128 34992 22282 35048
rect 22338 34992 22926 35048
rect 22982 34992 22987 35048
rect 17128 34990 22987 34992
rect 13905 34987 13971 34990
rect 8385 34914 8451 34917
rect 9949 34914 10015 34917
rect 8385 34912 10015 34914
rect 0 34778 800 34868
rect 8385 34856 8390 34912
rect 8446 34856 9954 34912
rect 10010 34856 10015 34912
rect 8385 34854 10015 34856
rect 8385 34851 8451 34854
rect 9949 34851 10015 34854
rect 10593 34914 10659 34917
rect 10726 34914 10732 34916
rect 10593 34912 10732 34914
rect 10593 34856 10598 34912
rect 10654 34856 10732 34912
rect 10593 34854 10732 34856
rect 10593 34851 10659 34854
rect 10726 34852 10732 34854
rect 10796 34852 10802 34916
rect 10869 34914 10935 34917
rect 17128 34914 17188 34990
rect 22277 34987 22343 34990
rect 22921 34987 22987 34990
rect 10869 34912 17188 34914
rect 10869 34856 10874 34912
rect 10930 34856 17188 34912
rect 10869 34854 17188 34856
rect 17309 34914 17375 34917
rect 18413 34914 18479 34917
rect 17309 34912 18479 34914
rect 17309 34856 17314 34912
rect 17370 34856 18418 34912
rect 18474 34856 18479 34912
rect 17309 34854 18479 34856
rect 10869 34851 10935 34854
rect 17309 34851 17375 34854
rect 18413 34851 18479 34854
rect 20161 34914 20227 34917
rect 20805 34914 20871 34917
rect 20161 34912 20871 34914
rect 20161 34856 20166 34912
rect 20222 34856 20810 34912
rect 20866 34856 20871 34912
rect 20161 34854 20871 34856
rect 20161 34851 20227 34854
rect 20805 34851 20871 34854
rect 21265 34914 21331 34917
rect 24761 34914 24827 34917
rect 21265 34912 24827 34914
rect 21265 34856 21270 34912
rect 21326 34856 24766 34912
rect 24822 34856 24827 34912
rect 21265 34854 24827 34856
rect 21265 34851 21331 34854
rect 24761 34851 24827 34854
rect 10208 34848 10528 34849
rect 10208 34784 10216 34848
rect 10280 34784 10296 34848
rect 10360 34784 10376 34848
rect 10440 34784 10456 34848
rect 10520 34784 10528 34848
rect 10208 34783 10528 34784
rect 19472 34848 19792 34849
rect 19472 34784 19480 34848
rect 19544 34784 19560 34848
rect 19624 34784 19640 34848
rect 19704 34784 19720 34848
rect 19784 34784 19792 34848
rect 19472 34783 19792 34784
rect 2773 34778 2839 34781
rect 0 34776 2839 34778
rect 0 34720 2778 34776
rect 2834 34720 2839 34776
rect 0 34718 2839 34720
rect 0 34628 800 34718
rect 2773 34715 2839 34718
rect 9806 34716 9812 34780
rect 9876 34778 9882 34780
rect 10041 34778 10107 34781
rect 11462 34778 11468 34780
rect 9876 34776 10107 34778
rect 9876 34720 10046 34776
rect 10102 34720 10107 34776
rect 10918 34744 11468 34778
rect 9876 34718 10107 34720
rect 9876 34716 9882 34718
rect 10041 34715 10107 34718
rect 10734 34718 11468 34744
rect 10734 34684 10978 34718
rect 11462 34716 11468 34718
rect 11532 34716 11538 34780
rect 12198 34716 12204 34780
rect 12268 34778 12274 34780
rect 16113 34778 16179 34781
rect 12268 34776 16179 34778
rect 12268 34720 16118 34776
rect 16174 34720 16179 34776
rect 12268 34718 16179 34720
rect 12268 34716 12274 34718
rect 16113 34715 16179 34718
rect 16481 34778 16547 34781
rect 18781 34778 18847 34781
rect 16481 34776 18847 34778
rect 16481 34720 16486 34776
rect 16542 34720 18786 34776
rect 18842 34720 18847 34776
rect 16481 34718 18847 34720
rect 16481 34715 16547 34718
rect 18781 34715 18847 34718
rect 20529 34778 20595 34781
rect 25589 34778 25655 34781
rect 20529 34776 25655 34778
rect 20529 34720 20534 34776
rect 20590 34720 25594 34776
rect 25650 34720 25655 34776
rect 20529 34718 25655 34720
rect 20529 34715 20595 34718
rect 25589 34715 25655 34718
rect 25865 34778 25931 34781
rect 29200 34778 30000 34868
rect 25865 34776 30000 34778
rect 25865 34720 25870 34776
rect 25926 34720 30000 34776
rect 25865 34718 30000 34720
rect 25865 34715 25931 34718
rect 10734 34676 10794 34684
rect 7097 34642 7163 34645
rect 7230 34642 7236 34644
rect 7097 34640 7236 34642
rect 7097 34584 7102 34640
rect 7158 34584 7236 34640
rect 7097 34582 7236 34584
rect 7097 34579 7163 34582
rect 7230 34580 7236 34582
rect 7300 34580 7306 34644
rect 7557 34642 7623 34645
rect 10182 34642 10794 34676
rect 7557 34640 10794 34642
rect 7557 34584 7562 34640
rect 7618 34616 10794 34640
rect 11237 34642 11303 34645
rect 15101 34642 15167 34645
rect 20805 34642 20871 34645
rect 11237 34640 20871 34642
rect 7618 34584 10242 34616
rect 7557 34582 10242 34584
rect 11237 34584 11242 34640
rect 11298 34584 15106 34640
rect 15162 34584 20810 34640
rect 20866 34584 20871 34640
rect 11237 34582 20871 34584
rect 7557 34579 7623 34582
rect 11237 34579 11303 34582
rect 15101 34579 15167 34582
rect 20805 34579 20871 34582
rect 22185 34640 22251 34645
rect 22185 34584 22190 34640
rect 22246 34584 22251 34640
rect 22185 34579 22251 34584
rect 24669 34642 24735 34645
rect 24945 34642 25011 34645
rect 24669 34640 25011 34642
rect 24669 34584 24674 34640
rect 24730 34584 24950 34640
rect 25006 34584 25011 34640
rect 29200 34628 30000 34718
rect 24669 34582 25011 34584
rect 24669 34579 24735 34582
rect 24945 34579 25011 34582
rect 9305 34506 9371 34509
rect 11973 34506 12039 34509
rect 9305 34504 12039 34506
rect 9305 34448 9310 34504
rect 9366 34448 11978 34504
rect 12034 34448 12039 34504
rect 9305 34446 12039 34448
rect 9305 34443 9371 34446
rect 11973 34443 12039 34446
rect 12249 34506 12315 34509
rect 18045 34506 18111 34509
rect 12249 34504 18111 34506
rect 12249 34448 12254 34504
rect 12310 34448 18050 34504
rect 18106 34448 18111 34504
rect 12249 34446 18111 34448
rect 12249 34443 12315 34446
rect 18045 34443 18111 34446
rect 18229 34506 18295 34509
rect 22188 34506 22248 34579
rect 18229 34504 22248 34506
rect 18229 34448 18234 34504
rect 18290 34448 22248 34504
rect 18229 34446 22248 34448
rect 18229 34443 18295 34446
rect 8753 34370 8819 34373
rect 13997 34370 14063 34373
rect 8753 34368 14063 34370
rect 8753 34312 8758 34368
rect 8814 34312 14002 34368
rect 14058 34312 14063 34368
rect 8753 34310 14063 34312
rect 8753 34307 8819 34310
rect 13997 34307 14063 34310
rect 15377 34370 15443 34373
rect 19057 34370 19123 34373
rect 15377 34368 19123 34370
rect 15377 34312 15382 34368
rect 15438 34312 19062 34368
rect 19118 34312 19123 34368
rect 15377 34310 19123 34312
rect 15377 34307 15443 34310
rect 19057 34307 19123 34310
rect 19333 34370 19399 34373
rect 19926 34370 19932 34372
rect 19333 34368 19932 34370
rect 19333 34312 19338 34368
rect 19394 34312 19932 34368
rect 19333 34310 19932 34312
rect 19333 34307 19399 34310
rect 19926 34308 19932 34310
rect 19996 34308 20002 34372
rect 20897 34370 20963 34373
rect 21030 34370 21036 34372
rect 20897 34368 21036 34370
rect 20897 34312 20902 34368
rect 20958 34312 21036 34368
rect 20897 34310 21036 34312
rect 20897 34307 20963 34310
rect 21030 34308 21036 34310
rect 21100 34308 21106 34372
rect 21173 34370 21239 34373
rect 23197 34370 23263 34373
rect 23657 34370 23723 34373
rect 21173 34368 23723 34370
rect 21173 34312 21178 34368
rect 21234 34312 23202 34368
rect 23258 34312 23662 34368
rect 23718 34312 23723 34368
rect 21173 34310 23723 34312
rect 21173 34307 21239 34310
rect 23197 34307 23263 34310
rect 23657 34307 23723 34310
rect 5576 34304 5896 34305
rect 5576 34240 5584 34304
rect 5648 34240 5664 34304
rect 5728 34240 5744 34304
rect 5808 34240 5824 34304
rect 5888 34240 5896 34304
rect 5576 34239 5896 34240
rect 14840 34304 15160 34305
rect 14840 34240 14848 34304
rect 14912 34240 14928 34304
rect 14992 34240 15008 34304
rect 15072 34240 15088 34304
rect 15152 34240 15160 34304
rect 14840 34239 15160 34240
rect 24104 34304 24424 34305
rect 24104 34240 24112 34304
rect 24176 34240 24192 34304
rect 24256 34240 24272 34304
rect 24336 34240 24352 34304
rect 24416 34240 24424 34304
rect 24104 34239 24424 34240
rect 8477 34234 8543 34237
rect 10910 34234 10916 34236
rect 8477 34232 10916 34234
rect 0 34098 800 34188
rect 8477 34176 8482 34232
rect 8538 34176 10916 34232
rect 8477 34174 10916 34176
rect 8477 34171 8543 34174
rect 10910 34172 10916 34174
rect 10980 34172 10986 34236
rect 11053 34234 11119 34237
rect 11053 34232 11944 34234
rect 11053 34176 11058 34232
rect 11114 34176 11944 34232
rect 11053 34174 11944 34176
rect 11053 34171 11119 34174
rect 2773 34098 2839 34101
rect 0 34096 2839 34098
rect 0 34040 2778 34096
rect 2834 34040 2839 34096
rect 0 34038 2839 34040
rect 0 33948 800 34038
rect 2773 34035 2839 34038
rect 7557 34098 7623 34101
rect 10726 34098 10732 34100
rect 7557 34096 10732 34098
rect 7557 34040 7562 34096
rect 7618 34040 10732 34096
rect 7557 34038 10732 34040
rect 7557 34035 7623 34038
rect 10726 34036 10732 34038
rect 10796 34036 10802 34100
rect 10869 34098 10935 34101
rect 11697 34098 11763 34101
rect 10869 34096 11763 34098
rect 10869 34040 10874 34096
rect 10930 34040 11702 34096
rect 11758 34040 11763 34096
rect 10869 34038 11763 34040
rect 11884 34098 11944 34174
rect 12014 34172 12020 34236
rect 12084 34234 12090 34236
rect 13905 34234 13971 34237
rect 12084 34232 13971 34234
rect 12084 34176 13910 34232
rect 13966 34176 13971 34232
rect 12084 34174 13971 34176
rect 12084 34172 12090 34174
rect 13905 34171 13971 34174
rect 14089 34234 14155 34237
rect 14641 34234 14707 34237
rect 14089 34232 14707 34234
rect 14089 34176 14094 34232
rect 14150 34176 14646 34232
rect 14702 34176 14707 34232
rect 14089 34174 14707 34176
rect 14089 34171 14155 34174
rect 14641 34171 14707 34174
rect 16430 34172 16436 34236
rect 16500 34234 16506 34236
rect 17861 34234 17927 34237
rect 23381 34234 23447 34237
rect 26325 34234 26391 34237
rect 16500 34232 23447 34234
rect 16500 34176 17866 34232
rect 17922 34176 23386 34232
rect 23442 34176 23447 34232
rect 16500 34174 23447 34176
rect 16500 34172 16506 34174
rect 17861 34171 17927 34174
rect 23381 34171 23447 34174
rect 24534 34232 26391 34234
rect 24534 34176 26330 34232
rect 26386 34176 26391 34232
rect 24534 34174 26391 34176
rect 15193 34098 15259 34101
rect 21173 34098 21239 34101
rect 11884 34038 15026 34098
rect 10869 34035 10935 34038
rect 11697 34035 11763 34038
rect 8477 33962 8543 33965
rect 9673 33962 9739 33965
rect 10409 33962 10475 33965
rect 12249 33962 12315 33965
rect 8477 33960 9739 33962
rect 8477 33904 8482 33960
rect 8538 33904 9678 33960
rect 9734 33904 9739 33960
rect 10182 33960 10475 33962
rect 10182 33928 10414 33960
rect 8477 33902 9739 33904
rect 8477 33899 8543 33902
rect 9673 33899 9739 33902
rect 9998 33904 10414 33928
rect 10470 33904 10475 33960
rect 9998 33902 10475 33904
rect 9998 33868 10242 33902
rect 10409 33899 10475 33902
rect 10596 33960 12315 33962
rect 10596 33904 12254 33960
rect 12310 33904 12315 33960
rect 10596 33902 12315 33904
rect 9998 33860 10058 33868
rect 9814 33829 10058 33860
rect 10596 33829 10656 33902
rect 12249 33899 12315 33902
rect 12382 33900 12388 33964
rect 12452 33962 12458 33964
rect 14549 33962 14615 33965
rect 12452 33960 14615 33962
rect 12452 33904 14554 33960
rect 14610 33904 14615 33960
rect 12452 33902 14615 33904
rect 14966 33962 15026 34038
rect 15193 34096 21239 34098
rect 15193 34040 15198 34096
rect 15254 34040 21178 34096
rect 21234 34040 21239 34096
rect 15193 34038 21239 34040
rect 15193 34035 15259 34038
rect 21173 34035 21239 34038
rect 21357 34098 21423 34101
rect 24534 34098 24594 34174
rect 26325 34171 26391 34174
rect 21357 34096 24594 34098
rect 21357 34040 21362 34096
rect 21418 34040 24594 34096
rect 21357 34038 24594 34040
rect 26141 34098 26207 34101
rect 29200 34098 30000 34188
rect 26141 34096 30000 34098
rect 26141 34040 26146 34096
rect 26202 34040 30000 34096
rect 26141 34038 30000 34040
rect 21357 34035 21423 34038
rect 26141 34035 26207 34038
rect 26509 33962 26575 33965
rect 14966 33960 26575 33962
rect 14966 33904 26514 33960
rect 26570 33904 26575 33960
rect 29200 33948 30000 34038
rect 14966 33902 26575 33904
rect 12452 33900 12458 33902
rect 14549 33899 14615 33902
rect 26509 33899 26575 33902
rect 9622 33764 9628 33828
rect 9692 33826 9698 33828
rect 9765 33826 10058 33829
rect 9692 33824 10058 33826
rect 9692 33768 9770 33824
rect 9826 33800 10058 33824
rect 10593 33824 10659 33829
rect 9826 33768 9874 33800
rect 9692 33766 9874 33768
rect 10593 33768 10598 33824
rect 10654 33768 10659 33824
rect 9692 33764 9698 33766
rect 9765 33763 9831 33766
rect 10593 33763 10659 33768
rect 10961 33826 11027 33829
rect 19333 33826 19399 33829
rect 10961 33824 19399 33826
rect 10961 33768 10966 33824
rect 11022 33768 19338 33824
rect 19394 33768 19399 33824
rect 10961 33766 19399 33768
rect 10961 33763 11027 33766
rect 19333 33763 19399 33766
rect 10208 33760 10528 33761
rect 10208 33696 10216 33760
rect 10280 33696 10296 33760
rect 10360 33696 10376 33760
rect 10440 33696 10456 33760
rect 10520 33696 10528 33760
rect 10208 33695 10528 33696
rect 19472 33760 19792 33761
rect 19472 33696 19480 33760
rect 19544 33696 19560 33760
rect 19624 33696 19640 33760
rect 19704 33696 19720 33760
rect 19784 33696 19792 33760
rect 19472 33695 19792 33696
rect 8937 33690 9003 33693
rect 10041 33690 10107 33693
rect 8937 33688 10107 33690
rect 8937 33632 8942 33688
rect 8998 33632 10046 33688
rect 10102 33632 10107 33688
rect 8937 33630 10107 33632
rect 8937 33627 9003 33630
rect 10041 33627 10107 33630
rect 10593 33690 10659 33693
rect 12985 33690 13051 33693
rect 10593 33688 13051 33690
rect 10593 33632 10598 33688
rect 10654 33632 12990 33688
rect 13046 33632 13051 33688
rect 10593 33630 13051 33632
rect 10593 33627 10659 33630
rect 12985 33627 13051 33630
rect 13118 33628 13124 33692
rect 13188 33690 13194 33692
rect 18689 33690 18755 33693
rect 13188 33688 18755 33690
rect 13188 33632 18694 33688
rect 18750 33632 18755 33688
rect 13188 33630 18755 33632
rect 13188 33628 13194 33630
rect 18689 33627 18755 33630
rect 8109 33554 8175 33557
rect 10409 33554 10475 33557
rect 8109 33552 10475 33554
rect 0 33418 800 33508
rect 8109 33496 8114 33552
rect 8170 33496 10414 33552
rect 10470 33496 10475 33552
rect 8109 33494 10475 33496
rect 8109 33491 8175 33494
rect 10409 33491 10475 33494
rect 11421 33554 11487 33557
rect 13813 33554 13879 33557
rect 11421 33552 13879 33554
rect 11421 33496 11426 33552
rect 11482 33496 13818 33552
rect 13874 33496 13879 33552
rect 11421 33494 13879 33496
rect 11421 33491 11487 33494
rect 13813 33491 13879 33494
rect 14406 33492 14412 33556
rect 14476 33554 14482 33556
rect 21357 33554 21423 33557
rect 14476 33552 21423 33554
rect 14476 33496 21362 33552
rect 21418 33496 21423 33552
rect 14476 33494 21423 33496
rect 14476 33492 14482 33494
rect 21357 33491 21423 33494
rect 1393 33418 1459 33421
rect 0 33416 1459 33418
rect 0 33360 1398 33416
rect 1454 33360 1459 33416
rect 0 33358 1459 33360
rect 0 33268 800 33358
rect 1393 33355 1459 33358
rect 10041 33418 10107 33421
rect 10596 33418 11116 33452
rect 13905 33418 13971 33421
rect 15101 33418 15167 33421
rect 10041 33416 13784 33418
rect 10041 33360 10046 33416
rect 10102 33392 13784 33416
rect 10102 33360 10656 33392
rect 10041 33358 10656 33360
rect 11056 33358 13784 33392
rect 10041 33355 10107 33358
rect 7557 33282 7623 33285
rect 10317 33282 10383 33285
rect 7557 33280 10383 33282
rect 7557 33224 7562 33280
rect 7618 33224 10322 33280
rect 10378 33224 10383 33280
rect 7557 33222 10383 33224
rect 7557 33219 7623 33222
rect 10317 33219 10383 33222
rect 10910 33220 10916 33284
rect 10980 33282 10986 33284
rect 11053 33282 11119 33285
rect 11462 33282 11468 33284
rect 10980 33280 11468 33282
rect 10980 33224 11058 33280
rect 11114 33224 11468 33280
rect 10980 33222 11468 33224
rect 10980 33220 10986 33222
rect 11053 33219 11119 33222
rect 11462 33220 11468 33222
rect 11532 33220 11538 33284
rect 11646 33220 11652 33284
rect 11716 33282 11722 33284
rect 12985 33282 13051 33285
rect 11716 33280 13051 33282
rect 11716 33224 12990 33280
rect 13046 33224 13051 33280
rect 11716 33222 13051 33224
rect 11716 33220 11722 33222
rect 12985 33219 13051 33222
rect 13261 33282 13327 33285
rect 13486 33282 13492 33284
rect 13261 33280 13492 33282
rect 13261 33224 13266 33280
rect 13322 33224 13492 33280
rect 13261 33222 13492 33224
rect 13261 33219 13327 33222
rect 13486 33220 13492 33222
rect 13556 33220 13562 33284
rect 13724 33282 13784 33358
rect 13905 33416 15167 33418
rect 13905 33360 13910 33416
rect 13966 33360 15106 33416
rect 15162 33360 15167 33416
rect 13905 33358 15167 33360
rect 13905 33355 13971 33358
rect 15101 33355 15167 33358
rect 15561 33418 15627 33421
rect 26325 33418 26391 33421
rect 15561 33416 26391 33418
rect 15561 33360 15566 33416
rect 15622 33360 26330 33416
rect 26386 33360 26391 33416
rect 15561 33358 26391 33360
rect 15561 33355 15627 33358
rect 26325 33355 26391 33358
rect 28165 33418 28231 33421
rect 29200 33418 30000 33508
rect 28165 33416 30000 33418
rect 28165 33360 28170 33416
rect 28226 33360 30000 33416
rect 28165 33358 30000 33360
rect 28165 33355 28231 33358
rect 14641 33282 14707 33285
rect 13724 33280 14707 33282
rect 13724 33224 14646 33280
rect 14702 33224 14707 33280
rect 13724 33222 14707 33224
rect 14641 33219 14707 33222
rect 17309 33282 17375 33285
rect 23473 33282 23539 33285
rect 17309 33280 23539 33282
rect 17309 33224 17314 33280
rect 17370 33224 23478 33280
rect 23534 33224 23539 33280
rect 29200 33268 30000 33358
rect 17309 33222 23539 33224
rect 17309 33219 17375 33222
rect 23473 33219 23539 33222
rect 5576 33216 5896 33217
rect 5576 33152 5584 33216
rect 5648 33152 5664 33216
rect 5728 33152 5744 33216
rect 5808 33152 5824 33216
rect 5888 33152 5896 33216
rect 5576 33151 5896 33152
rect 14840 33216 15160 33217
rect 14840 33152 14848 33216
rect 14912 33152 14928 33216
rect 14992 33152 15008 33216
rect 15072 33152 15088 33216
rect 15152 33152 15160 33216
rect 14840 33151 15160 33152
rect 24104 33216 24424 33217
rect 24104 33152 24112 33216
rect 24176 33152 24192 33216
rect 24256 33152 24272 33216
rect 24336 33152 24352 33216
rect 24416 33152 24424 33216
rect 24104 33151 24424 33152
rect 9397 33146 9463 33149
rect 9806 33146 9812 33148
rect 9397 33144 9812 33146
rect 9397 33088 9402 33144
rect 9458 33088 9812 33144
rect 9397 33086 9812 33088
rect 9397 33083 9463 33086
rect 9806 33084 9812 33086
rect 9876 33146 9882 33148
rect 10869 33146 10935 33149
rect 14457 33146 14523 33149
rect 9876 33144 14523 33146
rect 9876 33088 10874 33144
rect 10930 33088 14462 33144
rect 14518 33088 14523 33144
rect 9876 33086 14523 33088
rect 9876 33084 9882 33086
rect 10869 33083 10935 33086
rect 14457 33083 14523 33086
rect 18045 33146 18111 33149
rect 22461 33146 22527 33149
rect 18045 33144 22527 33146
rect 18045 33088 18050 33144
rect 18106 33088 22466 33144
rect 22522 33088 22527 33144
rect 18045 33086 22527 33088
rect 18045 33083 18111 33086
rect 22461 33083 22527 33086
rect 9765 33010 9831 33013
rect 12566 33010 12572 33012
rect 9765 33008 12572 33010
rect 9765 32952 9770 33008
rect 9826 32952 12572 33008
rect 9765 32950 12572 32952
rect 9765 32947 9831 32950
rect 12566 32948 12572 32950
rect 12636 32948 12642 33012
rect 12709 33010 12775 33013
rect 18413 33010 18479 33013
rect 12709 33008 18479 33010
rect 12709 32952 12714 33008
rect 12770 32952 18418 33008
rect 18474 32952 18479 33008
rect 12709 32950 18479 32952
rect 12709 32947 12775 32950
rect 18413 32947 18479 32950
rect 18689 33010 18755 33013
rect 20897 33010 20963 33013
rect 23933 33010 23999 33013
rect 18689 33008 23999 33010
rect 18689 32952 18694 33008
rect 18750 32952 20902 33008
rect 20958 32952 23938 33008
rect 23994 32952 23999 33008
rect 18689 32950 23999 32952
rect 18689 32947 18755 32950
rect 20897 32947 20963 32950
rect 23933 32947 23999 32950
rect 9673 32874 9739 32877
rect 11053 32874 11119 32877
rect 13537 32874 13603 32877
rect 9673 32872 10978 32874
rect 0 32738 800 32828
rect 9673 32816 9678 32872
rect 9734 32816 10978 32872
rect 9673 32814 10978 32816
rect 9673 32811 9739 32814
rect 2865 32738 2931 32741
rect 0 32736 2931 32738
rect 0 32680 2870 32736
rect 2926 32680 2931 32736
rect 0 32678 2931 32680
rect 0 32588 800 32678
rect 2865 32675 2931 32678
rect 10208 32672 10528 32673
rect 10208 32608 10216 32672
rect 10280 32608 10296 32672
rect 10360 32608 10376 32672
rect 10440 32608 10456 32672
rect 10520 32608 10528 32672
rect 10208 32607 10528 32608
rect 10918 32602 10978 32814
rect 11053 32872 13603 32874
rect 11053 32816 11058 32872
rect 11114 32816 13542 32872
rect 13598 32816 13603 32872
rect 11053 32814 13603 32816
rect 11053 32811 11119 32814
rect 13537 32811 13603 32814
rect 13721 32874 13787 32877
rect 22553 32874 22619 32877
rect 13721 32872 22619 32874
rect 13721 32816 13726 32872
rect 13782 32816 22558 32872
rect 22614 32816 22619 32872
rect 13721 32814 22619 32816
rect 13721 32811 13787 32814
rect 22553 32811 22619 32814
rect 23105 32874 23171 32877
rect 25773 32874 25839 32877
rect 23105 32872 25839 32874
rect 23105 32816 23110 32872
rect 23166 32816 25778 32872
rect 25834 32816 25839 32872
rect 23105 32814 25839 32816
rect 23105 32811 23171 32814
rect 25773 32811 25839 32814
rect 11237 32738 11303 32741
rect 11789 32738 11855 32741
rect 11237 32736 11855 32738
rect 11237 32680 11242 32736
rect 11298 32680 11794 32736
rect 11850 32680 11855 32736
rect 11237 32678 11855 32680
rect 11237 32675 11303 32678
rect 11789 32675 11855 32678
rect 12249 32738 12315 32741
rect 19333 32738 19399 32741
rect 12249 32736 19399 32738
rect 12249 32680 12254 32736
rect 12310 32680 19338 32736
rect 19394 32680 19399 32736
rect 12249 32678 19399 32680
rect 12249 32675 12315 32678
rect 19333 32675 19399 32678
rect 28165 32738 28231 32741
rect 29200 32738 30000 32828
rect 28165 32736 30000 32738
rect 28165 32680 28170 32736
rect 28226 32680 30000 32736
rect 28165 32678 30000 32680
rect 28165 32675 28231 32678
rect 19472 32672 19792 32673
rect 19472 32608 19480 32672
rect 19544 32608 19560 32672
rect 19624 32608 19640 32672
rect 19704 32608 19720 32672
rect 19784 32608 19792 32672
rect 19472 32607 19792 32608
rect 13353 32602 13419 32605
rect 10918 32600 13419 32602
rect 10918 32544 13358 32600
rect 13414 32544 13419 32600
rect 10918 32542 13419 32544
rect 13353 32539 13419 32542
rect 13486 32540 13492 32604
rect 13556 32602 13562 32604
rect 17309 32602 17375 32605
rect 13556 32600 17375 32602
rect 13556 32544 17314 32600
rect 17370 32544 17375 32600
rect 13556 32542 17375 32544
rect 13556 32540 13562 32542
rect 17309 32539 17375 32542
rect 22093 32602 22159 32605
rect 25037 32602 25103 32605
rect 22093 32600 25103 32602
rect 22093 32544 22098 32600
rect 22154 32544 25042 32600
rect 25098 32544 25103 32600
rect 29200 32588 30000 32678
rect 22093 32542 25103 32544
rect 22093 32539 22159 32542
rect 25037 32539 25103 32542
rect 9765 32466 9831 32469
rect 17493 32466 17559 32469
rect 9765 32464 17559 32466
rect 9765 32408 9770 32464
rect 9826 32408 17498 32464
rect 17554 32408 17559 32464
rect 9765 32406 17559 32408
rect 9765 32403 9831 32406
rect 17493 32403 17559 32406
rect 19333 32466 19399 32469
rect 26141 32466 26207 32469
rect 19333 32464 26207 32466
rect 19333 32408 19338 32464
rect 19394 32408 26146 32464
rect 26202 32408 26207 32464
rect 19333 32406 26207 32408
rect 19333 32403 19399 32406
rect 26141 32403 26207 32406
rect 8661 32330 8727 32333
rect 22093 32330 22159 32333
rect 26969 32330 27035 32333
rect 8661 32328 22159 32330
rect 8661 32272 8666 32328
rect 8722 32272 22098 32328
rect 22154 32272 22159 32328
rect 8661 32270 22159 32272
rect 8661 32267 8727 32270
rect 22093 32267 22159 32270
rect 23982 32328 27035 32330
rect 23982 32272 26974 32328
rect 27030 32272 27035 32328
rect 23982 32270 27035 32272
rect 9121 32194 9187 32197
rect 11278 32194 11284 32196
rect 9121 32192 11284 32194
rect 0 31908 800 32148
rect 9121 32136 9126 32192
rect 9182 32136 11284 32192
rect 9121 32134 11284 32136
rect 9121 32131 9187 32134
rect 11278 32132 11284 32134
rect 11348 32132 11354 32196
rect 11462 32132 11468 32196
rect 11532 32194 11538 32196
rect 12525 32194 12591 32197
rect 13997 32194 14063 32197
rect 11532 32192 12591 32194
rect 11532 32136 12530 32192
rect 12586 32136 12591 32192
rect 11532 32134 12591 32136
rect 11532 32132 11538 32134
rect 12525 32131 12591 32134
rect 12942 32192 14063 32194
rect 12942 32136 14002 32192
rect 14058 32136 14063 32192
rect 12942 32134 14063 32136
rect 5576 32128 5896 32129
rect 5576 32064 5584 32128
rect 5648 32064 5664 32128
rect 5728 32064 5744 32128
rect 5808 32064 5824 32128
rect 5888 32064 5896 32128
rect 5576 32063 5896 32064
rect 9121 32058 9187 32061
rect 12942 32058 13002 32134
rect 13997 32131 14063 32134
rect 14273 32194 14339 32197
rect 14641 32194 14707 32197
rect 14273 32192 14707 32194
rect 14273 32136 14278 32192
rect 14334 32136 14646 32192
rect 14702 32136 14707 32192
rect 14273 32134 14707 32136
rect 14273 32131 14339 32134
rect 14641 32131 14707 32134
rect 19517 32194 19583 32197
rect 23982 32194 24042 32270
rect 26969 32267 27035 32270
rect 19517 32192 24042 32194
rect 19517 32136 19522 32192
rect 19578 32136 24042 32192
rect 19517 32134 24042 32136
rect 19517 32131 19583 32134
rect 14840 32128 15160 32129
rect 14840 32064 14848 32128
rect 14912 32064 14928 32128
rect 14992 32064 15008 32128
rect 15072 32064 15088 32128
rect 15152 32064 15160 32128
rect 14840 32063 15160 32064
rect 24104 32128 24424 32129
rect 24104 32064 24112 32128
rect 24176 32064 24192 32128
rect 24256 32064 24272 32128
rect 24336 32064 24352 32128
rect 24416 32064 24424 32128
rect 24104 32063 24424 32064
rect 15285 32058 15351 32061
rect 19241 32058 19307 32061
rect 9121 32056 13002 32058
rect 9121 32000 9126 32056
rect 9182 32000 13002 32056
rect 9121 31998 13002 32000
rect 13080 31998 14474 32058
rect 9121 31995 9187 31998
rect 9949 31922 10015 31925
rect 13080 31922 13140 31998
rect 9949 31920 13140 31922
rect 9949 31864 9954 31920
rect 10010 31864 13140 31920
rect 9949 31862 13140 31864
rect 9949 31859 10015 31862
rect 13302 31860 13308 31924
rect 13372 31922 13378 31924
rect 13445 31922 13511 31925
rect 13372 31920 13511 31922
rect 13372 31864 13450 31920
rect 13506 31864 13511 31920
rect 13372 31862 13511 31864
rect 13372 31860 13378 31862
rect 13445 31859 13511 31862
rect 13813 31922 13879 31925
rect 14273 31922 14339 31925
rect 13813 31920 14339 31922
rect 13813 31864 13818 31920
rect 13874 31864 14278 31920
rect 14334 31864 14339 31920
rect 13813 31862 14339 31864
rect 14414 31922 14474 31998
rect 15285 32056 19307 32058
rect 15285 32000 15290 32056
rect 15346 32000 19246 32056
rect 19302 32000 19307 32056
rect 15285 31998 19307 32000
rect 15285 31995 15351 31998
rect 19241 31995 19307 31998
rect 19926 31996 19932 32060
rect 19996 32058 20002 32060
rect 20345 32058 20411 32061
rect 19996 32056 20411 32058
rect 19996 32000 20350 32056
rect 20406 32000 20411 32056
rect 19996 31998 20411 32000
rect 19996 31996 20002 31998
rect 20345 31995 20411 31998
rect 28717 32058 28783 32061
rect 29200 32058 30000 32148
rect 28717 32056 30000 32058
rect 28717 32000 28722 32056
rect 28778 32000 30000 32056
rect 28717 31998 30000 32000
rect 28717 31995 28783 31998
rect 16481 31922 16547 31925
rect 26325 31922 26391 31925
rect 14414 31920 16547 31922
rect 14414 31864 16486 31920
rect 16542 31864 16547 31920
rect 14414 31862 16547 31864
rect 13813 31859 13879 31862
rect 14273 31859 14339 31862
rect 16481 31859 16547 31862
rect 16622 31920 26391 31922
rect 16622 31864 26330 31920
rect 26386 31864 26391 31920
rect 29200 31908 30000 31998
rect 16622 31862 26391 31864
rect 10777 31786 10843 31789
rect 11421 31786 11487 31789
rect 9998 31726 10656 31786
rect 9397 31650 9463 31653
rect 9998 31650 10058 31726
rect 9397 31648 10058 31650
rect 9397 31592 9402 31648
rect 9458 31592 10058 31648
rect 9397 31590 10058 31592
rect 9397 31587 9463 31590
rect 10208 31584 10528 31585
rect 10208 31520 10216 31584
rect 10280 31520 10296 31584
rect 10360 31520 10376 31584
rect 10440 31520 10456 31584
rect 10520 31520 10528 31584
rect 10208 31519 10528 31520
rect 8937 31514 9003 31517
rect 9857 31514 9923 31517
rect 8937 31512 9923 31514
rect 0 31378 800 31468
rect 8937 31456 8942 31512
rect 8998 31456 9862 31512
rect 9918 31456 9923 31512
rect 8937 31454 9923 31456
rect 10596 31514 10656 31726
rect 10777 31784 11487 31786
rect 10777 31728 10782 31784
rect 10838 31728 11426 31784
rect 11482 31728 11487 31784
rect 10777 31726 11487 31728
rect 10777 31723 10843 31726
rect 11421 31723 11487 31726
rect 11973 31786 12039 31789
rect 14825 31786 14891 31789
rect 11973 31784 14891 31786
rect 11973 31728 11978 31784
rect 12034 31728 14830 31784
rect 14886 31728 14891 31784
rect 11973 31726 14891 31728
rect 11973 31723 12039 31726
rect 14825 31723 14891 31726
rect 15193 31786 15259 31789
rect 16622 31786 16682 31862
rect 26325 31859 26391 31862
rect 15193 31784 16682 31786
rect 15193 31728 15198 31784
rect 15254 31728 16682 31784
rect 15193 31726 16682 31728
rect 15193 31723 15259 31726
rect 20110 31724 20116 31788
rect 20180 31786 20186 31788
rect 20529 31786 20595 31789
rect 20180 31784 20595 31786
rect 20180 31728 20534 31784
rect 20590 31728 20595 31784
rect 20180 31726 20595 31728
rect 20180 31724 20186 31726
rect 20529 31723 20595 31726
rect 23381 31786 23447 31789
rect 25129 31786 25195 31789
rect 23381 31784 25195 31786
rect 23381 31728 23386 31784
rect 23442 31728 25134 31784
rect 25190 31728 25195 31784
rect 23381 31726 25195 31728
rect 23381 31723 23447 31726
rect 25129 31723 25195 31726
rect 11278 31588 11284 31652
rect 11348 31650 11354 31652
rect 13813 31650 13879 31653
rect 11348 31648 13879 31650
rect 11348 31592 13818 31648
rect 13874 31592 13879 31648
rect 11348 31590 13879 31592
rect 11348 31588 11354 31590
rect 13813 31587 13879 31590
rect 13997 31650 14063 31653
rect 17493 31650 17559 31653
rect 13997 31648 17559 31650
rect 13997 31592 14002 31648
rect 14058 31592 17498 31648
rect 17554 31592 17559 31648
rect 13997 31590 17559 31592
rect 13997 31587 14063 31590
rect 17493 31587 17559 31590
rect 19472 31584 19792 31585
rect 19472 31520 19480 31584
rect 19544 31520 19560 31584
rect 19624 31520 19640 31584
rect 19704 31520 19720 31584
rect 19784 31520 19792 31584
rect 19472 31519 19792 31520
rect 10596 31454 17234 31514
rect 8937 31451 9003 31454
rect 9857 31451 9923 31454
rect 2773 31378 2839 31381
rect 0 31376 2839 31378
rect 0 31320 2778 31376
rect 2834 31320 2839 31376
rect 0 31318 2839 31320
rect 0 31228 800 31318
rect 2773 31315 2839 31318
rect 9949 31378 10015 31381
rect 13721 31378 13787 31381
rect 9949 31376 13787 31378
rect 9949 31320 9954 31376
rect 10010 31320 13726 31376
rect 13782 31320 13787 31376
rect 9949 31318 13787 31320
rect 9949 31315 10015 31318
rect 13721 31315 13787 31318
rect 13854 31316 13860 31380
rect 13924 31378 13930 31380
rect 15101 31378 15167 31381
rect 13924 31376 15167 31378
rect 13924 31320 15106 31376
rect 15162 31320 15167 31376
rect 13924 31318 15167 31320
rect 13924 31316 13930 31318
rect 15101 31315 15167 31318
rect 16297 31378 16363 31381
rect 16481 31378 16547 31381
rect 16297 31376 16547 31378
rect 16297 31320 16302 31376
rect 16358 31320 16486 31376
rect 16542 31320 16547 31376
rect 16297 31318 16547 31320
rect 17174 31378 17234 31454
rect 26417 31378 26483 31381
rect 17174 31376 26483 31378
rect 17174 31320 26422 31376
rect 26478 31320 26483 31376
rect 17174 31318 26483 31320
rect 16297 31315 16363 31318
rect 16481 31315 16547 31318
rect 26417 31315 26483 31318
rect 8109 31242 8175 31245
rect 15193 31242 15259 31245
rect 8109 31240 15259 31242
rect 8109 31184 8114 31240
rect 8170 31184 15198 31240
rect 15254 31184 15259 31240
rect 8109 31182 15259 31184
rect 8109 31179 8175 31182
rect 15193 31179 15259 31182
rect 16205 31242 16271 31245
rect 19149 31242 19215 31245
rect 16205 31240 19215 31242
rect 16205 31184 16210 31240
rect 16266 31184 19154 31240
rect 19210 31184 19215 31240
rect 29200 31228 30000 31468
rect 16205 31182 19215 31184
rect 16205 31179 16271 31182
rect 19149 31179 19215 31182
rect 9806 31044 9812 31108
rect 9876 31106 9882 31108
rect 10726 31106 10732 31108
rect 9876 31046 10732 31106
rect 9876 31044 9882 31046
rect 10726 31044 10732 31046
rect 10796 31044 10802 31108
rect 10869 31106 10935 31109
rect 11697 31106 11763 31109
rect 10869 31104 11763 31106
rect 10869 31048 10874 31104
rect 10930 31048 11702 31104
rect 11758 31048 11763 31104
rect 10869 31046 11763 31048
rect 10869 31043 10935 31046
rect 11697 31043 11763 31046
rect 11881 31106 11947 31109
rect 14641 31106 14707 31109
rect 11881 31104 14707 31106
rect 11881 31048 11886 31104
rect 11942 31048 14646 31104
rect 14702 31048 14707 31104
rect 11881 31046 14707 31048
rect 11881 31043 11947 31046
rect 14641 31043 14707 31046
rect 5576 31040 5896 31041
rect 5576 30976 5584 31040
rect 5648 30976 5664 31040
rect 5728 30976 5744 31040
rect 5808 30976 5824 31040
rect 5888 30976 5896 31040
rect 5576 30975 5896 30976
rect 14840 31040 15160 31041
rect 14840 30976 14848 31040
rect 14912 30976 14928 31040
rect 14992 30976 15008 31040
rect 15072 30976 15088 31040
rect 15152 30976 15160 31040
rect 14840 30975 15160 30976
rect 24104 31040 24424 31041
rect 24104 30976 24112 31040
rect 24176 30976 24192 31040
rect 24256 30976 24272 31040
rect 24336 30976 24352 31040
rect 24416 30976 24424 31040
rect 24104 30975 24424 30976
rect 9397 30970 9463 30973
rect 10910 30970 10916 30972
rect 9397 30968 10916 30970
rect 9397 30912 9402 30968
rect 9458 30912 10916 30968
rect 9397 30910 10916 30912
rect 9397 30907 9463 30910
rect 10910 30908 10916 30910
rect 10980 30908 10986 30972
rect 11421 30970 11487 30973
rect 12709 30970 12775 30973
rect 11421 30968 12775 30970
rect 11421 30912 11426 30968
rect 11482 30912 12714 30968
rect 12770 30912 12775 30968
rect 11421 30910 12775 30912
rect 11421 30907 11487 30910
rect 12709 30907 12775 30910
rect 12893 30970 12959 30973
rect 14457 30970 14523 30973
rect 12893 30968 14523 30970
rect 12893 30912 12898 30968
rect 12954 30912 14462 30968
rect 14518 30912 14523 30968
rect 12893 30910 14523 30912
rect 12893 30907 12959 30910
rect 14457 30907 14523 30910
rect 15469 30970 15535 30973
rect 17769 30970 17835 30973
rect 15469 30968 17835 30970
rect 15469 30912 15474 30968
rect 15530 30912 17774 30968
rect 17830 30912 17835 30968
rect 15469 30910 17835 30912
rect 15469 30907 15535 30910
rect 17769 30907 17835 30910
rect 8569 30834 8635 30837
rect 23289 30834 23355 30837
rect 8569 30832 23355 30834
rect 0 30548 800 30788
rect 8569 30776 8574 30832
rect 8630 30776 23294 30832
rect 23350 30776 23355 30832
rect 8569 30774 23355 30776
rect 8569 30771 8635 30774
rect 23289 30771 23355 30774
rect 9121 30698 9187 30701
rect 10777 30698 10843 30701
rect 12709 30698 12775 30701
rect 9121 30696 10656 30698
rect 9121 30640 9126 30696
rect 9182 30640 10656 30696
rect 9121 30638 10656 30640
rect 9121 30635 9187 30638
rect 8201 30562 8267 30565
rect 10041 30562 10107 30565
rect 8201 30560 10107 30562
rect 8201 30504 8206 30560
rect 8262 30504 10046 30560
rect 10102 30504 10107 30560
rect 8201 30502 10107 30504
rect 10596 30562 10656 30638
rect 10777 30696 12775 30698
rect 10777 30640 10782 30696
rect 10838 30640 12714 30696
rect 12770 30640 12775 30696
rect 10777 30638 12775 30640
rect 10777 30635 10843 30638
rect 12709 30635 12775 30638
rect 13077 30698 13143 30701
rect 19057 30698 19123 30701
rect 13077 30696 19123 30698
rect 13077 30640 13082 30696
rect 13138 30640 19062 30696
rect 19118 30640 19123 30696
rect 13077 30638 19123 30640
rect 13077 30635 13143 30638
rect 19057 30635 19123 30638
rect 19609 30698 19675 30701
rect 22461 30698 22527 30701
rect 19609 30696 22527 30698
rect 19609 30640 19614 30696
rect 19670 30640 22466 30696
rect 22522 30640 22527 30696
rect 19609 30638 22527 30640
rect 19609 30635 19675 30638
rect 22461 30635 22527 30638
rect 11881 30562 11947 30565
rect 10596 30560 11947 30562
rect 10596 30504 11886 30560
rect 11942 30504 11947 30560
rect 10596 30502 11947 30504
rect 8201 30499 8267 30502
rect 10041 30499 10107 30502
rect 11881 30499 11947 30502
rect 12341 30562 12407 30565
rect 14181 30562 14247 30565
rect 12341 30560 14247 30562
rect 12341 30504 12346 30560
rect 12402 30504 14186 30560
rect 14242 30504 14247 30560
rect 12341 30502 14247 30504
rect 12341 30499 12407 30502
rect 14181 30499 14247 30502
rect 14457 30562 14523 30565
rect 18873 30562 18939 30565
rect 14457 30560 18939 30562
rect 14457 30504 14462 30560
rect 14518 30504 18878 30560
rect 18934 30504 18939 30560
rect 29200 30548 30000 30788
rect 14457 30502 18939 30504
rect 14457 30499 14523 30502
rect 18873 30499 18939 30502
rect 10208 30496 10528 30497
rect 10208 30432 10216 30496
rect 10280 30432 10296 30496
rect 10360 30432 10376 30496
rect 10440 30432 10456 30496
rect 10520 30432 10528 30496
rect 10208 30431 10528 30432
rect 19472 30496 19792 30497
rect 19472 30432 19480 30496
rect 19544 30432 19560 30496
rect 19624 30432 19640 30496
rect 19704 30432 19720 30496
rect 19784 30432 19792 30496
rect 19472 30431 19792 30432
rect 9857 30426 9923 30429
rect 9990 30426 9996 30428
rect 9857 30424 9996 30426
rect 9857 30368 9862 30424
rect 9918 30368 9996 30424
rect 9857 30366 9996 30368
rect 9857 30363 9923 30366
rect 9990 30364 9996 30366
rect 10060 30364 10066 30428
rect 11697 30426 11763 30429
rect 13169 30426 13235 30429
rect 11697 30424 13235 30426
rect 11697 30368 11702 30424
rect 11758 30368 13174 30424
rect 13230 30368 13235 30424
rect 11697 30366 13235 30368
rect 11697 30363 11763 30366
rect 13169 30363 13235 30366
rect 13353 30426 13419 30429
rect 16941 30426 17007 30429
rect 13353 30424 17007 30426
rect 13353 30368 13358 30424
rect 13414 30368 16946 30424
rect 17002 30368 17007 30424
rect 13353 30366 17007 30368
rect 13353 30363 13419 30366
rect 16941 30363 17007 30366
rect 21357 30426 21423 30429
rect 26049 30426 26115 30429
rect 21357 30424 26115 30426
rect 21357 30368 21362 30424
rect 21418 30368 26054 30424
rect 26110 30368 26115 30424
rect 21357 30366 26115 30368
rect 21357 30363 21423 30366
rect 26049 30363 26115 30366
rect 26325 30426 26391 30429
rect 26550 30426 26556 30428
rect 26325 30424 26556 30426
rect 26325 30368 26330 30424
rect 26386 30368 26556 30424
rect 26325 30366 26556 30368
rect 26325 30363 26391 30366
rect 26550 30364 26556 30366
rect 26620 30364 26626 30428
rect 9489 30290 9555 30293
rect 16757 30290 16823 30293
rect 9489 30288 16823 30290
rect 9489 30232 9494 30288
rect 9550 30232 16762 30288
rect 16818 30232 16823 30288
rect 9489 30230 16823 30232
rect 9489 30227 9555 30230
rect 16757 30227 16823 30230
rect 16982 30228 16988 30292
rect 17052 30290 17058 30292
rect 21081 30290 21147 30293
rect 17052 30288 21147 30290
rect 17052 30232 21086 30288
rect 21142 30232 21147 30288
rect 17052 30230 21147 30232
rect 17052 30228 17058 30230
rect 21081 30227 21147 30230
rect 9949 30154 10015 30157
rect 12065 30154 12131 30157
rect 9949 30152 12131 30154
rect 0 30018 800 30108
rect 9949 30096 9954 30152
rect 10010 30096 12070 30152
rect 12126 30096 12131 30152
rect 9949 30094 12131 30096
rect 9949 30091 10015 30094
rect 12065 30091 12131 30094
rect 12198 30092 12204 30156
rect 12268 30154 12274 30156
rect 12433 30154 12499 30157
rect 12268 30152 12499 30154
rect 12268 30096 12438 30152
rect 12494 30096 12499 30152
rect 12268 30094 12499 30096
rect 12268 30092 12274 30094
rect 12433 30091 12499 30094
rect 12709 30154 12775 30157
rect 17125 30154 17191 30157
rect 12709 30152 17191 30154
rect 12709 30096 12714 30152
rect 12770 30096 17130 30152
rect 17186 30096 17191 30152
rect 12709 30094 17191 30096
rect 12709 30091 12775 30094
rect 17125 30091 17191 30094
rect 18413 30154 18479 30157
rect 19425 30154 19491 30157
rect 18413 30152 19491 30154
rect 18413 30096 18418 30152
rect 18474 30096 19430 30152
rect 19486 30096 19491 30152
rect 18413 30094 19491 30096
rect 18413 30091 18479 30094
rect 19425 30091 19491 30094
rect 19977 30154 20043 30157
rect 25957 30154 26023 30157
rect 19977 30152 26023 30154
rect 19977 30096 19982 30152
rect 20038 30096 25962 30152
rect 26018 30096 26023 30152
rect 19977 30094 26023 30096
rect 19977 30091 20043 30094
rect 25957 30091 26023 30094
rect 3877 30018 3943 30021
rect 0 30016 3943 30018
rect 0 29960 3882 30016
rect 3938 29960 3943 30016
rect 0 29958 3943 29960
rect 0 29868 800 29958
rect 3877 29955 3943 29958
rect 9305 30018 9371 30021
rect 14089 30020 14155 30021
rect 9305 30016 13186 30018
rect 9305 29960 9310 30016
rect 9366 29960 13186 30016
rect 9305 29958 13186 29960
rect 9305 29955 9371 29958
rect 5576 29952 5896 29953
rect 5576 29888 5584 29952
rect 5648 29888 5664 29952
rect 5728 29888 5744 29952
rect 5808 29888 5824 29952
rect 5888 29888 5896 29952
rect 5576 29887 5896 29888
rect 8569 29882 8635 29885
rect 12985 29882 13051 29885
rect 8569 29880 13051 29882
rect 8569 29824 8574 29880
rect 8630 29824 12990 29880
rect 13046 29824 13051 29880
rect 8569 29822 13051 29824
rect 8569 29819 8635 29822
rect 12985 29819 13051 29822
rect 8661 29746 8727 29749
rect 11513 29746 11579 29749
rect 12617 29746 12683 29749
rect 8661 29744 12683 29746
rect 8661 29688 8666 29744
rect 8722 29688 11518 29744
rect 11574 29688 12622 29744
rect 12678 29688 12683 29744
rect 8661 29686 12683 29688
rect 13126 29746 13186 29958
rect 14038 29956 14044 30020
rect 14108 30018 14155 30020
rect 15837 30018 15903 30021
rect 17769 30018 17835 30021
rect 20989 30018 21055 30021
rect 14108 30016 14200 30018
rect 14150 29960 14200 30016
rect 14108 29958 14200 29960
rect 15837 30016 21055 30018
rect 15837 29960 15842 30016
rect 15898 29960 17774 30016
rect 17830 29960 20994 30016
rect 21050 29960 21055 30016
rect 15837 29958 21055 29960
rect 14108 29956 14155 29958
rect 14089 29955 14155 29956
rect 15837 29955 15903 29958
rect 17769 29955 17835 29958
rect 20989 29955 21055 29958
rect 24945 30018 25011 30021
rect 29200 30018 30000 30108
rect 24945 30016 30000 30018
rect 24945 29960 24950 30016
rect 25006 29960 30000 30016
rect 24945 29958 30000 29960
rect 24945 29955 25011 29958
rect 14840 29952 15160 29953
rect 14840 29888 14848 29952
rect 14912 29888 14928 29952
rect 14992 29888 15008 29952
rect 15072 29888 15088 29952
rect 15152 29888 15160 29952
rect 14840 29887 15160 29888
rect 24104 29952 24424 29953
rect 24104 29888 24112 29952
rect 24176 29888 24192 29952
rect 24256 29888 24272 29952
rect 24336 29888 24352 29952
rect 24416 29888 24424 29952
rect 24104 29887 24424 29888
rect 13261 29882 13327 29885
rect 13445 29882 13511 29885
rect 14365 29882 14431 29885
rect 13261 29880 14431 29882
rect 13261 29824 13266 29880
rect 13322 29824 13450 29880
rect 13506 29824 14370 29880
rect 14426 29824 14431 29880
rect 13261 29822 14431 29824
rect 13261 29819 13327 29822
rect 13445 29819 13511 29822
rect 14365 29819 14431 29822
rect 15285 29882 15351 29885
rect 16798 29882 16804 29884
rect 15285 29880 16804 29882
rect 15285 29824 15290 29880
rect 15346 29824 16804 29880
rect 15285 29822 16804 29824
rect 15285 29819 15351 29822
rect 16798 29820 16804 29822
rect 16868 29820 16874 29884
rect 16941 29882 17007 29885
rect 23749 29882 23815 29885
rect 16941 29880 23815 29882
rect 16941 29824 16946 29880
rect 17002 29824 23754 29880
rect 23810 29824 23815 29880
rect 29200 29868 30000 29958
rect 16941 29822 23815 29824
rect 16941 29819 17007 29822
rect 23749 29819 23815 29822
rect 17493 29746 17559 29749
rect 17953 29746 18019 29749
rect 19241 29746 19307 29749
rect 13126 29744 18019 29746
rect 13126 29688 17498 29744
rect 17554 29688 17958 29744
rect 18014 29688 18019 29744
rect 13126 29686 18019 29688
rect 8661 29683 8727 29686
rect 11513 29683 11579 29686
rect 12617 29683 12683 29686
rect 17493 29683 17559 29686
rect 17953 29683 18019 29686
rect 18094 29744 19307 29746
rect 18094 29688 19246 29744
rect 19302 29688 19307 29744
rect 18094 29686 19307 29688
rect 8385 29610 8451 29613
rect 11973 29610 12039 29613
rect 8385 29608 12039 29610
rect 8385 29552 8390 29608
rect 8446 29552 11978 29608
rect 12034 29552 12039 29608
rect 8385 29550 12039 29552
rect 8385 29547 8451 29550
rect 11973 29547 12039 29550
rect 12249 29610 12315 29613
rect 12985 29610 13051 29613
rect 13445 29610 13511 29613
rect 12249 29608 13511 29610
rect 12249 29552 12254 29608
rect 12310 29552 12990 29608
rect 13046 29552 13450 29608
rect 13506 29552 13511 29608
rect 12249 29550 13511 29552
rect 12249 29547 12315 29550
rect 12985 29547 13051 29550
rect 13445 29547 13511 29550
rect 14457 29610 14523 29613
rect 18094 29610 18154 29686
rect 19241 29683 19307 29686
rect 21541 29746 21607 29749
rect 22185 29746 22251 29749
rect 21541 29744 22251 29746
rect 21541 29688 21546 29744
rect 21602 29688 22190 29744
rect 22246 29688 22251 29744
rect 21541 29686 22251 29688
rect 21541 29683 21607 29686
rect 22185 29683 22251 29686
rect 23289 29746 23355 29749
rect 25589 29746 25655 29749
rect 23289 29744 25655 29746
rect 23289 29688 23294 29744
rect 23350 29688 25594 29744
rect 25650 29688 25655 29744
rect 23289 29686 25655 29688
rect 23289 29683 23355 29686
rect 25589 29683 25655 29686
rect 14457 29608 18154 29610
rect 14457 29552 14462 29608
rect 14518 29552 18154 29608
rect 14457 29550 18154 29552
rect 19333 29610 19399 29613
rect 19926 29610 19932 29612
rect 19333 29608 19932 29610
rect 19333 29552 19338 29608
rect 19394 29552 19932 29608
rect 19333 29550 19932 29552
rect 14457 29547 14523 29550
rect 19333 29547 19399 29550
rect 19926 29548 19932 29550
rect 19996 29548 20002 29612
rect 21725 29610 21791 29613
rect 25129 29610 25195 29613
rect 21725 29608 25195 29610
rect 21725 29552 21730 29608
rect 21786 29552 25134 29608
rect 25190 29552 25195 29608
rect 21725 29550 25195 29552
rect 21725 29547 21791 29550
rect 25129 29547 25195 29550
rect 10869 29474 10935 29477
rect 11646 29474 11652 29476
rect 10869 29472 11652 29474
rect 0 29338 800 29428
rect 10869 29416 10874 29472
rect 10930 29416 11652 29472
rect 10869 29414 11652 29416
rect 10869 29411 10935 29414
rect 11646 29412 11652 29414
rect 11716 29412 11722 29476
rect 11789 29474 11855 29477
rect 12198 29474 12204 29476
rect 11789 29472 12204 29474
rect 11789 29416 11794 29472
rect 11850 29416 12204 29472
rect 11789 29414 12204 29416
rect 11789 29411 11855 29414
rect 12198 29412 12204 29414
rect 12268 29412 12274 29476
rect 12433 29474 12499 29477
rect 19057 29474 19123 29477
rect 12433 29472 19123 29474
rect 12433 29416 12438 29472
rect 12494 29416 19062 29472
rect 19118 29416 19123 29472
rect 12433 29414 19123 29416
rect 12433 29411 12499 29414
rect 19057 29411 19123 29414
rect 22093 29476 22159 29477
rect 22093 29472 22140 29476
rect 22204 29474 22210 29476
rect 23749 29474 23815 29477
rect 22204 29472 23815 29474
rect 22093 29416 22098 29472
rect 22204 29416 23754 29472
rect 23810 29416 23815 29472
rect 22093 29412 22140 29416
rect 22204 29414 23815 29416
rect 22204 29412 22210 29414
rect 22093 29411 22159 29412
rect 23749 29411 23815 29414
rect 10208 29408 10528 29409
rect 10208 29344 10216 29408
rect 10280 29344 10296 29408
rect 10360 29344 10376 29408
rect 10440 29344 10456 29408
rect 10520 29344 10528 29408
rect 10208 29343 10528 29344
rect 19472 29408 19792 29409
rect 19472 29344 19480 29408
rect 19544 29344 19560 29408
rect 19624 29344 19640 29408
rect 19704 29344 19720 29408
rect 19784 29344 19792 29408
rect 19472 29343 19792 29344
rect 2773 29338 2839 29341
rect 0 29336 2839 29338
rect 0 29280 2778 29336
rect 2834 29280 2839 29336
rect 0 29278 2839 29280
rect 0 29188 800 29278
rect 2773 29275 2839 29278
rect 9765 29340 9831 29341
rect 9765 29336 9812 29340
rect 9876 29338 9882 29340
rect 10593 29338 10659 29341
rect 15929 29338 15995 29341
rect 9765 29280 9770 29336
rect 9765 29276 9812 29280
rect 9876 29278 9922 29338
rect 10593 29336 15995 29338
rect 10593 29280 10598 29336
rect 10654 29280 15934 29336
rect 15990 29280 15995 29336
rect 10593 29278 15995 29280
rect 9876 29276 9882 29278
rect 9765 29275 9831 29276
rect 10593 29275 10659 29278
rect 15929 29275 15995 29278
rect 16849 29338 16915 29341
rect 18413 29338 18479 29341
rect 16849 29336 18479 29338
rect 16849 29280 16854 29336
rect 16910 29280 18418 29336
rect 18474 29280 18479 29336
rect 16849 29278 18479 29280
rect 16849 29275 16915 29278
rect 18413 29275 18479 29278
rect 21541 29338 21607 29341
rect 23657 29338 23723 29341
rect 21541 29336 23723 29338
rect 21541 29280 21546 29336
rect 21602 29280 23662 29336
rect 23718 29280 23723 29336
rect 21541 29278 23723 29280
rect 21541 29275 21607 29278
rect 23657 29275 23723 29278
rect 24577 29338 24643 29341
rect 26601 29338 26667 29341
rect 24577 29336 26667 29338
rect 24577 29280 24582 29336
rect 24638 29280 26606 29336
rect 26662 29280 26667 29336
rect 24577 29278 26667 29280
rect 24577 29275 24643 29278
rect 26601 29275 26667 29278
rect 28165 29338 28231 29341
rect 29200 29338 30000 29428
rect 28165 29336 30000 29338
rect 28165 29280 28170 29336
rect 28226 29280 30000 29336
rect 28165 29278 30000 29280
rect 28165 29275 28231 29278
rect 9397 29202 9463 29205
rect 12382 29202 12388 29204
rect 9397 29200 12388 29202
rect 9397 29144 9402 29200
rect 9458 29144 12388 29200
rect 9397 29142 12388 29144
rect 9397 29139 9463 29142
rect 12382 29140 12388 29142
rect 12452 29140 12458 29204
rect 12617 29202 12683 29205
rect 15193 29202 15259 29205
rect 12617 29200 15259 29202
rect 12617 29144 12622 29200
rect 12678 29144 15198 29200
rect 15254 29144 15259 29200
rect 12617 29142 15259 29144
rect 12617 29139 12683 29142
rect 15193 29139 15259 29142
rect 15469 29202 15535 29205
rect 24025 29202 24091 29205
rect 15469 29200 24091 29202
rect 15469 29144 15474 29200
rect 15530 29144 24030 29200
rect 24086 29144 24091 29200
rect 29200 29188 30000 29278
rect 15469 29142 24091 29144
rect 15469 29139 15535 29142
rect 24025 29139 24091 29142
rect 9121 29066 9187 29069
rect 11605 29066 11671 29069
rect 9121 29064 11671 29066
rect 9121 29008 9126 29064
rect 9182 29008 11610 29064
rect 11666 29008 11671 29064
rect 9121 29006 11671 29008
rect 9121 29003 9187 29006
rect 11605 29003 11671 29006
rect 11973 29066 12039 29069
rect 13077 29066 13143 29069
rect 18045 29066 18111 29069
rect 11973 29064 13143 29066
rect 11973 29008 11978 29064
rect 12034 29008 13082 29064
rect 13138 29008 13143 29064
rect 11973 29006 13143 29008
rect 11973 29003 12039 29006
rect 13077 29003 13143 29006
rect 13356 29064 18111 29066
rect 13356 29008 18050 29064
rect 18106 29008 18111 29064
rect 13356 29006 18111 29008
rect 9121 28930 9187 28933
rect 12433 28930 12499 28933
rect 9121 28928 12499 28930
rect 9121 28872 9126 28928
rect 9182 28872 12438 28928
rect 12494 28872 12499 28928
rect 9121 28870 12499 28872
rect 9121 28867 9187 28870
rect 12433 28867 12499 28870
rect 12566 28868 12572 28932
rect 12636 28930 12642 28932
rect 13356 28930 13416 29006
rect 18045 29003 18111 29006
rect 18454 29004 18460 29068
rect 18524 29066 18530 29068
rect 21909 29066 21975 29069
rect 18524 29064 21975 29066
rect 18524 29008 21914 29064
rect 21970 29008 21975 29064
rect 18524 29006 21975 29008
rect 18524 29004 18530 29006
rect 21909 29003 21975 29006
rect 22093 29066 22159 29069
rect 23105 29066 23171 29069
rect 22093 29064 23171 29066
rect 22093 29008 22098 29064
rect 22154 29008 23110 29064
rect 23166 29008 23171 29064
rect 22093 29006 23171 29008
rect 22093 29003 22159 29006
rect 23105 29003 23171 29006
rect 12636 28870 13416 28930
rect 15285 28930 15351 28933
rect 17585 28930 17651 28933
rect 20110 28930 20116 28932
rect 15285 28928 20116 28930
rect 15285 28872 15290 28928
rect 15346 28872 17590 28928
rect 17646 28872 20116 28928
rect 15285 28870 20116 28872
rect 12636 28868 12642 28870
rect 15285 28867 15351 28870
rect 17585 28867 17651 28870
rect 20110 28868 20116 28870
rect 20180 28868 20186 28932
rect 20989 28930 21055 28933
rect 23381 28930 23447 28933
rect 20989 28928 23447 28930
rect 20989 28872 20994 28928
rect 21050 28872 23386 28928
rect 23442 28872 23447 28928
rect 20989 28870 23447 28872
rect 20989 28867 21055 28870
rect 23381 28867 23447 28870
rect 5576 28864 5896 28865
rect 5576 28800 5584 28864
rect 5648 28800 5664 28864
rect 5728 28800 5744 28864
rect 5808 28800 5824 28864
rect 5888 28800 5896 28864
rect 5576 28799 5896 28800
rect 14840 28864 15160 28865
rect 14840 28800 14848 28864
rect 14912 28800 14928 28864
rect 14992 28800 15008 28864
rect 15072 28800 15088 28864
rect 15152 28800 15160 28864
rect 14840 28799 15160 28800
rect 24104 28864 24424 28865
rect 24104 28800 24112 28864
rect 24176 28800 24192 28864
rect 24256 28800 24272 28864
rect 24336 28800 24352 28864
rect 24416 28800 24424 28864
rect 24104 28799 24424 28800
rect 9949 28794 10015 28797
rect 10501 28794 10567 28797
rect 9949 28792 10567 28794
rect 0 28508 800 28748
rect 9949 28736 9954 28792
rect 10010 28736 10506 28792
rect 10562 28736 10567 28792
rect 9949 28734 10567 28736
rect 9949 28731 10015 28734
rect 10501 28731 10567 28734
rect 11053 28794 11119 28797
rect 14181 28794 14247 28797
rect 11053 28792 14247 28794
rect 11053 28736 11058 28792
rect 11114 28736 14186 28792
rect 14242 28736 14247 28792
rect 11053 28734 14247 28736
rect 11053 28731 11119 28734
rect 14181 28731 14247 28734
rect 15285 28794 15351 28797
rect 19333 28794 19399 28797
rect 15285 28792 19399 28794
rect 15285 28736 15290 28792
rect 15346 28736 19338 28792
rect 19394 28736 19399 28792
rect 15285 28734 19399 28736
rect 15285 28731 15351 28734
rect 19333 28731 19399 28734
rect 19885 28794 19951 28797
rect 20805 28794 20871 28797
rect 19885 28792 20871 28794
rect 19885 28736 19890 28792
rect 19946 28736 20810 28792
rect 20866 28736 20871 28792
rect 19885 28734 20871 28736
rect 19885 28731 19951 28734
rect 20805 28731 20871 28734
rect 10041 28658 10107 28661
rect 12433 28658 12499 28661
rect 10041 28656 12499 28658
rect 10041 28600 10046 28656
rect 10102 28600 12438 28656
rect 12494 28600 12499 28656
rect 10041 28598 12499 28600
rect 10041 28595 10107 28598
rect 12433 28595 12499 28598
rect 12617 28658 12683 28661
rect 16757 28658 16823 28661
rect 16941 28660 17007 28661
rect 16941 28658 16988 28660
rect 12617 28656 16823 28658
rect 12617 28600 12622 28656
rect 12678 28600 16762 28656
rect 16818 28600 16823 28656
rect 12617 28598 16823 28600
rect 16896 28656 16988 28658
rect 16896 28600 16946 28656
rect 16896 28598 16988 28600
rect 12617 28595 12683 28598
rect 16757 28595 16823 28598
rect 16941 28596 16988 28598
rect 17052 28596 17058 28660
rect 19793 28658 19859 28661
rect 19926 28658 19932 28660
rect 19793 28656 19932 28658
rect 19793 28600 19798 28656
rect 19854 28600 19932 28656
rect 19793 28598 19932 28600
rect 16941 28595 17007 28596
rect 19793 28595 19859 28598
rect 19926 28596 19932 28598
rect 19996 28596 20002 28660
rect 9029 28522 9095 28525
rect 11053 28522 11119 28525
rect 12617 28522 12683 28525
rect 9029 28520 10978 28522
rect 9029 28464 9034 28520
rect 9090 28464 10978 28520
rect 9029 28462 10978 28464
rect 9029 28459 9095 28462
rect 10918 28386 10978 28462
rect 11053 28520 12683 28522
rect 11053 28464 11058 28520
rect 11114 28464 12622 28520
rect 12678 28464 12683 28520
rect 11053 28462 12683 28464
rect 11053 28459 11119 28462
rect 12617 28459 12683 28462
rect 12893 28522 12959 28525
rect 18413 28522 18479 28525
rect 19057 28522 19123 28525
rect 12893 28520 19123 28522
rect 12893 28464 12898 28520
rect 12954 28464 18418 28520
rect 18474 28464 19062 28520
rect 19118 28464 19123 28520
rect 12893 28462 19123 28464
rect 12893 28459 12959 28462
rect 18413 28459 18479 28462
rect 19057 28459 19123 28462
rect 19701 28522 19767 28525
rect 22093 28522 22159 28525
rect 22829 28522 22895 28525
rect 19701 28520 19994 28522
rect 19701 28464 19706 28520
rect 19762 28464 19994 28520
rect 19701 28462 19994 28464
rect 19701 28459 19767 28462
rect 17401 28386 17467 28389
rect 10918 28384 17467 28386
rect 10918 28328 17406 28384
rect 17462 28328 17467 28384
rect 10918 28326 17467 28328
rect 17401 28323 17467 28326
rect 10208 28320 10528 28321
rect 10208 28256 10216 28320
rect 10280 28256 10296 28320
rect 10360 28256 10376 28320
rect 10440 28256 10456 28320
rect 10520 28256 10528 28320
rect 10208 28255 10528 28256
rect 19472 28320 19792 28321
rect 19472 28256 19480 28320
rect 19544 28256 19560 28320
rect 19624 28256 19640 28320
rect 19704 28256 19720 28320
rect 19784 28256 19792 28320
rect 19472 28255 19792 28256
rect 10777 28250 10843 28253
rect 17125 28250 17191 28253
rect 10777 28248 17191 28250
rect 10777 28192 10782 28248
rect 10838 28192 17130 28248
rect 17186 28192 17191 28248
rect 10777 28190 17191 28192
rect 19934 28250 19994 28462
rect 22093 28520 22895 28522
rect 22093 28464 22098 28520
rect 22154 28464 22834 28520
rect 22890 28464 22895 28520
rect 29200 28508 30000 28748
rect 22093 28462 22895 28464
rect 22093 28459 22159 28462
rect 22829 28459 22895 28462
rect 28073 28386 28139 28389
rect 21774 28384 28139 28386
rect 21774 28328 28078 28384
rect 28134 28328 28139 28384
rect 21774 28326 28139 28328
rect 20713 28250 20779 28253
rect 19934 28248 20779 28250
rect 19934 28192 20718 28248
rect 20774 28192 20779 28248
rect 19934 28190 20779 28192
rect 10777 28187 10843 28190
rect 17125 28187 17191 28190
rect 20713 28187 20779 28190
rect 8293 28114 8359 28117
rect 11329 28114 11395 28117
rect 8293 28112 11395 28114
rect 0 27828 800 28068
rect 8293 28056 8298 28112
rect 8354 28056 11334 28112
rect 11390 28056 11395 28112
rect 8293 28054 11395 28056
rect 8293 28051 8359 28054
rect 11329 28051 11395 28054
rect 11789 28114 11855 28117
rect 12433 28114 12499 28117
rect 11789 28112 12499 28114
rect 11789 28056 11794 28112
rect 11850 28056 12438 28112
rect 12494 28056 12499 28112
rect 11789 28054 12499 28056
rect 11789 28051 11855 28054
rect 12433 28051 12499 28054
rect 12617 28114 12683 28117
rect 16849 28114 16915 28117
rect 12617 28112 16915 28114
rect 12617 28056 12622 28112
rect 12678 28056 16854 28112
rect 16910 28056 16915 28112
rect 12617 28054 16915 28056
rect 12617 28051 12683 28054
rect 16849 28051 16915 28054
rect 20437 28114 20503 28117
rect 21774 28114 21834 28326
rect 28073 28323 28139 28326
rect 23473 28250 23539 28253
rect 24526 28250 24532 28252
rect 23473 28248 24532 28250
rect 23473 28192 23478 28248
rect 23534 28192 24532 28248
rect 23473 28190 24532 28192
rect 23473 28187 23539 28190
rect 24526 28188 24532 28190
rect 24596 28188 24602 28252
rect 20437 28112 21834 28114
rect 20437 28056 20442 28112
rect 20498 28056 21834 28112
rect 20437 28054 21834 28056
rect 21909 28114 21975 28117
rect 24945 28114 25011 28117
rect 21909 28112 25011 28114
rect 21909 28056 21914 28112
rect 21970 28056 24950 28112
rect 25006 28056 25011 28112
rect 21909 28054 25011 28056
rect 20437 28051 20503 28054
rect 21909 28051 21975 28054
rect 24945 28051 25011 28054
rect 10041 27978 10107 27981
rect 10593 27978 10659 27981
rect 10041 27976 10659 27978
rect 10041 27920 10046 27976
rect 10102 27920 10598 27976
rect 10654 27920 10659 27976
rect 10041 27918 10659 27920
rect 10041 27915 10107 27918
rect 10593 27915 10659 27918
rect 10869 27978 10935 27981
rect 11605 27978 11671 27981
rect 10869 27976 11671 27978
rect 10869 27920 10874 27976
rect 10930 27920 11610 27976
rect 11666 27920 11671 27976
rect 10869 27918 11671 27920
rect 10869 27915 10935 27918
rect 11605 27915 11671 27918
rect 11881 27978 11947 27981
rect 12525 27978 12591 27981
rect 11881 27976 12591 27978
rect 11881 27920 11886 27976
rect 11942 27920 12530 27976
rect 12586 27920 12591 27976
rect 11881 27918 12591 27920
rect 11881 27915 11947 27918
rect 12525 27915 12591 27918
rect 12750 27916 12756 27980
rect 12820 27978 12826 27980
rect 15377 27978 15443 27981
rect 12820 27976 15443 27978
rect 12820 27920 15382 27976
rect 15438 27920 15443 27976
rect 12820 27918 15443 27920
rect 12820 27916 12826 27918
rect 15377 27915 15443 27918
rect 20713 27978 20779 27981
rect 22277 27978 22343 27981
rect 20713 27976 22343 27978
rect 20713 27920 20718 27976
rect 20774 27920 22282 27976
rect 22338 27920 22343 27976
rect 20713 27918 22343 27920
rect 20713 27915 20779 27918
rect 22277 27915 22343 27918
rect 10133 27842 10199 27845
rect 14181 27842 14247 27845
rect 10133 27840 14247 27842
rect 10133 27784 10138 27840
rect 10194 27784 14186 27840
rect 14242 27784 14247 27840
rect 10133 27782 14247 27784
rect 10133 27779 10199 27782
rect 14181 27779 14247 27782
rect 16205 27842 16271 27845
rect 19241 27842 19307 27845
rect 16205 27840 19307 27842
rect 16205 27784 16210 27840
rect 16266 27784 19246 27840
rect 19302 27784 19307 27840
rect 16205 27782 19307 27784
rect 16205 27779 16271 27782
rect 19241 27779 19307 27782
rect 21725 27842 21791 27845
rect 22185 27842 22251 27845
rect 22553 27842 22619 27845
rect 21725 27840 22619 27842
rect 21725 27784 21730 27840
rect 21786 27784 22190 27840
rect 22246 27784 22558 27840
rect 22614 27784 22619 27840
rect 29200 27828 30000 28068
rect 21725 27782 22619 27784
rect 21725 27779 21791 27782
rect 22185 27779 22251 27782
rect 22553 27779 22619 27782
rect 5576 27776 5896 27777
rect 5576 27712 5584 27776
rect 5648 27712 5664 27776
rect 5728 27712 5744 27776
rect 5808 27712 5824 27776
rect 5888 27712 5896 27776
rect 5576 27711 5896 27712
rect 14840 27776 15160 27777
rect 14840 27712 14848 27776
rect 14912 27712 14928 27776
rect 14992 27712 15008 27776
rect 15072 27712 15088 27776
rect 15152 27712 15160 27776
rect 14840 27711 15160 27712
rect 24104 27776 24424 27777
rect 24104 27712 24112 27776
rect 24176 27712 24192 27776
rect 24256 27712 24272 27776
rect 24336 27712 24352 27776
rect 24416 27712 24424 27776
rect 24104 27711 24424 27712
rect 9581 27706 9647 27709
rect 14457 27706 14523 27709
rect 9581 27704 14523 27706
rect 9581 27648 9586 27704
rect 9642 27648 14462 27704
rect 14518 27648 14523 27704
rect 9581 27646 14523 27648
rect 9581 27643 9647 27646
rect 14457 27643 14523 27646
rect 16849 27706 16915 27709
rect 18597 27706 18663 27709
rect 22001 27706 22067 27709
rect 16849 27704 22067 27706
rect 16849 27648 16854 27704
rect 16910 27648 18602 27704
rect 18658 27648 22006 27704
rect 22062 27648 22067 27704
rect 16849 27646 22067 27648
rect 16849 27643 16915 27646
rect 18597 27643 18663 27646
rect 22001 27643 22067 27646
rect 26182 27644 26188 27708
rect 26252 27706 26258 27708
rect 26325 27706 26391 27709
rect 26252 27704 26391 27706
rect 26252 27648 26330 27704
rect 26386 27648 26391 27704
rect 26252 27646 26391 27648
rect 26252 27644 26258 27646
rect 26325 27643 26391 27646
rect 8937 27570 9003 27573
rect 16430 27570 16436 27572
rect 8937 27568 16436 27570
rect 8937 27512 8942 27568
rect 8998 27512 16436 27568
rect 8937 27510 16436 27512
rect 8937 27507 9003 27510
rect 16430 27508 16436 27510
rect 16500 27508 16506 27572
rect 17309 27570 17375 27573
rect 18137 27570 18203 27573
rect 17309 27568 18203 27570
rect 17309 27512 17314 27568
rect 17370 27512 18142 27568
rect 18198 27512 18203 27568
rect 17309 27510 18203 27512
rect 17309 27507 17375 27510
rect 18137 27507 18203 27510
rect 21725 27570 21791 27573
rect 24485 27570 24551 27573
rect 21725 27568 24551 27570
rect 21725 27512 21730 27568
rect 21786 27512 24490 27568
rect 24546 27512 24551 27568
rect 21725 27510 24551 27512
rect 21725 27507 21791 27510
rect 24485 27507 24551 27510
rect 9489 27434 9555 27437
rect 13261 27434 13327 27437
rect 18873 27434 18939 27437
rect 26049 27434 26115 27437
rect 9489 27432 13186 27434
rect 0 27148 800 27388
rect 9489 27376 9494 27432
rect 9550 27376 13186 27432
rect 9489 27374 13186 27376
rect 9489 27371 9555 27374
rect 10961 27298 11027 27301
rect 12249 27298 12315 27301
rect 10961 27296 12315 27298
rect 10961 27240 10966 27296
rect 11022 27240 12254 27296
rect 12310 27240 12315 27296
rect 10961 27238 12315 27240
rect 10961 27235 11027 27238
rect 12249 27235 12315 27238
rect 12433 27298 12499 27301
rect 12985 27298 13051 27301
rect 12433 27296 13051 27298
rect 12433 27240 12438 27296
rect 12494 27240 12990 27296
rect 13046 27240 13051 27296
rect 12433 27238 13051 27240
rect 13126 27298 13186 27374
rect 13261 27432 18939 27434
rect 13261 27376 13266 27432
rect 13322 27376 18878 27432
rect 18934 27376 18939 27432
rect 13261 27374 18939 27376
rect 13261 27371 13327 27374
rect 18873 27371 18939 27374
rect 19290 27432 26115 27434
rect 19290 27376 26054 27432
rect 26110 27376 26115 27432
rect 19290 27374 26115 27376
rect 13445 27298 13511 27301
rect 13126 27296 13511 27298
rect 13126 27240 13450 27296
rect 13506 27240 13511 27296
rect 13126 27238 13511 27240
rect 12433 27235 12499 27238
rect 12985 27235 13051 27238
rect 13445 27235 13511 27238
rect 13629 27298 13695 27301
rect 17401 27298 17467 27301
rect 13629 27296 17467 27298
rect 13629 27240 13634 27296
rect 13690 27240 17406 27296
rect 17462 27240 17467 27296
rect 13629 27238 17467 27240
rect 13629 27235 13695 27238
rect 17401 27235 17467 27238
rect 17953 27298 18019 27301
rect 18413 27298 18479 27301
rect 17953 27296 18479 27298
rect 17953 27240 17958 27296
rect 18014 27240 18418 27296
rect 18474 27240 18479 27296
rect 17953 27238 18479 27240
rect 17953 27235 18019 27238
rect 18413 27235 18479 27238
rect 10208 27232 10528 27233
rect 10208 27168 10216 27232
rect 10280 27168 10296 27232
rect 10360 27168 10376 27232
rect 10440 27168 10456 27232
rect 10520 27168 10528 27232
rect 10208 27167 10528 27168
rect 11697 27162 11763 27165
rect 12750 27162 12756 27164
rect 11697 27160 12756 27162
rect 11697 27104 11702 27160
rect 11758 27104 12756 27160
rect 11697 27102 12756 27104
rect 11697 27099 11763 27102
rect 12750 27100 12756 27102
rect 12820 27100 12826 27164
rect 12934 27100 12940 27164
rect 13004 27162 13010 27164
rect 19290 27162 19350 27374
rect 26049 27371 26115 27374
rect 23105 27298 23171 27301
rect 25589 27298 25655 27301
rect 23105 27296 25655 27298
rect 23105 27240 23110 27296
rect 23166 27240 25594 27296
rect 25650 27240 25655 27296
rect 23105 27238 25655 27240
rect 23105 27235 23171 27238
rect 25589 27235 25655 27238
rect 28165 27298 28231 27301
rect 29200 27298 30000 27388
rect 28165 27296 30000 27298
rect 28165 27240 28170 27296
rect 28226 27240 30000 27296
rect 28165 27238 30000 27240
rect 28165 27235 28231 27238
rect 19472 27232 19792 27233
rect 19472 27168 19480 27232
rect 19544 27168 19560 27232
rect 19624 27168 19640 27232
rect 19704 27168 19720 27232
rect 19784 27168 19792 27232
rect 19472 27167 19792 27168
rect 13004 27102 19350 27162
rect 29200 27148 30000 27238
rect 13004 27100 13010 27102
rect 10777 27026 10843 27029
rect 24761 27026 24827 27029
rect 10777 27024 24827 27026
rect 10777 26968 10782 27024
rect 10838 26968 24766 27024
rect 24822 26968 24827 27024
rect 10777 26966 24827 26968
rect 10777 26963 10843 26966
rect 24761 26963 24827 26966
rect 9673 26890 9739 26893
rect 26325 26890 26391 26893
rect 9673 26888 26391 26890
rect 9673 26832 9678 26888
rect 9734 26832 26330 26888
rect 26386 26832 26391 26888
rect 9673 26830 26391 26832
rect 9673 26827 9739 26830
rect 26325 26827 26391 26830
rect 11789 26754 11855 26757
rect 15653 26754 15719 26757
rect 18137 26754 18203 26757
rect 11789 26752 13876 26754
rect 0 26468 800 26708
rect 11789 26696 11794 26752
rect 11850 26696 13876 26752
rect 11789 26694 13876 26696
rect 11789 26691 11855 26694
rect 5576 26688 5896 26689
rect 5576 26624 5584 26688
rect 5648 26624 5664 26688
rect 5728 26624 5744 26688
rect 5808 26624 5824 26688
rect 5888 26624 5896 26688
rect 5576 26623 5896 26624
rect 10225 26618 10291 26621
rect 10225 26616 13186 26618
rect 10225 26560 10230 26616
rect 10286 26560 13186 26616
rect 10225 26558 13186 26560
rect 10225 26555 10291 26558
rect 11329 26482 11395 26485
rect 12617 26482 12683 26485
rect 11329 26480 12683 26482
rect 11329 26424 11334 26480
rect 11390 26424 12622 26480
rect 12678 26424 12683 26480
rect 11329 26422 12683 26424
rect 11329 26419 11395 26422
rect 12617 26419 12683 26422
rect 9029 26346 9095 26349
rect 12934 26346 12940 26348
rect 9029 26344 12940 26346
rect 9029 26288 9034 26344
rect 9090 26288 12940 26344
rect 9029 26286 12940 26288
rect 9029 26283 9095 26286
rect 12934 26284 12940 26286
rect 13004 26284 13010 26348
rect 13126 26346 13186 26558
rect 13816 26482 13876 26694
rect 15653 26752 18203 26754
rect 15653 26696 15658 26752
rect 15714 26696 18142 26752
rect 18198 26696 18203 26752
rect 15653 26694 18203 26696
rect 15653 26691 15719 26694
rect 18137 26691 18203 26694
rect 19057 26754 19123 26757
rect 21633 26754 21699 26757
rect 19057 26752 21699 26754
rect 19057 26696 19062 26752
rect 19118 26696 21638 26752
rect 21694 26696 21699 26752
rect 19057 26694 21699 26696
rect 19057 26691 19123 26694
rect 21633 26691 21699 26694
rect 14840 26688 15160 26689
rect 14840 26624 14848 26688
rect 14912 26624 14928 26688
rect 14992 26624 15008 26688
rect 15072 26624 15088 26688
rect 15152 26624 15160 26688
rect 14840 26623 15160 26624
rect 24104 26688 24424 26689
rect 24104 26624 24112 26688
rect 24176 26624 24192 26688
rect 24256 26624 24272 26688
rect 24336 26624 24352 26688
rect 24416 26624 24424 26688
rect 24104 26623 24424 26624
rect 16941 26618 17007 26621
rect 18413 26618 18479 26621
rect 20253 26618 20319 26621
rect 16941 26616 20319 26618
rect 16941 26560 16946 26616
rect 17002 26560 18418 26616
rect 18474 26560 20258 26616
rect 20314 26560 20319 26616
rect 16941 26558 20319 26560
rect 16941 26555 17007 26558
rect 18413 26555 18479 26558
rect 20253 26555 20319 26558
rect 28165 26618 28231 26621
rect 29200 26618 30000 26708
rect 28165 26616 30000 26618
rect 28165 26560 28170 26616
rect 28226 26560 30000 26616
rect 28165 26558 30000 26560
rect 28165 26555 28231 26558
rect 18873 26482 18939 26485
rect 20161 26484 20227 26485
rect 13816 26480 18939 26482
rect 13816 26424 18878 26480
rect 18934 26424 18939 26480
rect 13816 26422 18939 26424
rect 18873 26419 18939 26422
rect 20110 26420 20116 26484
rect 20180 26482 20227 26484
rect 27429 26482 27495 26485
rect 20180 26480 27495 26482
rect 20222 26424 27434 26480
rect 27490 26424 27495 26480
rect 29200 26468 30000 26558
rect 20180 26422 27495 26424
rect 20180 26420 20227 26422
rect 20161 26419 20227 26420
rect 25408 26349 25468 26422
rect 27429 26419 27495 26422
rect 15377 26346 15443 26349
rect 13126 26344 15443 26346
rect 13126 26288 15382 26344
rect 15438 26288 15443 26344
rect 13126 26286 15443 26288
rect 15377 26283 15443 26286
rect 15561 26346 15627 26349
rect 16389 26346 16455 26349
rect 16573 26348 16639 26349
rect 16573 26346 16620 26348
rect 15561 26344 16455 26346
rect 15561 26288 15566 26344
rect 15622 26288 16394 26344
rect 16450 26288 16455 26344
rect 15561 26286 16455 26288
rect 16528 26344 16620 26346
rect 16528 26288 16578 26344
rect 16528 26286 16620 26288
rect 15561 26283 15627 26286
rect 16389 26283 16455 26286
rect 16573 26284 16620 26286
rect 16684 26284 16690 26348
rect 19701 26346 19767 26349
rect 23565 26346 23631 26349
rect 19701 26344 23631 26346
rect 19701 26288 19706 26344
rect 19762 26288 23570 26344
rect 23626 26288 23631 26344
rect 19701 26286 23631 26288
rect 16573 26283 16639 26284
rect 19701 26283 19767 26286
rect 23565 26283 23631 26286
rect 25405 26344 25471 26349
rect 25405 26288 25410 26344
rect 25466 26288 25471 26344
rect 25405 26283 25471 26288
rect 12065 26210 12131 26213
rect 17953 26210 18019 26213
rect 12065 26208 18019 26210
rect 12065 26152 12070 26208
rect 12126 26152 17958 26208
rect 18014 26152 18019 26208
rect 12065 26150 18019 26152
rect 12065 26147 12131 26150
rect 17953 26147 18019 26150
rect 10208 26144 10528 26145
rect 10208 26080 10216 26144
rect 10280 26080 10296 26144
rect 10360 26080 10376 26144
rect 10440 26080 10456 26144
rect 10520 26080 10528 26144
rect 10208 26079 10528 26080
rect 19472 26144 19792 26145
rect 19472 26080 19480 26144
rect 19544 26080 19560 26144
rect 19624 26080 19640 26144
rect 19704 26080 19720 26144
rect 19784 26080 19792 26144
rect 19472 26079 19792 26080
rect 10685 26074 10751 26077
rect 16573 26074 16639 26077
rect 10685 26072 16639 26074
rect 0 25788 800 26028
rect 10685 26016 10690 26072
rect 10746 26016 16578 26072
rect 16634 26016 16639 26072
rect 10685 26014 16639 26016
rect 10685 26011 10751 26014
rect 16573 26011 16639 26014
rect 20069 26074 20135 26077
rect 23473 26074 23539 26077
rect 20069 26072 23539 26074
rect 20069 26016 20074 26072
rect 20130 26016 23478 26072
rect 23534 26016 23539 26072
rect 20069 26014 23539 26016
rect 20069 26011 20135 26014
rect 23473 26011 23539 26014
rect 11053 25938 11119 25941
rect 12801 25938 12867 25941
rect 13813 25938 13879 25941
rect 11053 25936 13879 25938
rect 11053 25880 11058 25936
rect 11114 25880 12806 25936
rect 12862 25880 13818 25936
rect 13874 25880 13879 25936
rect 11053 25878 13879 25880
rect 11053 25875 11119 25878
rect 12801 25875 12867 25878
rect 13813 25875 13879 25878
rect 14222 25876 14228 25940
rect 14292 25938 14298 25940
rect 21081 25938 21147 25941
rect 26417 25938 26483 25941
rect 14292 25936 21147 25938
rect 14292 25880 21086 25936
rect 21142 25880 21147 25936
rect 14292 25878 21147 25880
rect 14292 25876 14298 25878
rect 21081 25875 21147 25878
rect 22326 25936 26483 25938
rect 22326 25880 26422 25936
rect 26478 25880 26483 25936
rect 22326 25878 26483 25880
rect 11145 25802 11211 25805
rect 14549 25802 14615 25805
rect 11145 25800 14615 25802
rect 11145 25744 11150 25800
rect 11206 25744 14554 25800
rect 14610 25744 14615 25800
rect 11145 25742 14615 25744
rect 11145 25739 11211 25742
rect 14549 25739 14615 25742
rect 15469 25802 15535 25805
rect 19149 25802 19215 25805
rect 15469 25800 19215 25802
rect 15469 25744 15474 25800
rect 15530 25744 19154 25800
rect 19210 25744 19215 25800
rect 15469 25742 19215 25744
rect 15469 25739 15535 25742
rect 19149 25739 19215 25742
rect 10777 25666 10843 25669
rect 14641 25666 14707 25669
rect 10777 25664 14707 25666
rect 10777 25608 10782 25664
rect 10838 25608 14646 25664
rect 14702 25608 14707 25664
rect 10777 25606 14707 25608
rect 10777 25603 10843 25606
rect 14641 25603 14707 25606
rect 15285 25666 15351 25669
rect 16021 25666 16087 25669
rect 15285 25664 16087 25666
rect 15285 25608 15290 25664
rect 15346 25608 16026 25664
rect 16082 25608 16087 25664
rect 15285 25606 16087 25608
rect 15285 25603 15351 25606
rect 16021 25603 16087 25606
rect 17217 25666 17283 25669
rect 19926 25666 19932 25668
rect 17217 25664 19932 25666
rect 17217 25608 17222 25664
rect 17278 25608 19932 25664
rect 17217 25606 19932 25608
rect 17217 25603 17283 25606
rect 19926 25604 19932 25606
rect 19996 25666 20002 25668
rect 20069 25666 20135 25669
rect 22326 25666 22386 25878
rect 26417 25875 26483 25878
rect 28165 25938 28231 25941
rect 29200 25938 30000 26028
rect 28165 25936 30000 25938
rect 28165 25880 28170 25936
rect 28226 25880 30000 25936
rect 28165 25878 30000 25880
rect 28165 25875 28231 25878
rect 22461 25802 22527 25805
rect 22461 25800 22754 25802
rect 22461 25744 22466 25800
rect 22522 25744 22754 25800
rect 29200 25788 30000 25878
rect 22461 25742 22754 25744
rect 22461 25739 22527 25742
rect 19996 25664 22386 25666
rect 19996 25608 20074 25664
rect 20130 25608 22386 25664
rect 19996 25606 22386 25608
rect 22694 25666 22754 25742
rect 22921 25666 22987 25669
rect 22694 25664 22987 25666
rect 22694 25608 22926 25664
rect 22982 25608 22987 25664
rect 22694 25606 22987 25608
rect 19996 25604 20002 25606
rect 20069 25603 20135 25606
rect 22921 25603 22987 25606
rect 5576 25600 5896 25601
rect 5576 25536 5584 25600
rect 5648 25536 5664 25600
rect 5728 25536 5744 25600
rect 5808 25536 5824 25600
rect 5888 25536 5896 25600
rect 5576 25535 5896 25536
rect 14840 25600 15160 25601
rect 14840 25536 14848 25600
rect 14912 25536 14928 25600
rect 14992 25536 15008 25600
rect 15072 25536 15088 25600
rect 15152 25536 15160 25600
rect 14840 25535 15160 25536
rect 24104 25600 24424 25601
rect 24104 25536 24112 25600
rect 24176 25536 24192 25600
rect 24256 25536 24272 25600
rect 24336 25536 24352 25600
rect 24416 25536 24424 25600
rect 24104 25535 24424 25536
rect 11053 25530 11119 25533
rect 12525 25530 12591 25533
rect 16982 25530 16988 25532
rect 11053 25528 12591 25530
rect 11053 25472 11058 25528
rect 11114 25472 12530 25528
rect 12586 25472 12591 25528
rect 11053 25470 12591 25472
rect 11053 25467 11119 25470
rect 12525 25467 12591 25470
rect 15288 25470 16988 25530
rect 10593 25394 10659 25397
rect 15288 25394 15348 25470
rect 16982 25468 16988 25470
rect 17052 25468 17058 25532
rect 10593 25392 15348 25394
rect 0 25108 800 25348
rect 10593 25336 10598 25392
rect 10654 25336 15348 25392
rect 10593 25334 15348 25336
rect 15561 25394 15627 25397
rect 19149 25394 19215 25397
rect 15561 25392 19215 25394
rect 15561 25336 15566 25392
rect 15622 25336 19154 25392
rect 19210 25336 19215 25392
rect 15561 25334 19215 25336
rect 10593 25331 10659 25334
rect 15561 25331 15627 25334
rect 19149 25331 19215 25334
rect 19885 25394 19951 25397
rect 23657 25396 23723 25397
rect 23606 25394 23612 25396
rect 19885 25392 23612 25394
rect 23676 25392 23723 25396
rect 19885 25336 19890 25392
rect 19946 25336 23612 25392
rect 23718 25336 23723 25392
rect 19885 25334 23612 25336
rect 19885 25331 19951 25334
rect 23606 25332 23612 25334
rect 23676 25332 23723 25336
rect 23657 25331 23723 25332
rect 10777 25258 10843 25261
rect 15745 25258 15811 25261
rect 10777 25256 15811 25258
rect 10777 25200 10782 25256
rect 10838 25200 15750 25256
rect 15806 25200 15811 25256
rect 10777 25198 15811 25200
rect 10777 25195 10843 25198
rect 15745 25195 15811 25198
rect 18638 25196 18644 25260
rect 18708 25258 18714 25260
rect 26325 25258 26391 25261
rect 18708 25256 26391 25258
rect 18708 25200 26330 25256
rect 26386 25200 26391 25256
rect 18708 25198 26391 25200
rect 18708 25196 18714 25198
rect 26325 25195 26391 25198
rect 28717 25258 28783 25261
rect 29200 25258 30000 25348
rect 28717 25256 30000 25258
rect 28717 25200 28722 25256
rect 28778 25200 30000 25256
rect 28717 25198 30000 25200
rect 28717 25195 28783 25198
rect 12617 25122 12683 25125
rect 16941 25122 17007 25125
rect 12617 25120 17007 25122
rect 12617 25064 12622 25120
rect 12678 25064 16946 25120
rect 17002 25064 17007 25120
rect 12617 25062 17007 25064
rect 12617 25059 12683 25062
rect 16941 25059 17007 25062
rect 19885 25122 19951 25125
rect 24526 25122 24532 25124
rect 19885 25120 24532 25122
rect 19885 25064 19890 25120
rect 19946 25064 24532 25120
rect 19885 25062 24532 25064
rect 19885 25059 19951 25062
rect 24526 25060 24532 25062
rect 24596 25060 24602 25124
rect 29200 25108 30000 25198
rect 10208 25056 10528 25057
rect 10208 24992 10216 25056
rect 10280 24992 10296 25056
rect 10360 24992 10376 25056
rect 10440 24992 10456 25056
rect 10520 24992 10528 25056
rect 10208 24991 10528 24992
rect 19472 25056 19792 25057
rect 19472 24992 19480 25056
rect 19544 24992 19560 25056
rect 19624 24992 19640 25056
rect 19704 24992 19720 25056
rect 19784 24992 19792 25056
rect 19472 24991 19792 24992
rect 11053 24986 11119 24989
rect 12985 24986 13051 24989
rect 11053 24984 13051 24986
rect 11053 24928 11058 24984
rect 11114 24928 12990 24984
rect 13046 24928 13051 24984
rect 11053 24926 13051 24928
rect 11053 24923 11119 24926
rect 12985 24923 13051 24926
rect 13169 24986 13235 24989
rect 17125 24986 17191 24989
rect 13169 24984 17191 24986
rect 13169 24928 13174 24984
rect 13230 24928 17130 24984
rect 17186 24928 17191 24984
rect 13169 24926 17191 24928
rect 13169 24923 13235 24926
rect 17125 24923 17191 24926
rect 21633 24986 21699 24989
rect 26509 24986 26575 24989
rect 21633 24984 26575 24986
rect 21633 24928 21638 24984
rect 21694 24928 26514 24984
rect 26570 24928 26575 24984
rect 21633 24926 26575 24928
rect 21633 24923 21699 24926
rect 26509 24923 26575 24926
rect 7833 24850 7899 24853
rect 13670 24850 13676 24852
rect 7833 24848 13676 24850
rect 7833 24792 7838 24848
rect 7894 24792 13676 24848
rect 7833 24790 13676 24792
rect 7833 24787 7899 24790
rect 13670 24788 13676 24790
rect 13740 24788 13746 24852
rect 13997 24850 14063 24853
rect 16113 24850 16179 24853
rect 13997 24848 16179 24850
rect 13997 24792 14002 24848
rect 14058 24792 16118 24848
rect 16174 24792 16179 24848
rect 13997 24790 16179 24792
rect 13997 24787 14063 24790
rect 16113 24787 16179 24790
rect 18137 24850 18203 24853
rect 20253 24850 20319 24853
rect 18137 24848 20319 24850
rect 18137 24792 18142 24848
rect 18198 24792 20258 24848
rect 20314 24792 20319 24848
rect 18137 24790 20319 24792
rect 18137 24787 18203 24790
rect 20253 24787 20319 24790
rect 20437 24850 20503 24853
rect 26141 24850 26207 24853
rect 20437 24848 26207 24850
rect 20437 24792 20442 24848
rect 20498 24792 26146 24848
rect 26202 24792 26207 24848
rect 20437 24790 26207 24792
rect 20437 24787 20503 24790
rect 26141 24787 26207 24790
rect 12065 24714 12131 24717
rect 14181 24714 14247 24717
rect 12065 24712 14247 24714
rect 12065 24656 12070 24712
rect 12126 24656 14186 24712
rect 14242 24656 14247 24712
rect 12065 24654 14247 24656
rect 12065 24651 12131 24654
rect 14181 24651 14247 24654
rect 14733 24714 14799 24717
rect 23013 24714 23079 24717
rect 23657 24714 23723 24717
rect 14733 24712 23723 24714
rect 14733 24656 14738 24712
rect 14794 24656 23018 24712
rect 23074 24656 23662 24712
rect 23718 24656 23723 24712
rect 14733 24654 23723 24656
rect 14733 24651 14799 24654
rect 23013 24651 23079 24654
rect 23657 24651 23723 24654
rect 11513 24578 11579 24581
rect 14641 24578 14707 24581
rect 11513 24576 14707 24578
rect 11513 24520 11518 24576
rect 11574 24520 14646 24576
rect 14702 24520 14707 24576
rect 11513 24518 14707 24520
rect 11513 24515 11579 24518
rect 14641 24515 14707 24518
rect 15377 24578 15443 24581
rect 15837 24578 15903 24581
rect 15377 24576 15903 24578
rect 15377 24520 15382 24576
rect 15438 24520 15842 24576
rect 15898 24520 15903 24576
rect 15377 24518 15903 24520
rect 15377 24515 15443 24518
rect 15837 24515 15903 24518
rect 16021 24578 16087 24581
rect 20989 24578 21055 24581
rect 16021 24576 21055 24578
rect 16021 24520 16026 24576
rect 16082 24520 20994 24576
rect 21050 24520 21055 24576
rect 16021 24518 21055 24520
rect 16021 24515 16087 24518
rect 20989 24515 21055 24518
rect 28165 24578 28231 24581
rect 29200 24578 30000 24668
rect 28165 24576 30000 24578
rect 28165 24520 28170 24576
rect 28226 24520 30000 24576
rect 28165 24518 30000 24520
rect 28165 24515 28231 24518
rect 5576 24512 5896 24513
rect 5576 24448 5584 24512
rect 5648 24448 5664 24512
rect 5728 24448 5744 24512
rect 5808 24448 5824 24512
rect 5888 24448 5896 24512
rect 5576 24447 5896 24448
rect 14840 24512 15160 24513
rect 14840 24448 14848 24512
rect 14912 24448 14928 24512
rect 14992 24448 15008 24512
rect 15072 24448 15088 24512
rect 15152 24448 15160 24512
rect 14840 24447 15160 24448
rect 24104 24512 24424 24513
rect 24104 24448 24112 24512
rect 24176 24448 24192 24512
rect 24256 24448 24272 24512
rect 24336 24448 24352 24512
rect 24416 24448 24424 24512
rect 24104 24447 24424 24448
rect 13077 24442 13143 24445
rect 14641 24442 14707 24445
rect 13077 24440 14707 24442
rect 13077 24384 13082 24440
rect 13138 24384 14646 24440
rect 14702 24384 14707 24440
rect 13077 24382 14707 24384
rect 13077 24379 13143 24382
rect 14641 24379 14707 24382
rect 15285 24442 15351 24445
rect 15929 24442 15995 24445
rect 15285 24440 15995 24442
rect 15285 24384 15290 24440
rect 15346 24384 15934 24440
rect 15990 24384 15995 24440
rect 15285 24382 15995 24384
rect 15285 24379 15351 24382
rect 15929 24379 15995 24382
rect 16113 24442 16179 24445
rect 19333 24442 19399 24445
rect 16113 24440 19399 24442
rect 16113 24384 16118 24440
rect 16174 24384 19338 24440
rect 19394 24384 19399 24440
rect 29200 24428 30000 24518
rect 16113 24382 19399 24384
rect 16113 24379 16179 24382
rect 19333 24379 19399 24382
rect 12893 24306 12959 24309
rect 20621 24306 20687 24309
rect 12893 24304 20687 24306
rect 12893 24248 12898 24304
rect 12954 24248 20626 24304
rect 20682 24248 20687 24304
rect 12893 24246 20687 24248
rect 12893 24243 12959 24246
rect 20621 24243 20687 24246
rect 20805 24306 20871 24309
rect 25221 24306 25287 24309
rect 20805 24304 25287 24306
rect 20805 24248 20810 24304
rect 20866 24248 25226 24304
rect 25282 24248 25287 24304
rect 20805 24246 25287 24248
rect 20805 24243 20871 24246
rect 25221 24243 25287 24246
rect 13261 24170 13327 24173
rect 14222 24170 14228 24172
rect 13261 24168 14228 24170
rect 13261 24112 13266 24168
rect 13322 24112 14228 24168
rect 13261 24110 14228 24112
rect 13261 24107 13327 24110
rect 14222 24108 14228 24110
rect 14292 24108 14298 24172
rect 14365 24170 14431 24173
rect 22185 24170 22251 24173
rect 24945 24170 25011 24173
rect 14365 24168 25011 24170
rect 14365 24112 14370 24168
rect 14426 24112 22190 24168
rect 22246 24112 24950 24168
rect 25006 24112 25011 24168
rect 14365 24110 25011 24112
rect 14365 24107 14431 24110
rect 22185 24107 22251 24110
rect 24945 24107 25011 24110
rect 10685 24034 10751 24037
rect 18229 24034 18295 24037
rect 10685 24032 18295 24034
rect 0 23748 800 23988
rect 10685 23976 10690 24032
rect 10746 23976 18234 24032
rect 18290 23976 18295 24032
rect 10685 23974 18295 23976
rect 10685 23971 10751 23974
rect 18229 23971 18295 23974
rect 18413 24034 18479 24037
rect 18781 24034 18847 24037
rect 23473 24034 23539 24037
rect 18413 24032 18847 24034
rect 18413 23976 18418 24032
rect 18474 23976 18786 24032
rect 18842 23976 18847 24032
rect 18413 23974 18847 23976
rect 18413 23971 18479 23974
rect 18781 23971 18847 23974
rect 21774 24032 23539 24034
rect 21774 23976 23478 24032
rect 23534 23976 23539 24032
rect 21774 23974 23539 23976
rect 10208 23968 10528 23969
rect 10208 23904 10216 23968
rect 10280 23904 10296 23968
rect 10360 23904 10376 23968
rect 10440 23904 10456 23968
rect 10520 23904 10528 23968
rect 10208 23903 10528 23904
rect 19472 23968 19792 23969
rect 19472 23904 19480 23968
rect 19544 23904 19560 23968
rect 19624 23904 19640 23968
rect 19704 23904 19720 23968
rect 19784 23904 19792 23968
rect 19472 23903 19792 23904
rect 10777 23898 10843 23901
rect 15009 23898 15075 23901
rect 10777 23896 15075 23898
rect 10777 23840 10782 23896
rect 10838 23840 15014 23896
rect 15070 23840 15075 23896
rect 10777 23838 15075 23840
rect 10777 23835 10843 23838
rect 15009 23835 15075 23838
rect 15193 23898 15259 23901
rect 15510 23898 15516 23900
rect 15193 23896 15516 23898
rect 15193 23840 15198 23896
rect 15254 23840 15516 23896
rect 15193 23838 15516 23840
rect 15193 23835 15259 23838
rect 15510 23836 15516 23838
rect 15580 23836 15586 23900
rect 15837 23898 15903 23901
rect 18781 23898 18847 23901
rect 15837 23896 18847 23898
rect 15837 23840 15842 23896
rect 15898 23840 18786 23896
rect 18842 23840 18847 23896
rect 15837 23838 18847 23840
rect 15837 23835 15903 23838
rect 18781 23835 18847 23838
rect 11421 23762 11487 23765
rect 12433 23762 12499 23765
rect 14733 23762 14799 23765
rect 11421 23760 14799 23762
rect 11421 23704 11426 23760
rect 11482 23704 12438 23760
rect 12494 23704 14738 23760
rect 14794 23704 14799 23760
rect 11421 23702 14799 23704
rect 11421 23699 11487 23702
rect 12433 23699 12499 23702
rect 14733 23699 14799 23702
rect 14917 23762 14983 23765
rect 21774 23762 21834 23974
rect 23473 23971 23539 23974
rect 24301 24034 24367 24037
rect 24853 24034 24919 24037
rect 24301 24032 24919 24034
rect 24301 23976 24306 24032
rect 24362 23976 24858 24032
rect 24914 23976 24919 24032
rect 24301 23974 24919 23976
rect 24301 23971 24367 23974
rect 24853 23971 24919 23974
rect 22645 23898 22711 23901
rect 24669 23898 24735 23901
rect 22645 23896 24735 23898
rect 22645 23840 22650 23896
rect 22706 23840 24674 23896
rect 24730 23840 24735 23896
rect 22645 23838 24735 23840
rect 22645 23835 22711 23838
rect 24669 23835 24735 23838
rect 14917 23760 21834 23762
rect 14917 23704 14922 23760
rect 14978 23704 21834 23760
rect 14917 23702 21834 23704
rect 21909 23762 21975 23765
rect 28625 23762 28691 23765
rect 21909 23760 28691 23762
rect 21909 23704 21914 23760
rect 21970 23704 28630 23760
rect 28686 23704 28691 23760
rect 29200 23748 30000 23988
rect 21909 23702 28691 23704
rect 14917 23699 14983 23702
rect 21909 23699 21975 23702
rect 28625 23699 28691 23702
rect 13905 23626 13971 23629
rect 13905 23624 15348 23626
rect 13905 23568 13910 23624
rect 13966 23568 15348 23624
rect 13905 23566 15348 23568
rect 13905 23563 13971 23566
rect 7230 23428 7236 23492
rect 7300 23490 7306 23492
rect 14406 23490 14412 23492
rect 7300 23430 14412 23490
rect 7300 23428 7306 23430
rect 14406 23428 14412 23430
rect 14476 23428 14482 23492
rect 15288 23490 15348 23566
rect 15510 23564 15516 23628
rect 15580 23626 15586 23628
rect 22369 23626 22435 23629
rect 15580 23624 22435 23626
rect 15580 23568 22374 23624
rect 22430 23568 22435 23624
rect 15580 23566 22435 23568
rect 15580 23564 15586 23566
rect 22369 23563 22435 23566
rect 22645 23490 22711 23493
rect 15288 23488 22711 23490
rect 15288 23432 22650 23488
rect 22706 23432 22711 23488
rect 15288 23430 22711 23432
rect 22645 23427 22711 23430
rect 26325 23492 26391 23493
rect 26325 23488 26372 23492
rect 26436 23490 26442 23492
rect 26325 23432 26330 23488
rect 26325 23428 26372 23432
rect 26436 23430 26482 23490
rect 26436 23428 26442 23430
rect 26325 23427 26391 23428
rect 5576 23424 5896 23425
rect 5576 23360 5584 23424
rect 5648 23360 5664 23424
rect 5728 23360 5744 23424
rect 5808 23360 5824 23424
rect 5888 23360 5896 23424
rect 5576 23359 5896 23360
rect 14840 23424 15160 23425
rect 14840 23360 14848 23424
rect 14912 23360 14928 23424
rect 14992 23360 15008 23424
rect 15072 23360 15088 23424
rect 15152 23360 15160 23424
rect 14840 23359 15160 23360
rect 24104 23424 24424 23425
rect 24104 23360 24112 23424
rect 24176 23360 24192 23424
rect 24256 23360 24272 23424
rect 24336 23360 24352 23424
rect 24416 23360 24424 23424
rect 24104 23359 24424 23360
rect 10317 23354 10383 23357
rect 14641 23354 14707 23357
rect 10317 23352 14707 23354
rect 0 23218 800 23308
rect 10317 23296 10322 23352
rect 10378 23296 14646 23352
rect 14702 23296 14707 23352
rect 10317 23294 14707 23296
rect 10317 23291 10383 23294
rect 14641 23291 14707 23294
rect 15273 23354 15339 23357
rect 16941 23354 17007 23357
rect 15273 23352 17007 23354
rect 15273 23296 15278 23352
rect 15334 23296 16946 23352
rect 17002 23296 17007 23352
rect 15273 23294 17007 23296
rect 15273 23291 15339 23294
rect 16941 23291 17007 23294
rect 18321 23354 18387 23357
rect 19701 23354 19767 23357
rect 18321 23352 19767 23354
rect 18321 23296 18326 23352
rect 18382 23296 19706 23352
rect 19762 23296 19767 23352
rect 18321 23294 19767 23296
rect 18321 23291 18387 23294
rect 19701 23291 19767 23294
rect 21633 23354 21699 23357
rect 22553 23354 22619 23357
rect 21633 23352 22619 23354
rect 21633 23296 21638 23352
rect 21694 23296 22558 23352
rect 22614 23296 22619 23352
rect 21633 23294 22619 23296
rect 21633 23291 21699 23294
rect 22553 23291 22619 23294
rect 2773 23218 2839 23221
rect 0 23216 2839 23218
rect 0 23160 2778 23216
rect 2834 23160 2839 23216
rect 0 23158 2839 23160
rect 0 23068 800 23158
rect 2773 23155 2839 23158
rect 10225 23218 10291 23221
rect 14181 23218 14247 23221
rect 10225 23216 14247 23218
rect 10225 23160 10230 23216
rect 10286 23160 14186 23216
rect 14242 23160 14247 23216
rect 10225 23158 14247 23160
rect 10225 23155 10291 23158
rect 14181 23155 14247 23158
rect 14457 23218 14523 23221
rect 16941 23218 17007 23221
rect 18137 23218 18203 23221
rect 14457 23216 18203 23218
rect 14457 23160 14462 23216
rect 14518 23160 16946 23216
rect 17002 23160 18142 23216
rect 18198 23160 18203 23216
rect 14457 23158 18203 23160
rect 14457 23155 14523 23158
rect 16941 23155 17007 23158
rect 18137 23155 18203 23158
rect 18321 23218 18387 23221
rect 18597 23218 18663 23221
rect 18321 23216 18663 23218
rect 18321 23160 18326 23216
rect 18382 23160 18602 23216
rect 18658 23160 18663 23216
rect 18321 23158 18663 23160
rect 18321 23155 18387 23158
rect 18597 23155 18663 23158
rect 19793 23218 19859 23221
rect 20805 23218 20871 23221
rect 19793 23216 20871 23218
rect 19793 23160 19798 23216
rect 19854 23160 20810 23216
rect 20866 23160 20871 23216
rect 19793 23158 20871 23160
rect 19793 23155 19859 23158
rect 20805 23155 20871 23158
rect 12157 23082 12223 23085
rect 12617 23082 12683 23085
rect 21081 23082 21147 23085
rect 12157 23080 21147 23082
rect 12157 23024 12162 23080
rect 12218 23024 12622 23080
rect 12678 23024 21086 23080
rect 21142 23024 21147 23080
rect 12157 23022 21147 23024
rect 22556 23082 22616 23291
rect 25681 23218 25747 23221
rect 29200 23218 30000 23308
rect 25681 23216 30000 23218
rect 25681 23160 25686 23216
rect 25742 23160 30000 23216
rect 25681 23158 30000 23160
rect 25681 23155 25747 23158
rect 23657 23082 23723 23085
rect 22556 23080 23723 23082
rect 22556 23024 23662 23080
rect 23718 23024 23723 23080
rect 22556 23022 23723 23024
rect 12157 23019 12223 23022
rect 12617 23019 12683 23022
rect 21081 23019 21147 23022
rect 23657 23019 23723 23022
rect 24526 23020 24532 23084
rect 24596 23082 24602 23084
rect 24669 23082 24735 23085
rect 24596 23080 24735 23082
rect 24596 23024 24674 23080
rect 24730 23024 24735 23080
rect 29200 23068 30000 23158
rect 24596 23022 24735 23024
rect 24596 23020 24602 23022
rect 24669 23019 24735 23022
rect 14181 22946 14247 22949
rect 16757 22946 16823 22949
rect 14181 22944 16823 22946
rect 14181 22888 14186 22944
rect 14242 22888 16762 22944
rect 16818 22888 16823 22944
rect 14181 22886 16823 22888
rect 14181 22883 14247 22886
rect 16757 22883 16823 22886
rect 17677 22946 17743 22949
rect 19057 22946 19123 22949
rect 17677 22944 19123 22946
rect 17677 22888 17682 22944
rect 17738 22888 19062 22944
rect 19118 22888 19123 22944
rect 17677 22886 19123 22888
rect 17677 22883 17743 22886
rect 19057 22883 19123 22886
rect 10208 22880 10528 22881
rect 10208 22816 10216 22880
rect 10280 22816 10296 22880
rect 10360 22816 10376 22880
rect 10440 22816 10456 22880
rect 10520 22816 10528 22880
rect 10208 22815 10528 22816
rect 19472 22880 19792 22881
rect 19472 22816 19480 22880
rect 19544 22816 19560 22880
rect 19624 22816 19640 22880
rect 19704 22816 19720 22880
rect 19784 22816 19792 22880
rect 19472 22815 19792 22816
rect 11329 22810 11395 22813
rect 13721 22810 13787 22813
rect 17769 22810 17835 22813
rect 11329 22808 17835 22810
rect 11329 22752 11334 22808
rect 11390 22752 13726 22808
rect 13782 22752 17774 22808
rect 17830 22752 17835 22808
rect 11329 22750 17835 22752
rect 11329 22747 11395 22750
rect 13721 22747 13787 22750
rect 17769 22747 17835 22750
rect 23749 22810 23815 22813
rect 26969 22810 27035 22813
rect 23749 22808 27035 22810
rect 23749 22752 23754 22808
rect 23810 22752 26974 22808
rect 27030 22752 27035 22808
rect 23749 22750 27035 22752
rect 23749 22747 23815 22750
rect 26969 22747 27035 22750
rect 11973 22674 12039 22677
rect 15745 22674 15811 22677
rect 17953 22674 18019 22677
rect 11973 22672 18019 22674
rect 0 22388 800 22628
rect 11973 22616 11978 22672
rect 12034 22616 15750 22672
rect 15806 22616 17958 22672
rect 18014 22616 18019 22672
rect 11973 22614 18019 22616
rect 11973 22611 12039 22614
rect 15745 22611 15811 22614
rect 17953 22611 18019 22614
rect 18505 22674 18571 22677
rect 20989 22674 21055 22677
rect 18505 22672 21055 22674
rect 18505 22616 18510 22672
rect 18566 22616 20994 22672
rect 21050 22616 21055 22672
rect 18505 22614 21055 22616
rect 18505 22611 18571 22614
rect 20989 22611 21055 22614
rect 23657 22674 23723 22677
rect 24945 22674 25011 22677
rect 25313 22674 25379 22677
rect 23657 22672 25379 22674
rect 23657 22616 23662 22672
rect 23718 22616 24950 22672
rect 25006 22616 25318 22672
rect 25374 22616 25379 22672
rect 23657 22614 25379 22616
rect 23657 22611 23723 22614
rect 24945 22611 25011 22614
rect 25313 22611 25379 22614
rect 13261 22538 13327 22541
rect 19609 22538 19675 22541
rect 13261 22536 19675 22538
rect 13261 22480 13266 22536
rect 13322 22480 19614 22536
rect 19670 22480 19675 22536
rect 13261 22478 19675 22480
rect 13261 22475 13327 22478
rect 19609 22475 19675 22478
rect 19793 22538 19859 22541
rect 24669 22538 24735 22541
rect 19793 22536 24735 22538
rect 19793 22480 19798 22536
rect 19854 22480 24674 22536
rect 24730 22480 24735 22536
rect 19793 22478 24735 22480
rect 19793 22475 19859 22478
rect 24669 22475 24735 22478
rect 28165 22538 28231 22541
rect 29200 22538 30000 22628
rect 28165 22536 30000 22538
rect 28165 22480 28170 22536
rect 28226 22480 30000 22536
rect 28165 22478 30000 22480
rect 28165 22475 28231 22478
rect 15285 22402 15351 22405
rect 18045 22402 18111 22405
rect 15285 22400 18111 22402
rect 15285 22344 15290 22400
rect 15346 22344 18050 22400
rect 18106 22344 18111 22400
rect 29200 22388 30000 22478
rect 15285 22342 18111 22344
rect 15285 22339 15351 22342
rect 18045 22339 18111 22342
rect 5576 22336 5896 22337
rect 5576 22272 5584 22336
rect 5648 22272 5664 22336
rect 5728 22272 5744 22336
rect 5808 22272 5824 22336
rect 5888 22272 5896 22336
rect 5576 22271 5896 22272
rect 14840 22336 15160 22337
rect 14840 22272 14848 22336
rect 14912 22272 14928 22336
rect 14992 22272 15008 22336
rect 15072 22272 15088 22336
rect 15152 22272 15160 22336
rect 14840 22271 15160 22272
rect 24104 22336 24424 22337
rect 24104 22272 24112 22336
rect 24176 22272 24192 22336
rect 24256 22272 24272 22336
rect 24336 22272 24352 22336
rect 24416 22272 24424 22336
rect 24104 22271 24424 22272
rect 15469 22266 15535 22269
rect 16481 22266 16547 22269
rect 17493 22266 17559 22269
rect 15469 22264 16547 22266
rect 15469 22208 15474 22264
rect 15530 22208 16486 22264
rect 16542 22208 16547 22264
rect 15469 22206 16547 22208
rect 15469 22203 15535 22206
rect 16481 22203 16547 22206
rect 16760 22264 17559 22266
rect 16760 22208 17498 22264
rect 17554 22208 17559 22264
rect 16760 22206 17559 22208
rect 12249 22130 12315 22133
rect 16760 22130 16820 22206
rect 17493 22203 17559 22206
rect 12249 22128 16820 22130
rect 12249 22072 12254 22128
rect 12310 22072 16820 22128
rect 12249 22070 16820 22072
rect 19609 22130 19675 22133
rect 19926 22130 19932 22132
rect 19609 22128 19932 22130
rect 19609 22072 19614 22128
rect 19670 22072 19932 22128
rect 19609 22070 19932 22072
rect 12249 22067 12315 22070
rect 19609 22067 19675 22070
rect 19926 22068 19932 22070
rect 19996 22068 20002 22132
rect 20069 22130 20135 22133
rect 23657 22132 23723 22133
rect 22134 22130 22140 22132
rect 20069 22128 22140 22130
rect 20069 22072 20074 22128
rect 20130 22072 22140 22128
rect 20069 22070 22140 22072
rect 20069 22067 20135 22070
rect 22134 22068 22140 22070
rect 22204 22068 22210 22132
rect 23606 22068 23612 22132
rect 23676 22130 23723 22132
rect 23676 22128 23768 22130
rect 23718 22072 23768 22128
rect 23676 22070 23768 22072
rect 23676 22068 23723 22070
rect 23657 22067 23723 22068
rect 13353 21994 13419 21997
rect 14181 21994 14247 21997
rect 15469 21994 15535 21997
rect 13353 21992 15535 21994
rect 0 21708 800 21948
rect 13353 21936 13358 21992
rect 13414 21936 14186 21992
rect 14242 21936 15474 21992
rect 15530 21936 15535 21992
rect 13353 21934 15535 21936
rect 13353 21931 13419 21934
rect 14181 21931 14247 21934
rect 15469 21931 15535 21934
rect 16021 21994 16087 21997
rect 18321 21994 18387 21997
rect 21357 21994 21423 21997
rect 16021 21992 18387 21994
rect 16021 21936 16026 21992
rect 16082 21936 18326 21992
rect 18382 21936 18387 21992
rect 16021 21934 18387 21936
rect 16021 21931 16087 21934
rect 18321 21931 18387 21934
rect 19198 21992 21423 21994
rect 19198 21936 21362 21992
rect 21418 21936 21423 21992
rect 19198 21934 21423 21936
rect 13629 21858 13695 21861
rect 16024 21858 16084 21931
rect 13629 21856 16084 21858
rect 13629 21800 13634 21856
rect 13690 21800 16084 21856
rect 13629 21798 16084 21800
rect 16573 21858 16639 21861
rect 19198 21858 19258 21934
rect 21357 21931 21423 21934
rect 16573 21856 19258 21858
rect 16573 21800 16578 21856
rect 16634 21800 19258 21856
rect 16573 21798 19258 21800
rect 26141 21858 26207 21861
rect 29200 21858 30000 21948
rect 26141 21856 30000 21858
rect 26141 21800 26146 21856
rect 26202 21800 30000 21856
rect 26141 21798 30000 21800
rect 13629 21795 13695 21798
rect 16573 21795 16639 21798
rect 26141 21795 26207 21798
rect 10208 21792 10528 21793
rect 10208 21728 10216 21792
rect 10280 21728 10296 21792
rect 10360 21728 10376 21792
rect 10440 21728 10456 21792
rect 10520 21728 10528 21792
rect 10208 21727 10528 21728
rect 19472 21792 19792 21793
rect 19472 21728 19480 21792
rect 19544 21728 19560 21792
rect 19624 21728 19640 21792
rect 19704 21728 19720 21792
rect 19784 21728 19792 21792
rect 19472 21727 19792 21728
rect 11237 21722 11303 21725
rect 14733 21722 14799 21725
rect 11237 21720 14799 21722
rect 11237 21664 11242 21720
rect 11298 21664 14738 21720
rect 14794 21664 14799 21720
rect 11237 21662 14799 21664
rect 11237 21659 11303 21662
rect 14733 21659 14799 21662
rect 14917 21722 14983 21725
rect 16113 21722 16179 21725
rect 16573 21722 16639 21725
rect 14917 21720 16639 21722
rect 14917 21664 14922 21720
rect 14978 21664 16118 21720
rect 16174 21664 16578 21720
rect 16634 21664 16639 21720
rect 14917 21662 16639 21664
rect 14917 21659 14983 21662
rect 16113 21659 16179 21662
rect 16573 21659 16639 21662
rect 16757 21722 16823 21725
rect 18505 21722 18571 21725
rect 16757 21720 18571 21722
rect 16757 21664 16762 21720
rect 16818 21664 18510 21720
rect 18566 21664 18571 21720
rect 29200 21708 30000 21798
rect 16757 21662 18571 21664
rect 16757 21659 16823 21662
rect 18505 21659 18571 21662
rect 14365 21586 14431 21589
rect 22921 21586 22987 21589
rect 14365 21584 22987 21586
rect 14365 21528 14370 21584
rect 14426 21528 22926 21584
rect 22982 21528 22987 21584
rect 14365 21526 22987 21528
rect 14365 21523 14431 21526
rect 22921 21523 22987 21526
rect 12617 21450 12683 21453
rect 19926 21450 19932 21452
rect 12617 21448 19932 21450
rect 12617 21392 12622 21448
rect 12678 21392 19932 21448
rect 12617 21390 19932 21392
rect 12617 21387 12683 21390
rect 19926 21388 19932 21390
rect 19996 21388 20002 21452
rect 16021 21314 16087 21317
rect 19149 21314 19215 21317
rect 16021 21312 19215 21314
rect 0 21028 800 21268
rect 16021 21256 16026 21312
rect 16082 21256 19154 21312
rect 19210 21256 19215 21312
rect 16021 21254 19215 21256
rect 16021 21251 16087 21254
rect 19149 21251 19215 21254
rect 5576 21248 5896 21249
rect 5576 21184 5584 21248
rect 5648 21184 5664 21248
rect 5728 21184 5744 21248
rect 5808 21184 5824 21248
rect 5888 21184 5896 21248
rect 5576 21183 5896 21184
rect 14840 21248 15160 21249
rect 14840 21184 14848 21248
rect 14912 21184 14928 21248
rect 14992 21184 15008 21248
rect 15072 21184 15088 21248
rect 15152 21184 15160 21248
rect 14840 21183 15160 21184
rect 24104 21248 24424 21249
rect 24104 21184 24112 21248
rect 24176 21184 24192 21248
rect 24256 21184 24272 21248
rect 24336 21184 24352 21248
rect 24416 21184 24424 21248
rect 24104 21183 24424 21184
rect 16573 21178 16639 21181
rect 22369 21178 22435 21181
rect 16573 21176 22435 21178
rect 16573 21120 16578 21176
rect 16634 21120 22374 21176
rect 22430 21120 22435 21176
rect 16573 21118 22435 21120
rect 16573 21115 16639 21118
rect 22369 21115 22435 21118
rect 24577 21178 24643 21181
rect 24853 21178 24919 21181
rect 24577 21176 24919 21178
rect 24577 21120 24582 21176
rect 24638 21120 24858 21176
rect 24914 21120 24919 21176
rect 24577 21118 24919 21120
rect 24577 21115 24643 21118
rect 24853 21115 24919 21118
rect 28165 21178 28231 21181
rect 29200 21178 30000 21268
rect 28165 21176 30000 21178
rect 28165 21120 28170 21176
rect 28226 21120 30000 21176
rect 28165 21118 30000 21120
rect 28165 21115 28231 21118
rect 13905 21042 13971 21045
rect 15377 21042 15443 21045
rect 13905 21040 15443 21042
rect 13905 20984 13910 21040
rect 13966 20984 15382 21040
rect 15438 20984 15443 21040
rect 13905 20982 15443 20984
rect 13905 20979 13971 20982
rect 15377 20979 15443 20982
rect 15745 21042 15811 21045
rect 22737 21042 22803 21045
rect 15745 21040 22803 21042
rect 15745 20984 15750 21040
rect 15806 20984 22742 21040
rect 22798 20984 22803 21040
rect 29200 21028 30000 21118
rect 15745 20982 22803 20984
rect 15745 20979 15811 20982
rect 22737 20979 22803 20982
rect 12065 20906 12131 20909
rect 14825 20906 14891 20909
rect 12065 20904 14891 20906
rect 12065 20848 12070 20904
rect 12126 20848 14830 20904
rect 14886 20848 14891 20904
rect 12065 20846 14891 20848
rect 12065 20843 12131 20846
rect 14825 20843 14891 20846
rect 16982 20844 16988 20908
rect 17052 20906 17058 20908
rect 17769 20906 17835 20909
rect 22185 20906 22251 20909
rect 17052 20904 17835 20906
rect 17052 20848 17774 20904
rect 17830 20848 17835 20904
rect 17052 20846 17835 20848
rect 17052 20844 17058 20846
rect 17769 20843 17835 20846
rect 19290 20904 22251 20906
rect 19290 20848 22190 20904
rect 22246 20848 22251 20904
rect 19290 20846 22251 20848
rect 12985 20770 13051 20773
rect 18505 20770 18571 20773
rect 19290 20770 19350 20846
rect 22185 20843 22251 20846
rect 12985 20768 19350 20770
rect 12985 20712 12990 20768
rect 13046 20712 18510 20768
rect 18566 20712 19350 20768
rect 12985 20710 19350 20712
rect 12985 20707 13051 20710
rect 18505 20707 18571 20710
rect 10208 20704 10528 20705
rect 10208 20640 10216 20704
rect 10280 20640 10296 20704
rect 10360 20640 10376 20704
rect 10440 20640 10456 20704
rect 10520 20640 10528 20704
rect 10208 20639 10528 20640
rect 19472 20704 19792 20705
rect 19472 20640 19480 20704
rect 19544 20640 19560 20704
rect 19624 20640 19640 20704
rect 19704 20640 19720 20704
rect 19784 20640 19792 20704
rect 19472 20639 19792 20640
rect 13261 20634 13327 20637
rect 18873 20634 18939 20637
rect 13261 20632 18939 20634
rect 0 20348 800 20588
rect 13261 20576 13266 20632
rect 13322 20576 18878 20632
rect 18934 20576 18939 20632
rect 13261 20574 18939 20576
rect 13261 20571 13327 20574
rect 18873 20571 18939 20574
rect 10869 20498 10935 20501
rect 13629 20498 13695 20501
rect 16614 20498 16620 20500
rect 10869 20496 16620 20498
rect 10869 20440 10874 20496
rect 10930 20440 13634 20496
rect 13690 20440 16620 20496
rect 10869 20438 16620 20440
rect 10869 20435 10935 20438
rect 13629 20435 13695 20438
rect 16614 20436 16620 20438
rect 16684 20498 16690 20500
rect 21817 20498 21883 20501
rect 16684 20496 21883 20498
rect 16684 20440 21822 20496
rect 21878 20440 21883 20496
rect 16684 20438 21883 20440
rect 16684 20436 16690 20438
rect 21817 20435 21883 20438
rect 12157 20362 12223 20365
rect 22645 20362 22711 20365
rect 12157 20360 22711 20362
rect 12157 20304 12162 20360
rect 12218 20304 22650 20360
rect 22706 20304 22711 20360
rect 29200 20348 30000 20588
rect 12157 20302 22711 20304
rect 12157 20299 12223 20302
rect 22645 20299 22711 20302
rect 5576 20160 5896 20161
rect 5576 20096 5584 20160
rect 5648 20096 5664 20160
rect 5728 20096 5744 20160
rect 5808 20096 5824 20160
rect 5888 20096 5896 20160
rect 5576 20095 5896 20096
rect 14840 20160 15160 20161
rect 14840 20096 14848 20160
rect 14912 20096 14928 20160
rect 14992 20096 15008 20160
rect 15072 20096 15088 20160
rect 15152 20096 15160 20160
rect 14840 20095 15160 20096
rect 24104 20160 24424 20161
rect 24104 20096 24112 20160
rect 24176 20096 24192 20160
rect 24256 20096 24272 20160
rect 24336 20096 24352 20160
rect 24416 20096 24424 20160
rect 24104 20095 24424 20096
rect 15101 19954 15167 19957
rect 16849 19954 16915 19957
rect 15101 19952 16915 19954
rect 0 19668 800 19908
rect 15101 19896 15106 19952
rect 15162 19896 16854 19952
rect 16910 19896 16915 19952
rect 15101 19894 16915 19896
rect 15101 19891 15167 19894
rect 16849 19891 16915 19894
rect 22134 19892 22140 19956
rect 22204 19954 22210 19956
rect 24301 19954 24367 19957
rect 27889 19954 27955 19957
rect 22204 19952 27955 19954
rect 22204 19896 24306 19952
rect 24362 19896 27894 19952
rect 27950 19896 27955 19952
rect 22204 19894 27955 19896
rect 22204 19892 22210 19894
rect 24301 19891 24367 19894
rect 27889 19891 27955 19894
rect 28165 19818 28231 19821
rect 29200 19818 30000 19908
rect 28165 19816 30000 19818
rect 28165 19760 28170 19816
rect 28226 19760 30000 19816
rect 28165 19758 30000 19760
rect 28165 19755 28231 19758
rect 15101 19682 15167 19685
rect 17033 19682 17099 19685
rect 15101 19680 17099 19682
rect 15101 19624 15106 19680
rect 15162 19624 17038 19680
rect 17094 19624 17099 19680
rect 29200 19668 30000 19758
rect 15101 19622 17099 19624
rect 15101 19619 15167 19622
rect 17033 19619 17099 19622
rect 10208 19616 10528 19617
rect 10208 19552 10216 19616
rect 10280 19552 10296 19616
rect 10360 19552 10376 19616
rect 10440 19552 10456 19616
rect 10520 19552 10528 19616
rect 10208 19551 10528 19552
rect 19472 19616 19792 19617
rect 19472 19552 19480 19616
rect 19544 19552 19560 19616
rect 19624 19552 19640 19616
rect 19704 19552 19720 19616
rect 19784 19552 19792 19616
rect 19472 19551 19792 19552
rect 12433 19410 12499 19413
rect 16849 19410 16915 19413
rect 12433 19408 16915 19410
rect 12433 19352 12438 19408
rect 12494 19352 16854 19408
rect 16910 19352 16915 19408
rect 12433 19350 16915 19352
rect 12433 19347 12499 19350
rect 16849 19347 16915 19350
rect 0 18988 800 19228
rect 28165 19138 28231 19141
rect 29200 19138 30000 19228
rect 28165 19136 30000 19138
rect 28165 19080 28170 19136
rect 28226 19080 30000 19136
rect 28165 19078 30000 19080
rect 28165 19075 28231 19078
rect 5576 19072 5896 19073
rect 5576 19008 5584 19072
rect 5648 19008 5664 19072
rect 5728 19008 5744 19072
rect 5808 19008 5824 19072
rect 5888 19008 5896 19072
rect 5576 19007 5896 19008
rect 14840 19072 15160 19073
rect 14840 19008 14848 19072
rect 14912 19008 14928 19072
rect 14992 19008 15008 19072
rect 15072 19008 15088 19072
rect 15152 19008 15160 19072
rect 14840 19007 15160 19008
rect 24104 19072 24424 19073
rect 24104 19008 24112 19072
rect 24176 19008 24192 19072
rect 24256 19008 24272 19072
rect 24336 19008 24352 19072
rect 24416 19008 24424 19072
rect 24104 19007 24424 19008
rect 29200 18988 30000 19078
rect 25221 18866 25287 18869
rect 25497 18866 25563 18869
rect 25221 18864 25563 18866
rect 25221 18808 25226 18864
rect 25282 18808 25502 18864
rect 25558 18808 25563 18864
rect 25221 18806 25563 18808
rect 25221 18803 25287 18806
rect 25497 18803 25563 18806
rect 0 18308 800 18548
rect 10208 18528 10528 18529
rect 10208 18464 10216 18528
rect 10280 18464 10296 18528
rect 10360 18464 10376 18528
rect 10440 18464 10456 18528
rect 10520 18464 10528 18528
rect 10208 18463 10528 18464
rect 19472 18528 19792 18529
rect 19472 18464 19480 18528
rect 19544 18464 19560 18528
rect 19624 18464 19640 18528
rect 19704 18464 19720 18528
rect 19784 18464 19792 18528
rect 19472 18463 19792 18464
rect 28165 18458 28231 18461
rect 29200 18458 30000 18548
rect 28165 18456 30000 18458
rect 28165 18400 28170 18456
rect 28226 18400 30000 18456
rect 28165 18398 30000 18400
rect 28165 18395 28231 18398
rect 14181 18322 14247 18325
rect 18321 18322 18387 18325
rect 14181 18320 18387 18322
rect 14181 18264 14186 18320
rect 14242 18264 18326 18320
rect 18382 18264 18387 18320
rect 29200 18308 30000 18398
rect 14181 18262 18387 18264
rect 14181 18259 14247 18262
rect 18321 18259 18387 18262
rect 25037 18186 25103 18189
rect 25221 18186 25287 18189
rect 25037 18184 25287 18186
rect 25037 18128 25042 18184
rect 25098 18128 25226 18184
rect 25282 18128 25287 18184
rect 25037 18126 25287 18128
rect 25037 18123 25103 18126
rect 25221 18123 25287 18126
rect 5576 17984 5896 17985
rect 5576 17920 5584 17984
rect 5648 17920 5664 17984
rect 5728 17920 5744 17984
rect 5808 17920 5824 17984
rect 5888 17920 5896 17984
rect 5576 17919 5896 17920
rect 14840 17984 15160 17985
rect 14840 17920 14848 17984
rect 14912 17920 14928 17984
rect 14992 17920 15008 17984
rect 15072 17920 15088 17984
rect 15152 17920 15160 17984
rect 14840 17919 15160 17920
rect 24104 17984 24424 17985
rect 24104 17920 24112 17984
rect 24176 17920 24192 17984
rect 24256 17920 24272 17984
rect 24336 17920 24352 17984
rect 24416 17920 24424 17984
rect 24104 17919 24424 17920
rect 0 17778 800 17868
rect 2773 17778 2839 17781
rect 0 17776 2839 17778
rect 0 17720 2778 17776
rect 2834 17720 2839 17776
rect 0 17718 2839 17720
rect 0 17628 800 17718
rect 2773 17715 2839 17718
rect 7557 17778 7623 17781
rect 18454 17778 18460 17780
rect 7557 17776 18460 17778
rect 7557 17720 7562 17776
rect 7618 17720 18460 17776
rect 7557 17718 18460 17720
rect 7557 17715 7623 17718
rect 18454 17716 18460 17718
rect 18524 17716 18530 17780
rect 24301 17778 24367 17781
rect 26550 17778 26556 17780
rect 24301 17776 26556 17778
rect 24301 17720 24306 17776
rect 24362 17720 26556 17776
rect 24301 17718 26556 17720
rect 24301 17715 24367 17718
rect 26550 17716 26556 17718
rect 26620 17716 26626 17780
rect 10593 17642 10659 17645
rect 26366 17642 26372 17644
rect 10593 17640 26372 17642
rect 10593 17584 10598 17640
rect 10654 17584 26372 17640
rect 10593 17582 26372 17584
rect 10593 17579 10659 17582
rect 26366 17580 26372 17582
rect 26436 17580 26442 17644
rect 29200 17628 30000 17868
rect 10208 17440 10528 17441
rect 10208 17376 10216 17440
rect 10280 17376 10296 17440
rect 10360 17376 10376 17440
rect 10440 17376 10456 17440
rect 10520 17376 10528 17440
rect 10208 17375 10528 17376
rect 19472 17440 19792 17441
rect 19472 17376 19480 17440
rect 19544 17376 19560 17440
rect 19624 17376 19640 17440
rect 19704 17376 19720 17440
rect 19784 17376 19792 17440
rect 19472 17375 19792 17376
rect 0 17098 800 17188
rect 1853 17098 1919 17101
rect 0 17096 1919 17098
rect 0 17040 1858 17096
rect 1914 17040 1919 17096
rect 0 17038 1919 17040
rect 0 16948 800 17038
rect 1853 17035 1919 17038
rect 5576 16896 5896 16897
rect 5576 16832 5584 16896
rect 5648 16832 5664 16896
rect 5728 16832 5744 16896
rect 5808 16832 5824 16896
rect 5888 16832 5896 16896
rect 5576 16831 5896 16832
rect 14840 16896 15160 16897
rect 14840 16832 14848 16896
rect 14912 16832 14928 16896
rect 14992 16832 15008 16896
rect 15072 16832 15088 16896
rect 15152 16832 15160 16896
rect 14840 16831 15160 16832
rect 24104 16896 24424 16897
rect 24104 16832 24112 16896
rect 24176 16832 24192 16896
rect 24256 16832 24272 16896
rect 24336 16832 24352 16896
rect 24416 16832 24424 16896
rect 24104 16831 24424 16832
rect 22001 16690 22067 16693
rect 23197 16690 23263 16693
rect 22001 16688 23263 16690
rect 22001 16632 22006 16688
rect 22062 16632 23202 16688
rect 23258 16632 23263 16688
rect 22001 16630 23263 16632
rect 22001 16627 22067 16630
rect 23197 16627 23263 16630
rect 7741 16554 7807 16557
rect 26182 16554 26188 16556
rect 7741 16552 26188 16554
rect 0 16268 800 16508
rect 7741 16496 7746 16552
rect 7802 16496 26188 16552
rect 7741 16494 26188 16496
rect 7741 16491 7807 16494
rect 26182 16492 26188 16494
rect 26252 16492 26258 16556
rect 28165 16418 28231 16421
rect 29200 16418 30000 16508
rect 28165 16416 30000 16418
rect 28165 16360 28170 16416
rect 28226 16360 30000 16416
rect 28165 16358 30000 16360
rect 28165 16355 28231 16358
rect 10208 16352 10528 16353
rect 10208 16288 10216 16352
rect 10280 16288 10296 16352
rect 10360 16288 10376 16352
rect 10440 16288 10456 16352
rect 10520 16288 10528 16352
rect 10208 16287 10528 16288
rect 19472 16352 19792 16353
rect 19472 16288 19480 16352
rect 19544 16288 19560 16352
rect 19624 16288 19640 16352
rect 19704 16288 19720 16352
rect 19784 16288 19792 16352
rect 19472 16287 19792 16288
rect 29200 16268 30000 16358
rect 9581 16146 9647 16149
rect 18638 16146 18644 16148
rect 9581 16144 18644 16146
rect 9581 16088 9586 16144
rect 9642 16088 18644 16144
rect 9581 16086 18644 16088
rect 9581 16083 9647 16086
rect 18638 16084 18644 16086
rect 18708 16084 18714 16148
rect 0 15738 800 15828
rect 5576 15808 5896 15809
rect 5576 15744 5584 15808
rect 5648 15744 5664 15808
rect 5728 15744 5744 15808
rect 5808 15744 5824 15808
rect 5888 15744 5896 15808
rect 5576 15743 5896 15744
rect 14840 15808 15160 15809
rect 14840 15744 14848 15808
rect 14912 15744 14928 15808
rect 14992 15744 15008 15808
rect 15072 15744 15088 15808
rect 15152 15744 15160 15808
rect 14840 15743 15160 15744
rect 24104 15808 24424 15809
rect 24104 15744 24112 15808
rect 24176 15744 24192 15808
rect 24256 15744 24272 15808
rect 24336 15744 24352 15808
rect 24416 15744 24424 15808
rect 24104 15743 24424 15744
rect 2773 15738 2839 15741
rect 0 15736 2839 15738
rect 0 15680 2778 15736
rect 2834 15680 2839 15736
rect 0 15678 2839 15680
rect 0 15588 800 15678
rect 2773 15675 2839 15678
rect 26141 15738 26207 15741
rect 29200 15738 30000 15828
rect 26141 15736 30000 15738
rect 26141 15680 26146 15736
rect 26202 15680 30000 15736
rect 26141 15678 30000 15680
rect 26141 15675 26207 15678
rect 29200 15588 30000 15678
rect 10208 15264 10528 15265
rect 10208 15200 10216 15264
rect 10280 15200 10296 15264
rect 10360 15200 10376 15264
rect 10440 15200 10456 15264
rect 10520 15200 10528 15264
rect 10208 15199 10528 15200
rect 19472 15264 19792 15265
rect 19472 15200 19480 15264
rect 19544 15200 19560 15264
rect 19624 15200 19640 15264
rect 19704 15200 19720 15264
rect 19784 15200 19792 15264
rect 19472 15199 19792 15200
rect 0 14908 800 15148
rect 28165 15058 28231 15061
rect 29200 15058 30000 15148
rect 28165 15056 30000 15058
rect 28165 15000 28170 15056
rect 28226 15000 30000 15056
rect 28165 14998 30000 15000
rect 28165 14995 28231 14998
rect 29200 14908 30000 14998
rect 5576 14720 5896 14721
rect 5576 14656 5584 14720
rect 5648 14656 5664 14720
rect 5728 14656 5744 14720
rect 5808 14656 5824 14720
rect 5888 14656 5896 14720
rect 5576 14655 5896 14656
rect 14840 14720 15160 14721
rect 14840 14656 14848 14720
rect 14912 14656 14928 14720
rect 14992 14656 15008 14720
rect 15072 14656 15088 14720
rect 15152 14656 15160 14720
rect 14840 14655 15160 14656
rect 24104 14720 24424 14721
rect 24104 14656 24112 14720
rect 24176 14656 24192 14720
rect 24256 14656 24272 14720
rect 24336 14656 24352 14720
rect 24416 14656 24424 14720
rect 24104 14655 24424 14656
rect 0 14378 800 14468
rect 1853 14378 1919 14381
rect 0 14376 1919 14378
rect 0 14320 1858 14376
rect 1914 14320 1919 14376
rect 0 14318 1919 14320
rect 0 14228 800 14318
rect 1853 14315 1919 14318
rect 28165 14378 28231 14381
rect 29200 14378 30000 14468
rect 28165 14376 30000 14378
rect 28165 14320 28170 14376
rect 28226 14320 30000 14376
rect 28165 14318 30000 14320
rect 28165 14315 28231 14318
rect 29200 14228 30000 14318
rect 10208 14176 10528 14177
rect 10208 14112 10216 14176
rect 10280 14112 10296 14176
rect 10360 14112 10376 14176
rect 10440 14112 10456 14176
rect 10520 14112 10528 14176
rect 10208 14111 10528 14112
rect 19472 14176 19792 14177
rect 19472 14112 19480 14176
rect 19544 14112 19560 14176
rect 19624 14112 19640 14176
rect 19704 14112 19720 14176
rect 19784 14112 19792 14176
rect 19472 14111 19792 14112
rect 0 13548 800 13788
rect 5576 13632 5896 13633
rect 5576 13568 5584 13632
rect 5648 13568 5664 13632
rect 5728 13568 5744 13632
rect 5808 13568 5824 13632
rect 5888 13568 5896 13632
rect 5576 13567 5896 13568
rect 14840 13632 15160 13633
rect 14840 13568 14848 13632
rect 14912 13568 14928 13632
rect 14992 13568 15008 13632
rect 15072 13568 15088 13632
rect 15152 13568 15160 13632
rect 14840 13567 15160 13568
rect 24104 13632 24424 13633
rect 24104 13568 24112 13632
rect 24176 13568 24192 13632
rect 24256 13568 24272 13632
rect 24336 13568 24352 13632
rect 24416 13568 24424 13632
rect 24104 13567 24424 13568
rect 29200 13548 30000 13788
rect 0 13018 800 13108
rect 10208 13088 10528 13089
rect 10208 13024 10216 13088
rect 10280 13024 10296 13088
rect 10360 13024 10376 13088
rect 10440 13024 10456 13088
rect 10520 13024 10528 13088
rect 10208 13023 10528 13024
rect 19472 13088 19792 13089
rect 19472 13024 19480 13088
rect 19544 13024 19560 13088
rect 19624 13024 19640 13088
rect 19704 13024 19720 13088
rect 19784 13024 19792 13088
rect 19472 13023 19792 13024
rect 2773 13018 2839 13021
rect 0 13016 2839 13018
rect 0 12960 2778 13016
rect 2834 12960 2839 13016
rect 0 12958 2839 12960
rect 0 12868 800 12958
rect 2773 12955 2839 12958
rect 29200 12868 30000 13108
rect 5576 12544 5896 12545
rect 5576 12480 5584 12544
rect 5648 12480 5664 12544
rect 5728 12480 5744 12544
rect 5808 12480 5824 12544
rect 5888 12480 5896 12544
rect 5576 12479 5896 12480
rect 14840 12544 15160 12545
rect 14840 12480 14848 12544
rect 14912 12480 14928 12544
rect 14992 12480 15008 12544
rect 15072 12480 15088 12544
rect 15152 12480 15160 12544
rect 14840 12479 15160 12480
rect 24104 12544 24424 12545
rect 24104 12480 24112 12544
rect 24176 12480 24192 12544
rect 24256 12480 24272 12544
rect 24336 12480 24352 12544
rect 24416 12480 24424 12544
rect 24104 12479 24424 12480
rect 0 12338 800 12428
rect 2773 12338 2839 12341
rect 0 12336 2839 12338
rect 0 12280 2778 12336
rect 2834 12280 2839 12336
rect 0 12278 2839 12280
rect 0 12188 800 12278
rect 2773 12275 2839 12278
rect 29200 12188 30000 12428
rect 10208 12000 10528 12001
rect 10208 11936 10216 12000
rect 10280 11936 10296 12000
rect 10360 11936 10376 12000
rect 10440 11936 10456 12000
rect 10520 11936 10528 12000
rect 10208 11935 10528 11936
rect 19472 12000 19792 12001
rect 19472 11936 19480 12000
rect 19544 11936 19560 12000
rect 19624 11936 19640 12000
rect 19704 11936 19720 12000
rect 19784 11936 19792 12000
rect 19472 11935 19792 11936
rect 0 11508 800 11748
rect 27981 11658 28047 11661
rect 29200 11658 30000 11748
rect 27981 11656 30000 11658
rect 27981 11600 27986 11656
rect 28042 11600 30000 11656
rect 27981 11598 30000 11600
rect 27981 11595 28047 11598
rect 29200 11508 30000 11598
rect 5576 11456 5896 11457
rect 5576 11392 5584 11456
rect 5648 11392 5664 11456
rect 5728 11392 5744 11456
rect 5808 11392 5824 11456
rect 5888 11392 5896 11456
rect 5576 11391 5896 11392
rect 14840 11456 15160 11457
rect 14840 11392 14848 11456
rect 14912 11392 14928 11456
rect 14992 11392 15008 11456
rect 15072 11392 15088 11456
rect 15152 11392 15160 11456
rect 14840 11391 15160 11392
rect 24104 11456 24424 11457
rect 24104 11392 24112 11456
rect 24176 11392 24192 11456
rect 24256 11392 24272 11456
rect 24336 11392 24352 11456
rect 24416 11392 24424 11456
rect 24104 11391 24424 11392
rect 0 10978 800 11068
rect 1853 10978 1919 10981
rect 0 10976 1919 10978
rect 0 10920 1858 10976
rect 1914 10920 1919 10976
rect 0 10918 1919 10920
rect 0 10828 800 10918
rect 1853 10915 1919 10918
rect 28165 10978 28231 10981
rect 29200 10978 30000 11068
rect 28165 10976 30000 10978
rect 28165 10920 28170 10976
rect 28226 10920 30000 10976
rect 28165 10918 30000 10920
rect 28165 10915 28231 10918
rect 10208 10912 10528 10913
rect 10208 10848 10216 10912
rect 10280 10848 10296 10912
rect 10360 10848 10376 10912
rect 10440 10848 10456 10912
rect 10520 10848 10528 10912
rect 10208 10847 10528 10848
rect 19472 10912 19792 10913
rect 19472 10848 19480 10912
rect 19544 10848 19560 10912
rect 19624 10848 19640 10912
rect 19704 10848 19720 10912
rect 19784 10848 19792 10912
rect 19472 10847 19792 10848
rect 29200 10828 30000 10918
rect 0 10298 800 10388
rect 5576 10368 5896 10369
rect 5576 10304 5584 10368
rect 5648 10304 5664 10368
rect 5728 10304 5744 10368
rect 5808 10304 5824 10368
rect 5888 10304 5896 10368
rect 5576 10303 5896 10304
rect 14840 10368 15160 10369
rect 14840 10304 14848 10368
rect 14912 10304 14928 10368
rect 14992 10304 15008 10368
rect 15072 10304 15088 10368
rect 15152 10304 15160 10368
rect 14840 10303 15160 10304
rect 24104 10368 24424 10369
rect 24104 10304 24112 10368
rect 24176 10304 24192 10368
rect 24256 10304 24272 10368
rect 24336 10304 24352 10368
rect 24416 10304 24424 10368
rect 24104 10303 24424 10304
rect 2865 10298 2931 10301
rect 0 10296 2931 10298
rect 0 10240 2870 10296
rect 2926 10240 2931 10296
rect 0 10238 2931 10240
rect 0 10148 800 10238
rect 2865 10235 2931 10238
rect 29200 10148 30000 10388
rect 10208 9824 10528 9825
rect 10208 9760 10216 9824
rect 10280 9760 10296 9824
rect 10360 9760 10376 9824
rect 10440 9760 10456 9824
rect 10520 9760 10528 9824
rect 10208 9759 10528 9760
rect 19472 9824 19792 9825
rect 19472 9760 19480 9824
rect 19544 9760 19560 9824
rect 19624 9760 19640 9824
rect 19704 9760 19720 9824
rect 19784 9760 19792 9824
rect 19472 9759 19792 9760
rect 0 9468 800 9708
rect 28165 9618 28231 9621
rect 29200 9618 30000 9708
rect 28165 9616 30000 9618
rect 28165 9560 28170 9616
rect 28226 9560 30000 9616
rect 28165 9558 30000 9560
rect 28165 9555 28231 9558
rect 29200 9468 30000 9558
rect 5576 9280 5896 9281
rect 5576 9216 5584 9280
rect 5648 9216 5664 9280
rect 5728 9216 5744 9280
rect 5808 9216 5824 9280
rect 5888 9216 5896 9280
rect 5576 9215 5896 9216
rect 14840 9280 15160 9281
rect 14840 9216 14848 9280
rect 14912 9216 14928 9280
rect 14992 9216 15008 9280
rect 15072 9216 15088 9280
rect 15152 9216 15160 9280
rect 14840 9215 15160 9216
rect 24104 9280 24424 9281
rect 24104 9216 24112 9280
rect 24176 9216 24192 9280
rect 24256 9216 24272 9280
rect 24336 9216 24352 9280
rect 24416 9216 24424 9280
rect 24104 9215 24424 9216
rect 0 8788 800 9028
rect 29200 8788 30000 9028
rect 10208 8736 10528 8737
rect 10208 8672 10216 8736
rect 10280 8672 10296 8736
rect 10360 8672 10376 8736
rect 10440 8672 10456 8736
rect 10520 8672 10528 8736
rect 10208 8671 10528 8672
rect 19472 8736 19792 8737
rect 19472 8672 19480 8736
rect 19544 8672 19560 8736
rect 19624 8672 19640 8736
rect 19704 8672 19720 8736
rect 19784 8672 19792 8736
rect 19472 8671 19792 8672
rect 0 8258 800 8348
rect 2773 8258 2839 8261
rect 0 8256 2839 8258
rect 0 8200 2778 8256
rect 2834 8200 2839 8256
rect 0 8198 2839 8200
rect 0 8108 800 8198
rect 2773 8195 2839 8198
rect 5576 8192 5896 8193
rect 5576 8128 5584 8192
rect 5648 8128 5664 8192
rect 5728 8128 5744 8192
rect 5808 8128 5824 8192
rect 5888 8128 5896 8192
rect 5576 8127 5896 8128
rect 14840 8192 15160 8193
rect 14840 8128 14848 8192
rect 14912 8128 14928 8192
rect 14992 8128 15008 8192
rect 15072 8128 15088 8192
rect 15152 8128 15160 8192
rect 14840 8127 15160 8128
rect 24104 8192 24424 8193
rect 24104 8128 24112 8192
rect 24176 8128 24192 8192
rect 24256 8128 24272 8192
rect 24336 8128 24352 8192
rect 24416 8128 24424 8192
rect 24104 8127 24424 8128
rect 29200 8108 30000 8348
rect 0 7578 800 7668
rect 10208 7648 10528 7649
rect 10208 7584 10216 7648
rect 10280 7584 10296 7648
rect 10360 7584 10376 7648
rect 10440 7584 10456 7648
rect 10520 7584 10528 7648
rect 10208 7583 10528 7584
rect 19472 7648 19792 7649
rect 19472 7584 19480 7648
rect 19544 7584 19560 7648
rect 19624 7584 19640 7648
rect 19704 7584 19720 7648
rect 19784 7584 19792 7648
rect 19472 7583 19792 7584
rect 2773 7578 2839 7581
rect 0 7576 2839 7578
rect 0 7520 2778 7576
rect 2834 7520 2839 7576
rect 0 7518 2839 7520
rect 0 7428 800 7518
rect 2773 7515 2839 7518
rect 28165 7578 28231 7581
rect 29200 7578 30000 7668
rect 28165 7576 30000 7578
rect 28165 7520 28170 7576
rect 28226 7520 30000 7576
rect 28165 7518 30000 7520
rect 28165 7515 28231 7518
rect 29200 7428 30000 7518
rect 5576 7104 5896 7105
rect 5576 7040 5584 7104
rect 5648 7040 5664 7104
rect 5728 7040 5744 7104
rect 5808 7040 5824 7104
rect 5888 7040 5896 7104
rect 5576 7039 5896 7040
rect 14840 7104 15160 7105
rect 14840 7040 14848 7104
rect 14912 7040 14928 7104
rect 14992 7040 15008 7104
rect 15072 7040 15088 7104
rect 15152 7040 15160 7104
rect 14840 7039 15160 7040
rect 24104 7104 24424 7105
rect 24104 7040 24112 7104
rect 24176 7040 24192 7104
rect 24256 7040 24272 7104
rect 24336 7040 24352 7104
rect 24416 7040 24424 7104
rect 24104 7039 24424 7040
rect 0 6898 800 6988
rect 2865 6898 2931 6901
rect 0 6896 2931 6898
rect 0 6840 2870 6896
rect 2926 6840 2931 6896
rect 0 6838 2931 6840
rect 0 6748 800 6838
rect 2865 6835 2931 6838
rect 28165 6898 28231 6901
rect 29200 6898 30000 6988
rect 28165 6896 30000 6898
rect 28165 6840 28170 6896
rect 28226 6840 30000 6896
rect 28165 6838 30000 6840
rect 28165 6835 28231 6838
rect 29200 6748 30000 6838
rect 10208 6560 10528 6561
rect 10208 6496 10216 6560
rect 10280 6496 10296 6560
rect 10360 6496 10376 6560
rect 10440 6496 10456 6560
rect 10520 6496 10528 6560
rect 10208 6495 10528 6496
rect 19472 6560 19792 6561
rect 19472 6496 19480 6560
rect 19544 6496 19560 6560
rect 19624 6496 19640 6560
rect 19704 6496 19720 6560
rect 19784 6496 19792 6560
rect 19472 6495 19792 6496
rect 0 6068 800 6308
rect 28165 6218 28231 6221
rect 29200 6218 30000 6308
rect 28165 6216 30000 6218
rect 28165 6160 28170 6216
rect 28226 6160 30000 6216
rect 28165 6158 30000 6160
rect 28165 6155 28231 6158
rect 29200 6068 30000 6158
rect 5576 6016 5896 6017
rect 5576 5952 5584 6016
rect 5648 5952 5664 6016
rect 5728 5952 5744 6016
rect 5808 5952 5824 6016
rect 5888 5952 5896 6016
rect 5576 5951 5896 5952
rect 14840 6016 15160 6017
rect 14840 5952 14848 6016
rect 14912 5952 14928 6016
rect 14992 5952 15008 6016
rect 15072 5952 15088 6016
rect 15152 5952 15160 6016
rect 14840 5951 15160 5952
rect 24104 6016 24424 6017
rect 24104 5952 24112 6016
rect 24176 5952 24192 6016
rect 24256 5952 24272 6016
rect 24336 5952 24352 6016
rect 24416 5952 24424 6016
rect 24104 5951 24424 5952
rect 0 5538 800 5628
rect 1853 5538 1919 5541
rect 0 5536 1919 5538
rect 0 5480 1858 5536
rect 1914 5480 1919 5536
rect 0 5478 1919 5480
rect 0 5388 800 5478
rect 1853 5475 1919 5478
rect 10208 5472 10528 5473
rect 10208 5408 10216 5472
rect 10280 5408 10296 5472
rect 10360 5408 10376 5472
rect 10440 5408 10456 5472
rect 10520 5408 10528 5472
rect 10208 5407 10528 5408
rect 19472 5472 19792 5473
rect 19472 5408 19480 5472
rect 19544 5408 19560 5472
rect 19624 5408 19640 5472
rect 19704 5408 19720 5472
rect 19784 5408 19792 5472
rect 19472 5407 19792 5408
rect 29200 5388 30000 5628
rect 0 4858 800 4948
rect 5576 4928 5896 4929
rect 5576 4864 5584 4928
rect 5648 4864 5664 4928
rect 5728 4864 5744 4928
rect 5808 4864 5824 4928
rect 5888 4864 5896 4928
rect 5576 4863 5896 4864
rect 14840 4928 15160 4929
rect 14840 4864 14848 4928
rect 14912 4864 14928 4928
rect 14992 4864 15008 4928
rect 15072 4864 15088 4928
rect 15152 4864 15160 4928
rect 14840 4863 15160 4864
rect 24104 4928 24424 4929
rect 24104 4864 24112 4928
rect 24176 4864 24192 4928
rect 24256 4864 24272 4928
rect 24336 4864 24352 4928
rect 24416 4864 24424 4928
rect 24104 4863 24424 4864
rect 2773 4858 2839 4861
rect 0 4856 2839 4858
rect 0 4800 2778 4856
rect 2834 4800 2839 4856
rect 0 4798 2839 4800
rect 0 4708 800 4798
rect 2773 4795 2839 4798
rect 26049 4858 26115 4861
rect 29200 4858 30000 4948
rect 26049 4856 30000 4858
rect 26049 4800 26054 4856
rect 26110 4800 30000 4856
rect 26049 4798 30000 4800
rect 26049 4795 26115 4798
rect 29200 4708 30000 4798
rect 10208 4384 10528 4385
rect 10208 4320 10216 4384
rect 10280 4320 10296 4384
rect 10360 4320 10376 4384
rect 10440 4320 10456 4384
rect 10520 4320 10528 4384
rect 10208 4319 10528 4320
rect 19472 4384 19792 4385
rect 19472 4320 19480 4384
rect 19544 4320 19560 4384
rect 19624 4320 19640 4384
rect 19704 4320 19720 4384
rect 19784 4320 19792 4384
rect 19472 4319 19792 4320
rect 0 4178 800 4268
rect 4061 4178 4127 4181
rect 0 4176 4127 4178
rect 0 4120 4066 4176
rect 4122 4120 4127 4176
rect 0 4118 4127 4120
rect 0 4028 800 4118
rect 4061 4115 4127 4118
rect 26141 4178 26207 4181
rect 29200 4178 30000 4268
rect 26141 4176 30000 4178
rect 26141 4120 26146 4176
rect 26202 4120 30000 4176
rect 26141 4118 30000 4120
rect 26141 4115 26207 4118
rect 29200 4028 30000 4118
rect 5576 3840 5896 3841
rect 5576 3776 5584 3840
rect 5648 3776 5664 3840
rect 5728 3776 5744 3840
rect 5808 3776 5824 3840
rect 5888 3776 5896 3840
rect 5576 3775 5896 3776
rect 14840 3840 15160 3841
rect 14840 3776 14848 3840
rect 14912 3776 14928 3840
rect 14992 3776 15008 3840
rect 15072 3776 15088 3840
rect 15152 3776 15160 3840
rect 14840 3775 15160 3776
rect 24104 3840 24424 3841
rect 24104 3776 24112 3840
rect 24176 3776 24192 3840
rect 24256 3776 24272 3840
rect 24336 3776 24352 3840
rect 24416 3776 24424 3840
rect 24104 3775 24424 3776
rect 0 3498 800 3588
rect 2957 3498 3023 3501
rect 0 3496 3023 3498
rect 0 3440 2962 3496
rect 3018 3440 3023 3496
rect 0 3438 3023 3440
rect 0 3348 800 3438
rect 2957 3435 3023 3438
rect 27429 3498 27495 3501
rect 29200 3498 30000 3588
rect 27429 3496 30000 3498
rect 27429 3440 27434 3496
rect 27490 3440 30000 3496
rect 27429 3438 30000 3440
rect 27429 3435 27495 3438
rect 29200 3348 30000 3438
rect 10208 3296 10528 3297
rect 10208 3232 10216 3296
rect 10280 3232 10296 3296
rect 10360 3232 10376 3296
rect 10440 3232 10456 3296
rect 10520 3232 10528 3296
rect 10208 3231 10528 3232
rect 19472 3296 19792 3297
rect 19472 3232 19480 3296
rect 19544 3232 19560 3296
rect 19624 3232 19640 3296
rect 19704 3232 19720 3296
rect 19784 3232 19792 3296
rect 19472 3231 19792 3232
rect 0 2818 800 2908
rect 2773 2818 2839 2821
rect 0 2816 2839 2818
rect 0 2760 2778 2816
rect 2834 2760 2839 2816
rect 0 2758 2839 2760
rect 0 2668 800 2758
rect 2773 2755 2839 2758
rect 26141 2818 26207 2821
rect 29200 2818 30000 2908
rect 26141 2816 30000 2818
rect 26141 2760 26146 2816
rect 26202 2760 30000 2816
rect 26141 2758 30000 2760
rect 26141 2755 26207 2758
rect 5576 2752 5896 2753
rect 5576 2688 5584 2752
rect 5648 2688 5664 2752
rect 5728 2688 5744 2752
rect 5808 2688 5824 2752
rect 5888 2688 5896 2752
rect 5576 2687 5896 2688
rect 14840 2752 15160 2753
rect 14840 2688 14848 2752
rect 14912 2688 14928 2752
rect 14992 2688 15008 2752
rect 15072 2688 15088 2752
rect 15152 2688 15160 2752
rect 14840 2687 15160 2688
rect 24104 2752 24424 2753
rect 24104 2688 24112 2752
rect 24176 2688 24192 2752
rect 24256 2688 24272 2752
rect 24336 2688 24352 2752
rect 24416 2688 24424 2752
rect 24104 2687 24424 2688
rect 29200 2668 30000 2758
rect 0 2138 800 2228
rect 10208 2208 10528 2209
rect 10208 2144 10216 2208
rect 10280 2144 10296 2208
rect 10360 2144 10376 2208
rect 10440 2144 10456 2208
rect 10520 2144 10528 2208
rect 10208 2143 10528 2144
rect 19472 2208 19792 2209
rect 19472 2144 19480 2208
rect 19544 2144 19560 2208
rect 19624 2144 19640 2208
rect 19704 2144 19720 2208
rect 19784 2144 19792 2208
rect 19472 2143 19792 2144
rect 3233 2138 3299 2141
rect 0 2136 3299 2138
rect 0 2080 3238 2136
rect 3294 2080 3299 2136
rect 0 2078 3299 2080
rect 0 1988 800 2078
rect 3233 2075 3299 2078
rect 26049 2138 26115 2141
rect 29200 2138 30000 2228
rect 26049 2136 30000 2138
rect 26049 2080 26054 2136
rect 26110 2080 30000 2136
rect 26049 2078 30000 2080
rect 26049 2075 26115 2078
rect 29200 1988 30000 2078
rect 0 1458 800 1548
rect 3049 1458 3115 1461
rect 0 1456 3115 1458
rect 0 1400 3054 1456
rect 3110 1400 3115 1456
rect 0 1398 3115 1400
rect 0 1308 800 1398
rect 3049 1395 3115 1398
rect 29200 1308 30000 1548
rect 0 628 800 868
rect 29200 628 30000 868
rect 26141 98 26207 101
rect 29200 98 30000 188
rect 26141 96 30000 98
rect 26141 40 26146 96
rect 26202 40 30000 96
rect 26141 38 30000 40
rect 26141 35 26207 38
rect 29200 -52 30000 38
<< via3 >>
rect 5584 39740 5648 39744
rect 5584 39684 5588 39740
rect 5588 39684 5644 39740
rect 5644 39684 5648 39740
rect 5584 39680 5648 39684
rect 5664 39740 5728 39744
rect 5664 39684 5668 39740
rect 5668 39684 5724 39740
rect 5724 39684 5728 39740
rect 5664 39680 5728 39684
rect 5744 39740 5808 39744
rect 5744 39684 5748 39740
rect 5748 39684 5804 39740
rect 5804 39684 5808 39740
rect 5744 39680 5808 39684
rect 5824 39740 5888 39744
rect 5824 39684 5828 39740
rect 5828 39684 5884 39740
rect 5884 39684 5888 39740
rect 5824 39680 5888 39684
rect 14848 39740 14912 39744
rect 14848 39684 14852 39740
rect 14852 39684 14908 39740
rect 14908 39684 14912 39740
rect 14848 39680 14912 39684
rect 14928 39740 14992 39744
rect 14928 39684 14932 39740
rect 14932 39684 14988 39740
rect 14988 39684 14992 39740
rect 14928 39680 14992 39684
rect 15008 39740 15072 39744
rect 15008 39684 15012 39740
rect 15012 39684 15068 39740
rect 15068 39684 15072 39740
rect 15008 39680 15072 39684
rect 15088 39740 15152 39744
rect 15088 39684 15092 39740
rect 15092 39684 15148 39740
rect 15148 39684 15152 39740
rect 15088 39680 15152 39684
rect 24112 39740 24176 39744
rect 24112 39684 24116 39740
rect 24116 39684 24172 39740
rect 24172 39684 24176 39740
rect 24112 39680 24176 39684
rect 24192 39740 24256 39744
rect 24192 39684 24196 39740
rect 24196 39684 24252 39740
rect 24252 39684 24256 39740
rect 24192 39680 24256 39684
rect 24272 39740 24336 39744
rect 24272 39684 24276 39740
rect 24276 39684 24332 39740
rect 24332 39684 24336 39740
rect 24272 39680 24336 39684
rect 24352 39740 24416 39744
rect 24352 39684 24356 39740
rect 24356 39684 24412 39740
rect 24412 39684 24416 39740
rect 24352 39680 24416 39684
rect 7604 39612 7668 39676
rect 11468 39204 11532 39268
rect 10216 39196 10280 39200
rect 10216 39140 10220 39196
rect 10220 39140 10276 39196
rect 10276 39140 10280 39196
rect 10216 39136 10280 39140
rect 10296 39196 10360 39200
rect 10296 39140 10300 39196
rect 10300 39140 10356 39196
rect 10356 39140 10360 39196
rect 10296 39136 10360 39140
rect 10376 39196 10440 39200
rect 10376 39140 10380 39196
rect 10380 39140 10436 39196
rect 10436 39140 10440 39196
rect 10376 39136 10440 39140
rect 10456 39196 10520 39200
rect 10456 39140 10460 39196
rect 10460 39140 10516 39196
rect 10516 39140 10520 39196
rect 10456 39136 10520 39140
rect 19480 39196 19544 39200
rect 19480 39140 19484 39196
rect 19484 39140 19540 39196
rect 19540 39140 19544 39196
rect 19480 39136 19544 39140
rect 19560 39196 19624 39200
rect 19560 39140 19564 39196
rect 19564 39140 19620 39196
rect 19620 39140 19624 39196
rect 19560 39136 19624 39140
rect 19640 39196 19704 39200
rect 19640 39140 19644 39196
rect 19644 39140 19700 39196
rect 19700 39140 19704 39196
rect 19640 39136 19704 39140
rect 19720 39196 19784 39200
rect 19720 39140 19724 39196
rect 19724 39140 19780 39196
rect 19780 39140 19784 39196
rect 19720 39136 19784 39140
rect 9996 38660 10060 38724
rect 5584 38652 5648 38656
rect 5584 38596 5588 38652
rect 5588 38596 5644 38652
rect 5644 38596 5648 38652
rect 5584 38592 5648 38596
rect 5664 38652 5728 38656
rect 5664 38596 5668 38652
rect 5668 38596 5724 38652
rect 5724 38596 5728 38652
rect 5664 38592 5728 38596
rect 5744 38652 5808 38656
rect 5744 38596 5748 38652
rect 5748 38596 5804 38652
rect 5804 38596 5808 38652
rect 5744 38592 5808 38596
rect 5824 38652 5888 38656
rect 5824 38596 5828 38652
rect 5828 38596 5884 38652
rect 5884 38596 5888 38652
rect 5824 38592 5888 38596
rect 9260 38524 9324 38588
rect 12020 38524 12084 38588
rect 14848 38652 14912 38656
rect 14848 38596 14852 38652
rect 14852 38596 14908 38652
rect 14908 38596 14912 38652
rect 14848 38592 14912 38596
rect 14928 38652 14992 38656
rect 14928 38596 14932 38652
rect 14932 38596 14988 38652
rect 14988 38596 14992 38652
rect 14928 38592 14992 38596
rect 15008 38652 15072 38656
rect 15008 38596 15012 38652
rect 15012 38596 15068 38652
rect 15068 38596 15072 38652
rect 15008 38592 15072 38596
rect 15088 38652 15152 38656
rect 15088 38596 15092 38652
rect 15092 38596 15148 38652
rect 15148 38596 15152 38652
rect 15088 38592 15152 38596
rect 24112 38652 24176 38656
rect 24112 38596 24116 38652
rect 24116 38596 24172 38652
rect 24172 38596 24176 38652
rect 24112 38592 24176 38596
rect 24192 38652 24256 38656
rect 24192 38596 24196 38652
rect 24196 38596 24252 38652
rect 24252 38596 24256 38652
rect 24192 38592 24256 38596
rect 24272 38652 24336 38656
rect 24272 38596 24276 38652
rect 24276 38596 24332 38652
rect 24332 38596 24336 38652
rect 24272 38592 24336 38596
rect 24352 38652 24416 38656
rect 24352 38596 24356 38652
rect 24356 38596 24412 38652
rect 24412 38596 24416 38652
rect 24352 38592 24416 38596
rect 19932 38252 19996 38316
rect 10216 38108 10280 38112
rect 10216 38052 10220 38108
rect 10220 38052 10276 38108
rect 10276 38052 10280 38108
rect 10216 38048 10280 38052
rect 10296 38108 10360 38112
rect 10296 38052 10300 38108
rect 10300 38052 10356 38108
rect 10356 38052 10360 38108
rect 10296 38048 10360 38052
rect 10376 38108 10440 38112
rect 10376 38052 10380 38108
rect 10380 38052 10436 38108
rect 10436 38052 10440 38108
rect 10376 38048 10440 38052
rect 10456 38108 10520 38112
rect 10456 38052 10460 38108
rect 10460 38052 10516 38108
rect 10516 38052 10520 38108
rect 10456 38048 10520 38052
rect 19480 38108 19544 38112
rect 19480 38052 19484 38108
rect 19484 38052 19540 38108
rect 19540 38052 19544 38108
rect 19480 38048 19544 38052
rect 19560 38108 19624 38112
rect 19560 38052 19564 38108
rect 19564 38052 19620 38108
rect 19620 38052 19624 38108
rect 19560 38048 19624 38052
rect 19640 38108 19704 38112
rect 19640 38052 19644 38108
rect 19644 38052 19700 38108
rect 19700 38052 19704 38108
rect 19640 38048 19704 38052
rect 19720 38108 19784 38112
rect 19720 38052 19724 38108
rect 19724 38052 19780 38108
rect 19780 38052 19784 38108
rect 19720 38048 19784 38052
rect 10732 37980 10796 38044
rect 12204 37708 12268 37772
rect 5584 37564 5648 37568
rect 5584 37508 5588 37564
rect 5588 37508 5644 37564
rect 5644 37508 5648 37564
rect 5584 37504 5648 37508
rect 5664 37564 5728 37568
rect 5664 37508 5668 37564
rect 5668 37508 5724 37564
rect 5724 37508 5728 37564
rect 5664 37504 5728 37508
rect 5744 37564 5808 37568
rect 5744 37508 5748 37564
rect 5748 37508 5804 37564
rect 5804 37508 5808 37564
rect 5744 37504 5808 37508
rect 5824 37564 5888 37568
rect 5824 37508 5828 37564
rect 5828 37508 5884 37564
rect 5884 37508 5888 37564
rect 5824 37504 5888 37508
rect 14848 37564 14912 37568
rect 14848 37508 14852 37564
rect 14852 37508 14908 37564
rect 14908 37508 14912 37564
rect 14848 37504 14912 37508
rect 14928 37564 14992 37568
rect 14928 37508 14932 37564
rect 14932 37508 14988 37564
rect 14988 37508 14992 37564
rect 14928 37504 14992 37508
rect 15008 37564 15072 37568
rect 15008 37508 15012 37564
rect 15012 37508 15068 37564
rect 15068 37508 15072 37564
rect 15008 37504 15072 37508
rect 15088 37564 15152 37568
rect 15088 37508 15092 37564
rect 15092 37508 15148 37564
rect 15148 37508 15152 37564
rect 15088 37504 15152 37508
rect 24112 37564 24176 37568
rect 24112 37508 24116 37564
rect 24116 37508 24172 37564
rect 24172 37508 24176 37564
rect 24112 37504 24176 37508
rect 24192 37564 24256 37568
rect 24192 37508 24196 37564
rect 24196 37508 24252 37564
rect 24252 37508 24256 37564
rect 24192 37504 24256 37508
rect 24272 37564 24336 37568
rect 24272 37508 24276 37564
rect 24276 37508 24332 37564
rect 24332 37508 24336 37564
rect 24272 37504 24336 37508
rect 24352 37564 24416 37568
rect 24352 37508 24356 37564
rect 24356 37508 24412 37564
rect 24412 37508 24416 37564
rect 24352 37504 24416 37508
rect 19196 37300 19260 37364
rect 9628 37028 9692 37092
rect 11652 37028 11716 37092
rect 14044 37028 14108 37092
rect 10216 37020 10280 37024
rect 10216 36964 10220 37020
rect 10220 36964 10276 37020
rect 10276 36964 10280 37020
rect 10216 36960 10280 36964
rect 10296 37020 10360 37024
rect 10296 36964 10300 37020
rect 10300 36964 10356 37020
rect 10356 36964 10360 37020
rect 10296 36960 10360 36964
rect 10376 37020 10440 37024
rect 10376 36964 10380 37020
rect 10380 36964 10436 37020
rect 10436 36964 10440 37020
rect 10376 36960 10440 36964
rect 10456 37020 10520 37024
rect 10456 36964 10460 37020
rect 10460 36964 10516 37020
rect 10516 36964 10520 37020
rect 10456 36960 10520 36964
rect 10916 36756 10980 36820
rect 12204 36620 12268 36684
rect 5584 36476 5648 36480
rect 5584 36420 5588 36476
rect 5588 36420 5644 36476
rect 5644 36420 5648 36476
rect 5584 36416 5648 36420
rect 5664 36476 5728 36480
rect 5664 36420 5668 36476
rect 5668 36420 5724 36476
rect 5724 36420 5728 36476
rect 5664 36416 5728 36420
rect 5744 36476 5808 36480
rect 5744 36420 5748 36476
rect 5748 36420 5804 36476
rect 5804 36420 5808 36476
rect 5744 36416 5808 36420
rect 5824 36476 5888 36480
rect 5824 36420 5828 36476
rect 5828 36420 5884 36476
rect 5884 36420 5888 36476
rect 5824 36416 5888 36420
rect 11652 36348 11716 36412
rect 20116 37164 20180 37228
rect 19480 37020 19544 37024
rect 19480 36964 19484 37020
rect 19484 36964 19540 37020
rect 19540 36964 19544 37020
rect 19480 36960 19544 36964
rect 19560 37020 19624 37024
rect 19560 36964 19564 37020
rect 19564 36964 19620 37020
rect 19620 36964 19624 37020
rect 19560 36960 19624 36964
rect 19640 37020 19704 37024
rect 19640 36964 19644 37020
rect 19644 36964 19700 37020
rect 19700 36964 19704 37020
rect 19640 36960 19704 36964
rect 19720 37020 19784 37024
rect 19720 36964 19724 37020
rect 19724 36964 19780 37020
rect 19780 36964 19784 37020
rect 19720 36960 19784 36964
rect 19932 36892 19996 36956
rect 14848 36476 14912 36480
rect 14848 36420 14852 36476
rect 14852 36420 14908 36476
rect 14908 36420 14912 36476
rect 14848 36416 14912 36420
rect 14928 36476 14992 36480
rect 14928 36420 14932 36476
rect 14932 36420 14988 36476
rect 14988 36420 14992 36476
rect 14928 36416 14992 36420
rect 15008 36476 15072 36480
rect 15008 36420 15012 36476
rect 15012 36420 15068 36476
rect 15068 36420 15072 36476
rect 15008 36416 15072 36420
rect 15088 36476 15152 36480
rect 15088 36420 15092 36476
rect 15092 36420 15148 36476
rect 15148 36420 15152 36476
rect 15088 36416 15152 36420
rect 24112 36476 24176 36480
rect 24112 36420 24116 36476
rect 24116 36420 24172 36476
rect 24172 36420 24176 36476
rect 24112 36416 24176 36420
rect 24192 36476 24256 36480
rect 24192 36420 24196 36476
rect 24196 36420 24252 36476
rect 24252 36420 24256 36476
rect 24192 36416 24256 36420
rect 24272 36476 24336 36480
rect 24272 36420 24276 36476
rect 24276 36420 24332 36476
rect 24332 36420 24336 36476
rect 24272 36416 24336 36420
rect 24352 36476 24416 36480
rect 24352 36420 24356 36476
rect 24356 36420 24412 36476
rect 24412 36420 24416 36476
rect 24352 36416 24416 36420
rect 12204 36348 12268 36412
rect 9812 36272 9876 36276
rect 9812 36216 9826 36272
rect 9826 36216 9876 36272
rect 9812 36212 9876 36216
rect 12020 36212 12084 36276
rect 13860 36212 13924 36276
rect 11836 36076 11900 36140
rect 11468 35940 11532 36004
rect 18644 36076 18708 36140
rect 19196 35940 19260 36004
rect 10216 35932 10280 35936
rect 10216 35876 10220 35932
rect 10220 35876 10276 35932
rect 10276 35876 10280 35932
rect 10216 35872 10280 35876
rect 10296 35932 10360 35936
rect 10296 35876 10300 35932
rect 10300 35876 10356 35932
rect 10356 35876 10360 35932
rect 10296 35872 10360 35876
rect 10376 35932 10440 35936
rect 10376 35876 10380 35932
rect 10380 35876 10436 35932
rect 10436 35876 10440 35932
rect 10376 35872 10440 35876
rect 10456 35932 10520 35936
rect 10456 35876 10460 35932
rect 10460 35876 10516 35932
rect 10516 35876 10520 35932
rect 10456 35872 10520 35876
rect 19480 35932 19544 35936
rect 19480 35876 19484 35932
rect 19484 35876 19540 35932
rect 19540 35876 19544 35932
rect 19480 35872 19544 35876
rect 19560 35932 19624 35936
rect 19560 35876 19564 35932
rect 19564 35876 19620 35932
rect 19620 35876 19624 35932
rect 19560 35872 19624 35876
rect 19640 35932 19704 35936
rect 19640 35876 19644 35932
rect 19644 35876 19700 35932
rect 19700 35876 19704 35932
rect 19640 35872 19704 35876
rect 19720 35932 19784 35936
rect 19720 35876 19724 35932
rect 19724 35876 19780 35932
rect 19780 35876 19784 35932
rect 19720 35872 19784 35876
rect 12388 35804 12452 35868
rect 7604 35728 7668 35732
rect 7604 35672 7618 35728
rect 7618 35672 7668 35728
rect 7604 35668 7668 35672
rect 21036 35728 21100 35732
rect 21036 35672 21050 35728
rect 21050 35672 21100 35728
rect 21036 35668 21100 35672
rect 5584 35388 5648 35392
rect 5584 35332 5588 35388
rect 5588 35332 5644 35388
rect 5644 35332 5648 35388
rect 5584 35328 5648 35332
rect 5664 35388 5728 35392
rect 5664 35332 5668 35388
rect 5668 35332 5724 35388
rect 5724 35332 5728 35388
rect 5664 35328 5728 35332
rect 5744 35388 5808 35392
rect 5744 35332 5748 35388
rect 5748 35332 5804 35388
rect 5804 35332 5808 35388
rect 5744 35328 5808 35332
rect 5824 35388 5888 35392
rect 5824 35332 5828 35388
rect 5828 35332 5884 35388
rect 5884 35332 5888 35388
rect 5824 35328 5888 35332
rect 14848 35388 14912 35392
rect 14848 35332 14852 35388
rect 14852 35332 14908 35388
rect 14908 35332 14912 35388
rect 14848 35328 14912 35332
rect 14928 35388 14992 35392
rect 14928 35332 14932 35388
rect 14932 35332 14988 35388
rect 14988 35332 14992 35388
rect 14928 35328 14992 35332
rect 15008 35388 15072 35392
rect 15008 35332 15012 35388
rect 15012 35332 15068 35388
rect 15068 35332 15072 35388
rect 15008 35328 15072 35332
rect 15088 35388 15152 35392
rect 15088 35332 15092 35388
rect 15092 35332 15148 35388
rect 15148 35332 15152 35388
rect 15088 35328 15152 35332
rect 24112 35388 24176 35392
rect 24112 35332 24116 35388
rect 24116 35332 24172 35388
rect 24172 35332 24176 35388
rect 24112 35328 24176 35332
rect 24192 35388 24256 35392
rect 24192 35332 24196 35388
rect 24196 35332 24252 35388
rect 24252 35332 24256 35388
rect 24192 35328 24256 35332
rect 24272 35388 24336 35392
rect 24272 35332 24276 35388
rect 24276 35332 24332 35388
rect 24332 35332 24336 35388
rect 24272 35328 24336 35332
rect 24352 35388 24416 35392
rect 24352 35332 24356 35388
rect 24356 35332 24412 35388
rect 24412 35332 24416 35388
rect 24352 35328 24416 35332
rect 9260 35320 9324 35324
rect 9260 35264 9274 35320
rect 9274 35264 9324 35320
rect 9260 35260 9324 35264
rect 12020 35260 12084 35324
rect 9812 35124 9876 35188
rect 13492 34988 13556 35052
rect 18644 35124 18708 35188
rect 10732 34852 10796 34916
rect 10216 34844 10280 34848
rect 10216 34788 10220 34844
rect 10220 34788 10276 34844
rect 10276 34788 10280 34844
rect 10216 34784 10280 34788
rect 10296 34844 10360 34848
rect 10296 34788 10300 34844
rect 10300 34788 10356 34844
rect 10356 34788 10360 34844
rect 10296 34784 10360 34788
rect 10376 34844 10440 34848
rect 10376 34788 10380 34844
rect 10380 34788 10436 34844
rect 10436 34788 10440 34844
rect 10376 34784 10440 34788
rect 10456 34844 10520 34848
rect 10456 34788 10460 34844
rect 10460 34788 10516 34844
rect 10516 34788 10520 34844
rect 10456 34784 10520 34788
rect 19480 34844 19544 34848
rect 19480 34788 19484 34844
rect 19484 34788 19540 34844
rect 19540 34788 19544 34844
rect 19480 34784 19544 34788
rect 19560 34844 19624 34848
rect 19560 34788 19564 34844
rect 19564 34788 19620 34844
rect 19620 34788 19624 34844
rect 19560 34784 19624 34788
rect 19640 34844 19704 34848
rect 19640 34788 19644 34844
rect 19644 34788 19700 34844
rect 19700 34788 19704 34844
rect 19640 34784 19704 34788
rect 19720 34844 19784 34848
rect 19720 34788 19724 34844
rect 19724 34788 19780 34844
rect 19780 34788 19784 34844
rect 19720 34784 19784 34788
rect 9812 34716 9876 34780
rect 11468 34716 11532 34780
rect 12204 34716 12268 34780
rect 7236 34580 7300 34644
rect 19932 34308 19996 34372
rect 21036 34308 21100 34372
rect 5584 34300 5648 34304
rect 5584 34244 5588 34300
rect 5588 34244 5644 34300
rect 5644 34244 5648 34300
rect 5584 34240 5648 34244
rect 5664 34300 5728 34304
rect 5664 34244 5668 34300
rect 5668 34244 5724 34300
rect 5724 34244 5728 34300
rect 5664 34240 5728 34244
rect 5744 34300 5808 34304
rect 5744 34244 5748 34300
rect 5748 34244 5804 34300
rect 5804 34244 5808 34300
rect 5744 34240 5808 34244
rect 5824 34300 5888 34304
rect 5824 34244 5828 34300
rect 5828 34244 5884 34300
rect 5884 34244 5888 34300
rect 5824 34240 5888 34244
rect 14848 34300 14912 34304
rect 14848 34244 14852 34300
rect 14852 34244 14908 34300
rect 14908 34244 14912 34300
rect 14848 34240 14912 34244
rect 14928 34300 14992 34304
rect 14928 34244 14932 34300
rect 14932 34244 14988 34300
rect 14988 34244 14992 34300
rect 14928 34240 14992 34244
rect 15008 34300 15072 34304
rect 15008 34244 15012 34300
rect 15012 34244 15068 34300
rect 15068 34244 15072 34300
rect 15008 34240 15072 34244
rect 15088 34300 15152 34304
rect 15088 34244 15092 34300
rect 15092 34244 15148 34300
rect 15148 34244 15152 34300
rect 15088 34240 15152 34244
rect 24112 34300 24176 34304
rect 24112 34244 24116 34300
rect 24116 34244 24172 34300
rect 24172 34244 24176 34300
rect 24112 34240 24176 34244
rect 24192 34300 24256 34304
rect 24192 34244 24196 34300
rect 24196 34244 24252 34300
rect 24252 34244 24256 34300
rect 24192 34240 24256 34244
rect 24272 34300 24336 34304
rect 24272 34244 24276 34300
rect 24276 34244 24332 34300
rect 24332 34244 24336 34300
rect 24272 34240 24336 34244
rect 24352 34300 24416 34304
rect 24352 34244 24356 34300
rect 24356 34244 24412 34300
rect 24412 34244 24416 34300
rect 24352 34240 24416 34244
rect 10916 34172 10980 34236
rect 10732 34036 10796 34100
rect 12020 34172 12084 34236
rect 16436 34172 16500 34236
rect 12388 33900 12452 33964
rect 9628 33764 9692 33828
rect 10216 33756 10280 33760
rect 10216 33700 10220 33756
rect 10220 33700 10276 33756
rect 10276 33700 10280 33756
rect 10216 33696 10280 33700
rect 10296 33756 10360 33760
rect 10296 33700 10300 33756
rect 10300 33700 10356 33756
rect 10356 33700 10360 33756
rect 10296 33696 10360 33700
rect 10376 33756 10440 33760
rect 10376 33700 10380 33756
rect 10380 33700 10436 33756
rect 10436 33700 10440 33756
rect 10376 33696 10440 33700
rect 10456 33756 10520 33760
rect 10456 33700 10460 33756
rect 10460 33700 10516 33756
rect 10516 33700 10520 33756
rect 10456 33696 10520 33700
rect 19480 33756 19544 33760
rect 19480 33700 19484 33756
rect 19484 33700 19540 33756
rect 19540 33700 19544 33756
rect 19480 33696 19544 33700
rect 19560 33756 19624 33760
rect 19560 33700 19564 33756
rect 19564 33700 19620 33756
rect 19620 33700 19624 33756
rect 19560 33696 19624 33700
rect 19640 33756 19704 33760
rect 19640 33700 19644 33756
rect 19644 33700 19700 33756
rect 19700 33700 19704 33756
rect 19640 33696 19704 33700
rect 19720 33756 19784 33760
rect 19720 33700 19724 33756
rect 19724 33700 19780 33756
rect 19780 33700 19784 33756
rect 19720 33696 19784 33700
rect 13124 33628 13188 33692
rect 14412 33492 14476 33556
rect 10916 33220 10980 33284
rect 11468 33220 11532 33284
rect 11652 33220 11716 33284
rect 13492 33220 13556 33284
rect 5584 33212 5648 33216
rect 5584 33156 5588 33212
rect 5588 33156 5644 33212
rect 5644 33156 5648 33212
rect 5584 33152 5648 33156
rect 5664 33212 5728 33216
rect 5664 33156 5668 33212
rect 5668 33156 5724 33212
rect 5724 33156 5728 33212
rect 5664 33152 5728 33156
rect 5744 33212 5808 33216
rect 5744 33156 5748 33212
rect 5748 33156 5804 33212
rect 5804 33156 5808 33212
rect 5744 33152 5808 33156
rect 5824 33212 5888 33216
rect 5824 33156 5828 33212
rect 5828 33156 5884 33212
rect 5884 33156 5888 33212
rect 5824 33152 5888 33156
rect 14848 33212 14912 33216
rect 14848 33156 14852 33212
rect 14852 33156 14908 33212
rect 14908 33156 14912 33212
rect 14848 33152 14912 33156
rect 14928 33212 14992 33216
rect 14928 33156 14932 33212
rect 14932 33156 14988 33212
rect 14988 33156 14992 33212
rect 14928 33152 14992 33156
rect 15008 33212 15072 33216
rect 15008 33156 15012 33212
rect 15012 33156 15068 33212
rect 15068 33156 15072 33212
rect 15008 33152 15072 33156
rect 15088 33212 15152 33216
rect 15088 33156 15092 33212
rect 15092 33156 15148 33212
rect 15148 33156 15152 33212
rect 15088 33152 15152 33156
rect 24112 33212 24176 33216
rect 24112 33156 24116 33212
rect 24116 33156 24172 33212
rect 24172 33156 24176 33212
rect 24112 33152 24176 33156
rect 24192 33212 24256 33216
rect 24192 33156 24196 33212
rect 24196 33156 24252 33212
rect 24252 33156 24256 33212
rect 24192 33152 24256 33156
rect 24272 33212 24336 33216
rect 24272 33156 24276 33212
rect 24276 33156 24332 33212
rect 24332 33156 24336 33212
rect 24272 33152 24336 33156
rect 24352 33212 24416 33216
rect 24352 33156 24356 33212
rect 24356 33156 24412 33212
rect 24412 33156 24416 33212
rect 24352 33152 24416 33156
rect 9812 33084 9876 33148
rect 12572 32948 12636 33012
rect 10216 32668 10280 32672
rect 10216 32612 10220 32668
rect 10220 32612 10276 32668
rect 10276 32612 10280 32668
rect 10216 32608 10280 32612
rect 10296 32668 10360 32672
rect 10296 32612 10300 32668
rect 10300 32612 10356 32668
rect 10356 32612 10360 32668
rect 10296 32608 10360 32612
rect 10376 32668 10440 32672
rect 10376 32612 10380 32668
rect 10380 32612 10436 32668
rect 10436 32612 10440 32668
rect 10376 32608 10440 32612
rect 10456 32668 10520 32672
rect 10456 32612 10460 32668
rect 10460 32612 10516 32668
rect 10516 32612 10520 32668
rect 10456 32608 10520 32612
rect 19480 32668 19544 32672
rect 19480 32612 19484 32668
rect 19484 32612 19540 32668
rect 19540 32612 19544 32668
rect 19480 32608 19544 32612
rect 19560 32668 19624 32672
rect 19560 32612 19564 32668
rect 19564 32612 19620 32668
rect 19620 32612 19624 32668
rect 19560 32608 19624 32612
rect 19640 32668 19704 32672
rect 19640 32612 19644 32668
rect 19644 32612 19700 32668
rect 19700 32612 19704 32668
rect 19640 32608 19704 32612
rect 19720 32668 19784 32672
rect 19720 32612 19724 32668
rect 19724 32612 19780 32668
rect 19780 32612 19784 32668
rect 19720 32608 19784 32612
rect 13492 32540 13556 32604
rect 11284 32132 11348 32196
rect 11468 32132 11532 32196
rect 5584 32124 5648 32128
rect 5584 32068 5588 32124
rect 5588 32068 5644 32124
rect 5644 32068 5648 32124
rect 5584 32064 5648 32068
rect 5664 32124 5728 32128
rect 5664 32068 5668 32124
rect 5668 32068 5724 32124
rect 5724 32068 5728 32124
rect 5664 32064 5728 32068
rect 5744 32124 5808 32128
rect 5744 32068 5748 32124
rect 5748 32068 5804 32124
rect 5804 32068 5808 32124
rect 5744 32064 5808 32068
rect 5824 32124 5888 32128
rect 5824 32068 5828 32124
rect 5828 32068 5884 32124
rect 5884 32068 5888 32124
rect 5824 32064 5888 32068
rect 14848 32124 14912 32128
rect 14848 32068 14852 32124
rect 14852 32068 14908 32124
rect 14908 32068 14912 32124
rect 14848 32064 14912 32068
rect 14928 32124 14992 32128
rect 14928 32068 14932 32124
rect 14932 32068 14988 32124
rect 14988 32068 14992 32124
rect 14928 32064 14992 32068
rect 15008 32124 15072 32128
rect 15008 32068 15012 32124
rect 15012 32068 15068 32124
rect 15068 32068 15072 32124
rect 15008 32064 15072 32068
rect 15088 32124 15152 32128
rect 15088 32068 15092 32124
rect 15092 32068 15148 32124
rect 15148 32068 15152 32124
rect 15088 32064 15152 32068
rect 24112 32124 24176 32128
rect 24112 32068 24116 32124
rect 24116 32068 24172 32124
rect 24172 32068 24176 32124
rect 24112 32064 24176 32068
rect 24192 32124 24256 32128
rect 24192 32068 24196 32124
rect 24196 32068 24252 32124
rect 24252 32068 24256 32124
rect 24192 32064 24256 32068
rect 24272 32124 24336 32128
rect 24272 32068 24276 32124
rect 24276 32068 24332 32124
rect 24332 32068 24336 32124
rect 24272 32064 24336 32068
rect 24352 32124 24416 32128
rect 24352 32068 24356 32124
rect 24356 32068 24412 32124
rect 24412 32068 24416 32124
rect 24352 32064 24416 32068
rect 13308 31860 13372 31924
rect 19932 31996 19996 32060
rect 10216 31580 10280 31584
rect 10216 31524 10220 31580
rect 10220 31524 10276 31580
rect 10276 31524 10280 31580
rect 10216 31520 10280 31524
rect 10296 31580 10360 31584
rect 10296 31524 10300 31580
rect 10300 31524 10356 31580
rect 10356 31524 10360 31580
rect 10296 31520 10360 31524
rect 10376 31580 10440 31584
rect 10376 31524 10380 31580
rect 10380 31524 10436 31580
rect 10436 31524 10440 31580
rect 10376 31520 10440 31524
rect 10456 31580 10520 31584
rect 10456 31524 10460 31580
rect 10460 31524 10516 31580
rect 10516 31524 10520 31580
rect 10456 31520 10520 31524
rect 20116 31724 20180 31788
rect 11284 31588 11348 31652
rect 19480 31580 19544 31584
rect 19480 31524 19484 31580
rect 19484 31524 19540 31580
rect 19540 31524 19544 31580
rect 19480 31520 19544 31524
rect 19560 31580 19624 31584
rect 19560 31524 19564 31580
rect 19564 31524 19620 31580
rect 19620 31524 19624 31580
rect 19560 31520 19624 31524
rect 19640 31580 19704 31584
rect 19640 31524 19644 31580
rect 19644 31524 19700 31580
rect 19700 31524 19704 31580
rect 19640 31520 19704 31524
rect 19720 31580 19784 31584
rect 19720 31524 19724 31580
rect 19724 31524 19780 31580
rect 19780 31524 19784 31580
rect 19720 31520 19784 31524
rect 13860 31316 13924 31380
rect 9812 31044 9876 31108
rect 10732 31044 10796 31108
rect 5584 31036 5648 31040
rect 5584 30980 5588 31036
rect 5588 30980 5644 31036
rect 5644 30980 5648 31036
rect 5584 30976 5648 30980
rect 5664 31036 5728 31040
rect 5664 30980 5668 31036
rect 5668 30980 5724 31036
rect 5724 30980 5728 31036
rect 5664 30976 5728 30980
rect 5744 31036 5808 31040
rect 5744 30980 5748 31036
rect 5748 30980 5804 31036
rect 5804 30980 5808 31036
rect 5744 30976 5808 30980
rect 5824 31036 5888 31040
rect 5824 30980 5828 31036
rect 5828 30980 5884 31036
rect 5884 30980 5888 31036
rect 5824 30976 5888 30980
rect 14848 31036 14912 31040
rect 14848 30980 14852 31036
rect 14852 30980 14908 31036
rect 14908 30980 14912 31036
rect 14848 30976 14912 30980
rect 14928 31036 14992 31040
rect 14928 30980 14932 31036
rect 14932 30980 14988 31036
rect 14988 30980 14992 31036
rect 14928 30976 14992 30980
rect 15008 31036 15072 31040
rect 15008 30980 15012 31036
rect 15012 30980 15068 31036
rect 15068 30980 15072 31036
rect 15008 30976 15072 30980
rect 15088 31036 15152 31040
rect 15088 30980 15092 31036
rect 15092 30980 15148 31036
rect 15148 30980 15152 31036
rect 15088 30976 15152 30980
rect 24112 31036 24176 31040
rect 24112 30980 24116 31036
rect 24116 30980 24172 31036
rect 24172 30980 24176 31036
rect 24112 30976 24176 30980
rect 24192 31036 24256 31040
rect 24192 30980 24196 31036
rect 24196 30980 24252 31036
rect 24252 30980 24256 31036
rect 24192 30976 24256 30980
rect 24272 31036 24336 31040
rect 24272 30980 24276 31036
rect 24276 30980 24332 31036
rect 24332 30980 24336 31036
rect 24272 30976 24336 30980
rect 24352 31036 24416 31040
rect 24352 30980 24356 31036
rect 24356 30980 24412 31036
rect 24412 30980 24416 31036
rect 24352 30976 24416 30980
rect 10916 30908 10980 30972
rect 10216 30492 10280 30496
rect 10216 30436 10220 30492
rect 10220 30436 10276 30492
rect 10276 30436 10280 30492
rect 10216 30432 10280 30436
rect 10296 30492 10360 30496
rect 10296 30436 10300 30492
rect 10300 30436 10356 30492
rect 10356 30436 10360 30492
rect 10296 30432 10360 30436
rect 10376 30492 10440 30496
rect 10376 30436 10380 30492
rect 10380 30436 10436 30492
rect 10436 30436 10440 30492
rect 10376 30432 10440 30436
rect 10456 30492 10520 30496
rect 10456 30436 10460 30492
rect 10460 30436 10516 30492
rect 10516 30436 10520 30492
rect 10456 30432 10520 30436
rect 19480 30492 19544 30496
rect 19480 30436 19484 30492
rect 19484 30436 19540 30492
rect 19540 30436 19544 30492
rect 19480 30432 19544 30436
rect 19560 30492 19624 30496
rect 19560 30436 19564 30492
rect 19564 30436 19620 30492
rect 19620 30436 19624 30492
rect 19560 30432 19624 30436
rect 19640 30492 19704 30496
rect 19640 30436 19644 30492
rect 19644 30436 19700 30492
rect 19700 30436 19704 30492
rect 19640 30432 19704 30436
rect 19720 30492 19784 30496
rect 19720 30436 19724 30492
rect 19724 30436 19780 30492
rect 19780 30436 19784 30492
rect 19720 30432 19784 30436
rect 9996 30364 10060 30428
rect 26556 30364 26620 30428
rect 16988 30228 17052 30292
rect 12204 30092 12268 30156
rect 5584 29948 5648 29952
rect 5584 29892 5588 29948
rect 5588 29892 5644 29948
rect 5644 29892 5648 29948
rect 5584 29888 5648 29892
rect 5664 29948 5728 29952
rect 5664 29892 5668 29948
rect 5668 29892 5724 29948
rect 5724 29892 5728 29948
rect 5664 29888 5728 29892
rect 5744 29948 5808 29952
rect 5744 29892 5748 29948
rect 5748 29892 5804 29948
rect 5804 29892 5808 29948
rect 5744 29888 5808 29892
rect 5824 29948 5888 29952
rect 5824 29892 5828 29948
rect 5828 29892 5884 29948
rect 5884 29892 5888 29948
rect 5824 29888 5888 29892
rect 14044 30016 14108 30020
rect 14044 29960 14094 30016
rect 14094 29960 14108 30016
rect 14044 29956 14108 29960
rect 14848 29948 14912 29952
rect 14848 29892 14852 29948
rect 14852 29892 14908 29948
rect 14908 29892 14912 29948
rect 14848 29888 14912 29892
rect 14928 29948 14992 29952
rect 14928 29892 14932 29948
rect 14932 29892 14988 29948
rect 14988 29892 14992 29948
rect 14928 29888 14992 29892
rect 15008 29948 15072 29952
rect 15008 29892 15012 29948
rect 15012 29892 15068 29948
rect 15068 29892 15072 29948
rect 15008 29888 15072 29892
rect 15088 29948 15152 29952
rect 15088 29892 15092 29948
rect 15092 29892 15148 29948
rect 15148 29892 15152 29948
rect 15088 29888 15152 29892
rect 24112 29948 24176 29952
rect 24112 29892 24116 29948
rect 24116 29892 24172 29948
rect 24172 29892 24176 29948
rect 24112 29888 24176 29892
rect 24192 29948 24256 29952
rect 24192 29892 24196 29948
rect 24196 29892 24252 29948
rect 24252 29892 24256 29948
rect 24192 29888 24256 29892
rect 24272 29948 24336 29952
rect 24272 29892 24276 29948
rect 24276 29892 24332 29948
rect 24332 29892 24336 29948
rect 24272 29888 24336 29892
rect 24352 29948 24416 29952
rect 24352 29892 24356 29948
rect 24356 29892 24412 29948
rect 24412 29892 24416 29948
rect 24352 29888 24416 29892
rect 16804 29820 16868 29884
rect 19932 29548 19996 29612
rect 11652 29412 11716 29476
rect 12204 29412 12268 29476
rect 22140 29472 22204 29476
rect 22140 29416 22154 29472
rect 22154 29416 22204 29472
rect 22140 29412 22204 29416
rect 10216 29404 10280 29408
rect 10216 29348 10220 29404
rect 10220 29348 10276 29404
rect 10276 29348 10280 29404
rect 10216 29344 10280 29348
rect 10296 29404 10360 29408
rect 10296 29348 10300 29404
rect 10300 29348 10356 29404
rect 10356 29348 10360 29404
rect 10296 29344 10360 29348
rect 10376 29404 10440 29408
rect 10376 29348 10380 29404
rect 10380 29348 10436 29404
rect 10436 29348 10440 29404
rect 10376 29344 10440 29348
rect 10456 29404 10520 29408
rect 10456 29348 10460 29404
rect 10460 29348 10516 29404
rect 10516 29348 10520 29404
rect 10456 29344 10520 29348
rect 19480 29404 19544 29408
rect 19480 29348 19484 29404
rect 19484 29348 19540 29404
rect 19540 29348 19544 29404
rect 19480 29344 19544 29348
rect 19560 29404 19624 29408
rect 19560 29348 19564 29404
rect 19564 29348 19620 29404
rect 19620 29348 19624 29404
rect 19560 29344 19624 29348
rect 19640 29404 19704 29408
rect 19640 29348 19644 29404
rect 19644 29348 19700 29404
rect 19700 29348 19704 29404
rect 19640 29344 19704 29348
rect 19720 29404 19784 29408
rect 19720 29348 19724 29404
rect 19724 29348 19780 29404
rect 19780 29348 19784 29404
rect 19720 29344 19784 29348
rect 9812 29336 9876 29340
rect 9812 29280 9826 29336
rect 9826 29280 9876 29336
rect 9812 29276 9876 29280
rect 12388 29140 12452 29204
rect 12572 28868 12636 28932
rect 18460 29004 18524 29068
rect 20116 28868 20180 28932
rect 5584 28860 5648 28864
rect 5584 28804 5588 28860
rect 5588 28804 5644 28860
rect 5644 28804 5648 28860
rect 5584 28800 5648 28804
rect 5664 28860 5728 28864
rect 5664 28804 5668 28860
rect 5668 28804 5724 28860
rect 5724 28804 5728 28860
rect 5664 28800 5728 28804
rect 5744 28860 5808 28864
rect 5744 28804 5748 28860
rect 5748 28804 5804 28860
rect 5804 28804 5808 28860
rect 5744 28800 5808 28804
rect 5824 28860 5888 28864
rect 5824 28804 5828 28860
rect 5828 28804 5884 28860
rect 5884 28804 5888 28860
rect 5824 28800 5888 28804
rect 14848 28860 14912 28864
rect 14848 28804 14852 28860
rect 14852 28804 14908 28860
rect 14908 28804 14912 28860
rect 14848 28800 14912 28804
rect 14928 28860 14992 28864
rect 14928 28804 14932 28860
rect 14932 28804 14988 28860
rect 14988 28804 14992 28860
rect 14928 28800 14992 28804
rect 15008 28860 15072 28864
rect 15008 28804 15012 28860
rect 15012 28804 15068 28860
rect 15068 28804 15072 28860
rect 15008 28800 15072 28804
rect 15088 28860 15152 28864
rect 15088 28804 15092 28860
rect 15092 28804 15148 28860
rect 15148 28804 15152 28860
rect 15088 28800 15152 28804
rect 24112 28860 24176 28864
rect 24112 28804 24116 28860
rect 24116 28804 24172 28860
rect 24172 28804 24176 28860
rect 24112 28800 24176 28804
rect 24192 28860 24256 28864
rect 24192 28804 24196 28860
rect 24196 28804 24252 28860
rect 24252 28804 24256 28860
rect 24192 28800 24256 28804
rect 24272 28860 24336 28864
rect 24272 28804 24276 28860
rect 24276 28804 24332 28860
rect 24332 28804 24336 28860
rect 24272 28800 24336 28804
rect 24352 28860 24416 28864
rect 24352 28804 24356 28860
rect 24356 28804 24412 28860
rect 24412 28804 24416 28860
rect 24352 28800 24416 28804
rect 16988 28656 17052 28660
rect 16988 28600 17002 28656
rect 17002 28600 17052 28656
rect 16988 28596 17052 28600
rect 19932 28596 19996 28660
rect 10216 28316 10280 28320
rect 10216 28260 10220 28316
rect 10220 28260 10276 28316
rect 10276 28260 10280 28316
rect 10216 28256 10280 28260
rect 10296 28316 10360 28320
rect 10296 28260 10300 28316
rect 10300 28260 10356 28316
rect 10356 28260 10360 28316
rect 10296 28256 10360 28260
rect 10376 28316 10440 28320
rect 10376 28260 10380 28316
rect 10380 28260 10436 28316
rect 10436 28260 10440 28316
rect 10376 28256 10440 28260
rect 10456 28316 10520 28320
rect 10456 28260 10460 28316
rect 10460 28260 10516 28316
rect 10516 28260 10520 28316
rect 10456 28256 10520 28260
rect 19480 28316 19544 28320
rect 19480 28260 19484 28316
rect 19484 28260 19540 28316
rect 19540 28260 19544 28316
rect 19480 28256 19544 28260
rect 19560 28316 19624 28320
rect 19560 28260 19564 28316
rect 19564 28260 19620 28316
rect 19620 28260 19624 28316
rect 19560 28256 19624 28260
rect 19640 28316 19704 28320
rect 19640 28260 19644 28316
rect 19644 28260 19700 28316
rect 19700 28260 19704 28316
rect 19640 28256 19704 28260
rect 19720 28316 19784 28320
rect 19720 28260 19724 28316
rect 19724 28260 19780 28316
rect 19780 28260 19784 28316
rect 19720 28256 19784 28260
rect 24532 28188 24596 28252
rect 12756 27916 12820 27980
rect 5584 27772 5648 27776
rect 5584 27716 5588 27772
rect 5588 27716 5644 27772
rect 5644 27716 5648 27772
rect 5584 27712 5648 27716
rect 5664 27772 5728 27776
rect 5664 27716 5668 27772
rect 5668 27716 5724 27772
rect 5724 27716 5728 27772
rect 5664 27712 5728 27716
rect 5744 27772 5808 27776
rect 5744 27716 5748 27772
rect 5748 27716 5804 27772
rect 5804 27716 5808 27772
rect 5744 27712 5808 27716
rect 5824 27772 5888 27776
rect 5824 27716 5828 27772
rect 5828 27716 5884 27772
rect 5884 27716 5888 27772
rect 5824 27712 5888 27716
rect 14848 27772 14912 27776
rect 14848 27716 14852 27772
rect 14852 27716 14908 27772
rect 14908 27716 14912 27772
rect 14848 27712 14912 27716
rect 14928 27772 14992 27776
rect 14928 27716 14932 27772
rect 14932 27716 14988 27772
rect 14988 27716 14992 27772
rect 14928 27712 14992 27716
rect 15008 27772 15072 27776
rect 15008 27716 15012 27772
rect 15012 27716 15068 27772
rect 15068 27716 15072 27772
rect 15008 27712 15072 27716
rect 15088 27772 15152 27776
rect 15088 27716 15092 27772
rect 15092 27716 15148 27772
rect 15148 27716 15152 27772
rect 15088 27712 15152 27716
rect 24112 27772 24176 27776
rect 24112 27716 24116 27772
rect 24116 27716 24172 27772
rect 24172 27716 24176 27772
rect 24112 27712 24176 27716
rect 24192 27772 24256 27776
rect 24192 27716 24196 27772
rect 24196 27716 24252 27772
rect 24252 27716 24256 27772
rect 24192 27712 24256 27716
rect 24272 27772 24336 27776
rect 24272 27716 24276 27772
rect 24276 27716 24332 27772
rect 24332 27716 24336 27772
rect 24272 27712 24336 27716
rect 24352 27772 24416 27776
rect 24352 27716 24356 27772
rect 24356 27716 24412 27772
rect 24412 27716 24416 27772
rect 24352 27712 24416 27716
rect 26188 27644 26252 27708
rect 16436 27508 16500 27572
rect 10216 27228 10280 27232
rect 10216 27172 10220 27228
rect 10220 27172 10276 27228
rect 10276 27172 10280 27228
rect 10216 27168 10280 27172
rect 10296 27228 10360 27232
rect 10296 27172 10300 27228
rect 10300 27172 10356 27228
rect 10356 27172 10360 27228
rect 10296 27168 10360 27172
rect 10376 27228 10440 27232
rect 10376 27172 10380 27228
rect 10380 27172 10436 27228
rect 10436 27172 10440 27228
rect 10376 27168 10440 27172
rect 10456 27228 10520 27232
rect 10456 27172 10460 27228
rect 10460 27172 10516 27228
rect 10516 27172 10520 27228
rect 10456 27168 10520 27172
rect 12756 27100 12820 27164
rect 12940 27100 13004 27164
rect 19480 27228 19544 27232
rect 19480 27172 19484 27228
rect 19484 27172 19540 27228
rect 19540 27172 19544 27228
rect 19480 27168 19544 27172
rect 19560 27228 19624 27232
rect 19560 27172 19564 27228
rect 19564 27172 19620 27228
rect 19620 27172 19624 27228
rect 19560 27168 19624 27172
rect 19640 27228 19704 27232
rect 19640 27172 19644 27228
rect 19644 27172 19700 27228
rect 19700 27172 19704 27228
rect 19640 27168 19704 27172
rect 19720 27228 19784 27232
rect 19720 27172 19724 27228
rect 19724 27172 19780 27228
rect 19780 27172 19784 27228
rect 19720 27168 19784 27172
rect 5584 26684 5648 26688
rect 5584 26628 5588 26684
rect 5588 26628 5644 26684
rect 5644 26628 5648 26684
rect 5584 26624 5648 26628
rect 5664 26684 5728 26688
rect 5664 26628 5668 26684
rect 5668 26628 5724 26684
rect 5724 26628 5728 26684
rect 5664 26624 5728 26628
rect 5744 26684 5808 26688
rect 5744 26628 5748 26684
rect 5748 26628 5804 26684
rect 5804 26628 5808 26684
rect 5744 26624 5808 26628
rect 5824 26684 5888 26688
rect 5824 26628 5828 26684
rect 5828 26628 5884 26684
rect 5884 26628 5888 26684
rect 5824 26624 5888 26628
rect 12940 26284 13004 26348
rect 14848 26684 14912 26688
rect 14848 26628 14852 26684
rect 14852 26628 14908 26684
rect 14908 26628 14912 26684
rect 14848 26624 14912 26628
rect 14928 26684 14992 26688
rect 14928 26628 14932 26684
rect 14932 26628 14988 26684
rect 14988 26628 14992 26684
rect 14928 26624 14992 26628
rect 15008 26684 15072 26688
rect 15008 26628 15012 26684
rect 15012 26628 15068 26684
rect 15068 26628 15072 26684
rect 15008 26624 15072 26628
rect 15088 26684 15152 26688
rect 15088 26628 15092 26684
rect 15092 26628 15148 26684
rect 15148 26628 15152 26684
rect 15088 26624 15152 26628
rect 24112 26684 24176 26688
rect 24112 26628 24116 26684
rect 24116 26628 24172 26684
rect 24172 26628 24176 26684
rect 24112 26624 24176 26628
rect 24192 26684 24256 26688
rect 24192 26628 24196 26684
rect 24196 26628 24252 26684
rect 24252 26628 24256 26684
rect 24192 26624 24256 26628
rect 24272 26684 24336 26688
rect 24272 26628 24276 26684
rect 24276 26628 24332 26684
rect 24332 26628 24336 26684
rect 24272 26624 24336 26628
rect 24352 26684 24416 26688
rect 24352 26628 24356 26684
rect 24356 26628 24412 26684
rect 24412 26628 24416 26684
rect 24352 26624 24416 26628
rect 20116 26480 20180 26484
rect 20116 26424 20166 26480
rect 20166 26424 20180 26480
rect 20116 26420 20180 26424
rect 16620 26344 16684 26348
rect 16620 26288 16634 26344
rect 16634 26288 16684 26344
rect 16620 26284 16684 26288
rect 10216 26140 10280 26144
rect 10216 26084 10220 26140
rect 10220 26084 10276 26140
rect 10276 26084 10280 26140
rect 10216 26080 10280 26084
rect 10296 26140 10360 26144
rect 10296 26084 10300 26140
rect 10300 26084 10356 26140
rect 10356 26084 10360 26140
rect 10296 26080 10360 26084
rect 10376 26140 10440 26144
rect 10376 26084 10380 26140
rect 10380 26084 10436 26140
rect 10436 26084 10440 26140
rect 10376 26080 10440 26084
rect 10456 26140 10520 26144
rect 10456 26084 10460 26140
rect 10460 26084 10516 26140
rect 10516 26084 10520 26140
rect 10456 26080 10520 26084
rect 19480 26140 19544 26144
rect 19480 26084 19484 26140
rect 19484 26084 19540 26140
rect 19540 26084 19544 26140
rect 19480 26080 19544 26084
rect 19560 26140 19624 26144
rect 19560 26084 19564 26140
rect 19564 26084 19620 26140
rect 19620 26084 19624 26140
rect 19560 26080 19624 26084
rect 19640 26140 19704 26144
rect 19640 26084 19644 26140
rect 19644 26084 19700 26140
rect 19700 26084 19704 26140
rect 19640 26080 19704 26084
rect 19720 26140 19784 26144
rect 19720 26084 19724 26140
rect 19724 26084 19780 26140
rect 19780 26084 19784 26140
rect 19720 26080 19784 26084
rect 14228 25876 14292 25940
rect 19932 25604 19996 25668
rect 5584 25596 5648 25600
rect 5584 25540 5588 25596
rect 5588 25540 5644 25596
rect 5644 25540 5648 25596
rect 5584 25536 5648 25540
rect 5664 25596 5728 25600
rect 5664 25540 5668 25596
rect 5668 25540 5724 25596
rect 5724 25540 5728 25596
rect 5664 25536 5728 25540
rect 5744 25596 5808 25600
rect 5744 25540 5748 25596
rect 5748 25540 5804 25596
rect 5804 25540 5808 25596
rect 5744 25536 5808 25540
rect 5824 25596 5888 25600
rect 5824 25540 5828 25596
rect 5828 25540 5884 25596
rect 5884 25540 5888 25596
rect 5824 25536 5888 25540
rect 14848 25596 14912 25600
rect 14848 25540 14852 25596
rect 14852 25540 14908 25596
rect 14908 25540 14912 25596
rect 14848 25536 14912 25540
rect 14928 25596 14992 25600
rect 14928 25540 14932 25596
rect 14932 25540 14988 25596
rect 14988 25540 14992 25596
rect 14928 25536 14992 25540
rect 15008 25596 15072 25600
rect 15008 25540 15012 25596
rect 15012 25540 15068 25596
rect 15068 25540 15072 25596
rect 15008 25536 15072 25540
rect 15088 25596 15152 25600
rect 15088 25540 15092 25596
rect 15092 25540 15148 25596
rect 15148 25540 15152 25596
rect 15088 25536 15152 25540
rect 24112 25596 24176 25600
rect 24112 25540 24116 25596
rect 24116 25540 24172 25596
rect 24172 25540 24176 25596
rect 24112 25536 24176 25540
rect 24192 25596 24256 25600
rect 24192 25540 24196 25596
rect 24196 25540 24252 25596
rect 24252 25540 24256 25596
rect 24192 25536 24256 25540
rect 24272 25596 24336 25600
rect 24272 25540 24276 25596
rect 24276 25540 24332 25596
rect 24332 25540 24336 25596
rect 24272 25536 24336 25540
rect 24352 25596 24416 25600
rect 24352 25540 24356 25596
rect 24356 25540 24412 25596
rect 24412 25540 24416 25596
rect 24352 25536 24416 25540
rect 16988 25468 17052 25532
rect 23612 25392 23676 25396
rect 23612 25336 23662 25392
rect 23662 25336 23676 25392
rect 23612 25332 23676 25336
rect 18644 25196 18708 25260
rect 24532 25060 24596 25124
rect 10216 25052 10280 25056
rect 10216 24996 10220 25052
rect 10220 24996 10276 25052
rect 10276 24996 10280 25052
rect 10216 24992 10280 24996
rect 10296 25052 10360 25056
rect 10296 24996 10300 25052
rect 10300 24996 10356 25052
rect 10356 24996 10360 25052
rect 10296 24992 10360 24996
rect 10376 25052 10440 25056
rect 10376 24996 10380 25052
rect 10380 24996 10436 25052
rect 10436 24996 10440 25052
rect 10376 24992 10440 24996
rect 10456 25052 10520 25056
rect 10456 24996 10460 25052
rect 10460 24996 10516 25052
rect 10516 24996 10520 25052
rect 10456 24992 10520 24996
rect 19480 25052 19544 25056
rect 19480 24996 19484 25052
rect 19484 24996 19540 25052
rect 19540 24996 19544 25052
rect 19480 24992 19544 24996
rect 19560 25052 19624 25056
rect 19560 24996 19564 25052
rect 19564 24996 19620 25052
rect 19620 24996 19624 25052
rect 19560 24992 19624 24996
rect 19640 25052 19704 25056
rect 19640 24996 19644 25052
rect 19644 24996 19700 25052
rect 19700 24996 19704 25052
rect 19640 24992 19704 24996
rect 19720 25052 19784 25056
rect 19720 24996 19724 25052
rect 19724 24996 19780 25052
rect 19780 24996 19784 25052
rect 19720 24992 19784 24996
rect 13676 24788 13740 24852
rect 5584 24508 5648 24512
rect 5584 24452 5588 24508
rect 5588 24452 5644 24508
rect 5644 24452 5648 24508
rect 5584 24448 5648 24452
rect 5664 24508 5728 24512
rect 5664 24452 5668 24508
rect 5668 24452 5724 24508
rect 5724 24452 5728 24508
rect 5664 24448 5728 24452
rect 5744 24508 5808 24512
rect 5744 24452 5748 24508
rect 5748 24452 5804 24508
rect 5804 24452 5808 24508
rect 5744 24448 5808 24452
rect 5824 24508 5888 24512
rect 5824 24452 5828 24508
rect 5828 24452 5884 24508
rect 5884 24452 5888 24508
rect 5824 24448 5888 24452
rect 14848 24508 14912 24512
rect 14848 24452 14852 24508
rect 14852 24452 14908 24508
rect 14908 24452 14912 24508
rect 14848 24448 14912 24452
rect 14928 24508 14992 24512
rect 14928 24452 14932 24508
rect 14932 24452 14988 24508
rect 14988 24452 14992 24508
rect 14928 24448 14992 24452
rect 15008 24508 15072 24512
rect 15008 24452 15012 24508
rect 15012 24452 15068 24508
rect 15068 24452 15072 24508
rect 15008 24448 15072 24452
rect 15088 24508 15152 24512
rect 15088 24452 15092 24508
rect 15092 24452 15148 24508
rect 15148 24452 15152 24508
rect 15088 24448 15152 24452
rect 24112 24508 24176 24512
rect 24112 24452 24116 24508
rect 24116 24452 24172 24508
rect 24172 24452 24176 24508
rect 24112 24448 24176 24452
rect 24192 24508 24256 24512
rect 24192 24452 24196 24508
rect 24196 24452 24252 24508
rect 24252 24452 24256 24508
rect 24192 24448 24256 24452
rect 24272 24508 24336 24512
rect 24272 24452 24276 24508
rect 24276 24452 24332 24508
rect 24332 24452 24336 24508
rect 24272 24448 24336 24452
rect 24352 24508 24416 24512
rect 24352 24452 24356 24508
rect 24356 24452 24412 24508
rect 24412 24452 24416 24508
rect 24352 24448 24416 24452
rect 14228 24108 14292 24172
rect 10216 23964 10280 23968
rect 10216 23908 10220 23964
rect 10220 23908 10276 23964
rect 10276 23908 10280 23964
rect 10216 23904 10280 23908
rect 10296 23964 10360 23968
rect 10296 23908 10300 23964
rect 10300 23908 10356 23964
rect 10356 23908 10360 23964
rect 10296 23904 10360 23908
rect 10376 23964 10440 23968
rect 10376 23908 10380 23964
rect 10380 23908 10436 23964
rect 10436 23908 10440 23964
rect 10376 23904 10440 23908
rect 10456 23964 10520 23968
rect 10456 23908 10460 23964
rect 10460 23908 10516 23964
rect 10516 23908 10520 23964
rect 10456 23904 10520 23908
rect 19480 23964 19544 23968
rect 19480 23908 19484 23964
rect 19484 23908 19540 23964
rect 19540 23908 19544 23964
rect 19480 23904 19544 23908
rect 19560 23964 19624 23968
rect 19560 23908 19564 23964
rect 19564 23908 19620 23964
rect 19620 23908 19624 23964
rect 19560 23904 19624 23908
rect 19640 23964 19704 23968
rect 19640 23908 19644 23964
rect 19644 23908 19700 23964
rect 19700 23908 19704 23964
rect 19640 23904 19704 23908
rect 19720 23964 19784 23968
rect 19720 23908 19724 23964
rect 19724 23908 19780 23964
rect 19780 23908 19784 23964
rect 19720 23904 19784 23908
rect 15516 23836 15580 23900
rect 7236 23428 7300 23492
rect 14412 23428 14476 23492
rect 15516 23564 15580 23628
rect 26372 23488 26436 23492
rect 26372 23432 26386 23488
rect 26386 23432 26436 23488
rect 26372 23428 26436 23432
rect 5584 23420 5648 23424
rect 5584 23364 5588 23420
rect 5588 23364 5644 23420
rect 5644 23364 5648 23420
rect 5584 23360 5648 23364
rect 5664 23420 5728 23424
rect 5664 23364 5668 23420
rect 5668 23364 5724 23420
rect 5724 23364 5728 23420
rect 5664 23360 5728 23364
rect 5744 23420 5808 23424
rect 5744 23364 5748 23420
rect 5748 23364 5804 23420
rect 5804 23364 5808 23420
rect 5744 23360 5808 23364
rect 5824 23420 5888 23424
rect 5824 23364 5828 23420
rect 5828 23364 5884 23420
rect 5884 23364 5888 23420
rect 5824 23360 5888 23364
rect 14848 23420 14912 23424
rect 14848 23364 14852 23420
rect 14852 23364 14908 23420
rect 14908 23364 14912 23420
rect 14848 23360 14912 23364
rect 14928 23420 14992 23424
rect 14928 23364 14932 23420
rect 14932 23364 14988 23420
rect 14988 23364 14992 23420
rect 14928 23360 14992 23364
rect 15008 23420 15072 23424
rect 15008 23364 15012 23420
rect 15012 23364 15068 23420
rect 15068 23364 15072 23420
rect 15008 23360 15072 23364
rect 15088 23420 15152 23424
rect 15088 23364 15092 23420
rect 15092 23364 15148 23420
rect 15148 23364 15152 23420
rect 15088 23360 15152 23364
rect 24112 23420 24176 23424
rect 24112 23364 24116 23420
rect 24116 23364 24172 23420
rect 24172 23364 24176 23420
rect 24112 23360 24176 23364
rect 24192 23420 24256 23424
rect 24192 23364 24196 23420
rect 24196 23364 24252 23420
rect 24252 23364 24256 23420
rect 24192 23360 24256 23364
rect 24272 23420 24336 23424
rect 24272 23364 24276 23420
rect 24276 23364 24332 23420
rect 24332 23364 24336 23420
rect 24272 23360 24336 23364
rect 24352 23420 24416 23424
rect 24352 23364 24356 23420
rect 24356 23364 24412 23420
rect 24412 23364 24416 23420
rect 24352 23360 24416 23364
rect 24532 23020 24596 23084
rect 10216 22876 10280 22880
rect 10216 22820 10220 22876
rect 10220 22820 10276 22876
rect 10276 22820 10280 22876
rect 10216 22816 10280 22820
rect 10296 22876 10360 22880
rect 10296 22820 10300 22876
rect 10300 22820 10356 22876
rect 10356 22820 10360 22876
rect 10296 22816 10360 22820
rect 10376 22876 10440 22880
rect 10376 22820 10380 22876
rect 10380 22820 10436 22876
rect 10436 22820 10440 22876
rect 10376 22816 10440 22820
rect 10456 22876 10520 22880
rect 10456 22820 10460 22876
rect 10460 22820 10516 22876
rect 10516 22820 10520 22876
rect 10456 22816 10520 22820
rect 19480 22876 19544 22880
rect 19480 22820 19484 22876
rect 19484 22820 19540 22876
rect 19540 22820 19544 22876
rect 19480 22816 19544 22820
rect 19560 22876 19624 22880
rect 19560 22820 19564 22876
rect 19564 22820 19620 22876
rect 19620 22820 19624 22876
rect 19560 22816 19624 22820
rect 19640 22876 19704 22880
rect 19640 22820 19644 22876
rect 19644 22820 19700 22876
rect 19700 22820 19704 22876
rect 19640 22816 19704 22820
rect 19720 22876 19784 22880
rect 19720 22820 19724 22876
rect 19724 22820 19780 22876
rect 19780 22820 19784 22876
rect 19720 22816 19784 22820
rect 5584 22332 5648 22336
rect 5584 22276 5588 22332
rect 5588 22276 5644 22332
rect 5644 22276 5648 22332
rect 5584 22272 5648 22276
rect 5664 22332 5728 22336
rect 5664 22276 5668 22332
rect 5668 22276 5724 22332
rect 5724 22276 5728 22332
rect 5664 22272 5728 22276
rect 5744 22332 5808 22336
rect 5744 22276 5748 22332
rect 5748 22276 5804 22332
rect 5804 22276 5808 22332
rect 5744 22272 5808 22276
rect 5824 22332 5888 22336
rect 5824 22276 5828 22332
rect 5828 22276 5884 22332
rect 5884 22276 5888 22332
rect 5824 22272 5888 22276
rect 14848 22332 14912 22336
rect 14848 22276 14852 22332
rect 14852 22276 14908 22332
rect 14908 22276 14912 22332
rect 14848 22272 14912 22276
rect 14928 22332 14992 22336
rect 14928 22276 14932 22332
rect 14932 22276 14988 22332
rect 14988 22276 14992 22332
rect 14928 22272 14992 22276
rect 15008 22332 15072 22336
rect 15008 22276 15012 22332
rect 15012 22276 15068 22332
rect 15068 22276 15072 22332
rect 15008 22272 15072 22276
rect 15088 22332 15152 22336
rect 15088 22276 15092 22332
rect 15092 22276 15148 22332
rect 15148 22276 15152 22332
rect 15088 22272 15152 22276
rect 24112 22332 24176 22336
rect 24112 22276 24116 22332
rect 24116 22276 24172 22332
rect 24172 22276 24176 22332
rect 24112 22272 24176 22276
rect 24192 22332 24256 22336
rect 24192 22276 24196 22332
rect 24196 22276 24252 22332
rect 24252 22276 24256 22332
rect 24192 22272 24256 22276
rect 24272 22332 24336 22336
rect 24272 22276 24276 22332
rect 24276 22276 24332 22332
rect 24332 22276 24336 22332
rect 24272 22272 24336 22276
rect 24352 22332 24416 22336
rect 24352 22276 24356 22332
rect 24356 22276 24412 22332
rect 24412 22276 24416 22332
rect 24352 22272 24416 22276
rect 19932 22068 19996 22132
rect 22140 22068 22204 22132
rect 23612 22128 23676 22132
rect 23612 22072 23662 22128
rect 23662 22072 23676 22128
rect 23612 22068 23676 22072
rect 10216 21788 10280 21792
rect 10216 21732 10220 21788
rect 10220 21732 10276 21788
rect 10276 21732 10280 21788
rect 10216 21728 10280 21732
rect 10296 21788 10360 21792
rect 10296 21732 10300 21788
rect 10300 21732 10356 21788
rect 10356 21732 10360 21788
rect 10296 21728 10360 21732
rect 10376 21788 10440 21792
rect 10376 21732 10380 21788
rect 10380 21732 10436 21788
rect 10436 21732 10440 21788
rect 10376 21728 10440 21732
rect 10456 21788 10520 21792
rect 10456 21732 10460 21788
rect 10460 21732 10516 21788
rect 10516 21732 10520 21788
rect 10456 21728 10520 21732
rect 19480 21788 19544 21792
rect 19480 21732 19484 21788
rect 19484 21732 19540 21788
rect 19540 21732 19544 21788
rect 19480 21728 19544 21732
rect 19560 21788 19624 21792
rect 19560 21732 19564 21788
rect 19564 21732 19620 21788
rect 19620 21732 19624 21788
rect 19560 21728 19624 21732
rect 19640 21788 19704 21792
rect 19640 21732 19644 21788
rect 19644 21732 19700 21788
rect 19700 21732 19704 21788
rect 19640 21728 19704 21732
rect 19720 21788 19784 21792
rect 19720 21732 19724 21788
rect 19724 21732 19780 21788
rect 19780 21732 19784 21788
rect 19720 21728 19784 21732
rect 19932 21388 19996 21452
rect 5584 21244 5648 21248
rect 5584 21188 5588 21244
rect 5588 21188 5644 21244
rect 5644 21188 5648 21244
rect 5584 21184 5648 21188
rect 5664 21244 5728 21248
rect 5664 21188 5668 21244
rect 5668 21188 5724 21244
rect 5724 21188 5728 21244
rect 5664 21184 5728 21188
rect 5744 21244 5808 21248
rect 5744 21188 5748 21244
rect 5748 21188 5804 21244
rect 5804 21188 5808 21244
rect 5744 21184 5808 21188
rect 5824 21244 5888 21248
rect 5824 21188 5828 21244
rect 5828 21188 5884 21244
rect 5884 21188 5888 21244
rect 5824 21184 5888 21188
rect 14848 21244 14912 21248
rect 14848 21188 14852 21244
rect 14852 21188 14908 21244
rect 14908 21188 14912 21244
rect 14848 21184 14912 21188
rect 14928 21244 14992 21248
rect 14928 21188 14932 21244
rect 14932 21188 14988 21244
rect 14988 21188 14992 21244
rect 14928 21184 14992 21188
rect 15008 21244 15072 21248
rect 15008 21188 15012 21244
rect 15012 21188 15068 21244
rect 15068 21188 15072 21244
rect 15008 21184 15072 21188
rect 15088 21244 15152 21248
rect 15088 21188 15092 21244
rect 15092 21188 15148 21244
rect 15148 21188 15152 21244
rect 15088 21184 15152 21188
rect 24112 21244 24176 21248
rect 24112 21188 24116 21244
rect 24116 21188 24172 21244
rect 24172 21188 24176 21244
rect 24112 21184 24176 21188
rect 24192 21244 24256 21248
rect 24192 21188 24196 21244
rect 24196 21188 24252 21244
rect 24252 21188 24256 21244
rect 24192 21184 24256 21188
rect 24272 21244 24336 21248
rect 24272 21188 24276 21244
rect 24276 21188 24332 21244
rect 24332 21188 24336 21244
rect 24272 21184 24336 21188
rect 24352 21244 24416 21248
rect 24352 21188 24356 21244
rect 24356 21188 24412 21244
rect 24412 21188 24416 21244
rect 24352 21184 24416 21188
rect 16988 20844 17052 20908
rect 10216 20700 10280 20704
rect 10216 20644 10220 20700
rect 10220 20644 10276 20700
rect 10276 20644 10280 20700
rect 10216 20640 10280 20644
rect 10296 20700 10360 20704
rect 10296 20644 10300 20700
rect 10300 20644 10356 20700
rect 10356 20644 10360 20700
rect 10296 20640 10360 20644
rect 10376 20700 10440 20704
rect 10376 20644 10380 20700
rect 10380 20644 10436 20700
rect 10436 20644 10440 20700
rect 10376 20640 10440 20644
rect 10456 20700 10520 20704
rect 10456 20644 10460 20700
rect 10460 20644 10516 20700
rect 10516 20644 10520 20700
rect 10456 20640 10520 20644
rect 19480 20700 19544 20704
rect 19480 20644 19484 20700
rect 19484 20644 19540 20700
rect 19540 20644 19544 20700
rect 19480 20640 19544 20644
rect 19560 20700 19624 20704
rect 19560 20644 19564 20700
rect 19564 20644 19620 20700
rect 19620 20644 19624 20700
rect 19560 20640 19624 20644
rect 19640 20700 19704 20704
rect 19640 20644 19644 20700
rect 19644 20644 19700 20700
rect 19700 20644 19704 20700
rect 19640 20640 19704 20644
rect 19720 20700 19784 20704
rect 19720 20644 19724 20700
rect 19724 20644 19780 20700
rect 19780 20644 19784 20700
rect 19720 20640 19784 20644
rect 16620 20436 16684 20500
rect 5584 20156 5648 20160
rect 5584 20100 5588 20156
rect 5588 20100 5644 20156
rect 5644 20100 5648 20156
rect 5584 20096 5648 20100
rect 5664 20156 5728 20160
rect 5664 20100 5668 20156
rect 5668 20100 5724 20156
rect 5724 20100 5728 20156
rect 5664 20096 5728 20100
rect 5744 20156 5808 20160
rect 5744 20100 5748 20156
rect 5748 20100 5804 20156
rect 5804 20100 5808 20156
rect 5744 20096 5808 20100
rect 5824 20156 5888 20160
rect 5824 20100 5828 20156
rect 5828 20100 5884 20156
rect 5884 20100 5888 20156
rect 5824 20096 5888 20100
rect 14848 20156 14912 20160
rect 14848 20100 14852 20156
rect 14852 20100 14908 20156
rect 14908 20100 14912 20156
rect 14848 20096 14912 20100
rect 14928 20156 14992 20160
rect 14928 20100 14932 20156
rect 14932 20100 14988 20156
rect 14988 20100 14992 20156
rect 14928 20096 14992 20100
rect 15008 20156 15072 20160
rect 15008 20100 15012 20156
rect 15012 20100 15068 20156
rect 15068 20100 15072 20156
rect 15008 20096 15072 20100
rect 15088 20156 15152 20160
rect 15088 20100 15092 20156
rect 15092 20100 15148 20156
rect 15148 20100 15152 20156
rect 15088 20096 15152 20100
rect 24112 20156 24176 20160
rect 24112 20100 24116 20156
rect 24116 20100 24172 20156
rect 24172 20100 24176 20156
rect 24112 20096 24176 20100
rect 24192 20156 24256 20160
rect 24192 20100 24196 20156
rect 24196 20100 24252 20156
rect 24252 20100 24256 20156
rect 24192 20096 24256 20100
rect 24272 20156 24336 20160
rect 24272 20100 24276 20156
rect 24276 20100 24332 20156
rect 24332 20100 24336 20156
rect 24272 20096 24336 20100
rect 24352 20156 24416 20160
rect 24352 20100 24356 20156
rect 24356 20100 24412 20156
rect 24412 20100 24416 20156
rect 24352 20096 24416 20100
rect 22140 19892 22204 19956
rect 10216 19612 10280 19616
rect 10216 19556 10220 19612
rect 10220 19556 10276 19612
rect 10276 19556 10280 19612
rect 10216 19552 10280 19556
rect 10296 19612 10360 19616
rect 10296 19556 10300 19612
rect 10300 19556 10356 19612
rect 10356 19556 10360 19612
rect 10296 19552 10360 19556
rect 10376 19612 10440 19616
rect 10376 19556 10380 19612
rect 10380 19556 10436 19612
rect 10436 19556 10440 19612
rect 10376 19552 10440 19556
rect 10456 19612 10520 19616
rect 10456 19556 10460 19612
rect 10460 19556 10516 19612
rect 10516 19556 10520 19612
rect 10456 19552 10520 19556
rect 19480 19612 19544 19616
rect 19480 19556 19484 19612
rect 19484 19556 19540 19612
rect 19540 19556 19544 19612
rect 19480 19552 19544 19556
rect 19560 19612 19624 19616
rect 19560 19556 19564 19612
rect 19564 19556 19620 19612
rect 19620 19556 19624 19612
rect 19560 19552 19624 19556
rect 19640 19612 19704 19616
rect 19640 19556 19644 19612
rect 19644 19556 19700 19612
rect 19700 19556 19704 19612
rect 19640 19552 19704 19556
rect 19720 19612 19784 19616
rect 19720 19556 19724 19612
rect 19724 19556 19780 19612
rect 19780 19556 19784 19612
rect 19720 19552 19784 19556
rect 5584 19068 5648 19072
rect 5584 19012 5588 19068
rect 5588 19012 5644 19068
rect 5644 19012 5648 19068
rect 5584 19008 5648 19012
rect 5664 19068 5728 19072
rect 5664 19012 5668 19068
rect 5668 19012 5724 19068
rect 5724 19012 5728 19068
rect 5664 19008 5728 19012
rect 5744 19068 5808 19072
rect 5744 19012 5748 19068
rect 5748 19012 5804 19068
rect 5804 19012 5808 19068
rect 5744 19008 5808 19012
rect 5824 19068 5888 19072
rect 5824 19012 5828 19068
rect 5828 19012 5884 19068
rect 5884 19012 5888 19068
rect 5824 19008 5888 19012
rect 14848 19068 14912 19072
rect 14848 19012 14852 19068
rect 14852 19012 14908 19068
rect 14908 19012 14912 19068
rect 14848 19008 14912 19012
rect 14928 19068 14992 19072
rect 14928 19012 14932 19068
rect 14932 19012 14988 19068
rect 14988 19012 14992 19068
rect 14928 19008 14992 19012
rect 15008 19068 15072 19072
rect 15008 19012 15012 19068
rect 15012 19012 15068 19068
rect 15068 19012 15072 19068
rect 15008 19008 15072 19012
rect 15088 19068 15152 19072
rect 15088 19012 15092 19068
rect 15092 19012 15148 19068
rect 15148 19012 15152 19068
rect 15088 19008 15152 19012
rect 24112 19068 24176 19072
rect 24112 19012 24116 19068
rect 24116 19012 24172 19068
rect 24172 19012 24176 19068
rect 24112 19008 24176 19012
rect 24192 19068 24256 19072
rect 24192 19012 24196 19068
rect 24196 19012 24252 19068
rect 24252 19012 24256 19068
rect 24192 19008 24256 19012
rect 24272 19068 24336 19072
rect 24272 19012 24276 19068
rect 24276 19012 24332 19068
rect 24332 19012 24336 19068
rect 24272 19008 24336 19012
rect 24352 19068 24416 19072
rect 24352 19012 24356 19068
rect 24356 19012 24412 19068
rect 24412 19012 24416 19068
rect 24352 19008 24416 19012
rect 10216 18524 10280 18528
rect 10216 18468 10220 18524
rect 10220 18468 10276 18524
rect 10276 18468 10280 18524
rect 10216 18464 10280 18468
rect 10296 18524 10360 18528
rect 10296 18468 10300 18524
rect 10300 18468 10356 18524
rect 10356 18468 10360 18524
rect 10296 18464 10360 18468
rect 10376 18524 10440 18528
rect 10376 18468 10380 18524
rect 10380 18468 10436 18524
rect 10436 18468 10440 18524
rect 10376 18464 10440 18468
rect 10456 18524 10520 18528
rect 10456 18468 10460 18524
rect 10460 18468 10516 18524
rect 10516 18468 10520 18524
rect 10456 18464 10520 18468
rect 19480 18524 19544 18528
rect 19480 18468 19484 18524
rect 19484 18468 19540 18524
rect 19540 18468 19544 18524
rect 19480 18464 19544 18468
rect 19560 18524 19624 18528
rect 19560 18468 19564 18524
rect 19564 18468 19620 18524
rect 19620 18468 19624 18524
rect 19560 18464 19624 18468
rect 19640 18524 19704 18528
rect 19640 18468 19644 18524
rect 19644 18468 19700 18524
rect 19700 18468 19704 18524
rect 19640 18464 19704 18468
rect 19720 18524 19784 18528
rect 19720 18468 19724 18524
rect 19724 18468 19780 18524
rect 19780 18468 19784 18524
rect 19720 18464 19784 18468
rect 5584 17980 5648 17984
rect 5584 17924 5588 17980
rect 5588 17924 5644 17980
rect 5644 17924 5648 17980
rect 5584 17920 5648 17924
rect 5664 17980 5728 17984
rect 5664 17924 5668 17980
rect 5668 17924 5724 17980
rect 5724 17924 5728 17980
rect 5664 17920 5728 17924
rect 5744 17980 5808 17984
rect 5744 17924 5748 17980
rect 5748 17924 5804 17980
rect 5804 17924 5808 17980
rect 5744 17920 5808 17924
rect 5824 17980 5888 17984
rect 5824 17924 5828 17980
rect 5828 17924 5884 17980
rect 5884 17924 5888 17980
rect 5824 17920 5888 17924
rect 14848 17980 14912 17984
rect 14848 17924 14852 17980
rect 14852 17924 14908 17980
rect 14908 17924 14912 17980
rect 14848 17920 14912 17924
rect 14928 17980 14992 17984
rect 14928 17924 14932 17980
rect 14932 17924 14988 17980
rect 14988 17924 14992 17980
rect 14928 17920 14992 17924
rect 15008 17980 15072 17984
rect 15008 17924 15012 17980
rect 15012 17924 15068 17980
rect 15068 17924 15072 17980
rect 15008 17920 15072 17924
rect 15088 17980 15152 17984
rect 15088 17924 15092 17980
rect 15092 17924 15148 17980
rect 15148 17924 15152 17980
rect 15088 17920 15152 17924
rect 24112 17980 24176 17984
rect 24112 17924 24116 17980
rect 24116 17924 24172 17980
rect 24172 17924 24176 17980
rect 24112 17920 24176 17924
rect 24192 17980 24256 17984
rect 24192 17924 24196 17980
rect 24196 17924 24252 17980
rect 24252 17924 24256 17980
rect 24192 17920 24256 17924
rect 24272 17980 24336 17984
rect 24272 17924 24276 17980
rect 24276 17924 24332 17980
rect 24332 17924 24336 17980
rect 24272 17920 24336 17924
rect 24352 17980 24416 17984
rect 24352 17924 24356 17980
rect 24356 17924 24412 17980
rect 24412 17924 24416 17980
rect 24352 17920 24416 17924
rect 18460 17716 18524 17780
rect 26556 17716 26620 17780
rect 26372 17580 26436 17644
rect 10216 17436 10280 17440
rect 10216 17380 10220 17436
rect 10220 17380 10276 17436
rect 10276 17380 10280 17436
rect 10216 17376 10280 17380
rect 10296 17436 10360 17440
rect 10296 17380 10300 17436
rect 10300 17380 10356 17436
rect 10356 17380 10360 17436
rect 10296 17376 10360 17380
rect 10376 17436 10440 17440
rect 10376 17380 10380 17436
rect 10380 17380 10436 17436
rect 10436 17380 10440 17436
rect 10376 17376 10440 17380
rect 10456 17436 10520 17440
rect 10456 17380 10460 17436
rect 10460 17380 10516 17436
rect 10516 17380 10520 17436
rect 10456 17376 10520 17380
rect 19480 17436 19544 17440
rect 19480 17380 19484 17436
rect 19484 17380 19540 17436
rect 19540 17380 19544 17436
rect 19480 17376 19544 17380
rect 19560 17436 19624 17440
rect 19560 17380 19564 17436
rect 19564 17380 19620 17436
rect 19620 17380 19624 17436
rect 19560 17376 19624 17380
rect 19640 17436 19704 17440
rect 19640 17380 19644 17436
rect 19644 17380 19700 17436
rect 19700 17380 19704 17436
rect 19640 17376 19704 17380
rect 19720 17436 19784 17440
rect 19720 17380 19724 17436
rect 19724 17380 19780 17436
rect 19780 17380 19784 17436
rect 19720 17376 19784 17380
rect 5584 16892 5648 16896
rect 5584 16836 5588 16892
rect 5588 16836 5644 16892
rect 5644 16836 5648 16892
rect 5584 16832 5648 16836
rect 5664 16892 5728 16896
rect 5664 16836 5668 16892
rect 5668 16836 5724 16892
rect 5724 16836 5728 16892
rect 5664 16832 5728 16836
rect 5744 16892 5808 16896
rect 5744 16836 5748 16892
rect 5748 16836 5804 16892
rect 5804 16836 5808 16892
rect 5744 16832 5808 16836
rect 5824 16892 5888 16896
rect 5824 16836 5828 16892
rect 5828 16836 5884 16892
rect 5884 16836 5888 16892
rect 5824 16832 5888 16836
rect 14848 16892 14912 16896
rect 14848 16836 14852 16892
rect 14852 16836 14908 16892
rect 14908 16836 14912 16892
rect 14848 16832 14912 16836
rect 14928 16892 14992 16896
rect 14928 16836 14932 16892
rect 14932 16836 14988 16892
rect 14988 16836 14992 16892
rect 14928 16832 14992 16836
rect 15008 16892 15072 16896
rect 15008 16836 15012 16892
rect 15012 16836 15068 16892
rect 15068 16836 15072 16892
rect 15008 16832 15072 16836
rect 15088 16892 15152 16896
rect 15088 16836 15092 16892
rect 15092 16836 15148 16892
rect 15148 16836 15152 16892
rect 15088 16832 15152 16836
rect 24112 16892 24176 16896
rect 24112 16836 24116 16892
rect 24116 16836 24172 16892
rect 24172 16836 24176 16892
rect 24112 16832 24176 16836
rect 24192 16892 24256 16896
rect 24192 16836 24196 16892
rect 24196 16836 24252 16892
rect 24252 16836 24256 16892
rect 24192 16832 24256 16836
rect 24272 16892 24336 16896
rect 24272 16836 24276 16892
rect 24276 16836 24332 16892
rect 24332 16836 24336 16892
rect 24272 16832 24336 16836
rect 24352 16892 24416 16896
rect 24352 16836 24356 16892
rect 24356 16836 24412 16892
rect 24412 16836 24416 16892
rect 24352 16832 24416 16836
rect 26188 16492 26252 16556
rect 10216 16348 10280 16352
rect 10216 16292 10220 16348
rect 10220 16292 10276 16348
rect 10276 16292 10280 16348
rect 10216 16288 10280 16292
rect 10296 16348 10360 16352
rect 10296 16292 10300 16348
rect 10300 16292 10356 16348
rect 10356 16292 10360 16348
rect 10296 16288 10360 16292
rect 10376 16348 10440 16352
rect 10376 16292 10380 16348
rect 10380 16292 10436 16348
rect 10436 16292 10440 16348
rect 10376 16288 10440 16292
rect 10456 16348 10520 16352
rect 10456 16292 10460 16348
rect 10460 16292 10516 16348
rect 10516 16292 10520 16348
rect 10456 16288 10520 16292
rect 19480 16348 19544 16352
rect 19480 16292 19484 16348
rect 19484 16292 19540 16348
rect 19540 16292 19544 16348
rect 19480 16288 19544 16292
rect 19560 16348 19624 16352
rect 19560 16292 19564 16348
rect 19564 16292 19620 16348
rect 19620 16292 19624 16348
rect 19560 16288 19624 16292
rect 19640 16348 19704 16352
rect 19640 16292 19644 16348
rect 19644 16292 19700 16348
rect 19700 16292 19704 16348
rect 19640 16288 19704 16292
rect 19720 16348 19784 16352
rect 19720 16292 19724 16348
rect 19724 16292 19780 16348
rect 19780 16292 19784 16348
rect 19720 16288 19784 16292
rect 18644 16084 18708 16148
rect 5584 15804 5648 15808
rect 5584 15748 5588 15804
rect 5588 15748 5644 15804
rect 5644 15748 5648 15804
rect 5584 15744 5648 15748
rect 5664 15804 5728 15808
rect 5664 15748 5668 15804
rect 5668 15748 5724 15804
rect 5724 15748 5728 15804
rect 5664 15744 5728 15748
rect 5744 15804 5808 15808
rect 5744 15748 5748 15804
rect 5748 15748 5804 15804
rect 5804 15748 5808 15804
rect 5744 15744 5808 15748
rect 5824 15804 5888 15808
rect 5824 15748 5828 15804
rect 5828 15748 5884 15804
rect 5884 15748 5888 15804
rect 5824 15744 5888 15748
rect 14848 15804 14912 15808
rect 14848 15748 14852 15804
rect 14852 15748 14908 15804
rect 14908 15748 14912 15804
rect 14848 15744 14912 15748
rect 14928 15804 14992 15808
rect 14928 15748 14932 15804
rect 14932 15748 14988 15804
rect 14988 15748 14992 15804
rect 14928 15744 14992 15748
rect 15008 15804 15072 15808
rect 15008 15748 15012 15804
rect 15012 15748 15068 15804
rect 15068 15748 15072 15804
rect 15008 15744 15072 15748
rect 15088 15804 15152 15808
rect 15088 15748 15092 15804
rect 15092 15748 15148 15804
rect 15148 15748 15152 15804
rect 15088 15744 15152 15748
rect 24112 15804 24176 15808
rect 24112 15748 24116 15804
rect 24116 15748 24172 15804
rect 24172 15748 24176 15804
rect 24112 15744 24176 15748
rect 24192 15804 24256 15808
rect 24192 15748 24196 15804
rect 24196 15748 24252 15804
rect 24252 15748 24256 15804
rect 24192 15744 24256 15748
rect 24272 15804 24336 15808
rect 24272 15748 24276 15804
rect 24276 15748 24332 15804
rect 24332 15748 24336 15804
rect 24272 15744 24336 15748
rect 24352 15804 24416 15808
rect 24352 15748 24356 15804
rect 24356 15748 24412 15804
rect 24412 15748 24416 15804
rect 24352 15744 24416 15748
rect 10216 15260 10280 15264
rect 10216 15204 10220 15260
rect 10220 15204 10276 15260
rect 10276 15204 10280 15260
rect 10216 15200 10280 15204
rect 10296 15260 10360 15264
rect 10296 15204 10300 15260
rect 10300 15204 10356 15260
rect 10356 15204 10360 15260
rect 10296 15200 10360 15204
rect 10376 15260 10440 15264
rect 10376 15204 10380 15260
rect 10380 15204 10436 15260
rect 10436 15204 10440 15260
rect 10376 15200 10440 15204
rect 10456 15260 10520 15264
rect 10456 15204 10460 15260
rect 10460 15204 10516 15260
rect 10516 15204 10520 15260
rect 10456 15200 10520 15204
rect 19480 15260 19544 15264
rect 19480 15204 19484 15260
rect 19484 15204 19540 15260
rect 19540 15204 19544 15260
rect 19480 15200 19544 15204
rect 19560 15260 19624 15264
rect 19560 15204 19564 15260
rect 19564 15204 19620 15260
rect 19620 15204 19624 15260
rect 19560 15200 19624 15204
rect 19640 15260 19704 15264
rect 19640 15204 19644 15260
rect 19644 15204 19700 15260
rect 19700 15204 19704 15260
rect 19640 15200 19704 15204
rect 19720 15260 19784 15264
rect 19720 15204 19724 15260
rect 19724 15204 19780 15260
rect 19780 15204 19784 15260
rect 19720 15200 19784 15204
rect 5584 14716 5648 14720
rect 5584 14660 5588 14716
rect 5588 14660 5644 14716
rect 5644 14660 5648 14716
rect 5584 14656 5648 14660
rect 5664 14716 5728 14720
rect 5664 14660 5668 14716
rect 5668 14660 5724 14716
rect 5724 14660 5728 14716
rect 5664 14656 5728 14660
rect 5744 14716 5808 14720
rect 5744 14660 5748 14716
rect 5748 14660 5804 14716
rect 5804 14660 5808 14716
rect 5744 14656 5808 14660
rect 5824 14716 5888 14720
rect 5824 14660 5828 14716
rect 5828 14660 5884 14716
rect 5884 14660 5888 14716
rect 5824 14656 5888 14660
rect 14848 14716 14912 14720
rect 14848 14660 14852 14716
rect 14852 14660 14908 14716
rect 14908 14660 14912 14716
rect 14848 14656 14912 14660
rect 14928 14716 14992 14720
rect 14928 14660 14932 14716
rect 14932 14660 14988 14716
rect 14988 14660 14992 14716
rect 14928 14656 14992 14660
rect 15008 14716 15072 14720
rect 15008 14660 15012 14716
rect 15012 14660 15068 14716
rect 15068 14660 15072 14716
rect 15008 14656 15072 14660
rect 15088 14716 15152 14720
rect 15088 14660 15092 14716
rect 15092 14660 15148 14716
rect 15148 14660 15152 14716
rect 15088 14656 15152 14660
rect 24112 14716 24176 14720
rect 24112 14660 24116 14716
rect 24116 14660 24172 14716
rect 24172 14660 24176 14716
rect 24112 14656 24176 14660
rect 24192 14716 24256 14720
rect 24192 14660 24196 14716
rect 24196 14660 24252 14716
rect 24252 14660 24256 14716
rect 24192 14656 24256 14660
rect 24272 14716 24336 14720
rect 24272 14660 24276 14716
rect 24276 14660 24332 14716
rect 24332 14660 24336 14716
rect 24272 14656 24336 14660
rect 24352 14716 24416 14720
rect 24352 14660 24356 14716
rect 24356 14660 24412 14716
rect 24412 14660 24416 14716
rect 24352 14656 24416 14660
rect 10216 14172 10280 14176
rect 10216 14116 10220 14172
rect 10220 14116 10276 14172
rect 10276 14116 10280 14172
rect 10216 14112 10280 14116
rect 10296 14172 10360 14176
rect 10296 14116 10300 14172
rect 10300 14116 10356 14172
rect 10356 14116 10360 14172
rect 10296 14112 10360 14116
rect 10376 14172 10440 14176
rect 10376 14116 10380 14172
rect 10380 14116 10436 14172
rect 10436 14116 10440 14172
rect 10376 14112 10440 14116
rect 10456 14172 10520 14176
rect 10456 14116 10460 14172
rect 10460 14116 10516 14172
rect 10516 14116 10520 14172
rect 10456 14112 10520 14116
rect 19480 14172 19544 14176
rect 19480 14116 19484 14172
rect 19484 14116 19540 14172
rect 19540 14116 19544 14172
rect 19480 14112 19544 14116
rect 19560 14172 19624 14176
rect 19560 14116 19564 14172
rect 19564 14116 19620 14172
rect 19620 14116 19624 14172
rect 19560 14112 19624 14116
rect 19640 14172 19704 14176
rect 19640 14116 19644 14172
rect 19644 14116 19700 14172
rect 19700 14116 19704 14172
rect 19640 14112 19704 14116
rect 19720 14172 19784 14176
rect 19720 14116 19724 14172
rect 19724 14116 19780 14172
rect 19780 14116 19784 14172
rect 19720 14112 19784 14116
rect 5584 13628 5648 13632
rect 5584 13572 5588 13628
rect 5588 13572 5644 13628
rect 5644 13572 5648 13628
rect 5584 13568 5648 13572
rect 5664 13628 5728 13632
rect 5664 13572 5668 13628
rect 5668 13572 5724 13628
rect 5724 13572 5728 13628
rect 5664 13568 5728 13572
rect 5744 13628 5808 13632
rect 5744 13572 5748 13628
rect 5748 13572 5804 13628
rect 5804 13572 5808 13628
rect 5744 13568 5808 13572
rect 5824 13628 5888 13632
rect 5824 13572 5828 13628
rect 5828 13572 5884 13628
rect 5884 13572 5888 13628
rect 5824 13568 5888 13572
rect 14848 13628 14912 13632
rect 14848 13572 14852 13628
rect 14852 13572 14908 13628
rect 14908 13572 14912 13628
rect 14848 13568 14912 13572
rect 14928 13628 14992 13632
rect 14928 13572 14932 13628
rect 14932 13572 14988 13628
rect 14988 13572 14992 13628
rect 14928 13568 14992 13572
rect 15008 13628 15072 13632
rect 15008 13572 15012 13628
rect 15012 13572 15068 13628
rect 15068 13572 15072 13628
rect 15008 13568 15072 13572
rect 15088 13628 15152 13632
rect 15088 13572 15092 13628
rect 15092 13572 15148 13628
rect 15148 13572 15152 13628
rect 15088 13568 15152 13572
rect 24112 13628 24176 13632
rect 24112 13572 24116 13628
rect 24116 13572 24172 13628
rect 24172 13572 24176 13628
rect 24112 13568 24176 13572
rect 24192 13628 24256 13632
rect 24192 13572 24196 13628
rect 24196 13572 24252 13628
rect 24252 13572 24256 13628
rect 24192 13568 24256 13572
rect 24272 13628 24336 13632
rect 24272 13572 24276 13628
rect 24276 13572 24332 13628
rect 24332 13572 24336 13628
rect 24272 13568 24336 13572
rect 24352 13628 24416 13632
rect 24352 13572 24356 13628
rect 24356 13572 24412 13628
rect 24412 13572 24416 13628
rect 24352 13568 24416 13572
rect 10216 13084 10280 13088
rect 10216 13028 10220 13084
rect 10220 13028 10276 13084
rect 10276 13028 10280 13084
rect 10216 13024 10280 13028
rect 10296 13084 10360 13088
rect 10296 13028 10300 13084
rect 10300 13028 10356 13084
rect 10356 13028 10360 13084
rect 10296 13024 10360 13028
rect 10376 13084 10440 13088
rect 10376 13028 10380 13084
rect 10380 13028 10436 13084
rect 10436 13028 10440 13084
rect 10376 13024 10440 13028
rect 10456 13084 10520 13088
rect 10456 13028 10460 13084
rect 10460 13028 10516 13084
rect 10516 13028 10520 13084
rect 10456 13024 10520 13028
rect 19480 13084 19544 13088
rect 19480 13028 19484 13084
rect 19484 13028 19540 13084
rect 19540 13028 19544 13084
rect 19480 13024 19544 13028
rect 19560 13084 19624 13088
rect 19560 13028 19564 13084
rect 19564 13028 19620 13084
rect 19620 13028 19624 13084
rect 19560 13024 19624 13028
rect 19640 13084 19704 13088
rect 19640 13028 19644 13084
rect 19644 13028 19700 13084
rect 19700 13028 19704 13084
rect 19640 13024 19704 13028
rect 19720 13084 19784 13088
rect 19720 13028 19724 13084
rect 19724 13028 19780 13084
rect 19780 13028 19784 13084
rect 19720 13024 19784 13028
rect 5584 12540 5648 12544
rect 5584 12484 5588 12540
rect 5588 12484 5644 12540
rect 5644 12484 5648 12540
rect 5584 12480 5648 12484
rect 5664 12540 5728 12544
rect 5664 12484 5668 12540
rect 5668 12484 5724 12540
rect 5724 12484 5728 12540
rect 5664 12480 5728 12484
rect 5744 12540 5808 12544
rect 5744 12484 5748 12540
rect 5748 12484 5804 12540
rect 5804 12484 5808 12540
rect 5744 12480 5808 12484
rect 5824 12540 5888 12544
rect 5824 12484 5828 12540
rect 5828 12484 5884 12540
rect 5884 12484 5888 12540
rect 5824 12480 5888 12484
rect 14848 12540 14912 12544
rect 14848 12484 14852 12540
rect 14852 12484 14908 12540
rect 14908 12484 14912 12540
rect 14848 12480 14912 12484
rect 14928 12540 14992 12544
rect 14928 12484 14932 12540
rect 14932 12484 14988 12540
rect 14988 12484 14992 12540
rect 14928 12480 14992 12484
rect 15008 12540 15072 12544
rect 15008 12484 15012 12540
rect 15012 12484 15068 12540
rect 15068 12484 15072 12540
rect 15008 12480 15072 12484
rect 15088 12540 15152 12544
rect 15088 12484 15092 12540
rect 15092 12484 15148 12540
rect 15148 12484 15152 12540
rect 15088 12480 15152 12484
rect 24112 12540 24176 12544
rect 24112 12484 24116 12540
rect 24116 12484 24172 12540
rect 24172 12484 24176 12540
rect 24112 12480 24176 12484
rect 24192 12540 24256 12544
rect 24192 12484 24196 12540
rect 24196 12484 24252 12540
rect 24252 12484 24256 12540
rect 24192 12480 24256 12484
rect 24272 12540 24336 12544
rect 24272 12484 24276 12540
rect 24276 12484 24332 12540
rect 24332 12484 24336 12540
rect 24272 12480 24336 12484
rect 24352 12540 24416 12544
rect 24352 12484 24356 12540
rect 24356 12484 24412 12540
rect 24412 12484 24416 12540
rect 24352 12480 24416 12484
rect 10216 11996 10280 12000
rect 10216 11940 10220 11996
rect 10220 11940 10276 11996
rect 10276 11940 10280 11996
rect 10216 11936 10280 11940
rect 10296 11996 10360 12000
rect 10296 11940 10300 11996
rect 10300 11940 10356 11996
rect 10356 11940 10360 11996
rect 10296 11936 10360 11940
rect 10376 11996 10440 12000
rect 10376 11940 10380 11996
rect 10380 11940 10436 11996
rect 10436 11940 10440 11996
rect 10376 11936 10440 11940
rect 10456 11996 10520 12000
rect 10456 11940 10460 11996
rect 10460 11940 10516 11996
rect 10516 11940 10520 11996
rect 10456 11936 10520 11940
rect 19480 11996 19544 12000
rect 19480 11940 19484 11996
rect 19484 11940 19540 11996
rect 19540 11940 19544 11996
rect 19480 11936 19544 11940
rect 19560 11996 19624 12000
rect 19560 11940 19564 11996
rect 19564 11940 19620 11996
rect 19620 11940 19624 11996
rect 19560 11936 19624 11940
rect 19640 11996 19704 12000
rect 19640 11940 19644 11996
rect 19644 11940 19700 11996
rect 19700 11940 19704 11996
rect 19640 11936 19704 11940
rect 19720 11996 19784 12000
rect 19720 11940 19724 11996
rect 19724 11940 19780 11996
rect 19780 11940 19784 11996
rect 19720 11936 19784 11940
rect 5584 11452 5648 11456
rect 5584 11396 5588 11452
rect 5588 11396 5644 11452
rect 5644 11396 5648 11452
rect 5584 11392 5648 11396
rect 5664 11452 5728 11456
rect 5664 11396 5668 11452
rect 5668 11396 5724 11452
rect 5724 11396 5728 11452
rect 5664 11392 5728 11396
rect 5744 11452 5808 11456
rect 5744 11396 5748 11452
rect 5748 11396 5804 11452
rect 5804 11396 5808 11452
rect 5744 11392 5808 11396
rect 5824 11452 5888 11456
rect 5824 11396 5828 11452
rect 5828 11396 5884 11452
rect 5884 11396 5888 11452
rect 5824 11392 5888 11396
rect 14848 11452 14912 11456
rect 14848 11396 14852 11452
rect 14852 11396 14908 11452
rect 14908 11396 14912 11452
rect 14848 11392 14912 11396
rect 14928 11452 14992 11456
rect 14928 11396 14932 11452
rect 14932 11396 14988 11452
rect 14988 11396 14992 11452
rect 14928 11392 14992 11396
rect 15008 11452 15072 11456
rect 15008 11396 15012 11452
rect 15012 11396 15068 11452
rect 15068 11396 15072 11452
rect 15008 11392 15072 11396
rect 15088 11452 15152 11456
rect 15088 11396 15092 11452
rect 15092 11396 15148 11452
rect 15148 11396 15152 11452
rect 15088 11392 15152 11396
rect 24112 11452 24176 11456
rect 24112 11396 24116 11452
rect 24116 11396 24172 11452
rect 24172 11396 24176 11452
rect 24112 11392 24176 11396
rect 24192 11452 24256 11456
rect 24192 11396 24196 11452
rect 24196 11396 24252 11452
rect 24252 11396 24256 11452
rect 24192 11392 24256 11396
rect 24272 11452 24336 11456
rect 24272 11396 24276 11452
rect 24276 11396 24332 11452
rect 24332 11396 24336 11452
rect 24272 11392 24336 11396
rect 24352 11452 24416 11456
rect 24352 11396 24356 11452
rect 24356 11396 24412 11452
rect 24412 11396 24416 11452
rect 24352 11392 24416 11396
rect 10216 10908 10280 10912
rect 10216 10852 10220 10908
rect 10220 10852 10276 10908
rect 10276 10852 10280 10908
rect 10216 10848 10280 10852
rect 10296 10908 10360 10912
rect 10296 10852 10300 10908
rect 10300 10852 10356 10908
rect 10356 10852 10360 10908
rect 10296 10848 10360 10852
rect 10376 10908 10440 10912
rect 10376 10852 10380 10908
rect 10380 10852 10436 10908
rect 10436 10852 10440 10908
rect 10376 10848 10440 10852
rect 10456 10908 10520 10912
rect 10456 10852 10460 10908
rect 10460 10852 10516 10908
rect 10516 10852 10520 10908
rect 10456 10848 10520 10852
rect 19480 10908 19544 10912
rect 19480 10852 19484 10908
rect 19484 10852 19540 10908
rect 19540 10852 19544 10908
rect 19480 10848 19544 10852
rect 19560 10908 19624 10912
rect 19560 10852 19564 10908
rect 19564 10852 19620 10908
rect 19620 10852 19624 10908
rect 19560 10848 19624 10852
rect 19640 10908 19704 10912
rect 19640 10852 19644 10908
rect 19644 10852 19700 10908
rect 19700 10852 19704 10908
rect 19640 10848 19704 10852
rect 19720 10908 19784 10912
rect 19720 10852 19724 10908
rect 19724 10852 19780 10908
rect 19780 10852 19784 10908
rect 19720 10848 19784 10852
rect 5584 10364 5648 10368
rect 5584 10308 5588 10364
rect 5588 10308 5644 10364
rect 5644 10308 5648 10364
rect 5584 10304 5648 10308
rect 5664 10364 5728 10368
rect 5664 10308 5668 10364
rect 5668 10308 5724 10364
rect 5724 10308 5728 10364
rect 5664 10304 5728 10308
rect 5744 10364 5808 10368
rect 5744 10308 5748 10364
rect 5748 10308 5804 10364
rect 5804 10308 5808 10364
rect 5744 10304 5808 10308
rect 5824 10364 5888 10368
rect 5824 10308 5828 10364
rect 5828 10308 5884 10364
rect 5884 10308 5888 10364
rect 5824 10304 5888 10308
rect 14848 10364 14912 10368
rect 14848 10308 14852 10364
rect 14852 10308 14908 10364
rect 14908 10308 14912 10364
rect 14848 10304 14912 10308
rect 14928 10364 14992 10368
rect 14928 10308 14932 10364
rect 14932 10308 14988 10364
rect 14988 10308 14992 10364
rect 14928 10304 14992 10308
rect 15008 10364 15072 10368
rect 15008 10308 15012 10364
rect 15012 10308 15068 10364
rect 15068 10308 15072 10364
rect 15008 10304 15072 10308
rect 15088 10364 15152 10368
rect 15088 10308 15092 10364
rect 15092 10308 15148 10364
rect 15148 10308 15152 10364
rect 15088 10304 15152 10308
rect 24112 10364 24176 10368
rect 24112 10308 24116 10364
rect 24116 10308 24172 10364
rect 24172 10308 24176 10364
rect 24112 10304 24176 10308
rect 24192 10364 24256 10368
rect 24192 10308 24196 10364
rect 24196 10308 24252 10364
rect 24252 10308 24256 10364
rect 24192 10304 24256 10308
rect 24272 10364 24336 10368
rect 24272 10308 24276 10364
rect 24276 10308 24332 10364
rect 24332 10308 24336 10364
rect 24272 10304 24336 10308
rect 24352 10364 24416 10368
rect 24352 10308 24356 10364
rect 24356 10308 24412 10364
rect 24412 10308 24416 10364
rect 24352 10304 24416 10308
rect 10216 9820 10280 9824
rect 10216 9764 10220 9820
rect 10220 9764 10276 9820
rect 10276 9764 10280 9820
rect 10216 9760 10280 9764
rect 10296 9820 10360 9824
rect 10296 9764 10300 9820
rect 10300 9764 10356 9820
rect 10356 9764 10360 9820
rect 10296 9760 10360 9764
rect 10376 9820 10440 9824
rect 10376 9764 10380 9820
rect 10380 9764 10436 9820
rect 10436 9764 10440 9820
rect 10376 9760 10440 9764
rect 10456 9820 10520 9824
rect 10456 9764 10460 9820
rect 10460 9764 10516 9820
rect 10516 9764 10520 9820
rect 10456 9760 10520 9764
rect 19480 9820 19544 9824
rect 19480 9764 19484 9820
rect 19484 9764 19540 9820
rect 19540 9764 19544 9820
rect 19480 9760 19544 9764
rect 19560 9820 19624 9824
rect 19560 9764 19564 9820
rect 19564 9764 19620 9820
rect 19620 9764 19624 9820
rect 19560 9760 19624 9764
rect 19640 9820 19704 9824
rect 19640 9764 19644 9820
rect 19644 9764 19700 9820
rect 19700 9764 19704 9820
rect 19640 9760 19704 9764
rect 19720 9820 19784 9824
rect 19720 9764 19724 9820
rect 19724 9764 19780 9820
rect 19780 9764 19784 9820
rect 19720 9760 19784 9764
rect 5584 9276 5648 9280
rect 5584 9220 5588 9276
rect 5588 9220 5644 9276
rect 5644 9220 5648 9276
rect 5584 9216 5648 9220
rect 5664 9276 5728 9280
rect 5664 9220 5668 9276
rect 5668 9220 5724 9276
rect 5724 9220 5728 9276
rect 5664 9216 5728 9220
rect 5744 9276 5808 9280
rect 5744 9220 5748 9276
rect 5748 9220 5804 9276
rect 5804 9220 5808 9276
rect 5744 9216 5808 9220
rect 5824 9276 5888 9280
rect 5824 9220 5828 9276
rect 5828 9220 5884 9276
rect 5884 9220 5888 9276
rect 5824 9216 5888 9220
rect 14848 9276 14912 9280
rect 14848 9220 14852 9276
rect 14852 9220 14908 9276
rect 14908 9220 14912 9276
rect 14848 9216 14912 9220
rect 14928 9276 14992 9280
rect 14928 9220 14932 9276
rect 14932 9220 14988 9276
rect 14988 9220 14992 9276
rect 14928 9216 14992 9220
rect 15008 9276 15072 9280
rect 15008 9220 15012 9276
rect 15012 9220 15068 9276
rect 15068 9220 15072 9276
rect 15008 9216 15072 9220
rect 15088 9276 15152 9280
rect 15088 9220 15092 9276
rect 15092 9220 15148 9276
rect 15148 9220 15152 9276
rect 15088 9216 15152 9220
rect 24112 9276 24176 9280
rect 24112 9220 24116 9276
rect 24116 9220 24172 9276
rect 24172 9220 24176 9276
rect 24112 9216 24176 9220
rect 24192 9276 24256 9280
rect 24192 9220 24196 9276
rect 24196 9220 24252 9276
rect 24252 9220 24256 9276
rect 24192 9216 24256 9220
rect 24272 9276 24336 9280
rect 24272 9220 24276 9276
rect 24276 9220 24332 9276
rect 24332 9220 24336 9276
rect 24272 9216 24336 9220
rect 24352 9276 24416 9280
rect 24352 9220 24356 9276
rect 24356 9220 24412 9276
rect 24412 9220 24416 9276
rect 24352 9216 24416 9220
rect 10216 8732 10280 8736
rect 10216 8676 10220 8732
rect 10220 8676 10276 8732
rect 10276 8676 10280 8732
rect 10216 8672 10280 8676
rect 10296 8732 10360 8736
rect 10296 8676 10300 8732
rect 10300 8676 10356 8732
rect 10356 8676 10360 8732
rect 10296 8672 10360 8676
rect 10376 8732 10440 8736
rect 10376 8676 10380 8732
rect 10380 8676 10436 8732
rect 10436 8676 10440 8732
rect 10376 8672 10440 8676
rect 10456 8732 10520 8736
rect 10456 8676 10460 8732
rect 10460 8676 10516 8732
rect 10516 8676 10520 8732
rect 10456 8672 10520 8676
rect 19480 8732 19544 8736
rect 19480 8676 19484 8732
rect 19484 8676 19540 8732
rect 19540 8676 19544 8732
rect 19480 8672 19544 8676
rect 19560 8732 19624 8736
rect 19560 8676 19564 8732
rect 19564 8676 19620 8732
rect 19620 8676 19624 8732
rect 19560 8672 19624 8676
rect 19640 8732 19704 8736
rect 19640 8676 19644 8732
rect 19644 8676 19700 8732
rect 19700 8676 19704 8732
rect 19640 8672 19704 8676
rect 19720 8732 19784 8736
rect 19720 8676 19724 8732
rect 19724 8676 19780 8732
rect 19780 8676 19784 8732
rect 19720 8672 19784 8676
rect 5584 8188 5648 8192
rect 5584 8132 5588 8188
rect 5588 8132 5644 8188
rect 5644 8132 5648 8188
rect 5584 8128 5648 8132
rect 5664 8188 5728 8192
rect 5664 8132 5668 8188
rect 5668 8132 5724 8188
rect 5724 8132 5728 8188
rect 5664 8128 5728 8132
rect 5744 8188 5808 8192
rect 5744 8132 5748 8188
rect 5748 8132 5804 8188
rect 5804 8132 5808 8188
rect 5744 8128 5808 8132
rect 5824 8188 5888 8192
rect 5824 8132 5828 8188
rect 5828 8132 5884 8188
rect 5884 8132 5888 8188
rect 5824 8128 5888 8132
rect 14848 8188 14912 8192
rect 14848 8132 14852 8188
rect 14852 8132 14908 8188
rect 14908 8132 14912 8188
rect 14848 8128 14912 8132
rect 14928 8188 14992 8192
rect 14928 8132 14932 8188
rect 14932 8132 14988 8188
rect 14988 8132 14992 8188
rect 14928 8128 14992 8132
rect 15008 8188 15072 8192
rect 15008 8132 15012 8188
rect 15012 8132 15068 8188
rect 15068 8132 15072 8188
rect 15008 8128 15072 8132
rect 15088 8188 15152 8192
rect 15088 8132 15092 8188
rect 15092 8132 15148 8188
rect 15148 8132 15152 8188
rect 15088 8128 15152 8132
rect 24112 8188 24176 8192
rect 24112 8132 24116 8188
rect 24116 8132 24172 8188
rect 24172 8132 24176 8188
rect 24112 8128 24176 8132
rect 24192 8188 24256 8192
rect 24192 8132 24196 8188
rect 24196 8132 24252 8188
rect 24252 8132 24256 8188
rect 24192 8128 24256 8132
rect 24272 8188 24336 8192
rect 24272 8132 24276 8188
rect 24276 8132 24332 8188
rect 24332 8132 24336 8188
rect 24272 8128 24336 8132
rect 24352 8188 24416 8192
rect 24352 8132 24356 8188
rect 24356 8132 24412 8188
rect 24412 8132 24416 8188
rect 24352 8128 24416 8132
rect 10216 7644 10280 7648
rect 10216 7588 10220 7644
rect 10220 7588 10276 7644
rect 10276 7588 10280 7644
rect 10216 7584 10280 7588
rect 10296 7644 10360 7648
rect 10296 7588 10300 7644
rect 10300 7588 10356 7644
rect 10356 7588 10360 7644
rect 10296 7584 10360 7588
rect 10376 7644 10440 7648
rect 10376 7588 10380 7644
rect 10380 7588 10436 7644
rect 10436 7588 10440 7644
rect 10376 7584 10440 7588
rect 10456 7644 10520 7648
rect 10456 7588 10460 7644
rect 10460 7588 10516 7644
rect 10516 7588 10520 7644
rect 10456 7584 10520 7588
rect 19480 7644 19544 7648
rect 19480 7588 19484 7644
rect 19484 7588 19540 7644
rect 19540 7588 19544 7644
rect 19480 7584 19544 7588
rect 19560 7644 19624 7648
rect 19560 7588 19564 7644
rect 19564 7588 19620 7644
rect 19620 7588 19624 7644
rect 19560 7584 19624 7588
rect 19640 7644 19704 7648
rect 19640 7588 19644 7644
rect 19644 7588 19700 7644
rect 19700 7588 19704 7644
rect 19640 7584 19704 7588
rect 19720 7644 19784 7648
rect 19720 7588 19724 7644
rect 19724 7588 19780 7644
rect 19780 7588 19784 7644
rect 19720 7584 19784 7588
rect 5584 7100 5648 7104
rect 5584 7044 5588 7100
rect 5588 7044 5644 7100
rect 5644 7044 5648 7100
rect 5584 7040 5648 7044
rect 5664 7100 5728 7104
rect 5664 7044 5668 7100
rect 5668 7044 5724 7100
rect 5724 7044 5728 7100
rect 5664 7040 5728 7044
rect 5744 7100 5808 7104
rect 5744 7044 5748 7100
rect 5748 7044 5804 7100
rect 5804 7044 5808 7100
rect 5744 7040 5808 7044
rect 5824 7100 5888 7104
rect 5824 7044 5828 7100
rect 5828 7044 5884 7100
rect 5884 7044 5888 7100
rect 5824 7040 5888 7044
rect 14848 7100 14912 7104
rect 14848 7044 14852 7100
rect 14852 7044 14908 7100
rect 14908 7044 14912 7100
rect 14848 7040 14912 7044
rect 14928 7100 14992 7104
rect 14928 7044 14932 7100
rect 14932 7044 14988 7100
rect 14988 7044 14992 7100
rect 14928 7040 14992 7044
rect 15008 7100 15072 7104
rect 15008 7044 15012 7100
rect 15012 7044 15068 7100
rect 15068 7044 15072 7100
rect 15008 7040 15072 7044
rect 15088 7100 15152 7104
rect 15088 7044 15092 7100
rect 15092 7044 15148 7100
rect 15148 7044 15152 7100
rect 15088 7040 15152 7044
rect 24112 7100 24176 7104
rect 24112 7044 24116 7100
rect 24116 7044 24172 7100
rect 24172 7044 24176 7100
rect 24112 7040 24176 7044
rect 24192 7100 24256 7104
rect 24192 7044 24196 7100
rect 24196 7044 24252 7100
rect 24252 7044 24256 7100
rect 24192 7040 24256 7044
rect 24272 7100 24336 7104
rect 24272 7044 24276 7100
rect 24276 7044 24332 7100
rect 24332 7044 24336 7100
rect 24272 7040 24336 7044
rect 24352 7100 24416 7104
rect 24352 7044 24356 7100
rect 24356 7044 24412 7100
rect 24412 7044 24416 7100
rect 24352 7040 24416 7044
rect 10216 6556 10280 6560
rect 10216 6500 10220 6556
rect 10220 6500 10276 6556
rect 10276 6500 10280 6556
rect 10216 6496 10280 6500
rect 10296 6556 10360 6560
rect 10296 6500 10300 6556
rect 10300 6500 10356 6556
rect 10356 6500 10360 6556
rect 10296 6496 10360 6500
rect 10376 6556 10440 6560
rect 10376 6500 10380 6556
rect 10380 6500 10436 6556
rect 10436 6500 10440 6556
rect 10376 6496 10440 6500
rect 10456 6556 10520 6560
rect 10456 6500 10460 6556
rect 10460 6500 10516 6556
rect 10516 6500 10520 6556
rect 10456 6496 10520 6500
rect 19480 6556 19544 6560
rect 19480 6500 19484 6556
rect 19484 6500 19540 6556
rect 19540 6500 19544 6556
rect 19480 6496 19544 6500
rect 19560 6556 19624 6560
rect 19560 6500 19564 6556
rect 19564 6500 19620 6556
rect 19620 6500 19624 6556
rect 19560 6496 19624 6500
rect 19640 6556 19704 6560
rect 19640 6500 19644 6556
rect 19644 6500 19700 6556
rect 19700 6500 19704 6556
rect 19640 6496 19704 6500
rect 19720 6556 19784 6560
rect 19720 6500 19724 6556
rect 19724 6500 19780 6556
rect 19780 6500 19784 6556
rect 19720 6496 19784 6500
rect 5584 6012 5648 6016
rect 5584 5956 5588 6012
rect 5588 5956 5644 6012
rect 5644 5956 5648 6012
rect 5584 5952 5648 5956
rect 5664 6012 5728 6016
rect 5664 5956 5668 6012
rect 5668 5956 5724 6012
rect 5724 5956 5728 6012
rect 5664 5952 5728 5956
rect 5744 6012 5808 6016
rect 5744 5956 5748 6012
rect 5748 5956 5804 6012
rect 5804 5956 5808 6012
rect 5744 5952 5808 5956
rect 5824 6012 5888 6016
rect 5824 5956 5828 6012
rect 5828 5956 5884 6012
rect 5884 5956 5888 6012
rect 5824 5952 5888 5956
rect 14848 6012 14912 6016
rect 14848 5956 14852 6012
rect 14852 5956 14908 6012
rect 14908 5956 14912 6012
rect 14848 5952 14912 5956
rect 14928 6012 14992 6016
rect 14928 5956 14932 6012
rect 14932 5956 14988 6012
rect 14988 5956 14992 6012
rect 14928 5952 14992 5956
rect 15008 6012 15072 6016
rect 15008 5956 15012 6012
rect 15012 5956 15068 6012
rect 15068 5956 15072 6012
rect 15008 5952 15072 5956
rect 15088 6012 15152 6016
rect 15088 5956 15092 6012
rect 15092 5956 15148 6012
rect 15148 5956 15152 6012
rect 15088 5952 15152 5956
rect 24112 6012 24176 6016
rect 24112 5956 24116 6012
rect 24116 5956 24172 6012
rect 24172 5956 24176 6012
rect 24112 5952 24176 5956
rect 24192 6012 24256 6016
rect 24192 5956 24196 6012
rect 24196 5956 24252 6012
rect 24252 5956 24256 6012
rect 24192 5952 24256 5956
rect 24272 6012 24336 6016
rect 24272 5956 24276 6012
rect 24276 5956 24332 6012
rect 24332 5956 24336 6012
rect 24272 5952 24336 5956
rect 24352 6012 24416 6016
rect 24352 5956 24356 6012
rect 24356 5956 24412 6012
rect 24412 5956 24416 6012
rect 24352 5952 24416 5956
rect 10216 5468 10280 5472
rect 10216 5412 10220 5468
rect 10220 5412 10276 5468
rect 10276 5412 10280 5468
rect 10216 5408 10280 5412
rect 10296 5468 10360 5472
rect 10296 5412 10300 5468
rect 10300 5412 10356 5468
rect 10356 5412 10360 5468
rect 10296 5408 10360 5412
rect 10376 5468 10440 5472
rect 10376 5412 10380 5468
rect 10380 5412 10436 5468
rect 10436 5412 10440 5468
rect 10376 5408 10440 5412
rect 10456 5468 10520 5472
rect 10456 5412 10460 5468
rect 10460 5412 10516 5468
rect 10516 5412 10520 5468
rect 10456 5408 10520 5412
rect 19480 5468 19544 5472
rect 19480 5412 19484 5468
rect 19484 5412 19540 5468
rect 19540 5412 19544 5468
rect 19480 5408 19544 5412
rect 19560 5468 19624 5472
rect 19560 5412 19564 5468
rect 19564 5412 19620 5468
rect 19620 5412 19624 5468
rect 19560 5408 19624 5412
rect 19640 5468 19704 5472
rect 19640 5412 19644 5468
rect 19644 5412 19700 5468
rect 19700 5412 19704 5468
rect 19640 5408 19704 5412
rect 19720 5468 19784 5472
rect 19720 5412 19724 5468
rect 19724 5412 19780 5468
rect 19780 5412 19784 5468
rect 19720 5408 19784 5412
rect 5584 4924 5648 4928
rect 5584 4868 5588 4924
rect 5588 4868 5644 4924
rect 5644 4868 5648 4924
rect 5584 4864 5648 4868
rect 5664 4924 5728 4928
rect 5664 4868 5668 4924
rect 5668 4868 5724 4924
rect 5724 4868 5728 4924
rect 5664 4864 5728 4868
rect 5744 4924 5808 4928
rect 5744 4868 5748 4924
rect 5748 4868 5804 4924
rect 5804 4868 5808 4924
rect 5744 4864 5808 4868
rect 5824 4924 5888 4928
rect 5824 4868 5828 4924
rect 5828 4868 5884 4924
rect 5884 4868 5888 4924
rect 5824 4864 5888 4868
rect 14848 4924 14912 4928
rect 14848 4868 14852 4924
rect 14852 4868 14908 4924
rect 14908 4868 14912 4924
rect 14848 4864 14912 4868
rect 14928 4924 14992 4928
rect 14928 4868 14932 4924
rect 14932 4868 14988 4924
rect 14988 4868 14992 4924
rect 14928 4864 14992 4868
rect 15008 4924 15072 4928
rect 15008 4868 15012 4924
rect 15012 4868 15068 4924
rect 15068 4868 15072 4924
rect 15008 4864 15072 4868
rect 15088 4924 15152 4928
rect 15088 4868 15092 4924
rect 15092 4868 15148 4924
rect 15148 4868 15152 4924
rect 15088 4864 15152 4868
rect 24112 4924 24176 4928
rect 24112 4868 24116 4924
rect 24116 4868 24172 4924
rect 24172 4868 24176 4924
rect 24112 4864 24176 4868
rect 24192 4924 24256 4928
rect 24192 4868 24196 4924
rect 24196 4868 24252 4924
rect 24252 4868 24256 4924
rect 24192 4864 24256 4868
rect 24272 4924 24336 4928
rect 24272 4868 24276 4924
rect 24276 4868 24332 4924
rect 24332 4868 24336 4924
rect 24272 4864 24336 4868
rect 24352 4924 24416 4928
rect 24352 4868 24356 4924
rect 24356 4868 24412 4924
rect 24412 4868 24416 4924
rect 24352 4864 24416 4868
rect 10216 4380 10280 4384
rect 10216 4324 10220 4380
rect 10220 4324 10276 4380
rect 10276 4324 10280 4380
rect 10216 4320 10280 4324
rect 10296 4380 10360 4384
rect 10296 4324 10300 4380
rect 10300 4324 10356 4380
rect 10356 4324 10360 4380
rect 10296 4320 10360 4324
rect 10376 4380 10440 4384
rect 10376 4324 10380 4380
rect 10380 4324 10436 4380
rect 10436 4324 10440 4380
rect 10376 4320 10440 4324
rect 10456 4380 10520 4384
rect 10456 4324 10460 4380
rect 10460 4324 10516 4380
rect 10516 4324 10520 4380
rect 10456 4320 10520 4324
rect 19480 4380 19544 4384
rect 19480 4324 19484 4380
rect 19484 4324 19540 4380
rect 19540 4324 19544 4380
rect 19480 4320 19544 4324
rect 19560 4380 19624 4384
rect 19560 4324 19564 4380
rect 19564 4324 19620 4380
rect 19620 4324 19624 4380
rect 19560 4320 19624 4324
rect 19640 4380 19704 4384
rect 19640 4324 19644 4380
rect 19644 4324 19700 4380
rect 19700 4324 19704 4380
rect 19640 4320 19704 4324
rect 19720 4380 19784 4384
rect 19720 4324 19724 4380
rect 19724 4324 19780 4380
rect 19780 4324 19784 4380
rect 19720 4320 19784 4324
rect 5584 3836 5648 3840
rect 5584 3780 5588 3836
rect 5588 3780 5644 3836
rect 5644 3780 5648 3836
rect 5584 3776 5648 3780
rect 5664 3836 5728 3840
rect 5664 3780 5668 3836
rect 5668 3780 5724 3836
rect 5724 3780 5728 3836
rect 5664 3776 5728 3780
rect 5744 3836 5808 3840
rect 5744 3780 5748 3836
rect 5748 3780 5804 3836
rect 5804 3780 5808 3836
rect 5744 3776 5808 3780
rect 5824 3836 5888 3840
rect 5824 3780 5828 3836
rect 5828 3780 5884 3836
rect 5884 3780 5888 3836
rect 5824 3776 5888 3780
rect 14848 3836 14912 3840
rect 14848 3780 14852 3836
rect 14852 3780 14908 3836
rect 14908 3780 14912 3836
rect 14848 3776 14912 3780
rect 14928 3836 14992 3840
rect 14928 3780 14932 3836
rect 14932 3780 14988 3836
rect 14988 3780 14992 3836
rect 14928 3776 14992 3780
rect 15008 3836 15072 3840
rect 15008 3780 15012 3836
rect 15012 3780 15068 3836
rect 15068 3780 15072 3836
rect 15008 3776 15072 3780
rect 15088 3836 15152 3840
rect 15088 3780 15092 3836
rect 15092 3780 15148 3836
rect 15148 3780 15152 3836
rect 15088 3776 15152 3780
rect 24112 3836 24176 3840
rect 24112 3780 24116 3836
rect 24116 3780 24172 3836
rect 24172 3780 24176 3836
rect 24112 3776 24176 3780
rect 24192 3836 24256 3840
rect 24192 3780 24196 3836
rect 24196 3780 24252 3836
rect 24252 3780 24256 3836
rect 24192 3776 24256 3780
rect 24272 3836 24336 3840
rect 24272 3780 24276 3836
rect 24276 3780 24332 3836
rect 24332 3780 24336 3836
rect 24272 3776 24336 3780
rect 24352 3836 24416 3840
rect 24352 3780 24356 3836
rect 24356 3780 24412 3836
rect 24412 3780 24416 3836
rect 24352 3776 24416 3780
rect 10216 3292 10280 3296
rect 10216 3236 10220 3292
rect 10220 3236 10276 3292
rect 10276 3236 10280 3292
rect 10216 3232 10280 3236
rect 10296 3292 10360 3296
rect 10296 3236 10300 3292
rect 10300 3236 10356 3292
rect 10356 3236 10360 3292
rect 10296 3232 10360 3236
rect 10376 3292 10440 3296
rect 10376 3236 10380 3292
rect 10380 3236 10436 3292
rect 10436 3236 10440 3292
rect 10376 3232 10440 3236
rect 10456 3292 10520 3296
rect 10456 3236 10460 3292
rect 10460 3236 10516 3292
rect 10516 3236 10520 3292
rect 10456 3232 10520 3236
rect 19480 3292 19544 3296
rect 19480 3236 19484 3292
rect 19484 3236 19540 3292
rect 19540 3236 19544 3292
rect 19480 3232 19544 3236
rect 19560 3292 19624 3296
rect 19560 3236 19564 3292
rect 19564 3236 19620 3292
rect 19620 3236 19624 3292
rect 19560 3232 19624 3236
rect 19640 3292 19704 3296
rect 19640 3236 19644 3292
rect 19644 3236 19700 3292
rect 19700 3236 19704 3292
rect 19640 3232 19704 3236
rect 19720 3292 19784 3296
rect 19720 3236 19724 3292
rect 19724 3236 19780 3292
rect 19780 3236 19784 3292
rect 19720 3232 19784 3236
rect 5584 2748 5648 2752
rect 5584 2692 5588 2748
rect 5588 2692 5644 2748
rect 5644 2692 5648 2748
rect 5584 2688 5648 2692
rect 5664 2748 5728 2752
rect 5664 2692 5668 2748
rect 5668 2692 5724 2748
rect 5724 2692 5728 2748
rect 5664 2688 5728 2692
rect 5744 2748 5808 2752
rect 5744 2692 5748 2748
rect 5748 2692 5804 2748
rect 5804 2692 5808 2748
rect 5744 2688 5808 2692
rect 5824 2748 5888 2752
rect 5824 2692 5828 2748
rect 5828 2692 5884 2748
rect 5884 2692 5888 2748
rect 5824 2688 5888 2692
rect 14848 2748 14912 2752
rect 14848 2692 14852 2748
rect 14852 2692 14908 2748
rect 14908 2692 14912 2748
rect 14848 2688 14912 2692
rect 14928 2748 14992 2752
rect 14928 2692 14932 2748
rect 14932 2692 14988 2748
rect 14988 2692 14992 2748
rect 14928 2688 14992 2692
rect 15008 2748 15072 2752
rect 15008 2692 15012 2748
rect 15012 2692 15068 2748
rect 15068 2692 15072 2748
rect 15008 2688 15072 2692
rect 15088 2748 15152 2752
rect 15088 2692 15092 2748
rect 15092 2692 15148 2748
rect 15148 2692 15152 2748
rect 15088 2688 15152 2692
rect 24112 2748 24176 2752
rect 24112 2692 24116 2748
rect 24116 2692 24172 2748
rect 24172 2692 24176 2748
rect 24112 2688 24176 2692
rect 24192 2748 24256 2752
rect 24192 2692 24196 2748
rect 24196 2692 24252 2748
rect 24252 2692 24256 2748
rect 24192 2688 24256 2692
rect 24272 2748 24336 2752
rect 24272 2692 24276 2748
rect 24276 2692 24332 2748
rect 24332 2692 24336 2748
rect 24272 2688 24336 2692
rect 24352 2748 24416 2752
rect 24352 2692 24356 2748
rect 24356 2692 24412 2748
rect 24412 2692 24416 2748
rect 24352 2688 24416 2692
rect 10216 2204 10280 2208
rect 10216 2148 10220 2204
rect 10220 2148 10276 2204
rect 10276 2148 10280 2204
rect 10216 2144 10280 2148
rect 10296 2204 10360 2208
rect 10296 2148 10300 2204
rect 10300 2148 10356 2204
rect 10356 2148 10360 2204
rect 10296 2144 10360 2148
rect 10376 2204 10440 2208
rect 10376 2148 10380 2204
rect 10380 2148 10436 2204
rect 10436 2148 10440 2204
rect 10376 2144 10440 2148
rect 10456 2204 10520 2208
rect 10456 2148 10460 2204
rect 10460 2148 10516 2204
rect 10516 2148 10520 2204
rect 10456 2144 10520 2148
rect 19480 2204 19544 2208
rect 19480 2148 19484 2204
rect 19484 2148 19540 2204
rect 19540 2148 19544 2204
rect 19480 2144 19544 2148
rect 19560 2204 19624 2208
rect 19560 2148 19564 2204
rect 19564 2148 19620 2204
rect 19620 2148 19624 2204
rect 19560 2144 19624 2148
rect 19640 2204 19704 2208
rect 19640 2148 19644 2204
rect 19644 2148 19700 2204
rect 19700 2148 19704 2204
rect 19640 2144 19704 2148
rect 19720 2204 19784 2208
rect 19720 2148 19724 2204
rect 19724 2148 19780 2204
rect 19780 2148 19784 2204
rect 19720 2144 19784 2148
<< metal4 >>
rect 5576 39744 5896 39760
rect 5576 39680 5584 39744
rect 5648 39680 5664 39744
rect 5728 39680 5744 39744
rect 5808 39680 5824 39744
rect 5888 39680 5896 39744
rect 5576 38656 5896 39680
rect 7603 39676 7669 39677
rect 7603 39612 7604 39676
rect 7668 39612 7669 39676
rect 7603 39611 7669 39612
rect 5576 38592 5584 38656
rect 5648 38592 5664 38656
rect 5728 38592 5744 38656
rect 5808 38592 5824 38656
rect 5888 38592 5896 38656
rect 5576 37568 5896 38592
rect 5576 37504 5584 37568
rect 5648 37504 5664 37568
rect 5728 37504 5744 37568
rect 5808 37504 5824 37568
rect 5888 37504 5896 37568
rect 5576 36480 5896 37504
rect 5576 36416 5584 36480
rect 5648 36416 5664 36480
rect 5728 36416 5744 36480
rect 5808 36416 5824 36480
rect 5888 36416 5896 36480
rect 5576 35392 5896 36416
rect 7606 35733 7666 39611
rect 10208 39200 10528 39760
rect 14840 39744 15160 39760
rect 14840 39680 14848 39744
rect 14912 39680 14928 39744
rect 14992 39680 15008 39744
rect 15072 39680 15088 39744
rect 15152 39680 15160 39744
rect 11467 39268 11533 39269
rect 11467 39204 11468 39268
rect 11532 39204 11533 39268
rect 11467 39203 11533 39204
rect 10208 39136 10216 39200
rect 10280 39136 10296 39200
rect 10360 39136 10376 39200
rect 10440 39136 10456 39200
rect 10520 39136 10528 39200
rect 9995 38724 10061 38725
rect 9995 38660 9996 38724
rect 10060 38660 10061 38724
rect 9995 38659 10061 38660
rect 9259 38588 9325 38589
rect 9259 38524 9260 38588
rect 9324 38524 9325 38588
rect 9259 38523 9325 38524
rect 7603 35732 7669 35733
rect 7603 35668 7604 35732
rect 7668 35668 7669 35732
rect 7603 35667 7669 35668
rect 5576 35328 5584 35392
rect 5648 35328 5664 35392
rect 5728 35328 5744 35392
rect 5808 35328 5824 35392
rect 5888 35328 5896 35392
rect 5576 34304 5896 35328
rect 9262 35325 9322 38523
rect 9627 37092 9693 37093
rect 9627 37028 9628 37092
rect 9692 37028 9693 37092
rect 9627 37027 9693 37028
rect 9259 35324 9325 35325
rect 9259 35260 9260 35324
rect 9324 35260 9325 35324
rect 9259 35259 9325 35260
rect 7235 34644 7301 34645
rect 7235 34580 7236 34644
rect 7300 34580 7301 34644
rect 7235 34579 7301 34580
rect 5576 34240 5584 34304
rect 5648 34240 5664 34304
rect 5728 34240 5744 34304
rect 5808 34240 5824 34304
rect 5888 34240 5896 34304
rect 5576 33216 5896 34240
rect 5576 33152 5584 33216
rect 5648 33152 5664 33216
rect 5728 33152 5744 33216
rect 5808 33152 5824 33216
rect 5888 33152 5896 33216
rect 5576 32128 5896 33152
rect 5576 32064 5584 32128
rect 5648 32064 5664 32128
rect 5728 32064 5744 32128
rect 5808 32064 5824 32128
rect 5888 32064 5896 32128
rect 5576 31040 5896 32064
rect 5576 30976 5584 31040
rect 5648 30976 5664 31040
rect 5728 30976 5744 31040
rect 5808 30976 5824 31040
rect 5888 30976 5896 31040
rect 5576 29952 5896 30976
rect 5576 29888 5584 29952
rect 5648 29888 5664 29952
rect 5728 29888 5744 29952
rect 5808 29888 5824 29952
rect 5888 29888 5896 29952
rect 5576 28864 5896 29888
rect 5576 28800 5584 28864
rect 5648 28800 5664 28864
rect 5728 28800 5744 28864
rect 5808 28800 5824 28864
rect 5888 28800 5896 28864
rect 5576 27776 5896 28800
rect 5576 27712 5584 27776
rect 5648 27712 5664 27776
rect 5728 27712 5744 27776
rect 5808 27712 5824 27776
rect 5888 27712 5896 27776
rect 5576 26688 5896 27712
rect 5576 26624 5584 26688
rect 5648 26624 5664 26688
rect 5728 26624 5744 26688
rect 5808 26624 5824 26688
rect 5888 26624 5896 26688
rect 5576 25600 5896 26624
rect 5576 25536 5584 25600
rect 5648 25536 5664 25600
rect 5728 25536 5744 25600
rect 5808 25536 5824 25600
rect 5888 25536 5896 25600
rect 5576 24512 5896 25536
rect 5576 24448 5584 24512
rect 5648 24448 5664 24512
rect 5728 24448 5744 24512
rect 5808 24448 5824 24512
rect 5888 24448 5896 24512
rect 5576 23424 5896 24448
rect 7238 23493 7298 34579
rect 9630 33829 9690 37027
rect 9811 36276 9877 36277
rect 9811 36212 9812 36276
rect 9876 36212 9877 36276
rect 9811 36211 9877 36212
rect 9814 35189 9874 36211
rect 9811 35188 9877 35189
rect 9811 35124 9812 35188
rect 9876 35124 9877 35188
rect 9811 35123 9877 35124
rect 9811 34780 9877 34781
rect 9811 34716 9812 34780
rect 9876 34716 9877 34780
rect 9811 34715 9877 34716
rect 9627 33828 9693 33829
rect 9627 33764 9628 33828
rect 9692 33764 9693 33828
rect 9627 33763 9693 33764
rect 9814 33149 9874 34715
rect 9811 33148 9877 33149
rect 9811 33084 9812 33148
rect 9876 33084 9877 33148
rect 9811 33083 9877 33084
rect 9811 31108 9877 31109
rect 9811 31044 9812 31108
rect 9876 31044 9877 31108
rect 9811 31043 9877 31044
rect 9814 29341 9874 31043
rect 9998 30429 10058 38659
rect 10208 38112 10528 39136
rect 10208 38048 10216 38112
rect 10280 38048 10296 38112
rect 10360 38048 10376 38112
rect 10440 38048 10456 38112
rect 10520 38048 10528 38112
rect 10208 37024 10528 38048
rect 10731 38044 10797 38045
rect 10731 37980 10732 38044
rect 10796 37980 10797 38044
rect 10731 37979 10797 37980
rect 10208 36960 10216 37024
rect 10280 36960 10296 37024
rect 10360 36960 10376 37024
rect 10440 36960 10456 37024
rect 10520 36960 10528 37024
rect 10208 35936 10528 36960
rect 10208 35872 10216 35936
rect 10280 35872 10296 35936
rect 10360 35872 10376 35936
rect 10440 35872 10456 35936
rect 10520 35872 10528 35936
rect 10208 34848 10528 35872
rect 10734 35322 10794 37979
rect 10915 36820 10981 36821
rect 10915 36756 10916 36820
rect 10980 36756 10981 36820
rect 10915 36755 10981 36756
rect 10208 34784 10216 34848
rect 10280 34784 10296 34848
rect 10360 34784 10376 34848
rect 10440 34784 10456 34848
rect 10520 34784 10528 34848
rect 10208 33760 10528 34784
rect 10208 33696 10216 33760
rect 10280 33696 10296 33760
rect 10360 33696 10376 33760
rect 10440 33696 10456 33760
rect 10520 33696 10528 33760
rect 10208 32672 10528 33696
rect 10596 35262 10794 35322
rect 10596 33554 10656 35262
rect 10731 34916 10797 34917
rect 10731 34852 10732 34916
rect 10796 34914 10797 34916
rect 10918 34914 10978 36755
rect 11470 36005 11530 39203
rect 14840 38656 15160 39680
rect 14840 38592 14848 38656
rect 14912 38592 14928 38656
rect 14992 38592 15008 38656
rect 15072 38592 15088 38656
rect 15152 38592 15160 38656
rect 12019 38588 12085 38589
rect 12019 38524 12020 38588
rect 12084 38524 12085 38588
rect 12019 38523 12085 38524
rect 12022 38450 12082 38523
rect 12022 38390 12266 38450
rect 12206 37773 12266 38390
rect 12203 37772 12269 37773
rect 12203 37708 12204 37772
rect 12268 37708 12269 37772
rect 12203 37707 12269 37708
rect 14840 37568 15160 38592
rect 14840 37504 14848 37568
rect 14912 37504 14928 37568
rect 14992 37504 15008 37568
rect 15072 37504 15088 37568
rect 15152 37504 15160 37568
rect 11651 37092 11717 37093
rect 11651 37028 11652 37092
rect 11716 37028 11717 37092
rect 11651 37027 11717 37028
rect 14043 37092 14109 37093
rect 14043 37028 14044 37092
rect 14108 37028 14109 37092
rect 14043 37027 14109 37028
rect 11654 36413 11714 37027
rect 12203 36684 12269 36685
rect 12203 36620 12204 36684
rect 12268 36620 12269 36684
rect 12203 36619 12269 36620
rect 12206 36413 12266 36619
rect 11651 36412 11717 36413
rect 11651 36348 11652 36412
rect 11716 36348 11717 36412
rect 11651 36347 11717 36348
rect 12203 36412 12269 36413
rect 12203 36348 12204 36412
rect 12268 36348 12269 36412
rect 12203 36347 12269 36348
rect 12019 36276 12085 36277
rect 12019 36212 12020 36276
rect 12084 36274 12085 36276
rect 13859 36276 13925 36277
rect 12084 36214 12266 36274
rect 12084 36212 12085 36214
rect 12019 36211 12085 36212
rect 11835 36140 11901 36141
rect 11835 36076 11836 36140
rect 11900 36076 11901 36140
rect 11835 36075 11901 36076
rect 11467 36004 11533 36005
rect 11467 35940 11468 36004
rect 11532 35940 11533 36004
rect 11467 35939 11533 35940
rect 11838 35050 11898 36075
rect 12206 36002 12266 36214
rect 13859 36212 13860 36276
rect 13924 36274 13925 36276
rect 14046 36274 14106 37027
rect 13924 36214 14106 36274
rect 13924 36212 13925 36214
rect 13859 36211 13925 36212
rect 12206 35942 13554 36002
rect 12387 35868 12453 35869
rect 12387 35866 12388 35868
rect 12022 35806 12388 35866
rect 12022 35325 12082 35806
rect 12387 35804 12388 35806
rect 12452 35804 12453 35868
rect 12387 35803 12453 35804
rect 12019 35324 12085 35325
rect 12019 35260 12020 35324
rect 12084 35260 12085 35324
rect 12019 35259 12085 35260
rect 13494 35053 13554 35942
rect 13491 35052 13557 35053
rect 11838 34990 12450 35050
rect 10796 34854 10978 34914
rect 10796 34852 10797 34854
rect 10731 34851 10797 34852
rect 11467 34780 11533 34781
rect 11467 34716 11468 34780
rect 11532 34716 11533 34780
rect 11467 34715 11533 34716
rect 12203 34780 12269 34781
rect 12203 34716 12204 34780
rect 12268 34716 12269 34780
rect 12203 34715 12269 34716
rect 11470 34642 11530 34715
rect 12206 34642 12266 34715
rect 11470 34582 12266 34642
rect 10915 34236 10981 34237
rect 10915 34172 10916 34236
rect 10980 34172 10981 34236
rect 12019 34236 12085 34237
rect 12019 34234 12020 34236
rect 10915 34171 10981 34172
rect 11838 34174 12020 34234
rect 10731 34100 10797 34101
rect 10731 34036 10732 34100
rect 10796 34036 10797 34100
rect 10918 34098 10978 34171
rect 10918 34038 11714 34098
rect 10731 34035 10797 34036
rect 10734 33690 10794 34035
rect 10734 33630 11162 33690
rect 10596 33494 10794 33554
rect 10208 32608 10216 32672
rect 10280 32608 10296 32672
rect 10360 32608 10376 32672
rect 10440 32608 10456 32672
rect 10520 32608 10528 32672
rect 10208 31584 10528 32608
rect 10208 31520 10216 31584
rect 10280 31520 10296 31584
rect 10360 31520 10376 31584
rect 10440 31520 10456 31584
rect 10520 31520 10528 31584
rect 10208 30496 10528 31520
rect 10734 31109 10794 33494
rect 10915 33284 10981 33285
rect 10915 33220 10916 33284
rect 10980 33220 10981 33284
rect 10915 33219 10981 33220
rect 10731 31108 10797 31109
rect 10731 31044 10732 31108
rect 10796 31044 10797 31108
rect 10731 31043 10797 31044
rect 10918 30973 10978 33219
rect 11102 32330 11162 33630
rect 11654 33285 11714 34038
rect 11467 33284 11533 33285
rect 11467 33220 11468 33284
rect 11532 33220 11533 33284
rect 11467 33219 11533 33220
rect 11651 33284 11717 33285
rect 11651 33220 11652 33284
rect 11716 33220 11717 33284
rect 11651 33219 11717 33220
rect 11470 33150 11530 33219
rect 11838 33150 11898 34174
rect 12019 34172 12020 34174
rect 12084 34172 12085 34236
rect 12019 34171 12085 34172
rect 12390 33965 12450 34990
rect 13491 34988 13492 35052
rect 13556 34988 13557 35052
rect 13491 34987 13557 34988
rect 12387 33964 12453 33965
rect 12387 33900 12388 33964
rect 12452 33900 12453 33964
rect 12387 33899 12453 33900
rect 13123 33692 13189 33693
rect 13123 33690 13124 33692
rect 11470 33090 11898 33150
rect 12574 33630 13124 33690
rect 12574 33013 12634 33630
rect 13123 33628 13124 33630
rect 13188 33628 13189 33692
rect 13123 33627 13189 33628
rect 13491 33284 13557 33285
rect 13491 33220 13492 33284
rect 13556 33220 13557 33284
rect 13491 33219 13557 33220
rect 12571 33012 12637 33013
rect 12571 32948 12572 33012
rect 12636 32948 12637 33012
rect 12571 32947 12637 32948
rect 13494 32605 13554 33219
rect 13491 32604 13557 32605
rect 13491 32540 13492 32604
rect 13556 32540 13557 32604
rect 13491 32539 13557 32540
rect 11102 32270 11530 32330
rect 11470 32197 11530 32270
rect 11283 32196 11349 32197
rect 11283 32132 11284 32196
rect 11348 32132 11349 32196
rect 11283 32131 11349 32132
rect 11467 32196 11533 32197
rect 11467 32132 11468 32196
rect 11532 32132 11533 32196
rect 11467 32131 11533 32132
rect 11286 31653 11346 32131
rect 13307 31924 13373 31925
rect 13307 31860 13308 31924
rect 13372 31860 13373 31924
rect 13307 31859 13373 31860
rect 11283 31652 11349 31653
rect 11283 31588 11284 31652
rect 11348 31588 11349 31652
rect 11283 31587 11349 31588
rect 10915 30972 10981 30973
rect 10915 30908 10916 30972
rect 10980 30908 10981 30972
rect 10915 30907 10981 30908
rect 10208 30432 10216 30496
rect 10280 30432 10296 30496
rect 10360 30432 10376 30496
rect 10440 30432 10456 30496
rect 10520 30432 10528 30496
rect 9995 30428 10061 30429
rect 9995 30364 9996 30428
rect 10060 30364 10061 30428
rect 9995 30363 10061 30364
rect 10208 29408 10528 30432
rect 13310 30290 13370 31859
rect 13859 31380 13925 31381
rect 13859 31316 13860 31380
rect 13924 31316 13925 31380
rect 13859 31315 13925 31316
rect 11654 30230 13370 30290
rect 11654 29477 11714 30230
rect 12203 30156 12269 30157
rect 12203 30092 12204 30156
rect 12268 30092 12269 30156
rect 12203 30091 12269 30092
rect 12206 29477 12266 30091
rect 11651 29476 11717 29477
rect 11651 29412 11652 29476
rect 11716 29412 11717 29476
rect 11651 29411 11717 29412
rect 12203 29476 12269 29477
rect 12203 29412 12204 29476
rect 12268 29412 12269 29476
rect 12203 29411 12269 29412
rect 10208 29344 10216 29408
rect 10280 29344 10296 29408
rect 10360 29344 10376 29408
rect 10440 29344 10456 29408
rect 10520 29344 10528 29408
rect 9811 29340 9877 29341
rect 9811 29276 9812 29340
rect 9876 29276 9877 29340
rect 9811 29275 9877 29276
rect 10208 28320 10528 29344
rect 12387 29204 12453 29205
rect 12387 29140 12388 29204
rect 12452 29140 12453 29204
rect 12387 29139 12453 29140
rect 12390 28930 12450 29139
rect 12571 28932 12637 28933
rect 12571 28930 12572 28932
rect 12390 28870 12572 28930
rect 12571 28868 12572 28870
rect 12636 28868 12637 28932
rect 13862 28930 13922 31315
rect 14046 30021 14106 36214
rect 14840 36480 15160 37504
rect 19472 39200 19792 39760
rect 19472 39136 19480 39200
rect 19544 39136 19560 39200
rect 19624 39136 19640 39200
rect 19704 39136 19720 39200
rect 19784 39136 19792 39200
rect 19472 38112 19792 39136
rect 24104 39744 24424 39760
rect 24104 39680 24112 39744
rect 24176 39680 24192 39744
rect 24256 39680 24272 39744
rect 24336 39680 24352 39744
rect 24416 39680 24424 39744
rect 24104 38656 24424 39680
rect 24104 38592 24112 38656
rect 24176 38592 24192 38656
rect 24256 38592 24272 38656
rect 24336 38592 24352 38656
rect 24416 38592 24424 38656
rect 19931 38316 19997 38317
rect 19931 38252 19932 38316
rect 19996 38252 19997 38316
rect 19931 38251 19997 38252
rect 19472 38048 19480 38112
rect 19544 38048 19560 38112
rect 19624 38048 19640 38112
rect 19704 38048 19720 38112
rect 19784 38048 19792 38112
rect 19195 37364 19261 37365
rect 19195 37300 19196 37364
rect 19260 37300 19261 37364
rect 19195 37299 19261 37300
rect 14840 36416 14848 36480
rect 14912 36416 14928 36480
rect 14992 36416 15008 36480
rect 15072 36416 15088 36480
rect 15152 36416 15160 36480
rect 14840 35392 15160 36416
rect 18643 36140 18709 36141
rect 18643 36076 18644 36140
rect 18708 36076 18709 36140
rect 18643 36075 18709 36076
rect 14840 35328 14848 35392
rect 14912 35328 14928 35392
rect 14992 35328 15008 35392
rect 15072 35328 15088 35392
rect 15152 35328 15160 35392
rect 14840 34304 15160 35328
rect 18646 35189 18706 36075
rect 19198 36005 19258 37299
rect 19472 37024 19792 38048
rect 19472 36960 19480 37024
rect 19544 36960 19560 37024
rect 19624 36960 19640 37024
rect 19704 36960 19720 37024
rect 19784 36960 19792 37024
rect 19195 36004 19261 36005
rect 19195 35940 19196 36004
rect 19260 35940 19261 36004
rect 19195 35939 19261 35940
rect 19472 35936 19792 36960
rect 19934 36957 19994 38251
rect 24104 37568 24424 38592
rect 24104 37504 24112 37568
rect 24176 37504 24192 37568
rect 24256 37504 24272 37568
rect 24336 37504 24352 37568
rect 24416 37504 24424 37568
rect 20115 37228 20181 37229
rect 20115 37164 20116 37228
rect 20180 37164 20181 37228
rect 20115 37163 20181 37164
rect 19931 36956 19997 36957
rect 19931 36892 19932 36956
rect 19996 36892 19997 36956
rect 19931 36891 19997 36892
rect 19472 35872 19480 35936
rect 19544 35872 19560 35936
rect 19624 35872 19640 35936
rect 19704 35872 19720 35936
rect 19784 35872 19792 35936
rect 18643 35188 18709 35189
rect 18643 35124 18644 35188
rect 18708 35124 18709 35188
rect 18643 35123 18709 35124
rect 14840 34240 14848 34304
rect 14912 34240 14928 34304
rect 14992 34240 15008 34304
rect 15072 34240 15088 34304
rect 15152 34240 15160 34304
rect 14411 33556 14477 33557
rect 14411 33492 14412 33556
rect 14476 33492 14477 33556
rect 14411 33491 14477 33492
rect 14043 30020 14109 30021
rect 14043 29956 14044 30020
rect 14108 29956 14109 30020
rect 14043 29955 14109 29956
rect 12571 28867 12637 28868
rect 13678 28870 13922 28930
rect 10208 28256 10216 28320
rect 10280 28256 10296 28320
rect 10360 28256 10376 28320
rect 10440 28256 10456 28320
rect 10520 28256 10528 28320
rect 10208 27232 10528 28256
rect 12755 27980 12821 27981
rect 12755 27916 12756 27980
rect 12820 27916 12821 27980
rect 12755 27915 12821 27916
rect 10208 27168 10216 27232
rect 10280 27168 10296 27232
rect 10360 27168 10376 27232
rect 10440 27168 10456 27232
rect 10520 27168 10528 27232
rect 10208 26144 10528 27168
rect 12758 27165 12818 27915
rect 12755 27164 12821 27165
rect 12755 27100 12756 27164
rect 12820 27100 12821 27164
rect 12755 27099 12821 27100
rect 12939 27164 13005 27165
rect 12939 27100 12940 27164
rect 13004 27100 13005 27164
rect 12939 27099 13005 27100
rect 12942 26349 13002 27099
rect 12939 26348 13005 26349
rect 12939 26284 12940 26348
rect 13004 26284 13005 26348
rect 12939 26283 13005 26284
rect 10208 26080 10216 26144
rect 10280 26080 10296 26144
rect 10360 26080 10376 26144
rect 10440 26080 10456 26144
rect 10520 26080 10528 26144
rect 10208 25056 10528 26080
rect 10208 24992 10216 25056
rect 10280 24992 10296 25056
rect 10360 24992 10376 25056
rect 10440 24992 10456 25056
rect 10520 24992 10528 25056
rect 10208 23968 10528 24992
rect 13678 24853 13738 28870
rect 14227 25940 14293 25941
rect 14227 25876 14228 25940
rect 14292 25876 14293 25940
rect 14227 25875 14293 25876
rect 13675 24852 13741 24853
rect 13675 24788 13676 24852
rect 13740 24788 13741 24852
rect 13675 24787 13741 24788
rect 14230 24173 14290 25875
rect 14227 24172 14293 24173
rect 14227 24108 14228 24172
rect 14292 24108 14293 24172
rect 14227 24107 14293 24108
rect 10208 23904 10216 23968
rect 10280 23904 10296 23968
rect 10360 23904 10376 23968
rect 10440 23904 10456 23968
rect 10520 23904 10528 23968
rect 7235 23492 7301 23493
rect 7235 23428 7236 23492
rect 7300 23428 7301 23492
rect 7235 23427 7301 23428
rect 5576 23360 5584 23424
rect 5648 23360 5664 23424
rect 5728 23360 5744 23424
rect 5808 23360 5824 23424
rect 5888 23360 5896 23424
rect 5576 22336 5896 23360
rect 5576 22272 5584 22336
rect 5648 22272 5664 22336
rect 5728 22272 5744 22336
rect 5808 22272 5824 22336
rect 5888 22272 5896 22336
rect 5576 21248 5896 22272
rect 5576 21184 5584 21248
rect 5648 21184 5664 21248
rect 5728 21184 5744 21248
rect 5808 21184 5824 21248
rect 5888 21184 5896 21248
rect 5576 20160 5896 21184
rect 5576 20096 5584 20160
rect 5648 20096 5664 20160
rect 5728 20096 5744 20160
rect 5808 20096 5824 20160
rect 5888 20096 5896 20160
rect 5576 19072 5896 20096
rect 5576 19008 5584 19072
rect 5648 19008 5664 19072
rect 5728 19008 5744 19072
rect 5808 19008 5824 19072
rect 5888 19008 5896 19072
rect 5576 17984 5896 19008
rect 5576 17920 5584 17984
rect 5648 17920 5664 17984
rect 5728 17920 5744 17984
rect 5808 17920 5824 17984
rect 5888 17920 5896 17984
rect 5576 16896 5896 17920
rect 5576 16832 5584 16896
rect 5648 16832 5664 16896
rect 5728 16832 5744 16896
rect 5808 16832 5824 16896
rect 5888 16832 5896 16896
rect 5576 15808 5896 16832
rect 5576 15744 5584 15808
rect 5648 15744 5664 15808
rect 5728 15744 5744 15808
rect 5808 15744 5824 15808
rect 5888 15744 5896 15808
rect 5576 14720 5896 15744
rect 5576 14656 5584 14720
rect 5648 14656 5664 14720
rect 5728 14656 5744 14720
rect 5808 14656 5824 14720
rect 5888 14656 5896 14720
rect 5576 13632 5896 14656
rect 5576 13568 5584 13632
rect 5648 13568 5664 13632
rect 5728 13568 5744 13632
rect 5808 13568 5824 13632
rect 5888 13568 5896 13632
rect 5576 12544 5896 13568
rect 5576 12480 5584 12544
rect 5648 12480 5664 12544
rect 5728 12480 5744 12544
rect 5808 12480 5824 12544
rect 5888 12480 5896 12544
rect 5576 11456 5896 12480
rect 5576 11392 5584 11456
rect 5648 11392 5664 11456
rect 5728 11392 5744 11456
rect 5808 11392 5824 11456
rect 5888 11392 5896 11456
rect 5576 10368 5896 11392
rect 5576 10304 5584 10368
rect 5648 10304 5664 10368
rect 5728 10304 5744 10368
rect 5808 10304 5824 10368
rect 5888 10304 5896 10368
rect 5576 9280 5896 10304
rect 5576 9216 5584 9280
rect 5648 9216 5664 9280
rect 5728 9216 5744 9280
rect 5808 9216 5824 9280
rect 5888 9216 5896 9280
rect 5576 8192 5896 9216
rect 5576 8128 5584 8192
rect 5648 8128 5664 8192
rect 5728 8128 5744 8192
rect 5808 8128 5824 8192
rect 5888 8128 5896 8192
rect 5576 7104 5896 8128
rect 5576 7040 5584 7104
rect 5648 7040 5664 7104
rect 5728 7040 5744 7104
rect 5808 7040 5824 7104
rect 5888 7040 5896 7104
rect 5576 6016 5896 7040
rect 5576 5952 5584 6016
rect 5648 5952 5664 6016
rect 5728 5952 5744 6016
rect 5808 5952 5824 6016
rect 5888 5952 5896 6016
rect 5576 4928 5896 5952
rect 5576 4864 5584 4928
rect 5648 4864 5664 4928
rect 5728 4864 5744 4928
rect 5808 4864 5824 4928
rect 5888 4864 5896 4928
rect 5576 3840 5896 4864
rect 5576 3776 5584 3840
rect 5648 3776 5664 3840
rect 5728 3776 5744 3840
rect 5808 3776 5824 3840
rect 5888 3776 5896 3840
rect 5576 2752 5896 3776
rect 5576 2688 5584 2752
rect 5648 2688 5664 2752
rect 5728 2688 5744 2752
rect 5808 2688 5824 2752
rect 5888 2688 5896 2752
rect 5576 2128 5896 2688
rect 10208 22880 10528 23904
rect 14414 23493 14474 33491
rect 14840 33216 15160 34240
rect 19472 34848 19792 35872
rect 19472 34784 19480 34848
rect 19544 34784 19560 34848
rect 19624 34784 19640 34848
rect 19704 34784 19720 34848
rect 19784 34784 19792 34848
rect 16435 34236 16501 34237
rect 16435 34172 16436 34236
rect 16500 34172 16501 34236
rect 16435 34171 16501 34172
rect 14840 33152 14848 33216
rect 14912 33152 14928 33216
rect 14992 33152 15008 33216
rect 15072 33152 15088 33216
rect 15152 33152 15160 33216
rect 14840 32128 15160 33152
rect 14840 32064 14848 32128
rect 14912 32064 14928 32128
rect 14992 32064 15008 32128
rect 15072 32064 15088 32128
rect 15152 32064 15160 32128
rect 14840 31040 15160 32064
rect 14840 30976 14848 31040
rect 14912 30976 14928 31040
rect 14992 30976 15008 31040
rect 15072 30976 15088 31040
rect 15152 30976 15160 31040
rect 14840 29952 15160 30976
rect 14840 29888 14848 29952
rect 14912 29888 14928 29952
rect 14992 29888 15008 29952
rect 15072 29888 15088 29952
rect 15152 29888 15160 29952
rect 14840 28864 15160 29888
rect 14840 28800 14848 28864
rect 14912 28800 14928 28864
rect 14992 28800 15008 28864
rect 15072 28800 15088 28864
rect 15152 28800 15160 28864
rect 14840 27776 15160 28800
rect 14840 27712 14848 27776
rect 14912 27712 14928 27776
rect 14992 27712 15008 27776
rect 15072 27712 15088 27776
rect 15152 27712 15160 27776
rect 14840 26688 15160 27712
rect 16438 27573 16498 34171
rect 19472 33760 19792 34784
rect 19934 34373 19994 36891
rect 19931 34372 19997 34373
rect 19931 34308 19932 34372
rect 19996 34308 19997 34372
rect 19931 34307 19997 34308
rect 19472 33696 19480 33760
rect 19544 33696 19560 33760
rect 19624 33696 19640 33760
rect 19704 33696 19720 33760
rect 19784 33696 19792 33760
rect 19472 32672 19792 33696
rect 19472 32608 19480 32672
rect 19544 32608 19560 32672
rect 19624 32608 19640 32672
rect 19704 32608 19720 32672
rect 19784 32608 19792 32672
rect 19472 31584 19792 32608
rect 19931 32060 19997 32061
rect 19931 31996 19932 32060
rect 19996 31996 19997 32060
rect 19931 31995 19997 31996
rect 19472 31520 19480 31584
rect 19544 31520 19560 31584
rect 19624 31520 19640 31584
rect 19704 31520 19720 31584
rect 19784 31520 19792 31584
rect 19472 30496 19792 31520
rect 19472 30432 19480 30496
rect 19544 30432 19560 30496
rect 19624 30432 19640 30496
rect 19704 30432 19720 30496
rect 19784 30432 19792 30496
rect 16987 30292 17053 30293
rect 16987 30228 16988 30292
rect 17052 30228 17053 30292
rect 16987 30227 17053 30228
rect 16803 29884 16869 29885
rect 16803 29820 16804 29884
rect 16868 29882 16869 29884
rect 16990 29882 17050 30227
rect 16868 29822 17050 29882
rect 16868 29820 16869 29822
rect 16803 29819 16869 29820
rect 19472 29408 19792 30432
rect 19934 29613 19994 31995
rect 20118 31789 20178 37163
rect 24104 36480 24424 37504
rect 24104 36416 24112 36480
rect 24176 36416 24192 36480
rect 24256 36416 24272 36480
rect 24336 36416 24352 36480
rect 24416 36416 24424 36480
rect 21035 35732 21101 35733
rect 21035 35668 21036 35732
rect 21100 35668 21101 35732
rect 21035 35667 21101 35668
rect 21038 34373 21098 35667
rect 24104 35392 24424 36416
rect 24104 35328 24112 35392
rect 24176 35328 24192 35392
rect 24256 35328 24272 35392
rect 24336 35328 24352 35392
rect 24416 35328 24424 35392
rect 21035 34372 21101 34373
rect 21035 34308 21036 34372
rect 21100 34308 21101 34372
rect 21035 34307 21101 34308
rect 24104 34304 24424 35328
rect 24104 34240 24112 34304
rect 24176 34240 24192 34304
rect 24256 34240 24272 34304
rect 24336 34240 24352 34304
rect 24416 34240 24424 34304
rect 24104 33216 24424 34240
rect 24104 33152 24112 33216
rect 24176 33152 24192 33216
rect 24256 33152 24272 33216
rect 24336 33152 24352 33216
rect 24416 33152 24424 33216
rect 24104 32128 24424 33152
rect 24104 32064 24112 32128
rect 24176 32064 24192 32128
rect 24256 32064 24272 32128
rect 24336 32064 24352 32128
rect 24416 32064 24424 32128
rect 20115 31788 20181 31789
rect 20115 31724 20116 31788
rect 20180 31724 20181 31788
rect 20115 31723 20181 31724
rect 24104 31040 24424 32064
rect 24104 30976 24112 31040
rect 24176 30976 24192 31040
rect 24256 30976 24272 31040
rect 24336 30976 24352 31040
rect 24416 30976 24424 31040
rect 24104 29952 24424 30976
rect 26555 30428 26621 30429
rect 26555 30364 26556 30428
rect 26620 30364 26621 30428
rect 26555 30363 26621 30364
rect 24104 29888 24112 29952
rect 24176 29888 24192 29952
rect 24256 29888 24272 29952
rect 24336 29888 24352 29952
rect 24416 29888 24424 29952
rect 19931 29612 19997 29613
rect 19931 29548 19932 29612
rect 19996 29548 19997 29612
rect 19931 29547 19997 29548
rect 22139 29476 22205 29477
rect 22139 29412 22140 29476
rect 22204 29412 22205 29476
rect 22139 29411 22205 29412
rect 19472 29344 19480 29408
rect 19544 29344 19560 29408
rect 19624 29344 19640 29408
rect 19704 29344 19720 29408
rect 19784 29344 19792 29408
rect 18459 29068 18525 29069
rect 18459 29004 18460 29068
rect 18524 29004 18525 29068
rect 18459 29003 18525 29004
rect 16987 28660 17053 28661
rect 16987 28596 16988 28660
rect 17052 28596 17053 28660
rect 16987 28595 17053 28596
rect 16435 27572 16501 27573
rect 16435 27508 16436 27572
rect 16500 27508 16501 27572
rect 16435 27507 16501 27508
rect 14840 26624 14848 26688
rect 14912 26624 14928 26688
rect 14992 26624 15008 26688
rect 15072 26624 15088 26688
rect 15152 26624 15160 26688
rect 14840 25600 15160 26624
rect 16619 26348 16685 26349
rect 16619 26284 16620 26348
rect 16684 26284 16685 26348
rect 16619 26283 16685 26284
rect 14840 25536 14848 25600
rect 14912 25536 14928 25600
rect 14992 25536 15008 25600
rect 15072 25536 15088 25600
rect 15152 25536 15160 25600
rect 14840 24512 15160 25536
rect 14840 24448 14848 24512
rect 14912 24448 14928 24512
rect 14992 24448 15008 24512
rect 15072 24448 15088 24512
rect 15152 24448 15160 24512
rect 14411 23492 14477 23493
rect 14411 23428 14412 23492
rect 14476 23428 14477 23492
rect 14411 23427 14477 23428
rect 10208 22816 10216 22880
rect 10280 22816 10296 22880
rect 10360 22816 10376 22880
rect 10440 22816 10456 22880
rect 10520 22816 10528 22880
rect 10208 21792 10528 22816
rect 10208 21728 10216 21792
rect 10280 21728 10296 21792
rect 10360 21728 10376 21792
rect 10440 21728 10456 21792
rect 10520 21728 10528 21792
rect 10208 20704 10528 21728
rect 10208 20640 10216 20704
rect 10280 20640 10296 20704
rect 10360 20640 10376 20704
rect 10440 20640 10456 20704
rect 10520 20640 10528 20704
rect 10208 19616 10528 20640
rect 10208 19552 10216 19616
rect 10280 19552 10296 19616
rect 10360 19552 10376 19616
rect 10440 19552 10456 19616
rect 10520 19552 10528 19616
rect 10208 18528 10528 19552
rect 10208 18464 10216 18528
rect 10280 18464 10296 18528
rect 10360 18464 10376 18528
rect 10440 18464 10456 18528
rect 10520 18464 10528 18528
rect 10208 17440 10528 18464
rect 10208 17376 10216 17440
rect 10280 17376 10296 17440
rect 10360 17376 10376 17440
rect 10440 17376 10456 17440
rect 10520 17376 10528 17440
rect 10208 16352 10528 17376
rect 10208 16288 10216 16352
rect 10280 16288 10296 16352
rect 10360 16288 10376 16352
rect 10440 16288 10456 16352
rect 10520 16288 10528 16352
rect 10208 15264 10528 16288
rect 10208 15200 10216 15264
rect 10280 15200 10296 15264
rect 10360 15200 10376 15264
rect 10440 15200 10456 15264
rect 10520 15200 10528 15264
rect 10208 14176 10528 15200
rect 10208 14112 10216 14176
rect 10280 14112 10296 14176
rect 10360 14112 10376 14176
rect 10440 14112 10456 14176
rect 10520 14112 10528 14176
rect 10208 13088 10528 14112
rect 10208 13024 10216 13088
rect 10280 13024 10296 13088
rect 10360 13024 10376 13088
rect 10440 13024 10456 13088
rect 10520 13024 10528 13088
rect 10208 12000 10528 13024
rect 10208 11936 10216 12000
rect 10280 11936 10296 12000
rect 10360 11936 10376 12000
rect 10440 11936 10456 12000
rect 10520 11936 10528 12000
rect 10208 10912 10528 11936
rect 10208 10848 10216 10912
rect 10280 10848 10296 10912
rect 10360 10848 10376 10912
rect 10440 10848 10456 10912
rect 10520 10848 10528 10912
rect 10208 9824 10528 10848
rect 10208 9760 10216 9824
rect 10280 9760 10296 9824
rect 10360 9760 10376 9824
rect 10440 9760 10456 9824
rect 10520 9760 10528 9824
rect 10208 8736 10528 9760
rect 10208 8672 10216 8736
rect 10280 8672 10296 8736
rect 10360 8672 10376 8736
rect 10440 8672 10456 8736
rect 10520 8672 10528 8736
rect 10208 7648 10528 8672
rect 10208 7584 10216 7648
rect 10280 7584 10296 7648
rect 10360 7584 10376 7648
rect 10440 7584 10456 7648
rect 10520 7584 10528 7648
rect 10208 6560 10528 7584
rect 10208 6496 10216 6560
rect 10280 6496 10296 6560
rect 10360 6496 10376 6560
rect 10440 6496 10456 6560
rect 10520 6496 10528 6560
rect 10208 5472 10528 6496
rect 10208 5408 10216 5472
rect 10280 5408 10296 5472
rect 10360 5408 10376 5472
rect 10440 5408 10456 5472
rect 10520 5408 10528 5472
rect 10208 4384 10528 5408
rect 10208 4320 10216 4384
rect 10280 4320 10296 4384
rect 10360 4320 10376 4384
rect 10440 4320 10456 4384
rect 10520 4320 10528 4384
rect 10208 3296 10528 4320
rect 10208 3232 10216 3296
rect 10280 3232 10296 3296
rect 10360 3232 10376 3296
rect 10440 3232 10456 3296
rect 10520 3232 10528 3296
rect 10208 2208 10528 3232
rect 10208 2144 10216 2208
rect 10280 2144 10296 2208
rect 10360 2144 10376 2208
rect 10440 2144 10456 2208
rect 10520 2144 10528 2208
rect 10208 2128 10528 2144
rect 14840 23424 15160 24448
rect 15515 23900 15581 23901
rect 15515 23836 15516 23900
rect 15580 23836 15581 23900
rect 15515 23835 15581 23836
rect 15518 23629 15578 23835
rect 15515 23628 15581 23629
rect 15515 23564 15516 23628
rect 15580 23564 15581 23628
rect 15515 23563 15581 23564
rect 14840 23360 14848 23424
rect 14912 23360 14928 23424
rect 14992 23360 15008 23424
rect 15072 23360 15088 23424
rect 15152 23360 15160 23424
rect 14840 22336 15160 23360
rect 14840 22272 14848 22336
rect 14912 22272 14928 22336
rect 14992 22272 15008 22336
rect 15072 22272 15088 22336
rect 15152 22272 15160 22336
rect 14840 21248 15160 22272
rect 14840 21184 14848 21248
rect 14912 21184 14928 21248
rect 14992 21184 15008 21248
rect 15072 21184 15088 21248
rect 15152 21184 15160 21248
rect 14840 20160 15160 21184
rect 16622 20501 16682 26283
rect 16990 25533 17050 28595
rect 16987 25532 17053 25533
rect 16987 25468 16988 25532
rect 17052 25468 17053 25532
rect 16987 25467 17053 25468
rect 16990 20909 17050 25467
rect 16987 20908 17053 20909
rect 16987 20844 16988 20908
rect 17052 20844 17053 20908
rect 16987 20843 17053 20844
rect 16619 20500 16685 20501
rect 16619 20436 16620 20500
rect 16684 20436 16685 20500
rect 16619 20435 16685 20436
rect 14840 20096 14848 20160
rect 14912 20096 14928 20160
rect 14992 20096 15008 20160
rect 15072 20096 15088 20160
rect 15152 20096 15160 20160
rect 14840 19072 15160 20096
rect 14840 19008 14848 19072
rect 14912 19008 14928 19072
rect 14992 19008 15008 19072
rect 15072 19008 15088 19072
rect 15152 19008 15160 19072
rect 14840 17984 15160 19008
rect 14840 17920 14848 17984
rect 14912 17920 14928 17984
rect 14992 17920 15008 17984
rect 15072 17920 15088 17984
rect 15152 17920 15160 17984
rect 14840 16896 15160 17920
rect 18462 17781 18522 29003
rect 19472 28320 19792 29344
rect 20115 28932 20181 28933
rect 20115 28868 20116 28932
rect 20180 28868 20181 28932
rect 20115 28867 20181 28868
rect 19931 28660 19997 28661
rect 19931 28596 19932 28660
rect 19996 28596 19997 28660
rect 19931 28595 19997 28596
rect 19472 28256 19480 28320
rect 19544 28256 19560 28320
rect 19624 28256 19640 28320
rect 19704 28256 19720 28320
rect 19784 28256 19792 28320
rect 19472 27232 19792 28256
rect 19472 27168 19480 27232
rect 19544 27168 19560 27232
rect 19624 27168 19640 27232
rect 19704 27168 19720 27232
rect 19784 27168 19792 27232
rect 19472 26144 19792 27168
rect 19472 26080 19480 26144
rect 19544 26080 19560 26144
rect 19624 26080 19640 26144
rect 19704 26080 19720 26144
rect 19784 26080 19792 26144
rect 18643 25260 18709 25261
rect 18643 25196 18644 25260
rect 18708 25196 18709 25260
rect 18643 25195 18709 25196
rect 18459 17780 18525 17781
rect 18459 17716 18460 17780
rect 18524 17716 18525 17780
rect 18459 17715 18525 17716
rect 14840 16832 14848 16896
rect 14912 16832 14928 16896
rect 14992 16832 15008 16896
rect 15072 16832 15088 16896
rect 15152 16832 15160 16896
rect 14840 15808 15160 16832
rect 18646 16149 18706 25195
rect 19472 25056 19792 26080
rect 19934 25669 19994 28595
rect 20118 26485 20178 28867
rect 20115 26484 20181 26485
rect 20115 26420 20116 26484
rect 20180 26420 20181 26484
rect 20115 26419 20181 26420
rect 19931 25668 19997 25669
rect 19931 25604 19932 25668
rect 19996 25604 19997 25668
rect 19931 25603 19997 25604
rect 19472 24992 19480 25056
rect 19544 24992 19560 25056
rect 19624 24992 19640 25056
rect 19704 24992 19720 25056
rect 19784 24992 19792 25056
rect 19472 23968 19792 24992
rect 19472 23904 19480 23968
rect 19544 23904 19560 23968
rect 19624 23904 19640 23968
rect 19704 23904 19720 23968
rect 19784 23904 19792 23968
rect 19472 22880 19792 23904
rect 19472 22816 19480 22880
rect 19544 22816 19560 22880
rect 19624 22816 19640 22880
rect 19704 22816 19720 22880
rect 19784 22816 19792 22880
rect 19472 21792 19792 22816
rect 22142 22133 22202 29411
rect 24104 28864 24424 29888
rect 24104 28800 24112 28864
rect 24176 28800 24192 28864
rect 24256 28800 24272 28864
rect 24336 28800 24352 28864
rect 24416 28800 24424 28864
rect 24104 27776 24424 28800
rect 24531 28252 24597 28253
rect 24531 28188 24532 28252
rect 24596 28188 24597 28252
rect 24531 28187 24597 28188
rect 24104 27712 24112 27776
rect 24176 27712 24192 27776
rect 24256 27712 24272 27776
rect 24336 27712 24352 27776
rect 24416 27712 24424 27776
rect 24104 26688 24424 27712
rect 24104 26624 24112 26688
rect 24176 26624 24192 26688
rect 24256 26624 24272 26688
rect 24336 26624 24352 26688
rect 24416 26624 24424 26688
rect 24104 25600 24424 26624
rect 24104 25536 24112 25600
rect 24176 25536 24192 25600
rect 24256 25536 24272 25600
rect 24336 25536 24352 25600
rect 24416 25536 24424 25600
rect 23611 25396 23677 25397
rect 23611 25332 23612 25396
rect 23676 25332 23677 25396
rect 23611 25331 23677 25332
rect 23614 22133 23674 25331
rect 24104 24512 24424 25536
rect 24534 25125 24594 28187
rect 26187 27708 26253 27709
rect 26187 27644 26188 27708
rect 26252 27644 26253 27708
rect 26187 27643 26253 27644
rect 24531 25124 24597 25125
rect 24531 25060 24532 25124
rect 24596 25060 24597 25124
rect 24531 25059 24597 25060
rect 24104 24448 24112 24512
rect 24176 24448 24192 24512
rect 24256 24448 24272 24512
rect 24336 24448 24352 24512
rect 24416 24448 24424 24512
rect 24104 23424 24424 24448
rect 24104 23360 24112 23424
rect 24176 23360 24192 23424
rect 24256 23360 24272 23424
rect 24336 23360 24352 23424
rect 24416 23360 24424 23424
rect 24104 22336 24424 23360
rect 24534 23085 24594 25059
rect 24531 23084 24597 23085
rect 24531 23020 24532 23084
rect 24596 23020 24597 23084
rect 24531 23019 24597 23020
rect 24104 22272 24112 22336
rect 24176 22272 24192 22336
rect 24256 22272 24272 22336
rect 24336 22272 24352 22336
rect 24416 22272 24424 22336
rect 19931 22132 19997 22133
rect 19931 22068 19932 22132
rect 19996 22068 19997 22132
rect 19931 22067 19997 22068
rect 22139 22132 22205 22133
rect 22139 22068 22140 22132
rect 22204 22068 22205 22132
rect 22139 22067 22205 22068
rect 23611 22132 23677 22133
rect 23611 22068 23612 22132
rect 23676 22068 23677 22132
rect 23611 22067 23677 22068
rect 19472 21728 19480 21792
rect 19544 21728 19560 21792
rect 19624 21728 19640 21792
rect 19704 21728 19720 21792
rect 19784 21728 19792 21792
rect 19472 20704 19792 21728
rect 19934 21453 19994 22067
rect 19931 21452 19997 21453
rect 19931 21388 19932 21452
rect 19996 21388 19997 21452
rect 19931 21387 19997 21388
rect 19472 20640 19480 20704
rect 19544 20640 19560 20704
rect 19624 20640 19640 20704
rect 19704 20640 19720 20704
rect 19784 20640 19792 20704
rect 19472 19616 19792 20640
rect 22142 19957 22202 22067
rect 24104 21248 24424 22272
rect 24104 21184 24112 21248
rect 24176 21184 24192 21248
rect 24256 21184 24272 21248
rect 24336 21184 24352 21248
rect 24416 21184 24424 21248
rect 24104 20160 24424 21184
rect 24104 20096 24112 20160
rect 24176 20096 24192 20160
rect 24256 20096 24272 20160
rect 24336 20096 24352 20160
rect 24416 20096 24424 20160
rect 22139 19956 22205 19957
rect 22139 19892 22140 19956
rect 22204 19892 22205 19956
rect 22139 19891 22205 19892
rect 19472 19552 19480 19616
rect 19544 19552 19560 19616
rect 19624 19552 19640 19616
rect 19704 19552 19720 19616
rect 19784 19552 19792 19616
rect 19472 18528 19792 19552
rect 19472 18464 19480 18528
rect 19544 18464 19560 18528
rect 19624 18464 19640 18528
rect 19704 18464 19720 18528
rect 19784 18464 19792 18528
rect 19472 17440 19792 18464
rect 19472 17376 19480 17440
rect 19544 17376 19560 17440
rect 19624 17376 19640 17440
rect 19704 17376 19720 17440
rect 19784 17376 19792 17440
rect 19472 16352 19792 17376
rect 19472 16288 19480 16352
rect 19544 16288 19560 16352
rect 19624 16288 19640 16352
rect 19704 16288 19720 16352
rect 19784 16288 19792 16352
rect 18643 16148 18709 16149
rect 18643 16084 18644 16148
rect 18708 16084 18709 16148
rect 18643 16083 18709 16084
rect 14840 15744 14848 15808
rect 14912 15744 14928 15808
rect 14992 15744 15008 15808
rect 15072 15744 15088 15808
rect 15152 15744 15160 15808
rect 14840 14720 15160 15744
rect 14840 14656 14848 14720
rect 14912 14656 14928 14720
rect 14992 14656 15008 14720
rect 15072 14656 15088 14720
rect 15152 14656 15160 14720
rect 14840 13632 15160 14656
rect 14840 13568 14848 13632
rect 14912 13568 14928 13632
rect 14992 13568 15008 13632
rect 15072 13568 15088 13632
rect 15152 13568 15160 13632
rect 14840 12544 15160 13568
rect 14840 12480 14848 12544
rect 14912 12480 14928 12544
rect 14992 12480 15008 12544
rect 15072 12480 15088 12544
rect 15152 12480 15160 12544
rect 14840 11456 15160 12480
rect 14840 11392 14848 11456
rect 14912 11392 14928 11456
rect 14992 11392 15008 11456
rect 15072 11392 15088 11456
rect 15152 11392 15160 11456
rect 14840 10368 15160 11392
rect 14840 10304 14848 10368
rect 14912 10304 14928 10368
rect 14992 10304 15008 10368
rect 15072 10304 15088 10368
rect 15152 10304 15160 10368
rect 14840 9280 15160 10304
rect 14840 9216 14848 9280
rect 14912 9216 14928 9280
rect 14992 9216 15008 9280
rect 15072 9216 15088 9280
rect 15152 9216 15160 9280
rect 14840 8192 15160 9216
rect 14840 8128 14848 8192
rect 14912 8128 14928 8192
rect 14992 8128 15008 8192
rect 15072 8128 15088 8192
rect 15152 8128 15160 8192
rect 14840 7104 15160 8128
rect 14840 7040 14848 7104
rect 14912 7040 14928 7104
rect 14992 7040 15008 7104
rect 15072 7040 15088 7104
rect 15152 7040 15160 7104
rect 14840 6016 15160 7040
rect 14840 5952 14848 6016
rect 14912 5952 14928 6016
rect 14992 5952 15008 6016
rect 15072 5952 15088 6016
rect 15152 5952 15160 6016
rect 14840 4928 15160 5952
rect 14840 4864 14848 4928
rect 14912 4864 14928 4928
rect 14992 4864 15008 4928
rect 15072 4864 15088 4928
rect 15152 4864 15160 4928
rect 14840 3840 15160 4864
rect 14840 3776 14848 3840
rect 14912 3776 14928 3840
rect 14992 3776 15008 3840
rect 15072 3776 15088 3840
rect 15152 3776 15160 3840
rect 14840 2752 15160 3776
rect 14840 2688 14848 2752
rect 14912 2688 14928 2752
rect 14992 2688 15008 2752
rect 15072 2688 15088 2752
rect 15152 2688 15160 2752
rect 14840 2128 15160 2688
rect 19472 15264 19792 16288
rect 19472 15200 19480 15264
rect 19544 15200 19560 15264
rect 19624 15200 19640 15264
rect 19704 15200 19720 15264
rect 19784 15200 19792 15264
rect 19472 14176 19792 15200
rect 19472 14112 19480 14176
rect 19544 14112 19560 14176
rect 19624 14112 19640 14176
rect 19704 14112 19720 14176
rect 19784 14112 19792 14176
rect 19472 13088 19792 14112
rect 19472 13024 19480 13088
rect 19544 13024 19560 13088
rect 19624 13024 19640 13088
rect 19704 13024 19720 13088
rect 19784 13024 19792 13088
rect 19472 12000 19792 13024
rect 19472 11936 19480 12000
rect 19544 11936 19560 12000
rect 19624 11936 19640 12000
rect 19704 11936 19720 12000
rect 19784 11936 19792 12000
rect 19472 10912 19792 11936
rect 19472 10848 19480 10912
rect 19544 10848 19560 10912
rect 19624 10848 19640 10912
rect 19704 10848 19720 10912
rect 19784 10848 19792 10912
rect 19472 9824 19792 10848
rect 19472 9760 19480 9824
rect 19544 9760 19560 9824
rect 19624 9760 19640 9824
rect 19704 9760 19720 9824
rect 19784 9760 19792 9824
rect 19472 8736 19792 9760
rect 19472 8672 19480 8736
rect 19544 8672 19560 8736
rect 19624 8672 19640 8736
rect 19704 8672 19720 8736
rect 19784 8672 19792 8736
rect 19472 7648 19792 8672
rect 19472 7584 19480 7648
rect 19544 7584 19560 7648
rect 19624 7584 19640 7648
rect 19704 7584 19720 7648
rect 19784 7584 19792 7648
rect 19472 6560 19792 7584
rect 19472 6496 19480 6560
rect 19544 6496 19560 6560
rect 19624 6496 19640 6560
rect 19704 6496 19720 6560
rect 19784 6496 19792 6560
rect 19472 5472 19792 6496
rect 19472 5408 19480 5472
rect 19544 5408 19560 5472
rect 19624 5408 19640 5472
rect 19704 5408 19720 5472
rect 19784 5408 19792 5472
rect 19472 4384 19792 5408
rect 19472 4320 19480 4384
rect 19544 4320 19560 4384
rect 19624 4320 19640 4384
rect 19704 4320 19720 4384
rect 19784 4320 19792 4384
rect 19472 3296 19792 4320
rect 19472 3232 19480 3296
rect 19544 3232 19560 3296
rect 19624 3232 19640 3296
rect 19704 3232 19720 3296
rect 19784 3232 19792 3296
rect 19472 2208 19792 3232
rect 19472 2144 19480 2208
rect 19544 2144 19560 2208
rect 19624 2144 19640 2208
rect 19704 2144 19720 2208
rect 19784 2144 19792 2208
rect 19472 2128 19792 2144
rect 24104 19072 24424 20096
rect 24104 19008 24112 19072
rect 24176 19008 24192 19072
rect 24256 19008 24272 19072
rect 24336 19008 24352 19072
rect 24416 19008 24424 19072
rect 24104 17984 24424 19008
rect 24104 17920 24112 17984
rect 24176 17920 24192 17984
rect 24256 17920 24272 17984
rect 24336 17920 24352 17984
rect 24416 17920 24424 17984
rect 24104 16896 24424 17920
rect 24104 16832 24112 16896
rect 24176 16832 24192 16896
rect 24256 16832 24272 16896
rect 24336 16832 24352 16896
rect 24416 16832 24424 16896
rect 24104 15808 24424 16832
rect 26190 16557 26250 27643
rect 26371 23492 26437 23493
rect 26371 23428 26372 23492
rect 26436 23428 26437 23492
rect 26371 23427 26437 23428
rect 26374 17645 26434 23427
rect 26558 17781 26618 30363
rect 26555 17780 26621 17781
rect 26555 17716 26556 17780
rect 26620 17716 26621 17780
rect 26555 17715 26621 17716
rect 26371 17644 26437 17645
rect 26371 17580 26372 17644
rect 26436 17580 26437 17644
rect 26371 17579 26437 17580
rect 26187 16556 26253 16557
rect 26187 16492 26188 16556
rect 26252 16492 26253 16556
rect 26187 16491 26253 16492
rect 24104 15744 24112 15808
rect 24176 15744 24192 15808
rect 24256 15744 24272 15808
rect 24336 15744 24352 15808
rect 24416 15744 24424 15808
rect 24104 14720 24424 15744
rect 24104 14656 24112 14720
rect 24176 14656 24192 14720
rect 24256 14656 24272 14720
rect 24336 14656 24352 14720
rect 24416 14656 24424 14720
rect 24104 13632 24424 14656
rect 24104 13568 24112 13632
rect 24176 13568 24192 13632
rect 24256 13568 24272 13632
rect 24336 13568 24352 13632
rect 24416 13568 24424 13632
rect 24104 12544 24424 13568
rect 24104 12480 24112 12544
rect 24176 12480 24192 12544
rect 24256 12480 24272 12544
rect 24336 12480 24352 12544
rect 24416 12480 24424 12544
rect 24104 11456 24424 12480
rect 24104 11392 24112 11456
rect 24176 11392 24192 11456
rect 24256 11392 24272 11456
rect 24336 11392 24352 11456
rect 24416 11392 24424 11456
rect 24104 10368 24424 11392
rect 24104 10304 24112 10368
rect 24176 10304 24192 10368
rect 24256 10304 24272 10368
rect 24336 10304 24352 10368
rect 24416 10304 24424 10368
rect 24104 9280 24424 10304
rect 24104 9216 24112 9280
rect 24176 9216 24192 9280
rect 24256 9216 24272 9280
rect 24336 9216 24352 9280
rect 24416 9216 24424 9280
rect 24104 8192 24424 9216
rect 24104 8128 24112 8192
rect 24176 8128 24192 8192
rect 24256 8128 24272 8192
rect 24336 8128 24352 8192
rect 24416 8128 24424 8192
rect 24104 7104 24424 8128
rect 24104 7040 24112 7104
rect 24176 7040 24192 7104
rect 24256 7040 24272 7104
rect 24336 7040 24352 7104
rect 24416 7040 24424 7104
rect 24104 6016 24424 7040
rect 24104 5952 24112 6016
rect 24176 5952 24192 6016
rect 24256 5952 24272 6016
rect 24336 5952 24352 6016
rect 24416 5952 24424 6016
rect 24104 4928 24424 5952
rect 24104 4864 24112 4928
rect 24176 4864 24192 4928
rect 24256 4864 24272 4928
rect 24336 4864 24352 4928
rect 24416 4864 24424 4928
rect 24104 3840 24424 4864
rect 24104 3776 24112 3840
rect 24176 3776 24192 3840
rect 24256 3776 24272 3840
rect 24336 3776 24352 3840
rect 24416 3776 24424 3840
rect 24104 2752 24424 3776
rect 24104 2688 24112 2752
rect 24176 2688 24192 2752
rect 24256 2688 24272 2752
rect 24336 2688 24352 2752
rect 24416 2688 24424 2752
rect 24104 2128 24424 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 7360 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1644511149
transform -1 0 7728 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1644511149
transform 1 0 26036 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1644511149
transform -1 0 9844 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1644511149
transform 1 0 11500 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1644511149
transform -1 0 28152 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1644511149
transform 1 0 5244 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1644511149
transform 1 0 19872 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1644511149
transform 1 0 23092 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52
timestamp 1644511149
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8280 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_107
timestamp 1644511149
transform 1 0 10948 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1644511149
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_113
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_120 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12144 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_132 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 13248 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_141 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_147
timestamp 1644511149
transform 1 0 14628 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_162
timestamp 1644511149
transform 1 0 16008 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_169
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_177
timestamp 1644511149
transform 1 0 17388 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_184
timestamp 1644511149
transform 1 0 18032 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_218
timestamp 1644511149
transform 1 0 21160 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1644511149
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_248
timestamp 1644511149
transform 1 0 23920 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_276
timestamp 1644511149
transform 1 0 26496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_284
timestamp 1644511149
transform 1 0 27232 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_293
timestamp 1644511149
transform 1 0 28060 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_1_3
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_9
timestamp 1644511149
transform 1 0 1932 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_34
timestamp 1644511149
transform 1 0 4232 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_41
timestamp 1644511149
transform 1 0 4876 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_45
timestamp 1644511149
transform 1 0 5244 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_49
timestamp 1644511149
transform 1 0 5612 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1644511149
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_57
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_84
timestamp 1644511149
transform 1 0 8832 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_92
timestamp 1644511149
transform 1 0 9568 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_96
timestamp 1644511149
transform 1 0 9936 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_108
timestamp 1644511149
transform 1 0 11040 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_136
timestamp 1644511149
transform 1 0 13616 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_163
timestamp 1644511149
transform 1 0 16100 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1644511149
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_169
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_177
timestamp 1644511149
transform 1 0 17388 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_182
timestamp 1644511149
transform 1 0 17848 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_189
timestamp 1644511149
transform 1 0 18492 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_214
timestamp 1644511149
transform 1 0 20792 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1644511149
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_225
timestamp 1644511149
transform 1 0 21804 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_247
timestamp 1644511149
transform 1 0 23828 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_276
timestamp 1644511149
transform 1 0 26496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_284
timestamp 1644511149
transform 1 0 27232 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_291
timestamp 1644511149
transform 1 0 27876 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_24
timestamp 1644511149
transform 1 0 3312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_32
timestamp 1644511149
transform 1 0 4048 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_38
timestamp 1644511149
transform 1 0 4600 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_42
timestamp 1644511149
transform 1 0 4968 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_67
timestamp 1644511149
transform 1 0 7268 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_74
timestamp 1644511149
transform 1 0 7912 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1644511149
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_85
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_108
timestamp 1644511149
transform 1 0 11040 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_114
timestamp 1644511149
transform 1 0 11592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_118
timestamp 1644511149
transform 1 0 11960 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_125
timestamp 1644511149
transform 1 0 12604 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_132
timestamp 1644511149
transform 1 0 13248 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_146
timestamp 1644511149
transform 1 0 14536 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_179
timestamp 1644511149
transform 1 0 17572 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_187
timestamp 1644511149
transform 1 0 18308 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_192
timestamp 1644511149
transform 1 0 18768 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_201
timestamp 1644511149
transform 1 0 19596 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_208
timestamp 1644511149
transform 1 0 20240 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_215
timestamp 1644511149
transform 1 0 20884 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_224
timestamp 1644511149
transform 1 0 21712 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_231
timestamp 1644511149
transform 1 0 22356 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_237
timestamp 1644511149
transform 1 0 22908 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_241
timestamp 1644511149
transform 1 0 23276 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_248
timestamp 1644511149
transform 1 0 23920 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_253
timestamp 1644511149
transform 1 0 24380 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_257
timestamp 1644511149
transform 1 0 24748 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_282
timestamp 1644511149
transform 1 0 27048 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_2_293
timestamp 1644511149
transform 1 0 28060 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_24
timestamp 1644511149
transform 1 0 3312 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_49
timestamp 1644511149
transform 1 0 5612 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1644511149
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_62
timestamp 1644511149
transform 1 0 6808 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_87
timestamp 1644511149
transform 1 0 9108 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_94
timestamp 1644511149
transform 1 0 9752 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_101
timestamp 1644511149
transform 1 0 10396 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_109
timestamp 1644511149
transform 1 0 11132 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_113
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_125
timestamp 1644511149
transform 1 0 12604 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_150
timestamp 1644511149
transform 1 0 14904 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1644511149
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1644511149
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_169
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_177
timestamp 1644511149
transform 1 0 17388 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_199
timestamp 1644511149
transform 1 0 19412 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_211
timestamp 1644511149
transform 1 0 20516 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1644511149
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_225
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_233
timestamp 1644511149
transform 1 0 22540 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_239
timestamp 1644511149
transform 1 0 23092 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_264
timestamp 1644511149
transform 1 0 25392 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_271
timestamp 1644511149
transform 1 0 26036 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1644511149
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_281
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_291
timestamp 1644511149
transform 1 0 27876 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_10
timestamp 1644511149
transform 1 0 2024 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_17
timestamp 1644511149
transform 1 0 2668 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_24
timestamp 1644511149
transform 1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_50
timestamp 1644511149
transform 1 0 5704 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_57
timestamp 1644511149
transform 1 0 6348 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_65
timestamp 1644511149
transform 1 0 7084 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_70
timestamp 1644511149
transform 1 0 7544 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1644511149
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1644511149
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_85
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_89
timestamp 1644511149
transform 1 0 9292 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_101
timestamp 1644511149
transform 1 0 10396 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_113
timestamp 1644511149
transform 1 0 11500 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_125
timestamp 1644511149
transform 1 0 12604 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_137
timestamp 1644511149
transform 1 0 13708 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_153
timestamp 1644511149
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_165
timestamp 1644511149
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_177
timestamp 1644511149
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1644511149
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1644511149
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_197
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_209
timestamp 1644511149
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_221
timestamp 1644511149
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_233
timestamp 1644511149
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_248
timestamp 1644511149
transform 1 0 23920 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_253
timestamp 1644511149
transform 1 0 24380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_263
timestamp 1644511149
transform 1 0 25300 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_270
timestamp 1644511149
transform 1 0 25944 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_295
timestamp 1644511149
transform 1 0 28244 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_6
timestamp 1644511149
transform 1 0 1656 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_31
timestamp 1644511149
transform 1 0 3956 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_38
timestamp 1644511149
transform 1 0 4600 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_45
timestamp 1644511149
transform 1 0 5244 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_52
timestamp 1644511149
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_60
timestamp 1644511149
transform 1 0 6624 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_67
timestamp 1644511149
transform 1 0 7268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_79
timestamp 1644511149
transform 1 0 8372 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_91
timestamp 1644511149
transform 1 0 9476 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_103
timestamp 1644511149
transform 1 0 10580 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1644511149
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_113
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_125
timestamp 1644511149
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_137
timestamp 1644511149
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_149
timestamp 1644511149
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1644511149
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1644511149
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_169
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_181
timestamp 1644511149
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_193
timestamp 1644511149
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_205
timestamp 1644511149
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1644511149
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1644511149
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_225
timestamp 1644511149
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_237
timestamp 1644511149
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_249
timestamp 1644511149
transform 1 0 24012 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_276
timestamp 1644511149
transform 1 0 26496 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_281
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_286
timestamp 1644511149
transform 1 0 27416 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_293
timestamp 1644511149
transform 1 0 28060 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp 1644511149
transform 1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_32
timestamp 1644511149
transform 1 0 4048 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_39
timestamp 1644511149
transform 1 0 4692 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_46
timestamp 1644511149
transform 1 0 5336 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_53
timestamp 1644511149
transform 1 0 5980 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_60
timestamp 1644511149
transform 1 0 6624 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_67
timestamp 1644511149
transform 1 0 7268 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_79
timestamp 1644511149
transform 1 0 8372 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1644511149
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_97
timestamp 1644511149
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_109
timestamp 1644511149
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_121
timestamp 1644511149
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1644511149
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1644511149
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_153
timestamp 1644511149
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_165
timestamp 1644511149
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_177
timestamp 1644511149
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1644511149
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1644511149
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_197
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_209
timestamp 1644511149
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_221
timestamp 1644511149
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_233
timestamp 1644511149
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1644511149
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1644511149
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_253
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_259
timestamp 1644511149
transform 1 0 24932 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_263
timestamp 1644511149
transform 1 0 25300 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_270
timestamp 1644511149
transform 1 0 25944 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_295
timestamp 1644511149
transform 1 0 28244 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_11
timestamp 1644511149
transform 1 0 2116 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_18
timestamp 1644511149
transform 1 0 2760 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_24
timestamp 1644511149
transform 1 0 3312 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_46
timestamp 1644511149
transform 1 0 5336 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1644511149
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1644511149
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_81
timestamp 1644511149
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1644511149
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1644511149
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1644511149
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_113
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_125
timestamp 1644511149
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_137
timestamp 1644511149
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_149
timestamp 1644511149
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1644511149
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1644511149
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_169
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_181
timestamp 1644511149
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_193
timestamp 1644511149
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_205
timestamp 1644511149
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1644511149
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1644511149
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_225
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_237
timestamp 1644511149
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_249
timestamp 1644511149
transform 1 0 24012 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_276
timestamp 1644511149
transform 1 0 26496 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_281
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_286
timestamp 1644511149
transform 1 0 27416 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_293
timestamp 1644511149
transform 1 0 28060 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_24
timestamp 1644511149
transform 1 0 3312 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_32
timestamp 1644511149
transform 1 0 4048 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_39
timestamp 1644511149
transform 1 0 4692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_51
timestamp 1644511149
transform 1 0 5796 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_63
timestamp 1644511149
transform 1 0 6900 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_75
timestamp 1644511149
transform 1 0 8004 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1644511149
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_97
timestamp 1644511149
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_109
timestamp 1644511149
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_121
timestamp 1644511149
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1644511149
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1644511149
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_153
timestamp 1644511149
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_165
timestamp 1644511149
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_177
timestamp 1644511149
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1644511149
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1644511149
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_197
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_209
timestamp 1644511149
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_221
timestamp 1644511149
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_233
timestamp 1644511149
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1644511149
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1644511149
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_253
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_265
timestamp 1644511149
transform 1 0 25484 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_273
timestamp 1644511149
transform 1 0 26220 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_295
timestamp 1644511149
transform 1 0 28244 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_30
timestamp 1644511149
transform 1 0 3864 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_37
timestamp 1644511149
transform 1 0 4508 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_49
timestamp 1644511149
transform 1 0 5612 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1644511149
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_69
timestamp 1644511149
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_81
timestamp 1644511149
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_93
timestamp 1644511149
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1644511149
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1644511149
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_113
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_125
timestamp 1644511149
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_137
timestamp 1644511149
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_149
timestamp 1644511149
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1644511149
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1644511149
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_181
timestamp 1644511149
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_193
timestamp 1644511149
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_205
timestamp 1644511149
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1644511149
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1644511149
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_225
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_237
timestamp 1644511149
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_249
timestamp 1644511149
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_261
timestamp 1644511149
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1644511149
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1644511149
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_281
timestamp 1644511149
transform 1 0 26956 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_285
timestamp 1644511149
transform 1 0 27324 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_292
timestamp 1644511149
transform 1 0 27968 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_298
timestamp 1644511149
transform 1 0 28520 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_24
timestamp 1644511149
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1644511149
transform 1 0 4048 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_44
timestamp 1644511149
transform 1 0 5152 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_56
timestamp 1644511149
transform 1 0 6256 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_68
timestamp 1644511149
transform 1 0 7360 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_80
timestamp 1644511149
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_97
timestamp 1644511149
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_109
timestamp 1644511149
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_121
timestamp 1644511149
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1644511149
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1644511149
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_153
timestamp 1644511149
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_165
timestamp 1644511149
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_177
timestamp 1644511149
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1644511149
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1644511149
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_197
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_209
timestamp 1644511149
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_221
timestamp 1644511149
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_233
timestamp 1644511149
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1644511149
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1644511149
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_253
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_265
timestamp 1644511149
transform 1 0 25484 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_273
timestamp 1644511149
transform 1 0 26220 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_295
timestamp 1644511149
transform 1 0 28244 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_7
timestamp 1644511149
transform 1 0 1748 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_11
timestamp 1644511149
transform 1 0 2116 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_18
timestamp 1644511149
transform 1 0 2760 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_25
timestamp 1644511149
transform 1 0 3404 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_37
timestamp 1644511149
transform 1 0 4508 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_49
timestamp 1644511149
transform 1 0 5612 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1644511149
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_69
timestamp 1644511149
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_81
timestamp 1644511149
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_93
timestamp 1644511149
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1644511149
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1644511149
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_113
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_125
timestamp 1644511149
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_137
timestamp 1644511149
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_149
timestamp 1644511149
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1644511149
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1644511149
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_169
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_181
timestamp 1644511149
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_193
timestamp 1644511149
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_205
timestamp 1644511149
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1644511149
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1644511149
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_225
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_237
timestamp 1644511149
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_249
timestamp 1644511149
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_261
timestamp 1644511149
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1644511149
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1644511149
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_281
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_285
timestamp 1644511149
transform 1 0 27324 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_292
timestamp 1644511149
transform 1 0 27968 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_298
timestamp 1644511149
transform 1 0 28520 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_24
timestamp 1644511149
transform 1 0 3312 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_41
timestamp 1644511149
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_53
timestamp 1644511149
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_65
timestamp 1644511149
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1644511149
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1644511149
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_85
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_97
timestamp 1644511149
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_109
timestamp 1644511149
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_121
timestamp 1644511149
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1644511149
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1644511149
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_153
timestamp 1644511149
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_165
timestamp 1644511149
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_177
timestamp 1644511149
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1644511149
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1644511149
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_197
timestamp 1644511149
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_209
timestamp 1644511149
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_221
timestamp 1644511149
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_233
timestamp 1644511149
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1644511149
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1644511149
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_253
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_265
timestamp 1644511149
transform 1 0 25484 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_273
timestamp 1644511149
transform 1 0 26220 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_295
timestamp 1644511149
transform 1 0 28244 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_8
timestamp 1644511149
transform 1 0 1840 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1644511149
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1644511149
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1644511149
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1644511149
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1644511149
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_69
timestamp 1644511149
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_81
timestamp 1644511149
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_93
timestamp 1644511149
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1644511149
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1644511149
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_113
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_125
timestamp 1644511149
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_137
timestamp 1644511149
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_149
timestamp 1644511149
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1644511149
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1644511149
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_169
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_181
timestamp 1644511149
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_193
timestamp 1644511149
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_205
timestamp 1644511149
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1644511149
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1644511149
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_225
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_237
timestamp 1644511149
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_249
timestamp 1644511149
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_261
timestamp 1644511149
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1644511149
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1644511149
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_281
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_285
timestamp 1644511149
transform 1 0 27324 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_292
timestamp 1644511149
transform 1 0 27968 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_298
timestamp 1644511149
transform 1 0 28520 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_3
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_7
timestamp 1644511149
transform 1 0 1748 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_11
timestamp 1644511149
transform 1 0 2116 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_23
timestamp 1644511149
transform 1 0 3220 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1644511149
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_53
timestamp 1644511149
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_65
timestamp 1644511149
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1644511149
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1644511149
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_97
timestamp 1644511149
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_109
timestamp 1644511149
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_121
timestamp 1644511149
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1644511149
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1644511149
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_153
timestamp 1644511149
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_165
timestamp 1644511149
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_177
timestamp 1644511149
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1644511149
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1644511149
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_197
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_209
timestamp 1644511149
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_221
timestamp 1644511149
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_233
timestamp 1644511149
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1644511149
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1644511149
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_253
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_265
timestamp 1644511149
transform 1 0 25484 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_273
timestamp 1644511149
transform 1 0 26220 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_295
timestamp 1644511149
transform 1 0 28244 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_3
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_25
timestamp 1644511149
transform 1 0 3404 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_37
timestamp 1644511149
transform 1 0 4508 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_49
timestamp 1644511149
transform 1 0 5612 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1644511149
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1644511149
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_81
timestamp 1644511149
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_93
timestamp 1644511149
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1644511149
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1644511149
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_113
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_125
timestamp 1644511149
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_137
timestamp 1644511149
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_149
timestamp 1644511149
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1644511149
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1644511149
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_169
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_181
timestamp 1644511149
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_193
timestamp 1644511149
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_205
timestamp 1644511149
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1644511149
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1644511149
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_225
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_237
timestamp 1644511149
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_249
timestamp 1644511149
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_261
timestamp 1644511149
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1644511149
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1644511149
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_281
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_286
timestamp 1644511149
transform 1 0 27416 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_293
timestamp 1644511149
transform 1 0 28060 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_24
timestamp 1644511149
transform 1 0 3312 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1644511149
transform 1 0 4048 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_44
timestamp 1644511149
transform 1 0 5152 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_56
timestamp 1644511149
transform 1 0 6256 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_68
timestamp 1644511149
transform 1 0 7360 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_80
timestamp 1644511149
transform 1 0 8464 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_85
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_97
timestamp 1644511149
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_109
timestamp 1644511149
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_121
timestamp 1644511149
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1644511149
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1644511149
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_141
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_153
timestamp 1644511149
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_165
timestamp 1644511149
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_177
timestamp 1644511149
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1644511149
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1644511149
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_197
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_209
timestamp 1644511149
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_221
timestamp 1644511149
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_233
timestamp 1644511149
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1644511149
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1644511149
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_253
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_265
timestamp 1644511149
transform 1 0 25484 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_273
timestamp 1644511149
transform 1 0 26220 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_295
timestamp 1644511149
transform 1 0 28244 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_3
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_10
timestamp 1644511149
transform 1 0 2024 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_17
timestamp 1644511149
transform 1 0 2668 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_24
timestamp 1644511149
transform 1 0 3312 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_36
timestamp 1644511149
transform 1 0 4416 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_48
timestamp 1644511149
transform 1 0 5520 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_69
timestamp 1644511149
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_81
timestamp 1644511149
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_93
timestamp 1644511149
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1644511149
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1644511149
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_113
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_125
timestamp 1644511149
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_137
timestamp 1644511149
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_149
timestamp 1644511149
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1644511149
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1644511149
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_169
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_181
timestamp 1644511149
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_193
timestamp 1644511149
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_205
timestamp 1644511149
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1644511149
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1644511149
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_225
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_237
timestamp 1644511149
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_249
timestamp 1644511149
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_261
timestamp 1644511149
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1644511149
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1644511149
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_281
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_287
timestamp 1644511149
transform 1 0 27508 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_295
timestamp 1644511149
transform 1 0 28244 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_24
timestamp 1644511149
transform 1 0 3312 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1644511149
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_53
timestamp 1644511149
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_65
timestamp 1644511149
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1644511149
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1644511149
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_85
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_97
timestamp 1644511149
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_109
timestamp 1644511149
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_121
timestamp 1644511149
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1644511149
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1644511149
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_153
timestamp 1644511149
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_165
timestamp 1644511149
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_177
timestamp 1644511149
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1644511149
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1644511149
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_197
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_209
timestamp 1644511149
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_221
timestamp 1644511149
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_233
timestamp 1644511149
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1644511149
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1644511149
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_253
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_265
timestamp 1644511149
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_277
timestamp 1644511149
transform 1 0 26588 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_283
timestamp 1644511149
transform 1 0 27140 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_287
timestamp 1644511149
transform 1 0 27508 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_294
timestamp 1644511149
transform 1 0 28152 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_298
timestamp 1644511149
transform 1 0 28520 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_24
timestamp 1644511149
transform 1 0 3312 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_36
timestamp 1644511149
transform 1 0 4416 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_48
timestamp 1644511149
transform 1 0 5520 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 1644511149
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_81
timestamp 1644511149
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_93
timestamp 1644511149
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1644511149
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1644511149
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_113
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_125
timestamp 1644511149
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_137
timestamp 1644511149
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_149
timestamp 1644511149
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1644511149
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1644511149
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_169
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_181
timestamp 1644511149
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_193
timestamp 1644511149
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_205
timestamp 1644511149
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1644511149
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1644511149
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_225
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_237
timestamp 1644511149
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_249
timestamp 1644511149
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_261
timestamp 1644511149
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_276
timestamp 1644511149
transform 1 0 26496 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_281
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_287
timestamp 1644511149
transform 1 0 27508 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_294
timestamp 1644511149
transform 1 0 28152 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_298
timestamp 1644511149
transform 1 0 28520 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_8
timestamp 1644511149
transform 1 0 1840 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_15
timestamp 1644511149
transform 1 0 2484 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_22
timestamp 1644511149
transform 1 0 3128 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1644511149
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 1644511149
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1644511149
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1644511149
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1644511149
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_97
timestamp 1644511149
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_109
timestamp 1644511149
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_121
timestamp 1644511149
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1644511149
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1644511149
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_153
timestamp 1644511149
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_165
timestamp 1644511149
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_177
timestamp 1644511149
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1644511149
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1644511149
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_197
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_209
timestamp 1644511149
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_221
timestamp 1644511149
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_233
timestamp 1644511149
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1644511149
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1644511149
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_253
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_261
timestamp 1644511149
transform 1 0 25116 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_267
timestamp 1644511149
transform 1 0 25668 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_274
timestamp 1644511149
transform 1 0 26312 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_282
timestamp 1644511149
transform 1 0 27048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_286
timestamp 1644511149
transform 1 0 27416 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_293
timestamp 1644511149
transform 1 0 28060 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_3
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_10
timestamp 1644511149
transform 1 0 2024 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_22
timestamp 1644511149
transform 1 0 3128 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_34
timestamp 1644511149
transform 1 0 4232 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_46
timestamp 1644511149
transform 1 0 5336 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1644511149
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_81
timestamp 1644511149
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_93
timestamp 1644511149
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1644511149
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1644511149
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_113
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_125
timestamp 1644511149
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_137
timestamp 1644511149
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_149
timestamp 1644511149
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1644511149
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1644511149
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_169
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_181
timestamp 1644511149
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_193
timestamp 1644511149
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_205
timestamp 1644511149
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1644511149
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1644511149
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_225
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_237
timestamp 1644511149
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_249
timestamp 1644511149
transform 1 0 24012 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_257
timestamp 1644511149
transform 1 0 24748 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_263
timestamp 1644511149
transform 1 0 25300 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_270
timestamp 1644511149
transform 1 0 25944 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_278
timestamp 1644511149
transform 1 0 26680 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_281
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_285
timestamp 1644511149
transform 1 0 27324 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_292
timestamp 1644511149
transform 1 0 27968 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_298
timestamp 1644511149
transform 1 0 28520 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_24
timestamp 1644511149
transform 1 0 3312 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1644511149
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_53
timestamp 1644511149
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_65
timestamp 1644511149
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1644511149
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1644511149
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_85
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_97
timestamp 1644511149
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_109
timestamp 1644511149
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_121
timestamp 1644511149
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1644511149
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1644511149
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_141
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_153
timestamp 1644511149
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_165
timestamp 1644511149
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_177
timestamp 1644511149
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1644511149
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1644511149
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_197
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_209
timestamp 1644511149
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_221
timestamp 1644511149
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_233
timestamp 1644511149
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_248
timestamp 1644511149
transform 1 0 23920 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_253
timestamp 1644511149
transform 1 0 24380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_257
timestamp 1644511149
transform 1 0 24748 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_261
timestamp 1644511149
transform 1 0 25116 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_265
timestamp 1644511149
transform 1 0 25484 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_269
timestamp 1644511149
transform 1 0 25852 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_273
timestamp 1644511149
transform 1 0 26220 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_295
timestamp 1644511149
transform 1 0 28244 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_8
timestamp 1644511149
transform 1 0 1840 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1644511149
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1644511149
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1644511149
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1644511149
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1644511149
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1644511149
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_81
timestamp 1644511149
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_93
timestamp 1644511149
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1644511149
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1644511149
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_113
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_125
timestamp 1644511149
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_137
timestamp 1644511149
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_149
timestamp 1644511149
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1644511149
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1644511149
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_169
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_181
timestamp 1644511149
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_193
timestamp 1644511149
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_205
timestamp 1644511149
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1644511149
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1644511149
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_225
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_237
timestamp 1644511149
transform 1 0 22908 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_248
timestamp 1644511149
transform 1 0 23920 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_255
timestamp 1644511149
transform 1 0 24564 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_262
timestamp 1644511149
transform 1 0 25208 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_269
timestamp 1644511149
transform 1 0 25852 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_276
timestamp 1644511149
transform 1 0 26496 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_281
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_285
timestamp 1644511149
transform 1 0 27324 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_293
timestamp 1644511149
transform 1 0 28060 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_24
timestamp 1644511149
transform 1 0 3312 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1644511149
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_53
timestamp 1644511149
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_65
timestamp 1644511149
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1644511149
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1644511149
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_85
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_97
timestamp 1644511149
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_109
timestamp 1644511149
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_121
timestamp 1644511149
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1644511149
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1644511149
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_153
timestamp 1644511149
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_165
timestamp 1644511149
transform 1 0 16284 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_173
timestamp 1644511149
transform 1 0 17020 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_177
timestamp 1644511149
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1644511149
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1644511149
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_197
timestamp 1644511149
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_209
timestamp 1644511149
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_221
timestamp 1644511149
transform 1 0 21436 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_229
timestamp 1644511149
transform 1 0 22172 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_233
timestamp 1644511149
transform 1 0 22540 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_240
timestamp 1644511149
transform 1 0 23184 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_248
timestamp 1644511149
transform 1 0 23920 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_257
timestamp 1644511149
transform 1 0 24748 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_265
timestamp 1644511149
transform 1 0 25484 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_273
timestamp 1644511149
transform 1 0 26220 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_295
timestamp 1644511149
transform 1 0 28244 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_6
timestamp 1644511149
transform 1 0 1656 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_18
timestamp 1644511149
transform 1 0 2760 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_30
timestamp 1644511149
transform 1 0 3864 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_42
timestamp 1644511149
transform 1 0 4968 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1644511149
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_69
timestamp 1644511149
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_81
timestamp 1644511149
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_93
timestamp 1644511149
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1644511149
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1644511149
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_113
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_125
timestamp 1644511149
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_137
timestamp 1644511149
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_149
timestamp 1644511149
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1644511149
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1644511149
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_175
timestamp 1644511149
transform 1 0 17204 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_183
timestamp 1644511149
transform 1 0 17940 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_189
timestamp 1644511149
transform 1 0 18492 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_201
timestamp 1644511149
transform 1 0 19596 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_205
timestamp 1644511149
transform 1 0 19964 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_209
timestamp 1644511149
transform 1 0 20332 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_213
timestamp 1644511149
transform 1 0 20700 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1644511149
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1644511149
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1644511149
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_230
timestamp 1644511149
transform 1 0 22264 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_237
timestamp 1644511149
transform 1 0 22908 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_245
timestamp 1644511149
transform 1 0 23644 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_253
timestamp 1644511149
transform 1 0 24380 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_276
timestamp 1644511149
transform 1 0 26496 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_281
timestamp 1644511149
transform 1 0 26956 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_289
timestamp 1644511149
transform 1 0 27692 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_297
timestamp 1644511149
transform 1 0 28428 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_3
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_9
timestamp 1644511149
transform 1 0 1932 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_16
timestamp 1644511149
transform 1 0 2576 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1644511149
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_53
timestamp 1644511149
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_65
timestamp 1644511149
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1644511149
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1644511149
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_85
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_97
timestamp 1644511149
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_109
timestamp 1644511149
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_121
timestamp 1644511149
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1644511149
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1644511149
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_153
timestamp 1644511149
transform 1 0 15180 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_161
timestamp 1644511149
transform 1 0 15916 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_165
timestamp 1644511149
transform 1 0 16284 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_185
timestamp 1644511149
transform 1 0 18124 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_192
timestamp 1644511149
transform 1 0 18768 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_197
timestamp 1644511149
transform 1 0 19228 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_201
timestamp 1644511149
transform 1 0 19596 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_206
timestamp 1644511149
transform 1 0 20056 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_213
timestamp 1644511149
transform 1 0 20700 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_224
timestamp 1644511149
transform 1 0 21712 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_232
timestamp 1644511149
transform 1 0 22448 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_240
timestamp 1644511149
transform 1 0 23184 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_247
timestamp 1644511149
transform 1 0 23828 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1644511149
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_253
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_270
timestamp 1644511149
transform 1 0 25944 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_295
timestamp 1644511149
transform 1 0 28244 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_24
timestamp 1644511149
transform 1 0 3312 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_36
timestamp 1644511149
transform 1 0 4416 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_48
timestamp 1644511149
transform 1 0 5520 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_69
timestamp 1644511149
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_81
timestamp 1644511149
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_93
timestamp 1644511149
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1644511149
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1644511149
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_113
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_125
timestamp 1644511149
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_137
timestamp 1644511149
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_149
timestamp 1644511149
transform 1 0 14812 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_157
timestamp 1644511149
transform 1 0 15548 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_164
timestamp 1644511149
transform 1 0 16192 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_179
timestamp 1644511149
transform 1 0 17572 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_199
timestamp 1644511149
transform 1 0 19412 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_219
timestamp 1644511149
transform 1 0 21252 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1644511149
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_241
timestamp 1644511149
transform 1 0 23276 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_261
timestamp 1644511149
transform 1 0 25116 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_270
timestamp 1644511149
transform 1 0 25944 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_278
timestamp 1644511149
transform 1 0 26680 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_286
timestamp 1644511149
transform 1 0 27416 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_294
timestamp 1644511149
transform 1 0 28152 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_298
timestamp 1644511149
transform 1 0 28520 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_24
timestamp 1644511149
transform 1 0 3312 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_41
timestamp 1644511149
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_53
timestamp 1644511149
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_65
timestamp 1644511149
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1644511149
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1644511149
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_85
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_97
timestamp 1644511149
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_109
timestamp 1644511149
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_121
timestamp 1644511149
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1644511149
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1644511149
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_141
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_156
timestamp 1644511149
transform 1 0 15456 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_176
timestamp 1644511149
transform 1 0 17296 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_190
timestamp 1644511149
transform 1 0 18584 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_202
timestamp 1644511149
transform 1 0 19688 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_211
timestamp 1644511149
transform 1 0 20516 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_215
timestamp 1644511149
transform 1 0 20884 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_232
timestamp 1644511149
transform 1 0 22448 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_240
timestamp 1644511149
transform 1 0 23184 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_248
timestamp 1644511149
transform 1 0 23920 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_269
timestamp 1644511149
transform 1 0 25852 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_273
timestamp 1644511149
transform 1 0 26220 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_295
timestamp 1644511149
transform 1 0 28244 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_3
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_9
timestamp 1644511149
transform 1 0 1932 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_16
timestamp 1644511149
transform 1 0 2576 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_28
timestamp 1644511149
transform 1 0 3680 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_40
timestamp 1644511149
transform 1 0 4784 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_52
timestamp 1644511149
transform 1 0 5888 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_69
timestamp 1644511149
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_81
timestamp 1644511149
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_93
timestamp 1644511149
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1644511149
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1644511149
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_113
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_125
timestamp 1644511149
transform 1 0 12604 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_133
timestamp 1644511149
transform 1 0 13340 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_139
timestamp 1644511149
transform 1 0 13892 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_159
timestamp 1644511149
transform 1 0 15732 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1644511149
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_172
timestamp 1644511149
transform 1 0 16928 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_185
timestamp 1644511149
transform 1 0 18124 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_197
timestamp 1644511149
transform 1 0 19228 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_219
timestamp 1644511149
transform 1 0 21252 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1644511149
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_231
timestamp 1644511149
transform 1 0 22356 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_240
timestamp 1644511149
transform 1 0 23184 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_248
timestamp 1644511149
transform 1 0 23920 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_256
timestamp 1644511149
transform 1 0 24656 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_276
timestamp 1644511149
transform 1 0 26496 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_287
timestamp 1644511149
transform 1 0 27508 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_295
timestamp 1644511149
transform 1 0 28244 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1644511149
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1644511149
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1644511149
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_53
timestamp 1644511149
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_65
timestamp 1644511149
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1644511149
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1644511149
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_97
timestamp 1644511149
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_109
timestamp 1644511149
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_121
timestamp 1644511149
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1644511149
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1644511149
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_141
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_147
timestamp 1644511149
transform 1 0 14628 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_158
timestamp 1644511149
transform 1 0 15640 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_168
timestamp 1644511149
transform 1 0 16560 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_179
timestamp 1644511149
transform 1 0 17572 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_187
timestamp 1644511149
transform 1 0 18308 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1644511149
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_202
timestamp 1644511149
transform 1 0 19688 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_211
timestamp 1644511149
transform 1 0 20516 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_219
timestamp 1644511149
transform 1 0 21252 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_223
timestamp 1644511149
transform 1 0 21620 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_228
timestamp 1644511149
transform 1 0 22080 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_236
timestamp 1644511149
transform 1 0 22816 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_248
timestamp 1644511149
transform 1 0 23920 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_253
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_257
timestamp 1644511149
transform 1 0 24748 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_265
timestamp 1644511149
transform 1 0 25484 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_273
timestamp 1644511149
transform 1 0 26220 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_295
timestamp 1644511149
transform 1 0 28244 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1644511149
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1644511149
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1644511149
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1644511149
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1644511149
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_69
timestamp 1644511149
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_81
timestamp 1644511149
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_93
timestamp 1644511149
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1644511149
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1644511149
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_113
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_125
timestamp 1644511149
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_137
timestamp 1644511149
transform 1 0 13708 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_148
timestamp 1644511149
transform 1 0 14720 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_159
timestamp 1644511149
transform 1 0 15732 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1644511149
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_176
timestamp 1644511149
transform 1 0 17296 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_183
timestamp 1644511149
transform 1 0 17940 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_194
timestamp 1644511149
transform 1 0 18952 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_207
timestamp 1644511149
transform 1 0 20148 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_213
timestamp 1644511149
transform 1 0 20700 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_218
timestamp 1644511149
transform 1 0 21160 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_225
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_229
timestamp 1644511149
transform 1 0 22172 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_240
timestamp 1644511149
transform 1 0 23184 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_251
timestamp 1644511149
transform 1 0 24196 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_259
timestamp 1644511149
transform 1 0 24932 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_276
timestamp 1644511149
transform 1 0 26496 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_287
timestamp 1644511149
transform 1 0 27508 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_295
timestamp 1644511149
transform 1 0 28244 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1644511149
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1644511149
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_41
timestamp 1644511149
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_53
timestamp 1644511149
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_65
timestamp 1644511149
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1644511149
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1644511149
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_85
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_97
timestamp 1644511149
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_109
timestamp 1644511149
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_121
timestamp 1644511149
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_136
timestamp 1644511149
transform 1 0 13616 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_141
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_148
timestamp 1644511149
transform 1 0 14720 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_159
timestamp 1644511149
transform 1 0 15732 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_181
timestamp 1644511149
transform 1 0 17756 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_192
timestamp 1644511149
transform 1 0 18768 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_197
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_215
timestamp 1644511149
transform 1 0 20884 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_235
timestamp 1644511149
transform 1 0 22724 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_246
timestamp 1644511149
transform 1 0 23736 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_269
timestamp 1644511149
transform 1 0 25852 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_273
timestamp 1644511149
transform 1 0 26220 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_295
timestamp 1644511149
transform 1 0 28244 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1644511149
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1644511149
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1644511149
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1644511149
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1644511149
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_57
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_69
timestamp 1644511149
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_81
timestamp 1644511149
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_93
timestamp 1644511149
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1644511149
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1644511149
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_113
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_125
timestamp 1644511149
transform 1 0 12604 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_149
timestamp 1644511149
transform 1 0 14812 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1644511149
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1644511149
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_177
timestamp 1644511149
transform 1 0 17388 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_185
timestamp 1644511149
transform 1 0 18124 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_203
timestamp 1644511149
transform 1 0 19780 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_213
timestamp 1644511149
transform 1 0 20700 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_220
timestamp 1644511149
transform 1 0 21344 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_230
timestamp 1644511149
transform 1 0 22264 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_234
timestamp 1644511149
transform 1 0 22632 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_242
timestamp 1644511149
transform 1 0 23368 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_250
timestamp 1644511149
transform 1 0 24104 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_259
timestamp 1644511149
transform 1 0 24932 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_272
timestamp 1644511149
transform 1 0 26128 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_33_289
timestamp 1644511149
transform 1 0 27692 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_297
timestamp 1644511149
transform 1 0 28428 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1644511149
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1644511149
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_41
timestamp 1644511149
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_53
timestamp 1644511149
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_65
timestamp 1644511149
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1644511149
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1644511149
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_85
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_97
timestamp 1644511149
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_109
timestamp 1644511149
transform 1 0 11132 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_117
timestamp 1644511149
transform 1 0 11868 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_122
timestamp 1644511149
transform 1 0 12328 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_129
timestamp 1644511149
transform 1 0 12972 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_136
timestamp 1644511149
transform 1 0 13616 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_145
timestamp 1644511149
transform 1 0 14444 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_157
timestamp 1644511149
transform 1 0 15548 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_163
timestamp 1644511149
transform 1 0 16100 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_172
timestamp 1644511149
transform 1 0 16928 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_184
timestamp 1644511149
transform 1 0 18032 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_192
timestamp 1644511149
transform 1 0 18768 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_197
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_208
timestamp 1644511149
transform 1 0 20240 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_228
timestamp 1644511149
transform 1 0 22080 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_236
timestamp 1644511149
transform 1 0 22816 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_246
timestamp 1644511149
transform 1 0 23736 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_34_253
timestamp 1644511149
transform 1 0 24380 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_34_266
timestamp 1644511149
transform 1 0 25576 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_295
timestamp 1644511149
transform 1 0 28244 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1644511149
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1644511149
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1644511149
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1644511149
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1644511149
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1644511149
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_57
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_69
timestamp 1644511149
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_81
timestamp 1644511149
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_93
timestamp 1644511149
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1644511149
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1644511149
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_113
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_119
timestamp 1644511149
transform 1 0 12052 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_126
timestamp 1644511149
transform 1 0 12696 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_134
timestamp 1644511149
transform 1 0 13432 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_142
timestamp 1644511149
transform 1 0 14168 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_154
timestamp 1644511149
transform 1 0 15272 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_163
timestamp 1644511149
transform 1 0 16100 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1644511149
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_169
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_179
timestamp 1644511149
transform 1 0 17572 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_190
timestamp 1644511149
transform 1 0 18584 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_200
timestamp 1644511149
transform 1 0 19504 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_208
timestamp 1644511149
transform 1 0 20240 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_214
timestamp 1644511149
transform 1 0 20792 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_222
timestamp 1644511149
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_231
timestamp 1644511149
transform 1 0 22356 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_251
timestamp 1644511149
transform 1 0 24196 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_276
timestamp 1644511149
transform 1 0 26496 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_287
timestamp 1644511149
transform 1 0 27508 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_295
timestamp 1644511149
transform 1 0 28244 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1644511149
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1644511149
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_41
timestamp 1644511149
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_53
timestamp 1644511149
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_65
timestamp 1644511149
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1644511149
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1644511149
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_85
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_97
timestamp 1644511149
transform 1 0 10028 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_105
timestamp 1644511149
transform 1 0 10764 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_111
timestamp 1644511149
transform 1 0 11316 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_115
timestamp 1644511149
transform 1 0 11684 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_120
timestamp 1644511149
transform 1 0 12144 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_128
timestamp 1644511149
transform 1 0 12880 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_136
timestamp 1644511149
transform 1 0 13616 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_141
timestamp 1644511149
transform 1 0 14076 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_149
timestamp 1644511149
transform 1 0 14812 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_158
timestamp 1644511149
transform 1 0 15640 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_166
timestamp 1644511149
transform 1 0 16376 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_175
timestamp 1644511149
transform 1 0 17204 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_179
timestamp 1644511149
transform 1 0 17572 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_186
timestamp 1644511149
transform 1 0 18216 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_194
timestamp 1644511149
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_202
timestamp 1644511149
transform 1 0 19688 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_218
timestamp 1644511149
transform 1 0 21160 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_240
timestamp 1644511149
transform 1 0 23184 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_248
timestamp 1644511149
transform 1 0 23920 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_261
timestamp 1644511149
transform 1 0 25116 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_270
timestamp 1644511149
transform 1 0 25944 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_295
timestamp 1644511149
transform 1 0 28244 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_3
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_11
timestamp 1644511149
transform 1 0 2116 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_17
timestamp 1644511149
transform 1 0 2668 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_29
timestamp 1644511149
transform 1 0 3772 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_41
timestamp 1644511149
transform 1 0 4876 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_53
timestamp 1644511149
transform 1 0 5980 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_57
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_69
timestamp 1644511149
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_81
timestamp 1644511149
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_93
timestamp 1644511149
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_108
timestamp 1644511149
transform 1 0 11040 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_113
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_117
timestamp 1644511149
transform 1 0 11868 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_121
timestamp 1644511149
transform 1 0 12236 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_128
timestamp 1644511149
transform 1 0 12880 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_136
timestamp 1644511149
transform 1 0 13616 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_144
timestamp 1644511149
transform 1 0 14352 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_154
timestamp 1644511149
transform 1 0 15272 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_158
timestamp 1644511149
transform 1 0 15640 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_164
timestamp 1644511149
transform 1 0 16192 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_172
timestamp 1644511149
transform 1 0 16928 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_183
timestamp 1644511149
transform 1 0 17940 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_189
timestamp 1644511149
transform 1 0 18492 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_206
timestamp 1644511149
transform 1 0 20056 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1644511149
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1644511149
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_231
timestamp 1644511149
transform 1 0 22356 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_245
timestamp 1644511149
transform 1 0 23644 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_256
timestamp 1644511149
transform 1 0 24656 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_276
timestamp 1644511149
transform 1 0 26496 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_288
timestamp 1644511149
transform 1 0 27600 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_295
timestamp 1644511149
transform 1 0 28244 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_24
timestamp 1644511149
transform 1 0 3312 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_41
timestamp 1644511149
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_53
timestamp 1644511149
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_65
timestamp 1644511149
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1644511149
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1644511149
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_85
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_97
timestamp 1644511149
transform 1 0 10028 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_103
timestamp 1644511149
transform 1 0 10580 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_107
timestamp 1644511149
transform 1 0 10948 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_114
timestamp 1644511149
transform 1 0 11592 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_121
timestamp 1644511149
transform 1 0 12236 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_128
timestamp 1644511149
transform 1 0 12880 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_136
timestamp 1644511149
transform 1 0 13616 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_157
timestamp 1644511149
transform 1 0 15548 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_171
timestamp 1644511149
transform 1 0 16836 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_182
timestamp 1644511149
transform 1 0 17848 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_192
timestamp 1644511149
transform 1 0 18768 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_201
timestamp 1644511149
transform 1 0 19596 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_221
timestamp 1644511149
transform 1 0 21436 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_225
timestamp 1644511149
transform 1 0 21804 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_232
timestamp 1644511149
transform 1 0 22448 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_240
timestamp 1644511149
transform 1 0 23184 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_248
timestamp 1644511149
transform 1 0 23920 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_257
timestamp 1644511149
transform 1 0 24748 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_269
timestamp 1644511149
transform 1 0 25852 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_273
timestamp 1644511149
transform 1 0 26220 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_295
timestamp 1644511149
transform 1 0 28244 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_3
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_10
timestamp 1644511149
transform 1 0 2024 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_22
timestamp 1644511149
transform 1 0 3128 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_34
timestamp 1644511149
transform 1 0 4232 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_46
timestamp 1644511149
transform 1 0 5336 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 1644511149
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_69
timestamp 1644511149
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_81
timestamp 1644511149
transform 1 0 8556 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_89
timestamp 1644511149
transform 1 0 9292 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_94
timestamp 1644511149
transform 1 0 9752 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_101
timestamp 1644511149
transform 1 0 10396 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_108
timestamp 1644511149
transform 1 0 11040 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_113
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_119
timestamp 1644511149
transform 1 0 12052 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_126
timestamp 1644511149
transform 1 0 12696 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_133
timestamp 1644511149
transform 1 0 13340 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_141
timestamp 1644511149
transform 1 0 14076 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_149
timestamp 1644511149
transform 1 0 14812 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_160
timestamp 1644511149
transform 1 0 15824 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_179
timestamp 1644511149
transform 1 0 17572 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_190
timestamp 1644511149
transform 1 0 18584 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_200
timestamp 1644511149
transform 1 0 19504 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_211
timestamp 1644511149
transform 1 0 20516 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_220
timestamp 1644511149
transform 1 0 21344 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_233
timestamp 1644511149
transform 1 0 22540 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_239
timestamp 1644511149
transform 1 0 23092 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_246
timestamp 1644511149
transform 1 0 23736 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_256
timestamp 1644511149
transform 1 0 24656 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_276
timestamp 1644511149
transform 1 0 26496 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_288
timestamp 1644511149
transform 1 0 27600 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_295
timestamp 1644511149
transform 1 0 28244 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1644511149
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1644511149
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1644511149
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_41
timestamp 1644511149
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_53
timestamp 1644511149
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_65
timestamp 1644511149
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1644511149
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1644511149
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_85
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_100
timestamp 1644511149
transform 1 0 10304 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_107
timestamp 1644511149
transform 1 0 10948 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_114
timestamp 1644511149
transform 1 0 11592 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_121
timestamp 1644511149
transform 1 0 12236 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_128
timestamp 1644511149
transform 1 0 12880 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_136
timestamp 1644511149
transform 1 0 13616 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_141
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_148
timestamp 1644511149
transform 1 0 14720 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_158
timestamp 1644511149
transform 1 0 15640 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_179
timestamp 1644511149
transform 1 0 17572 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_183
timestamp 1644511149
transform 1 0 17940 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_192
timestamp 1644511149
transform 1 0 18768 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_213
timestamp 1644511149
transform 1 0 20700 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_217
timestamp 1644511149
transform 1 0 21068 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_234
timestamp 1644511149
transform 1 0 22632 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1644511149
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1644511149
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_260
timestamp 1644511149
transform 1 0 25024 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_269
timestamp 1644511149
transform 1 0 25852 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_273
timestamp 1644511149
transform 1 0 26220 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_295
timestamp 1644511149
transform 1 0 28244 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1644511149
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1644511149
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1644511149
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1644511149
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1644511149
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_69
timestamp 1644511149
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_81
timestamp 1644511149
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_93
timestamp 1644511149
transform 1 0 9660 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_97
timestamp 1644511149
transform 1 0 10028 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_101
timestamp 1644511149
transform 1 0 10396 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_108
timestamp 1644511149
transform 1 0 11040 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_113
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_122
timestamp 1644511149
transform 1 0 12328 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_131
timestamp 1644511149
transform 1 0 13156 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_139
timestamp 1644511149
transform 1 0 13892 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_147
timestamp 1644511149
transform 1 0 14628 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_158
timestamp 1644511149
transform 1 0 15640 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_166
timestamp 1644511149
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_175
timestamp 1644511149
transform 1 0 17204 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_182
timestamp 1644511149
transform 1 0 17848 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_191
timestamp 1644511149
transform 1 0 18676 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_200
timestamp 1644511149
transform 1 0 19504 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_213
timestamp 1644511149
transform 1 0 20700 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_220
timestamp 1644511149
transform 1 0 21344 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_225
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_235
timestamp 1644511149
transform 1 0 22724 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_243
timestamp 1644511149
transform 1 0 23460 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_251
timestamp 1644511149
transform 1 0 24196 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_266
timestamp 1644511149
transform 1 0 25576 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_276
timestamp 1644511149
transform 1 0 26496 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_288
timestamp 1644511149
transform 1 0 27600 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_295
timestamp 1644511149
transform 1 0 28244 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1644511149
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1644511149
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_41
timestamp 1644511149
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_53
timestamp 1644511149
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_65
timestamp 1644511149
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1644511149
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1644511149
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_85
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_94
timestamp 1644511149
transform 1 0 9752 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_101
timestamp 1644511149
transform 1 0 10396 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_108
timestamp 1644511149
transform 1 0 11040 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_128
timestamp 1644511149
transform 1 0 12880 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_136
timestamp 1644511149
transform 1 0 13616 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_148
timestamp 1644511149
transform 1 0 14720 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_161
timestamp 1644511149
transform 1 0 15916 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_165
timestamp 1644511149
transform 1 0 16284 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_182
timestamp 1644511149
transform 1 0 17848 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_186
timestamp 1644511149
transform 1 0 18216 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_192
timestamp 1644511149
transform 1 0 18768 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_201
timestamp 1644511149
transform 1 0 19596 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_221
timestamp 1644511149
transform 1 0 21436 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_42_234
timestamp 1644511149
transform 1 0 22632 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_240
timestamp 1644511149
transform 1 0 23184 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_248
timestamp 1644511149
transform 1 0 23920 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_42_253
timestamp 1644511149
transform 1 0 24380 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_42_264
timestamp 1644511149
transform 1 0 25392 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_272
timestamp 1644511149
transform 1 0 26128 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_295
timestamp 1644511149
transform 1 0 28244 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1644511149
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1644511149
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_39
timestamp 1644511149
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1644511149
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1644511149
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_57
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_69
timestamp 1644511149
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_81
timestamp 1644511149
transform 1 0 8556 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_89
timestamp 1644511149
transform 1 0 9292 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_94
timestamp 1644511149
transform 1 0 9752 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_101
timestamp 1644511149
transform 1 0 10396 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_108
timestamp 1644511149
transform 1 0 11040 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_129
timestamp 1644511149
transform 1 0 12972 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_151
timestamp 1644511149
transform 1 0 14996 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_163
timestamp 1644511149
transform 1 0 16100 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1644511149
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_185
timestamp 1644511149
transform 1 0 18124 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_205
timestamp 1644511149
transform 1 0 19964 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_213
timestamp 1644511149
transform 1 0 20700 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_220
timestamp 1644511149
transform 1 0 21344 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_225
timestamp 1644511149
transform 1 0 21804 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_235
timestamp 1644511149
transform 1 0 22724 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_239
timestamp 1644511149
transform 1 0 23092 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_247
timestamp 1644511149
transform 1 0 23828 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_256
timestamp 1644511149
transform 1 0 24656 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_276
timestamp 1644511149
transform 1 0 26496 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_286
timestamp 1644511149
transform 1 0 27416 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_295
timestamp 1644511149
transform 1 0 28244 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1644511149
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1644511149
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_41
timestamp 1644511149
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_53
timestamp 1644511149
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_65
timestamp 1644511149
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1644511149
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1644511149
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_85
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_89
timestamp 1644511149
transform 1 0 9292 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_93
timestamp 1644511149
transform 1 0 9660 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_100
timestamp 1644511149
transform 1 0 10304 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_107
timestamp 1644511149
transform 1 0 10948 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_116
timestamp 1644511149
transform 1 0 11776 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_136
timestamp 1644511149
transform 1 0 13616 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_145
timestamp 1644511149
transform 1 0 14444 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_155
timestamp 1644511149
transform 1 0 15364 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_175
timestamp 1644511149
transform 1 0 17204 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_182
timestamp 1644511149
transform 1 0 17848 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_192
timestamp 1644511149
transform 1 0 18768 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_44_197
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_44_208
timestamp 1644511149
transform 1 0 20240 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_216
timestamp 1644511149
transform 1 0 20976 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_225
timestamp 1644511149
transform 1 0 21804 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_235
timestamp 1644511149
transform 1 0 22724 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_248
timestamp 1644511149
transform 1 0 23920 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_253
timestamp 1644511149
transform 1 0 24380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_260
timestamp 1644511149
transform 1 0 25024 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_270
timestamp 1644511149
transform 1 0 25944 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_295
timestamp 1644511149
transform 1 0 28244 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1644511149
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1644511149
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_27
timestamp 1644511149
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_39
timestamp 1644511149
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1644511149
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1644511149
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_69
timestamp 1644511149
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_81
timestamp 1644511149
transform 1 0 8556 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_87
timestamp 1644511149
transform 1 0 9108 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_94
timestamp 1644511149
transform 1 0 9752 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_101
timestamp 1644511149
transform 1 0 10396 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_108
timestamp 1644511149
transform 1 0 11040 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_45_113
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_121
timestamp 1644511149
transform 1 0 12236 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_132
timestamp 1644511149
transform 1 0 13248 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_142
timestamp 1644511149
transform 1 0 14168 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_148
timestamp 1644511149
transform 1 0 14720 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_155
timestamp 1644511149
transform 1 0 15364 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_164
timestamp 1644511149
transform 1 0 16192 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_169
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_176
timestamp 1644511149
transform 1 0 17296 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_187
timestamp 1644511149
transform 1 0 18308 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_194
timestamp 1644511149
transform 1 0 18952 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_214
timestamp 1644511149
transform 1 0 20792 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_222
timestamp 1644511149
transform 1 0 21528 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_232
timestamp 1644511149
transform 1 0 22448 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_240
timestamp 1644511149
transform 1 0 23184 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_260
timestamp 1644511149
transform 1 0 25024 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_270
timestamp 1644511149
transform 1 0 25944 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_278
timestamp 1644511149
transform 1 0 26680 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_281
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_291
timestamp 1644511149
transform 1 0 27876 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1644511149
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1644511149
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_41
timestamp 1644511149
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_53
timestamp 1644511149
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_65
timestamp 1644511149
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_80
timestamp 1644511149
transform 1 0 8464 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_85
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_92
timestamp 1644511149
transform 1 0 9568 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_99
timestamp 1644511149
transform 1 0 10212 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_106
timestamp 1644511149
transform 1 0 10856 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_126
timestamp 1644511149
transform 1 0 12696 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_136
timestamp 1644511149
transform 1 0 13616 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_157
timestamp 1644511149
transform 1 0 15548 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_181
timestamp 1644511149
transform 1 0 17756 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_192
timestamp 1644511149
transform 1 0 18768 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_197
timestamp 1644511149
transform 1 0 19228 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_221
timestamp 1644511149
transform 1 0 21436 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_227
timestamp 1644511149
transform 1 0 21988 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_234
timestamp 1644511149
transform 1 0 22632 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_238
timestamp 1644511149
transform 1 0 23000 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_244
timestamp 1644511149
transform 1 0 23552 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_253
timestamp 1644511149
transform 1 0 24380 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_270
timestamp 1644511149
transform 1 0 25944 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_295
timestamp 1644511149
transform 1 0 28244 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1644511149
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1644511149
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1644511149
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_39
timestamp 1644511149
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1644511149
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1644511149
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_69
timestamp 1644511149
transform 1 0 7452 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_47_80
timestamp 1644511149
transform 1 0 8464 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_88
timestamp 1644511149
transform 1 0 9200 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_92
timestamp 1644511149
transform 1 0 9568 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_99
timestamp 1644511149
transform 1 0 10212 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_108
timestamp 1644511149
transform 1 0 11040 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_113
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_117
timestamp 1644511149
transform 1 0 11868 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_123
timestamp 1644511149
transform 1 0 12420 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_129
timestamp 1644511149
transform 1 0 12972 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_138
timestamp 1644511149
transform 1 0 13800 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_158
timestamp 1644511149
transform 1 0 15640 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_166
timestamp 1644511149
transform 1 0 16376 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_169
timestamp 1644511149
transform 1 0 16652 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_173
timestamp 1644511149
transform 1 0 17020 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_190
timestamp 1644511149
transform 1 0 18584 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_210
timestamp 1644511149
transform 1 0 20424 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_214
timestamp 1644511149
transform 1 0 20792 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_220
timestamp 1644511149
transform 1 0 21344 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_228
timestamp 1644511149
transform 1 0 22080 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_248
timestamp 1644511149
transform 1 0 23920 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_256
timestamp 1644511149
transform 1 0 24656 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_276
timestamp 1644511149
transform 1 0 26496 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_287
timestamp 1644511149
transform 1 0 27508 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_295
timestamp 1644511149
transform 1 0 28244 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_3
timestamp 1644511149
transform 1 0 1380 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_48_8
timestamp 1644511149
transform 1 0 1840 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_20
timestamp 1644511149
transform 1 0 2944 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1644511149
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_53
timestamp 1644511149
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_65
timestamp 1644511149
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_80
timestamp 1644511149
transform 1 0 8464 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_48_85
timestamp 1644511149
transform 1 0 8924 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_91
timestamp 1644511149
transform 1 0 9476 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_98
timestamp 1644511149
transform 1 0 10120 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_106
timestamp 1644511149
transform 1 0 10856 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_126
timestamp 1644511149
transform 1 0 12696 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_136
timestamp 1644511149
transform 1 0 13616 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_144
timestamp 1644511149
transform 1 0 14352 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_153
timestamp 1644511149
transform 1 0 15180 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_159
timestamp 1644511149
transform 1 0 15732 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_165
timestamp 1644511149
transform 1 0 16284 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_179
timestamp 1644511149
transform 1 0 17572 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1644511149
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1644511149
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_197
timestamp 1644511149
transform 1 0 19228 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_206
timestamp 1644511149
transform 1 0 20056 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_220
timestamp 1644511149
transform 1 0 21344 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_240
timestamp 1644511149
transform 1 0 23184 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_248
timestamp 1644511149
transform 1 0 23920 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_269
timestamp 1644511149
transform 1 0 25852 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_273
timestamp 1644511149
transform 1 0 26220 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_295
timestamp 1644511149
transform 1 0 28244 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_24
timestamp 1644511149
transform 1 0 3312 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_36
timestamp 1644511149
transform 1 0 4416 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_48
timestamp 1644511149
transform 1 0 5520 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_69
timestamp 1644511149
transform 1 0 7452 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_73
timestamp 1644511149
transform 1 0 7820 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_80
timestamp 1644511149
transform 1 0 8464 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_87
timestamp 1644511149
transform 1 0 9108 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_94
timestamp 1644511149
transform 1 0 9752 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_101
timestamp 1644511149
transform 1 0 10396 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_108
timestamp 1644511149
transform 1 0 11040 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_49_113
timestamp 1644511149
transform 1 0 11500 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_120
timestamp 1644511149
transform 1 0 12144 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_140
timestamp 1644511149
transform 1 0 13984 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_148
timestamp 1644511149
transform 1 0 14720 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_154
timestamp 1644511149
transform 1 0 15272 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_164
timestamp 1644511149
transform 1 0 16192 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_173
timestamp 1644511149
transform 1 0 17020 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_193
timestamp 1644511149
transform 1 0 18860 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_201
timestamp 1644511149
transform 1 0 19596 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_218
timestamp 1644511149
transform 1 0 21160 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_49_225
timestamp 1644511149
transform 1 0 21804 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_233
timestamp 1644511149
transform 1 0 22540 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_237
timestamp 1644511149
transform 1 0 22908 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_248
timestamp 1644511149
transform 1 0 23920 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_268
timestamp 1644511149
transform 1 0 25760 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_276
timestamp 1644511149
transform 1 0 26496 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_287
timestamp 1644511149
transform 1 0 27508 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_295
timestamp 1644511149
transform 1 0 28244 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_6
timestamp 1644511149
transform 1 0 1656 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_18
timestamp 1644511149
transform 1 0 2760 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_26
timestamp 1644511149
transform 1 0 3496 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_29
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_41
timestamp 1644511149
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_53
timestamp 1644511149
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_65
timestamp 1644511149
transform 1 0 7084 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_69
timestamp 1644511149
transform 1 0 7452 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_73
timestamp 1644511149
transform 1 0 7820 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_80
timestamp 1644511149
transform 1 0 8464 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_50_85
timestamp 1644511149
transform 1 0 8924 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_91
timestamp 1644511149
transform 1 0 9476 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_95
timestamp 1644511149
transform 1 0 9844 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_100
timestamp 1644511149
transform 1 0 10304 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_107
timestamp 1644511149
transform 1 0 10948 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_116
timestamp 1644511149
transform 1 0 11776 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_136
timestamp 1644511149
transform 1 0 13616 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_144
timestamp 1644511149
transform 1 0 14352 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_164
timestamp 1644511149
transform 1 0 16192 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_184
timestamp 1644511149
transform 1 0 18032 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_192
timestamp 1644511149
transform 1 0 18768 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_202
timestamp 1644511149
transform 1 0 19688 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_208
timestamp 1644511149
transform 1 0 20240 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_230
timestamp 1644511149
transform 1 0 22264 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_238
timestamp 1644511149
transform 1 0 23000 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_248
timestamp 1644511149
transform 1 0 23920 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_253
timestamp 1644511149
transform 1 0 24380 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_270
timestamp 1644511149
transform 1 0 25944 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_295
timestamp 1644511149
transform 1 0 28244 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1644511149
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_15
timestamp 1644511149
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_27
timestamp 1644511149
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_39
timestamp 1644511149
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1644511149
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1644511149
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_57
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_64
timestamp 1644511149
transform 1 0 6992 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_68
timestamp 1644511149
transform 1 0 7360 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_78
timestamp 1644511149
transform 1 0 8280 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_85
timestamp 1644511149
transform 1 0 8924 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_92
timestamp 1644511149
transform 1 0 9568 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_100
timestamp 1644511149
transform 1 0 10304 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_108
timestamp 1644511149
transform 1 0 11040 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_129
timestamp 1644511149
transform 1 0 12972 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_136
timestamp 1644511149
transform 1 0 13616 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_156
timestamp 1644511149
transform 1 0 15456 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_164
timestamp 1644511149
transform 1 0 16192 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_169
timestamp 1644511149
transform 1 0 16652 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_173
timestamp 1644511149
transform 1 0 17020 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_190
timestamp 1644511149
transform 1 0 18584 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_210
timestamp 1644511149
transform 1 0 20424 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_220
timestamp 1644511149
transform 1 0 21344 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_241
timestamp 1644511149
transform 1 0 23276 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_255
timestamp 1644511149
transform 1 0 24564 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_261
timestamp 1644511149
transform 1 0 25116 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_271
timestamp 1644511149
transform 1 0 26036 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1644511149
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_290
timestamp 1644511149
transform 1 0 27784 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_298
timestamp 1644511149
transform 1 0 28520 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_3
timestamp 1644511149
transform 1 0 1380 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_11
timestamp 1644511149
transform 1 0 2116 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_15
timestamp 1644511149
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1644511149
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_29
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_41
timestamp 1644511149
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_53
timestamp 1644511149
transform 1 0 5980 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_61
timestamp 1644511149
transform 1 0 6716 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_66
timestamp 1644511149
transform 1 0 7176 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_73
timestamp 1644511149
transform 1 0 7820 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_80
timestamp 1644511149
transform 1 0 8464 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_52_85
timestamp 1644511149
transform 1 0 8924 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_91
timestamp 1644511149
transform 1 0 9476 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_100
timestamp 1644511149
transform 1 0 10304 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_109
timestamp 1644511149
transform 1 0 11132 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_118
timestamp 1644511149
transform 1 0 11960 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_127
timestamp 1644511149
transform 1 0 12788 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_136
timestamp 1644511149
transform 1 0 13616 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_146
timestamp 1644511149
transform 1 0 14536 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_155
timestamp 1644511149
transform 1 0 15364 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_159
timestamp 1644511149
transform 1 0 15732 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_167
timestamp 1644511149
transform 1 0 16468 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_179
timestamp 1644511149
transform 1 0 17572 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_192
timestamp 1644511149
transform 1 0 18768 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_197
timestamp 1644511149
transform 1 0 19228 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_201
timestamp 1644511149
transform 1 0 19596 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_208
timestamp 1644511149
transform 1 0 20240 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_212
timestamp 1644511149
transform 1 0 20608 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_229
timestamp 1644511149
transform 1 0 22172 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_52_242
timestamp 1644511149
transform 1 0 23368 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_250
timestamp 1644511149
transform 1 0 24104 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_258
timestamp 1644511149
transform 1 0 24840 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_270
timestamp 1644511149
transform 1 0 25944 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_295
timestamp 1644511149
transform 1 0 28244 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_53_3
timestamp 1644511149
transform 1 0 1380 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_27
timestamp 1644511149
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_39
timestamp 1644511149
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1644511149
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1644511149
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_57
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_62
timestamp 1644511149
transform 1 0 6808 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_69
timestamp 1644511149
transform 1 0 7452 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_76
timestamp 1644511149
transform 1 0 8096 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_83
timestamp 1644511149
transform 1 0 8740 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_90
timestamp 1644511149
transform 1 0 9384 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_99
timestamp 1644511149
transform 1 0 10212 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_108
timestamp 1644511149
transform 1 0 11040 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_117
timestamp 1644511149
transform 1 0 11868 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_126
timestamp 1644511149
transform 1 0 12696 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_135
timestamp 1644511149
transform 1 0 13524 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_144
timestamp 1644511149
transform 1 0 14352 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_164
timestamp 1644511149
transform 1 0 16192 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_175
timestamp 1644511149
transform 1 0 17204 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_179
timestamp 1644511149
transform 1 0 17572 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_196
timestamp 1644511149
transform 1 0 19136 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_220
timestamp 1644511149
transform 1 0 21344 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_225
timestamp 1644511149
transform 1 0 21804 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_232
timestamp 1644511149
transform 1 0 22448 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_243
timestamp 1644511149
transform 1 0 23460 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_256
timestamp 1644511149
transform 1 0 24656 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_276
timestamp 1644511149
transform 1 0 26496 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_287
timestamp 1644511149
transform 1 0 27508 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_295
timestamp 1644511149
transform 1 0 28244 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_3
timestamp 1644511149
transform 1 0 1380 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_8
timestamp 1644511149
transform 1 0 1840 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_15
timestamp 1644511149
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1644511149
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_29
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_41
timestamp 1644511149
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_53
timestamp 1644511149
transform 1 0 5980 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_57
timestamp 1644511149
transform 1 0 6348 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_64
timestamp 1644511149
transform 1 0 6992 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_73
timestamp 1644511149
transform 1 0 7820 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_80
timestamp 1644511149
transform 1 0 8464 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_85
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_89
timestamp 1644511149
transform 1 0 9292 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_93
timestamp 1644511149
transform 1 0 9660 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_102
timestamp 1644511149
transform 1 0 10488 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_111
timestamp 1644511149
transform 1 0 11316 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_131
timestamp 1644511149
transform 1 0 13156 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1644511149
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_157
timestamp 1644511149
transform 1 0 15548 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_163
timestamp 1644511149
transform 1 0 16100 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_180
timestamp 1644511149
transform 1 0 17664 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_186
timestamp 1644511149
transform 1 0 18216 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_192
timestamp 1644511149
transform 1 0 18768 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_197
timestamp 1644511149
transform 1 0 19228 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_210
timestamp 1644511149
transform 1 0 20424 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_220
timestamp 1644511149
transform 1 0 21344 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_230
timestamp 1644511149
transform 1 0 22264 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_238
timestamp 1644511149
transform 1 0 23000 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_248
timestamp 1644511149
transform 1 0 23920 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_253
timestamp 1644511149
transform 1 0 24380 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_270
timestamp 1644511149
transform 1 0 25944 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_295
timestamp 1644511149
transform 1 0 28244 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_3
timestamp 1644511149
transform 1 0 1380 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_25
timestamp 1644511149
transform 1 0 3404 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_37
timestamp 1644511149
transform 1 0 4508 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_49
timestamp 1644511149
transform 1 0 5612 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1644511149
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_65
timestamp 1644511149
transform 1 0 7084 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_70
timestamp 1644511149
transform 1 0 7544 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_77
timestamp 1644511149
transform 1 0 8188 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_84
timestamp 1644511149
transform 1 0 8832 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_91
timestamp 1644511149
transform 1 0 9476 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_99
timestamp 1644511149
transform 1 0 10212 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_108
timestamp 1644511149
transform 1 0 11040 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_129
timestamp 1644511149
transform 1 0 12972 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_139
timestamp 1644511149
transform 1 0 13892 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_159
timestamp 1644511149
transform 1 0 15732 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1644511149
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_55_169
timestamp 1644511149
transform 1 0 16652 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_177
timestamp 1644511149
transform 1 0 17388 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_185
timestamp 1644511149
transform 1 0 18124 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_202
timestamp 1644511149
transform 1 0 19688 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_210
timestamp 1644511149
transform 1 0 20424 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_220
timestamp 1644511149
transform 1 0 21344 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_241
timestamp 1644511149
transform 1 0 23276 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_261
timestamp 1644511149
transform 1 0 25116 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_272
timestamp 1644511149
transform 1 0 26128 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_288
timestamp 1644511149
transform 1 0 27600 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_295
timestamp 1644511149
transform 1 0 28244 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_6
timestamp 1644511149
transform 1 0 1656 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_18
timestamp 1644511149
transform 1 0 2760 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_26
timestamp 1644511149
transform 1 0 3496 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_29
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_41
timestamp 1644511149
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_53
timestamp 1644511149
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_65
timestamp 1644511149
transform 1 0 7084 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_69
timestamp 1644511149
transform 1 0 7452 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_73
timestamp 1644511149
transform 1 0 7820 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_80
timestamp 1644511149
transform 1 0 8464 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_85
timestamp 1644511149
transform 1 0 8924 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_94
timestamp 1644511149
transform 1 0 9752 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_103
timestamp 1644511149
transform 1 0 10580 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_123
timestamp 1644511149
transform 1 0 12420 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_134
timestamp 1644511149
transform 1 0 13432 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_56_149
timestamp 1644511149
transform 1 0 14812 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_157
timestamp 1644511149
transform 1 0 15548 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_174
timestamp 1644511149
transform 1 0 17112 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_182
timestamp 1644511149
transform 1 0 17848 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_192
timestamp 1644511149
transform 1 0 18768 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_202
timestamp 1644511149
transform 1 0 19688 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_215
timestamp 1644511149
transform 1 0 20884 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_235
timestamp 1644511149
transform 1 0 22724 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_246
timestamp 1644511149
transform 1 0 23736 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_253
timestamp 1644511149
transform 1 0 24380 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_262
timestamp 1644511149
transform 1 0 25208 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_270
timestamp 1644511149
transform 1 0 25944 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_295
timestamp 1644511149
transform 1 0 28244 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_7
timestamp 1644511149
transform 1 0 1748 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_14
timestamp 1644511149
transform 1 0 2392 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_26
timestamp 1644511149
transform 1 0 3496 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_38
timestamp 1644511149
transform 1 0 4600 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_50
timestamp 1644511149
transform 1 0 5704 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_69
timestamp 1644511149
transform 1 0 7452 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_73
timestamp 1644511149
transform 1 0 7820 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_80
timestamp 1644511149
transform 1 0 8464 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_87
timestamp 1644511149
transform 1 0 9108 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_94
timestamp 1644511149
transform 1 0 9752 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_101
timestamp 1644511149
transform 1 0 10396 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_108
timestamp 1644511149
transform 1 0 11040 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_113
timestamp 1644511149
transform 1 0 11500 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_117
timestamp 1644511149
transform 1 0 11868 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_123
timestamp 1644511149
transform 1 0 12420 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_130
timestamp 1644511149
transform 1 0 13064 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_150
timestamp 1644511149
transform 1 0 14904 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_164
timestamp 1644511149
transform 1 0 16192 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_169
timestamp 1644511149
transform 1 0 16652 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_191
timestamp 1644511149
transform 1 0 18676 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_199
timestamp 1644511149
transform 1 0 19412 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_219
timestamp 1644511149
transform 1 0 21252 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1644511149
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_233
timestamp 1644511149
transform 1 0 22540 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_241
timestamp 1644511149
transform 1 0 23276 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_250
timestamp 1644511149
transform 1 0 24104 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_254
timestamp 1644511149
transform 1 0 24472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_276
timestamp 1644511149
transform 1 0 26496 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_288
timestamp 1644511149
transform 1 0 27600 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_295
timestamp 1644511149
transform 1 0 28244 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_24
timestamp 1644511149
transform 1 0 3312 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1644511149
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_41
timestamp 1644511149
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_53
timestamp 1644511149
transform 1 0 5980 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_61
timestamp 1644511149
transform 1 0 6716 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_66
timestamp 1644511149
transform 1 0 7176 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_73
timestamp 1644511149
transform 1 0 7820 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_80
timestamp 1644511149
transform 1 0 8464 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_85
timestamp 1644511149
transform 1 0 8924 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_89
timestamp 1644511149
transform 1 0 9292 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_96
timestamp 1644511149
transform 1 0 9936 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_105
timestamp 1644511149
transform 1 0 10764 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_114
timestamp 1644511149
transform 1 0 11592 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_123
timestamp 1644511149
transform 1 0 12420 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_129
timestamp 1644511149
transform 1 0 12972 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_136
timestamp 1644511149
transform 1 0 13616 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_148
timestamp 1644511149
transform 1 0 14720 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_156
timestamp 1644511149
transform 1 0 15456 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_173
timestamp 1644511149
transform 1 0 17020 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_181
timestamp 1644511149
transform 1 0 17756 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_192
timestamp 1644511149
transform 1 0 18768 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_213
timestamp 1644511149
transform 1 0 20700 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_223
timestamp 1644511149
transform 1 0 21620 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_233
timestamp 1644511149
transform 1 0 22540 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_243
timestamp 1644511149
transform 1 0 23460 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1644511149
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_258
timestamp 1644511149
transform 1 0 24840 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_269
timestamp 1644511149
transform 1 0 25852 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_273
timestamp 1644511149
transform 1 0 26220 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_295
timestamp 1644511149
transform 1 0 28244 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_59_3
timestamp 1644511149
transform 1 0 1380 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_27
timestamp 1644511149
transform 1 0 3588 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_34
timestamp 1644511149
transform 1 0 4232 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_46
timestamp 1644511149
transform 1 0 5336 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_54
timestamp 1644511149
transform 1 0 6072 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_59_57
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_66
timestamp 1644511149
transform 1 0 7176 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_73
timestamp 1644511149
transform 1 0 7820 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_80
timestamp 1644511149
transform 1 0 8464 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_87
timestamp 1644511149
transform 1 0 9108 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_94
timestamp 1644511149
transform 1 0 9752 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_101
timestamp 1644511149
transform 1 0 10396 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_108
timestamp 1644511149
transform 1 0 11040 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_129
timestamp 1644511149
transform 1 0 12972 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_149
timestamp 1644511149
transform 1 0 14812 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_157
timestamp 1644511149
transform 1 0 15548 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_164
timestamp 1644511149
transform 1 0 16192 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_174
timestamp 1644511149
transform 1 0 17112 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_183
timestamp 1644511149
transform 1 0 17940 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_203
timestamp 1644511149
transform 1 0 19780 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_215
timestamp 1644511149
transform 1 0 20884 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1644511149
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_229
timestamp 1644511149
transform 1 0 22172 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_240
timestamp 1644511149
transform 1 0 23184 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_251
timestamp 1644511149
transform 1 0 24196 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_260
timestamp 1644511149
transform 1 0 25024 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_271
timestamp 1644511149
transform 1 0 26036 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1644511149
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_287
timestamp 1644511149
transform 1 0 27508 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_295
timestamp 1644511149
transform 1 0 28244 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_60_3
timestamp 1644511149
transform 1 0 1380 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_9
timestamp 1644511149
transform 1 0 1932 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_13
timestamp 1644511149
transform 1 0 2300 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_17
timestamp 1644511149
transform 1 0 2668 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_24
timestamp 1644511149
transform 1 0 3312 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_32
timestamp 1644511149
transform 1 0 4048 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_39
timestamp 1644511149
transform 1 0 4692 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_60_47
timestamp 1644511149
transform 1 0 5428 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_52
timestamp 1644511149
transform 1 0 5888 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_59
timestamp 1644511149
transform 1 0 6532 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_66
timestamp 1644511149
transform 1 0 7176 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_73
timestamp 1644511149
transform 1 0 7820 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_80
timestamp 1644511149
transform 1 0 8464 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_85
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_90
timestamp 1644511149
transform 1 0 9384 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_97
timestamp 1644511149
transform 1 0 10028 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_104
timestamp 1644511149
transform 1 0 10672 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_111
timestamp 1644511149
transform 1 0 11316 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_119
timestamp 1644511149
transform 1 0 12052 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_128
timestamp 1644511149
transform 1 0 12880 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_136
timestamp 1644511149
transform 1 0 13616 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_146
timestamp 1644511149
transform 1 0 14536 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_154
timestamp 1644511149
transform 1 0 15272 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_174
timestamp 1644511149
transform 1 0 17112 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_182
timestamp 1644511149
transform 1 0 17848 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_192
timestamp 1644511149
transform 1 0 18768 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_200
timestamp 1644511149
transform 1 0 19504 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_220
timestamp 1644511149
transform 1 0 21344 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_231
timestamp 1644511149
transform 1 0 22356 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_242
timestamp 1644511149
transform 1 0 23368 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_250
timestamp 1644511149
transform 1 0 24104 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_263
timestamp 1644511149
transform 1 0 25300 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_270
timestamp 1644511149
transform 1 0 25944 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_295
timestamp 1644511149
transform 1 0 28244 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_3
timestamp 1644511149
transform 1 0 1380 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_25
timestamp 1644511149
transform 1 0 3404 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_32
timestamp 1644511149
transform 1 0 4048 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_39
timestamp 1644511149
transform 1 0 4692 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_46
timestamp 1644511149
transform 1 0 5336 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_54
timestamp 1644511149
transform 1 0 6072 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_60
timestamp 1644511149
transform 1 0 6624 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_71
timestamp 1644511149
transform 1 0 7636 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_78
timestamp 1644511149
transform 1 0 8280 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_85
timestamp 1644511149
transform 1 0 8924 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_92
timestamp 1644511149
transform 1 0 9568 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_99
timestamp 1644511149
transform 1 0 10212 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_108
timestamp 1644511149
transform 1 0 11040 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_113
timestamp 1644511149
transform 1 0 11500 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_117
timestamp 1644511149
transform 1 0 11868 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_121
timestamp 1644511149
transform 1 0 12236 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_129
timestamp 1644511149
transform 1 0 12972 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_138
timestamp 1644511149
transform 1 0 13800 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_147
timestamp 1644511149
transform 1 0 14628 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_153
timestamp 1644511149
transform 1 0 15180 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_160
timestamp 1644511149
transform 1 0 15824 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_172
timestamp 1644511149
transform 1 0 16928 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_181
timestamp 1644511149
transform 1 0 17756 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_193
timestamp 1644511149
transform 1 0 18860 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_201
timestamp 1644511149
transform 1 0 19596 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_208
timestamp 1644511149
transform 1 0 20240 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_220
timestamp 1644511149
transform 1 0 21344 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_234
timestamp 1644511149
transform 1 0 22632 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_249
timestamp 1644511149
transform 1 0 24012 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_256
timestamp 1644511149
transform 1 0 24656 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_276
timestamp 1644511149
transform 1 0 26496 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_290
timestamp 1644511149
transform 1 0 27784 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_294
timestamp 1644511149
transform 1 0 28152 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_298
timestamp 1644511149
transform 1 0 28520 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_62_3
timestamp 1644511149
transform 1 0 1380 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_7
timestamp 1644511149
transform 1 0 1748 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_24
timestamp 1644511149
transform 1 0 3312 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_32
timestamp 1644511149
transform 1 0 4048 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_39
timestamp 1644511149
transform 1 0 4692 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_46
timestamp 1644511149
transform 1 0 5336 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_54
timestamp 1644511149
transform 1 0 6072 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_59
timestamp 1644511149
transform 1 0 6532 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_66
timestamp 1644511149
transform 1 0 7176 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_73
timestamp 1644511149
transform 1 0 7820 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_80
timestamp 1644511149
transform 1 0 8464 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_88
timestamp 1644511149
transform 1 0 9200 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_95
timestamp 1644511149
transform 1 0 9844 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_102
timestamp 1644511149
transform 1 0 10488 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_111
timestamp 1644511149
transform 1 0 11316 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_115
timestamp 1644511149
transform 1 0 11684 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_132
timestamp 1644511149
transform 1 0 13248 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_157
timestamp 1644511149
transform 1 0 15548 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_166
timestamp 1644511149
transform 1 0 16376 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_186
timestamp 1644511149
transform 1 0 18216 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_194
timestamp 1644511149
transform 1 0 18952 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_204
timestamp 1644511149
transform 1 0 19872 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_217
timestamp 1644511149
transform 1 0 21068 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_221
timestamp 1644511149
transform 1 0 21436 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_229
timestamp 1644511149
transform 1 0 22172 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_62_243
timestamp 1644511149
transform 1 0 23460 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1644511149
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_261
timestamp 1644511149
transform 1 0 25116 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_270
timestamp 1644511149
transform 1 0 25944 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_295
timestamp 1644511149
transform 1 0 28244 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_3
timestamp 1644511149
transform 1 0 1380 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_7
timestamp 1644511149
transform 1 0 1748 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_15
timestamp 1644511149
transform 1 0 2484 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_31
timestamp 1644511149
transform 1 0 3956 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_44
timestamp 1644511149
transform 1 0 5152 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1644511149
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1644511149
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_57
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_66
timestamp 1644511149
transform 1 0 7176 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_70
timestamp 1644511149
transform 1 0 7544 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_74
timestamp 1644511149
transform 1 0 7912 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_81
timestamp 1644511149
transform 1 0 8556 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_88
timestamp 1644511149
transform 1 0 9200 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_95
timestamp 1644511149
transform 1 0 9844 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_108
timestamp 1644511149
transform 1 0 11040 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_63_113
timestamp 1644511149
transform 1 0 11500 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_132
timestamp 1644511149
transform 1 0 13248 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_152
timestamp 1644511149
transform 1 0 15088 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_163
timestamp 1644511149
transform 1 0 16100 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1644511149
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_174
timestamp 1644511149
transform 1 0 17112 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_194
timestamp 1644511149
transform 1 0 18952 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_214
timestamp 1644511149
transform 1 0 20792 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_222
timestamp 1644511149
transform 1 0 21528 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_229
timestamp 1644511149
transform 1 0 22172 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_241
timestamp 1644511149
transform 1 0 23276 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_251
timestamp 1644511149
transform 1 0 24196 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_276
timestamp 1644511149
transform 1 0 26496 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_287
timestamp 1644511149
transform 1 0 27508 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_295
timestamp 1644511149
transform 1 0 28244 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_24
timestamp 1644511149
transform 1 0 3312 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_38
timestamp 1644511149
transform 1 0 4600 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_51
timestamp 1644511149
transform 1 0 5796 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_58
timestamp 1644511149
transform 1 0 6440 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_62
timestamp 1644511149
transform 1 0 6808 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_66
timestamp 1644511149
transform 1 0 7176 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_73
timestamp 1644511149
transform 1 0 7820 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_80
timestamp 1644511149
transform 1 0 8464 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_88
timestamp 1644511149
transform 1 0 9200 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_96
timestamp 1644511149
transform 1 0 9936 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_109
timestamp 1644511149
transform 1 0 11132 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_122
timestamp 1644511149
transform 1 0 12328 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1644511149
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1644511149
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_141
timestamp 1644511149
transform 1 0 14076 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_145
timestamp 1644511149
transform 1 0 14444 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_162
timestamp 1644511149
transform 1 0 16008 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_182
timestamp 1644511149
transform 1 0 17848 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_192
timestamp 1644511149
transform 1 0 18768 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_197
timestamp 1644511149
transform 1 0 19228 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_204
timestamp 1644511149
transform 1 0 19872 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_217
timestamp 1644511149
transform 1 0 21068 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_227
timestamp 1644511149
transform 1 0 21988 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_231
timestamp 1644511149
transform 1 0 22356 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_248
timestamp 1644511149
transform 1 0 23920 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_269
timestamp 1644511149
transform 1 0 25852 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_273
timestamp 1644511149
transform 1 0 26220 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_295
timestamp 1644511149
transform 1 0 28244 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_3
timestamp 1644511149
transform 1 0 1380 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_26
timestamp 1644511149
transform 1 0 3496 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1644511149
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1644511149
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_60
timestamp 1644511149
transform 1 0 6624 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_68
timestamp 1644511149
transform 1 0 7360 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_72
timestamp 1644511149
transform 1 0 7728 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_79
timestamp 1644511149
transform 1 0 8372 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_92
timestamp 1644511149
transform 1 0 9568 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_108
timestamp 1644511149
transform 1 0 11040 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_113
timestamp 1644511149
transform 1 0 11500 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_118
timestamp 1644511149
transform 1 0 11960 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_143
timestamp 1644511149
transform 1 0 14260 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_152
timestamp 1644511149
transform 1 0 15088 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_158
timestamp 1644511149
transform 1 0 15640 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_164
timestamp 1644511149
transform 1 0 16192 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_185
timestamp 1644511149
transform 1 0 18124 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_205
timestamp 1644511149
transform 1 0 19964 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_218
timestamp 1644511149
transform 1 0 21160 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_65_246
timestamp 1644511149
transform 1 0 23736 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_254
timestamp 1644511149
transform 1 0 24472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_276
timestamp 1644511149
transform 1 0 26496 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_287
timestamp 1644511149
transform 1 0 27508 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_295
timestamp 1644511149
transform 1 0 28244 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_24
timestamp 1644511149
transform 1 0 3312 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_66_29
timestamp 1644511149
transform 1 0 3772 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_66_35
timestamp 1644511149
transform 1 0 4324 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_60
timestamp 1644511149
transform 1 0 6624 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_68
timestamp 1644511149
transform 1 0 7360 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_73
timestamp 1644511149
transform 1 0 7820 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_80
timestamp 1644511149
transform 1 0 8464 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_85
timestamp 1644511149
transform 1 0 8924 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_89
timestamp 1644511149
transform 1 0 9292 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_96
timestamp 1644511149
transform 1 0 9936 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_121
timestamp 1644511149
transform 1 0 12236 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_129
timestamp 1644511149
transform 1 0 12972 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_66_134
timestamp 1644511149
transform 1 0 13432 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_66_141
timestamp 1644511149
transform 1 0 14076 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_146
timestamp 1644511149
transform 1 0 14536 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_153
timestamp 1644511149
transform 1 0 15180 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_178
timestamp 1644511149
transform 1 0 17480 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_187
timestamp 1644511149
transform 1 0 18308 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1644511149
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_202
timestamp 1644511149
transform 1 0 19688 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_206
timestamp 1644511149
transform 1 0 20056 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_228
timestamp 1644511149
transform 1 0 22080 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_237
timestamp 1644511149
transform 1 0 22908 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_241
timestamp 1644511149
transform 1 0 23276 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_248
timestamp 1644511149
transform 1 0 23920 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_261
timestamp 1644511149
transform 1 0 25116 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_270
timestamp 1644511149
transform 1 0 25944 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_295
timestamp 1644511149
transform 1 0 28244 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_3
timestamp 1644511149
transform 1 0 1380 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_25
timestamp 1644511149
transform 1 0 3404 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_50
timestamp 1644511149
transform 1 0 5704 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_67_60
timestamp 1644511149
transform 1 0 6624 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_67_69
timestamp 1644511149
transform 1 0 7452 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_76
timestamp 1644511149
transform 1 0 8096 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_83
timestamp 1644511149
transform 1 0 8740 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_90
timestamp 1644511149
transform 1 0 9384 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_97
timestamp 1644511149
transform 1 0 10028 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_104
timestamp 1644511149
transform 1 0 10672 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_113
timestamp 1644511149
transform 1 0 11500 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_118
timestamp 1644511149
transform 1 0 11960 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_125
timestamp 1644511149
transform 1 0 12604 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_150
timestamp 1644511149
transform 1 0 14904 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_156
timestamp 1644511149
transform 1 0 15456 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_160
timestamp 1644511149
transform 1 0 15824 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_67_174
timestamp 1644511149
transform 1 0 17112 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_199
timestamp 1644511149
transform 1 0 19412 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_208
timestamp 1644511149
transform 1 0 20240 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1644511149
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1644511149
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_225
timestamp 1644511149
transform 1 0 21804 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_229
timestamp 1644511149
transform 1 0 22172 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_251
timestamp 1644511149
transform 1 0 24196 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_276
timestamp 1644511149
transform 1 0 26496 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_286
timestamp 1644511149
transform 1 0 27416 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_290
timestamp 1644511149
transform 1 0 27784 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_295
timestamp 1644511149
transform 1 0 28244 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_3
timestamp 1644511149
transform 1 0 1380 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_10
timestamp 1644511149
transform 1 0 2024 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_17
timestamp 1644511149
transform 1 0 2668 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_24
timestamp 1644511149
transform 1 0 3312 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_50
timestamp 1644511149
transform 1 0 5704 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_68_57
timestamp 1644511149
transform 1 0 6348 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_68_66
timestamp 1644511149
transform 1 0 7176 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_73
timestamp 1644511149
transform 1 0 7820 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_80
timestamp 1644511149
transform 1 0 8464 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_85
timestamp 1644511149
transform 1 0 8924 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_68_94
timestamp 1644511149
transform 1 0 9752 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_101
timestamp 1644511149
transform 1 0 10396 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_108
timestamp 1644511149
transform 1 0 11040 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_113
timestamp 1644511149
transform 1 0 11500 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_135
timestamp 1644511149
transform 1 0 13524 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1644511149
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_141
timestamp 1644511149
transform 1 0 14076 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_164
timestamp 1644511149
transform 1 0 16192 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_172
timestamp 1644511149
transform 1 0 16928 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_179
timestamp 1644511149
transform 1 0 17572 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_188
timestamp 1644511149
transform 1 0 18400 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_197
timestamp 1644511149
transform 1 0 19228 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_220
timestamp 1644511149
transform 1 0 21344 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_225
timestamp 1644511149
transform 1 0 21804 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_248
timestamp 1644511149
transform 1 0 23920 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_253
timestamp 1644511149
transform 1 0 24380 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_276
timestamp 1644511149
transform 1 0 26496 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_281
timestamp 1644511149
transform 1 0 26956 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_289
timestamp 1644511149
transform 1 0 27692 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_297
timestamp 1644511149
transform 1 0 28428 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 28888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 28888 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 28888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 28888 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 28888 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 28888 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 28888 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 28888 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 28888 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 28888 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 28888 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 28888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 28888 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 28888 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 28888 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 28888 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 28888 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 28888 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 28888 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 28888 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 28888 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 28888 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 28888 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 28888 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 28888 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 28888 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 28888 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 28888 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 28888 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 28888 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 28888 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 28888 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 28888 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 28888 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 28888 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 28888 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 28888 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 28888 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 28888 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 28888 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 28888 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 28888 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 28888 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 28888 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 28888 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 28888 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 28888 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 28888 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 28888 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 28888 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 28888 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 28888 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 28888 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 28888 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 28888 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 28888 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 28888 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 28888 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 28888 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 28888 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 28888 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 28888 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 28888 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 28888 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 28888 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1644511149
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1644511149
transform -1 0 28888 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1644511149
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1644511149
transform -1 0 28888 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1644511149
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1644511149
transform -1 0 28888 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1644511149
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1644511149
transform -1 0 28888 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1644511149
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1644511149
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1644511149
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1644511149
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1644511149
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1644511149
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1644511149
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1644511149
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1644511149
transform 1 0 6256 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1644511149
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1644511149
transform 1 0 11408 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1644511149
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1644511149
transform 1 0 16560 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1644511149
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1644511149
transform 1 0 21712 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1644511149
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1644511149
transform 1 0 26864 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _0708_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19044 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _0709_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20792 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0710_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24748 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0711_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5336 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0712_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1748 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0713_
timestamp 1644511149
transform 1 0 14352 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0714_
timestamp 1644511149
transform 1 0 2484 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0715_
timestamp 1644511149
transform 1 0 24472 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0716_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27048 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0717_
timestamp 1644511149
transform 1 0 2392 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0718_
timestamp 1644511149
transform 1 0 27968 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0719_
timestamp 1644511149
transform 1 0 1748 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0720_
timestamp 1644511149
transform 1 0 1748 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0721_
timestamp 1644511149
transform 1 0 27968 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0722_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9568 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  _0723_
timestamp 1644511149
transform 1 0 10304 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0724_
timestamp 1644511149
transform 1 0 13156 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0725_
timestamp 1644511149
transform 1 0 15732 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0726_
timestamp 1644511149
transform 1 0 7636 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0727_
timestamp 1644511149
transform 1 0 27692 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0728_
timestamp 1644511149
transform 1 0 27048 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0729_
timestamp 1644511149
transform 1 0 8740 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0730_
timestamp 1644511149
transform 1 0 25668 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0731_
timestamp 1644511149
transform 1 0 27968 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0732_
timestamp 1644511149
transform 1 0 2392 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0733_
timestamp 1644511149
transform 1 0 27968 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0734_
timestamp 1644511149
transform 1 0 1840 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0735_
timestamp 1644511149
transform 1 0 10212 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0736_
timestamp 1644511149
transform 1 0 24380 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0737_
timestamp 1644511149
transform 1 0 15548 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0738_
timestamp 1644511149
transform 1 0 9660 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0739_
timestamp 1644511149
transform 1 0 27968 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0740_
timestamp 1644511149
transform 1 0 26220 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0741_
timestamp 1644511149
transform 1 0 11500 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0742_
timestamp 1644511149
transform 1 0 4600 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0743_
timestamp 1644511149
transform 1 0 19228 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0744_
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0745_
timestamp 1644511149
transform 1 0 17296 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0746_
timestamp 1644511149
transform 1 0 2392 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0747_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9936 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0748_
timestamp 1644511149
transform 1 0 4692 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0749_
timestamp 1644511149
transform 1 0 27692 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0750_
timestamp 1644511149
transform 1 0 2208 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0751_
timestamp 1644511149
transform 1 0 21804 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0752_
timestamp 1644511149
transform 1 0 10396 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0753_
timestamp 1644511149
transform 1 0 21804 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  _0754_
timestamp 1644511149
transform 1 0 20240 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0755_
timestamp 1644511149
transform 1 0 16652 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0756_
timestamp 1644511149
transform 1 0 1748 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0757_
timestamp 1644511149
transform 1 0 12972 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0758_
timestamp 1644511149
transform 1 0 1748 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0759_
timestamp 1644511149
transform 1 0 21068 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0760_
timestamp 1644511149
transform 1 0 21436 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0761_
timestamp 1644511149
transform 1 0 17572 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0762_
timestamp 1644511149
transform 1 0 18676 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0763_
timestamp 1644511149
transform 1 0 11960 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0764_
timestamp 1644511149
transform 1 0 14076 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0765_
timestamp 1644511149
transform 1 0 27784 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0766_
timestamp 1644511149
transform 1 0 20332 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0767_
timestamp 1644511149
transform 1 0 23000 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0768_
timestamp 1644511149
transform 1 0 1656 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0769_
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0770_
timestamp 1644511149
transform 1 0 16652 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0771_
timestamp 1644511149
transform 1 0 1564 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0772_
timestamp 1644511149
transform 1 0 19320 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0773_
timestamp 1644511149
transform 1 0 22080 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0774_
timestamp 1644511149
transform 1 0 21068 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0775_
timestamp 1644511149
transform 1 0 18216 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0776_
timestamp 1644511149
transform 1 0 14904 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0777_
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  _0778_
timestamp 1644511149
transform 1 0 20240 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0779_
timestamp 1644511149
transform 1 0 14260 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0780_
timestamp 1644511149
transform 1 0 27232 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0781_
timestamp 1644511149
transform 1 0 2116 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0782_
timestamp 1644511149
transform 1 0 11040 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0783_
timestamp 1644511149
transform 1 0 1840 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0784_
timestamp 1644511149
transform 1 0 2116 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  _0785_
timestamp 1644511149
transform 1 0 3772 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0786_
timestamp 1644511149
transform 1 0 12788 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0787_
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0788_
timestamp 1644511149
transform 1 0 4048 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0789_
timestamp 1644511149
transform 1 0 27784 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0790_
timestamp 1644511149
transform 1 0 11684 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0791_
timestamp 1644511149
transform 1 0 4324 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0792_
timestamp 1644511149
transform 1 0 27600 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0793_
timestamp 1644511149
transform 1 0 12328 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0794_
timestamp 1644511149
transform 1 0 17572 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0795_
timestamp 1644511149
transform 1 0 27140 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0796_
timestamp 1644511149
transform 1 0 2392 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0797_
timestamp 1644511149
transform 1 0 4968 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0798_
timestamp 1644511149
transform 1 0 25576 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0799_
timestamp 1644511149
transform 1 0 3036 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0800_
timestamp 1644511149
transform 1 0 27784 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0801_
timestamp 1644511149
transform 1 0 27048 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0802_
timestamp 1644511149
transform 1 0 2484 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0803_
timestamp 1644511149
transform 1 0 2852 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0804_
timestamp 1644511149
transform 1 0 17572 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0805_
timestamp 1644511149
transform 1 0 3772 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0806_
timestamp 1644511149
transform 1 0 2392 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0807_
timestamp 1644511149
transform 1 0 27692 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0808_
timestamp 1644511149
transform 1 0 7268 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0809_
timestamp 1644511149
transform 1 0 2484 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0810_
timestamp 1644511149
transform 1 0 9476 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0811_
timestamp 1644511149
transform 1 0 11684 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0812_
timestamp 1644511149
transform 1 0 6348 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0813_
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0814_
timestamp 1644511149
transform 1 0 1472 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0815_
timestamp 1644511149
transform 1 0 20056 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0816_
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0817_
timestamp 1644511149
transform 1 0 9660 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0818_
timestamp 1644511149
transform 1 0 10764 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0819_
timestamp 1644511149
transform 1 0 3772 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0820_
timestamp 1644511149
transform 1 0 14076 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0821_
timestamp 1644511149
transform 1 0 20516 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0822_
timestamp 1644511149
transform 1 0 27784 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0823_
timestamp 1644511149
transform 1 0 27784 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0824_
timestamp 1644511149
transform 1 0 2300 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0825_
timestamp 1644511149
transform 1 0 9752 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0826_
timestamp 1644511149
transform 1 0 27784 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0827_
timestamp 1644511149
transform 1 0 21068 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0828_
timestamp 1644511149
transform 1 0 9936 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0829_
timestamp 1644511149
transform 1 0 1656 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0830_
timestamp 1644511149
transform 1 0 1564 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0831_
timestamp 1644511149
transform 1 0 1564 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0832_
timestamp 1644511149
transform 1 0 1564 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0833_
timestamp 1644511149
transform 1 0 21712 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0834_
timestamp 1644511149
transform 1 0 13340 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0835_
timestamp 1644511149
transform 1 0 1656 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0836_
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0837_
timestamp 1644511149
transform 1 0 11868 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0838_
timestamp 1644511149
transform 1 0 3036 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0839_
timestamp 1644511149
transform 1 0 27140 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0840_
timestamp 1644511149
transform 1 0 19964 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0841_
timestamp 1644511149
transform 1 0 10396 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0842_
timestamp 1644511149
transform 1 0 10764 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0843_
timestamp 1644511149
transform 1 0 23552 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0844_
timestamp 1644511149
transform 1 0 18400 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _0845_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26956 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0846_
timestamp 1644511149
transform 1 0 25576 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0847_
timestamp 1644511149
transform 1 0 25668 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0848_
timestamp 1644511149
transform 1 0 24932 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0849_
timestamp 1644511149
transform 1 0 24840 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0850_
timestamp 1644511149
transform 1 0 23644 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0851_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24288 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0852_
timestamp 1644511149
transform 1 0 22632 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0853_
timestamp 1644511149
transform 1 0 17664 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0854_
timestamp 1644511149
transform 1 0 22816 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _0855_
timestamp 1644511149
transform 1 0 23092 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0856_
timestamp 1644511149
transform 1 0 12604 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0857_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21988 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0858_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22448 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0859_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22724 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0860_
timestamp 1644511149
transform 1 0 23552 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0861_
timestamp 1644511149
transform 1 0 23552 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0862_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23184 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0863_
timestamp 1644511149
transform 1 0 27876 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0864_
timestamp 1644511149
transform 1 0 24840 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0865_
timestamp 1644511149
transform 1 0 24104 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _0866_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25300 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0867_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26956 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0868_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25484 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0869_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27140 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0870_
timestamp 1644511149
transform 1 0 12604 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0871_
timestamp 1644511149
transform 1 0 11960 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0872_
timestamp 1644511149
transform 1 0 16652 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0873_
timestamp 1644511149
transform 1 0 16008 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0874_
timestamp 1644511149
transform 1 0 14352 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0875_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19228 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0876_
timestamp 1644511149
transform 1 0 14444 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0877_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17664 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _0878_
timestamp 1644511149
transform 1 0 18492 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0879_
timestamp 1644511149
transform 1 0 13616 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0880_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16928 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0881_
timestamp 1644511149
transform 1 0 17296 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0882_
timestamp 1644511149
transform 1 0 18492 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0883_
timestamp 1644511149
transform 1 0 18308 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0884_
timestamp 1644511149
transform 1 0 19320 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0885_
timestamp 1644511149
transform 1 0 19504 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _0886_
timestamp 1644511149
transform 1 0 20424 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0887_
timestamp 1644511149
transform 1 0 9936 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0888_
timestamp 1644511149
transform 1 0 24288 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a221oi_2  _0889_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20056 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0890_
timestamp 1644511149
transform 1 0 9384 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0891_
timestamp 1644511149
transform 1 0 9108 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0892_
timestamp 1644511149
transform 1 0 10212 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0893_
timestamp 1644511149
transform 1 0 10672 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0894_
timestamp 1644511149
transform 1 0 23368 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0895_
timestamp 1644511149
transform 1 0 10764 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0896_
timestamp 1644511149
transform 1 0 9200 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0897_
timestamp 1644511149
transform 1 0 8464 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0898_
timestamp 1644511149
transform 1 0 22724 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0899_
timestamp 1644511149
transform 1 0 23644 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__o22a_1  _0900_
timestamp 1644511149
transform 1 0 22816 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0901_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21896 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0902_
timestamp 1644511149
transform 1 0 23184 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0903_
timestamp 1644511149
transform 1 0 24012 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0904_
timestamp 1644511149
transform 1 0 25208 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0905_
timestamp 1644511149
transform 1 0 25208 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _0906_
timestamp 1644511149
transform 1 0 26956 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0907_
timestamp 1644511149
transform 1 0 19228 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a211oi_1  _0908_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26956 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0909_
timestamp 1644511149
transform 1 0 16652 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0910_
timestamp 1644511149
transform 1 0 22264 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _0911_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21436 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0912_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21712 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0913_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0914_
timestamp 1644511149
transform 1 0 22080 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0915_
timestamp 1644511149
transform 1 0 22724 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0916_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22448 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0917_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23368 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0918_
timestamp 1644511149
transform 1 0 27876 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0919_
timestamp 1644511149
transform 1 0 23276 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0920_
timestamp 1644511149
transform 1 0 22908 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0921_
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0922_
timestamp 1644511149
transform 1 0 23368 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0923_
timestamp 1644511149
transform 1 0 25116 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0924_
timestamp 1644511149
transform 1 0 25484 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0925_
timestamp 1644511149
transform 1 0 27784 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0926_
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0927_
timestamp 1644511149
transform 1 0 27876 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0928_
timestamp 1644511149
transform 1 0 26036 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0929_
timestamp 1644511149
transform 1 0 27876 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0930_
timestamp 1644511149
transform 1 0 26956 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0931_
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _0932_
timestamp 1644511149
transform 1 0 17112 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0933_
timestamp 1644511149
transform 1 0 26128 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0934_
timestamp 1644511149
transform 1 0 16836 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0935_
timestamp 1644511149
transform 1 0 15640 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0936_
timestamp 1644511149
transform 1 0 17940 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0937_
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0938_
timestamp 1644511149
transform 1 0 18124 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0939_
timestamp 1644511149
transform 1 0 20056 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0940_
timestamp 1644511149
transform 1 0 19688 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0941_
timestamp 1644511149
transform 1 0 20424 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0942_
timestamp 1644511149
transform 1 0 20056 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0943_
timestamp 1644511149
transform 1 0 20884 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0944_
timestamp 1644511149
transform 1 0 20056 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0945_
timestamp 1644511149
transform 1 0 27876 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0946_
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0947_
timestamp 1644511149
transform 1 0 13340 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0948_
timestamp 1644511149
transform 1 0 20148 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0949_
timestamp 1644511149
transform 1 0 20332 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0950_
timestamp 1644511149
transform 1 0 16652 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0951_
timestamp 1644511149
transform 1 0 22632 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0952_
timestamp 1644511149
transform 1 0 20792 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0953_
timestamp 1644511149
transform 1 0 20792 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0954_
timestamp 1644511149
transform 1 0 19228 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0955_
timestamp 1644511149
transform 1 0 21804 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0956_
timestamp 1644511149
transform 1 0 23000 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _0957_
timestamp 1644511149
transform 1 0 9844 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0958_
timestamp 1644511149
transform 1 0 27876 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0959_
timestamp 1644511149
transform 1 0 21988 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0960_
timestamp 1644511149
transform 1 0 27876 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0961_
timestamp 1644511149
transform 1 0 23092 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0962_
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0963_
timestamp 1644511149
transform 1 0 24380 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0964_
timestamp 1644511149
transform 1 0 25576 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0965_
timestamp 1644511149
transform 1 0 10028 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0966_
timestamp 1644511149
transform 1 0 24564 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0967_
timestamp 1644511149
transform 1 0 10120 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0968_
timestamp 1644511149
transform 1 0 25392 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0969_
timestamp 1644511149
transform 1 0 26956 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0970_
timestamp 1644511149
transform 1 0 10580 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0971_
timestamp 1644511149
transform 1 0 25392 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0972_
timestamp 1644511149
transform 1 0 27784 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0973_
timestamp 1644511149
transform 1 0 27876 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0974_
timestamp 1644511149
transform 1 0 10764 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0975_
timestamp 1644511149
transform 1 0 15824 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0976_
timestamp 1644511149
transform 1 0 26956 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0977_
timestamp 1644511149
transform 1 0 20424 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0978_
timestamp 1644511149
transform 1 0 20240 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0979_
timestamp 1644511149
transform 1 0 12604 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0980_
timestamp 1644511149
transform 1 0 22172 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0981_
timestamp 1644511149
transform 1 0 20792 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0982_
timestamp 1644511149
transform 1 0 20884 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0983_
timestamp 1644511149
transform 1 0 13064 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0984_
timestamp 1644511149
transform 1 0 21804 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0985_
timestamp 1644511149
transform 1 0 10764 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0986_
timestamp 1644511149
transform 1 0 23552 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0987_
timestamp 1644511149
transform 1 0 18400 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0988_
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0989_
timestamp 1644511149
transform 1 0 16008 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0990_
timestamp 1644511149
transform 1 0 27324 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__and4b_1  _0991_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21068 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0992_
timestamp 1644511149
transform 1 0 22080 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0993_
timestamp 1644511149
transform 1 0 14352 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0994_
timestamp 1644511149
transform 1 0 14444 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0995_
timestamp 1644511149
transform 1 0 12420 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _0996_
timestamp 1644511149
transform 1 0 21896 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0997_
timestamp 1644511149
transform 1 0 11776 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0998_
timestamp 1644511149
transform 1 0 20884 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0999_
timestamp 1644511149
transform 1 0 11960 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1000_
timestamp 1644511149
transform 1 0 21896 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1001_
timestamp 1644511149
transform 1 0 14260 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1002_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1003_
timestamp 1644511149
transform 1 0 21988 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1004_
timestamp 1644511149
transform 1 0 22172 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1005_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23000 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1006_
timestamp 1644511149
transform 1 0 25392 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1007_
timestamp 1644511149
transform 1 0 11960 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1008_
timestamp 1644511149
transform 1 0 23184 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1009_
timestamp 1644511149
transform 1 0 22908 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1010_
timestamp 1644511149
transform 1 0 11316 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1011_
timestamp 1644511149
transform 1 0 23184 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1012_
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1013_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23276 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1014_
timestamp 1644511149
transform 1 0 21804 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1015_
timestamp 1644511149
transform 1 0 23092 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1016_
timestamp 1644511149
transform 1 0 23644 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1017_
timestamp 1644511149
transform 1 0 24380 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1018_
timestamp 1644511149
transform 1 0 24012 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1019_
timestamp 1644511149
transform 1 0 24196 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1020_
timestamp 1644511149
transform 1 0 11868 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1021_
timestamp 1644511149
transform 1 0 24104 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1022_
timestamp 1644511149
transform 1 0 24380 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1023_
timestamp 1644511149
transform 1 0 24932 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1024_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25116 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1025_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1026_
timestamp 1644511149
transform 1 0 27692 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1027_
timestamp 1644511149
transform 1 0 14444 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1028_
timestamp 1644511149
transform 1 0 10764 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1029_
timestamp 1644511149
transform 1 0 20056 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1030_
timestamp 1644511149
transform 1 0 10672 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1031_
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1032_
timestamp 1644511149
transform 1 0 23276 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1033_
timestamp 1644511149
transform 1 0 24932 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1034_
timestamp 1644511149
transform 1 0 19596 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1035_
timestamp 1644511149
transform 1 0 24656 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1036_
timestamp 1644511149
transform 1 0 25944 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1037_
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1038_
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1039_
timestamp 1644511149
transform 1 0 13248 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1040_
timestamp 1644511149
transform 1 0 13708 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1041_
timestamp 1644511149
transform 1 0 14720 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1042_
timestamp 1644511149
transform 1 0 9936 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1043_
timestamp 1644511149
transform 1 0 11776 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1044_
timestamp 1644511149
transform 1 0 19228 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1045_
timestamp 1644511149
transform 1 0 9200 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1046_
timestamp 1644511149
transform 1 0 14812 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1047_
timestamp 1644511149
transform 1 0 14812 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1048_
timestamp 1644511149
transform 1 0 15732 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1049_
timestamp 1644511149
transform 1 0 10764 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1050_
timestamp 1644511149
transform 1 0 14996 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1051_
timestamp 1644511149
transform 1 0 13984 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1052_
timestamp 1644511149
transform 1 0 13800 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1053_
timestamp 1644511149
transform 1 0 13248 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1054_
timestamp 1644511149
transform 1 0 14720 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1055_
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__and4b_1  _1056_
timestamp 1644511149
transform 1 0 15364 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1057_
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1058_
timestamp 1644511149
transform 1 0 13248 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1059_
timestamp 1644511149
transform 1 0 13064 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1060_
timestamp 1644511149
transform 1 0 11316 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1061_
timestamp 1644511149
transform 1 0 15088 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1062_
timestamp 1644511149
transform 1 0 10764 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1063_
timestamp 1644511149
transform 1 0 15180 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1064_
timestamp 1644511149
transform 1 0 10120 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1065_
timestamp 1644511149
transform 1 0 16100 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1066_
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1067_
timestamp 1644511149
transform 1 0 15088 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1068_
timestamp 1644511149
transform 1 0 14812 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1069_
timestamp 1644511149
transform 1 0 15640 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1070_
timestamp 1644511149
transform 1 0 12696 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1071_
timestamp 1644511149
transform 1 0 14812 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1072_
timestamp 1644511149
transform 1 0 17480 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1073_
timestamp 1644511149
transform 1 0 14536 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1074_
timestamp 1644511149
transform 1 0 12420 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1075_
timestamp 1644511149
transform 1 0 14996 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1076_
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1077_
timestamp 1644511149
transform 1 0 15180 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1078_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15088 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1079_
timestamp 1644511149
transform 1 0 15180 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1080_
timestamp 1644511149
transform 1 0 14168 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1081_
timestamp 1644511149
transform 1 0 15088 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1082_
timestamp 1644511149
transform 1 0 16652 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1083_
timestamp 1644511149
transform 1 0 16744 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1084_
timestamp 1644511149
transform 1 0 13340 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1085_
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1086_
timestamp 1644511149
transform 1 0 16192 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1087_
timestamp 1644511149
transform 1 0 18124 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1088_
timestamp 1644511149
transform 1 0 17296 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1089_
timestamp 1644511149
transform 1 0 17940 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1090_
timestamp 1644511149
transform 1 0 12052 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _1091_
timestamp 1644511149
transform 1 0 18952 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1092_
timestamp 1644511149
transform 1 0 10672 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1093_
timestamp 1644511149
transform 1 0 15732 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1094_
timestamp 1644511149
transform 1 0 10764 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1095_
timestamp 1644511149
transform 1 0 17664 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1096_
timestamp 1644511149
transform 1 0 16928 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1097_
timestamp 1644511149
transform 1 0 17204 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1098_
timestamp 1644511149
transform 1 0 9476 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1099_
timestamp 1644511149
transform 1 0 18032 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1100_
timestamp 1644511149
transform 1 0 18216 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1101_
timestamp 1644511149
transform 1 0 17296 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1102_
timestamp 1644511149
transform 1 0 17940 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1103_
timestamp 1644511149
transform 1 0 11776 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _1104_
timestamp 1644511149
transform 1 0 18952 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1105_
timestamp 1644511149
transform 1 0 17296 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1106_
timestamp 1644511149
transform 1 0 9568 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1107_
timestamp 1644511149
transform 1 0 14904 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1108_
timestamp 1644511149
transform 1 0 9200 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1109_
timestamp 1644511149
transform 1 0 19688 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1110_
timestamp 1644511149
transform 1 0 21988 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1111_
timestamp 1644511149
transform 1 0 24564 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1112_
timestamp 1644511149
transform 1 0 9752 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1113_
timestamp 1644511149
transform 1 0 21528 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1114_
timestamp 1644511149
transform 1 0 27876 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1115_
timestamp 1644511149
transform 1 0 17388 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1116_
timestamp 1644511149
transform 1 0 17480 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1117_
timestamp 1644511149
transform 1 0 22908 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1118_
timestamp 1644511149
transform 1 0 27876 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__and4b_1  _1119_
timestamp 1644511149
transform 1 0 20608 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1120_
timestamp 1644511149
transform 1 0 23644 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1121_
timestamp 1644511149
transform 1 0 24380 0 1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1122_
timestamp 1644511149
transform 1 0 27324 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1123_
timestamp 1644511149
transform 1 0 10764 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1124_
timestamp 1644511149
transform 1 0 21804 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1125_
timestamp 1644511149
transform 1 0 10120 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1126_
timestamp 1644511149
transform 1 0 23092 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1127_
timestamp 1644511149
transform 1 0 9476 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1128_
timestamp 1644511149
transform 1 0 21804 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1129_
timestamp 1644511149
transform 1 0 21712 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1130_
timestamp 1644511149
transform 1 0 18216 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1131_
timestamp 1644511149
transform 1 0 22724 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1132_
timestamp 1644511149
transform 1 0 25484 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1133_
timestamp 1644511149
transform 1 0 9292 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1134_
timestamp 1644511149
transform 1 0 22724 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1135_
timestamp 1644511149
transform 1 0 22540 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1136_
timestamp 1644511149
transform 1 0 10120 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1137_
timestamp 1644511149
transform 1 0 23552 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1138_
timestamp 1644511149
transform 1 0 14904 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1139_
timestamp 1644511149
transform 1 0 24380 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1140_
timestamp 1644511149
transform 1 0 23368 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1141_
timestamp 1644511149
transform 1 0 23368 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1142_
timestamp 1644511149
transform 1 0 26956 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1143_
timestamp 1644511149
transform 1 0 22540 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1144_
timestamp 1644511149
transform 1 0 25484 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1145_
timestamp 1644511149
transform 1 0 9108 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1146_
timestamp 1644511149
transform 1 0 23460 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1147_
timestamp 1644511149
transform 1 0 22448 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1148_
timestamp 1644511149
transform 1 0 9568 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1149_
timestamp 1644511149
transform 1 0 24380 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1150_
timestamp 1644511149
transform 1 0 24380 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1151_
timestamp 1644511149
transform 1 0 25392 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1152_
timestamp 1644511149
transform 1 0 26956 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1153_
timestamp 1644511149
transform 1 0 26956 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1154_
timestamp 1644511149
transform 1 0 8924 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1155_
timestamp 1644511149
transform 1 0 27324 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1156_
timestamp 1644511149
transform 1 0 26956 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1157_
timestamp 1644511149
transform 1 0 9476 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1158_
timestamp 1644511149
transform 1 0 19228 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1159_
timestamp 1644511149
transform 1 0 9660 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1160_
timestamp 1644511149
transform 1 0 26956 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1161_
timestamp 1644511149
transform 1 0 25208 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1162_
timestamp 1644511149
transform 1 0 25484 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1163_
timestamp 1644511149
transform 1 0 8556 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1164_
timestamp 1644511149
transform 1 0 24472 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1165_
timestamp 1644511149
transform 1 0 26956 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1166_
timestamp 1644511149
transform 1 0 26956 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1167_
timestamp 1644511149
transform 1 0 26956 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1168_
timestamp 1644511149
transform 1 0 8188 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _1169_
timestamp 1644511149
transform 1 0 20792 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1170_
timestamp 1644511149
transform 1 0 10488 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1171_
timestamp 1644511149
transform 1 0 15824 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1172_
timestamp 1644511149
transform 1 0 9476 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1173_
timestamp 1644511149
transform 1 0 18308 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1174_
timestamp 1644511149
transform 1 0 9200 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1175_
timestamp 1644511149
transform 1 0 9292 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1176_
timestamp 1644511149
transform 1 0 16836 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1177_
timestamp 1644511149
transform 1 0 10120 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1178_
timestamp 1644511149
transform 1 0 18308 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1179_
timestamp 1644511149
transform 1 0 10672 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1180_
timestamp 1644511149
transform 1 0 18216 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1181_
timestamp 1644511149
transform 1 0 10120 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1182_
timestamp 1644511149
transform 1 0 19044 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1183_
timestamp 1644511149
transform 1 0 10120 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1184_
timestamp 1644511149
transform 1 0 19228 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1185_
timestamp 1644511149
transform 1 0 10028 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1186_
timestamp 1644511149
transform 1 0 9292 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1187_
timestamp 1644511149
transform 1 0 14812 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1188_
timestamp 1644511149
transform 1 0 9292 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1189_
timestamp 1644511149
transform 1 0 17480 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1190_
timestamp 1644511149
transform 1 0 9476 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1191_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17664 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1192_
timestamp 1644511149
transform 1 0 18308 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1193_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18216 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1194_
timestamp 1644511149
transform 1 0 17940 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1195_
timestamp 1644511149
transform 1 0 19504 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1196_
timestamp 1644511149
transform 1 0 18124 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1197_
timestamp 1644511149
transform 1 0 15916 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1198_
timestamp 1644511149
transform 1 0 8648 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1199_
timestamp 1644511149
transform 1 0 16652 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1200_
timestamp 1644511149
transform 1 0 9016 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1201_
timestamp 1644511149
transform 1 0 15732 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1202_
timestamp 1644511149
transform 1 0 8832 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1203_
timestamp 1644511149
transform 1 0 13892 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1204_
timestamp 1644511149
transform 1 0 8188 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1205_
timestamp 1644511149
transform 1 0 14076 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1206_
timestamp 1644511149
transform 1 0 7820 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1207_
timestamp 1644511149
transform 1 0 13248 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1208_
timestamp 1644511149
transform 1 0 8648 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1209_
timestamp 1644511149
transform 1 0 13156 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1210_
timestamp 1644511149
transform 1 0 8004 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1211_
timestamp 1644511149
transform 1 0 13064 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1212_
timestamp 1644511149
transform 1 0 8832 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1213_
timestamp 1644511149
transform 1 0 12328 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1214_
timestamp 1644511149
transform 1 0 8188 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1215_
timestamp 1644511149
transform 1 0 15824 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1216_
timestamp 1644511149
transform 1 0 16744 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1217_
timestamp 1644511149
transform 1 0 16652 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1218_
timestamp 1644511149
transform 1 0 15640 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1219_
timestamp 1644511149
transform 1 0 11500 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1220_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16836 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1221_
timestamp 1644511149
transform 1 0 10580 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1222_
timestamp 1644511149
transform 1 0 7544 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1223_
timestamp 1644511149
transform 1 0 12236 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1224_
timestamp 1644511149
transform 1 0 8188 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1225_
timestamp 1644511149
transform 1 0 11316 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1226_
timestamp 1644511149
transform 1 0 7544 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1227_
timestamp 1644511149
transform 1 0 8188 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1228_
timestamp 1644511149
transform 1 0 11960 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1229_
timestamp 1644511149
transform 1 0 8188 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1230_
timestamp 1644511149
transform 1 0 10580 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1231_
timestamp 1644511149
transform 1 0 8188 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1232_
timestamp 1644511149
transform 1 0 11868 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1233_
timestamp 1644511149
transform 1 0 9476 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1234_
timestamp 1644511149
transform 1 0 11316 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1235_
timestamp 1644511149
transform 1 0 10120 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1236_
timestamp 1644511149
transform 1 0 12696 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1237_
timestamp 1644511149
transform 1 0 9476 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1238_
timestamp 1644511149
transform 1 0 12604 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1239_
timestamp 1644511149
transform 1 0 11776 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1240_
timestamp 1644511149
transform 1 0 13064 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1241_
timestamp 1644511149
transform 1 0 13616 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1242_
timestamp 1644511149
transform 1 0 13064 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a41o_1  _1243_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 13064 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1244_
timestamp 1644511149
transform 1 0 12880 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1245_
timestamp 1644511149
transform 1 0 8924 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1246_
timestamp 1644511149
transform 1 0 8188 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1247_
timestamp 1644511149
transform 1 0 11960 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1248_
timestamp 1644511149
transform 1 0 7912 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1249_
timestamp 1644511149
transform 1 0 10580 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1250_
timestamp 1644511149
transform 1 0 7544 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1251_
timestamp 1644511149
transform 1 0 10580 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1252_
timestamp 1644511149
transform 1 0 8188 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1253_
timestamp 1644511149
transform 1 0 11960 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1254_
timestamp 1644511149
transform 1 0 8832 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1255_
timestamp 1644511149
transform 1 0 12420 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1256_
timestamp 1644511149
transform 1 0 8188 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1257_
timestamp 1644511149
transform 1 0 8188 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1258_
timestamp 1644511149
transform 1 0 14076 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1259_
timestamp 1644511149
transform 1 0 8188 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1260_
timestamp 1644511149
transform 1 0 14168 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1261_
timestamp 1644511149
transform 1 0 7544 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1262_
timestamp 1644511149
transform 1 0 14076 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1263_
timestamp 1644511149
transform 1 0 12788 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1264_
timestamp 1644511149
transform 1 0 13340 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1265_
timestamp 1644511149
transform 1 0 13064 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1266_
timestamp 1644511149
transform 1 0 10856 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1267_
timestamp 1644511149
transform 1 0 14076 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1268_
timestamp 1644511149
transform 1 0 10856 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1269_
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1270_
timestamp 1644511149
transform 1 0 13340 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1271_
timestamp 1644511149
transform 1 0 8188 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1272_
timestamp 1644511149
transform 1 0 14628 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1273_
timestamp 1644511149
transform 1 0 8188 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1274_
timestamp 1644511149
transform 1 0 16652 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1275_
timestamp 1644511149
transform 1 0 8004 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1276_
timestamp 1644511149
transform 1 0 15272 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1277_
timestamp 1644511149
transform 1 0 15732 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1278_
timestamp 1644511149
transform 1 0 8280 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1279_
timestamp 1644511149
transform 1 0 17848 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1280_
timestamp 1644511149
transform 1 0 9016 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1281_
timestamp 1644511149
transform 1 0 19228 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1282_
timestamp 1644511149
transform 1 0 8096 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1283_
timestamp 1644511149
transform 1 0 16652 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1284_
timestamp 1644511149
transform 1 0 7544 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1285_
timestamp 1644511149
transform 1 0 19228 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1286_
timestamp 1644511149
transform 1 0 15456 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1287_
timestamp 1644511149
transform 1 0 15272 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1288_
timestamp 1644511149
transform 1 0 18216 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1289_
timestamp 1644511149
transform 1 0 17940 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1290_
timestamp 1644511149
transform 1 0 18124 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1291_
timestamp 1644511149
transform 1 0 10672 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1292_
timestamp 1644511149
transform 1 0 6900 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1293_
timestamp 1644511149
transform 1 0 11132 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1294_
timestamp 1644511149
transform 1 0 7544 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1295_
timestamp 1644511149
transform 1 0 7176 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1296_
timestamp 1644511149
transform 1 0 10304 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1297_
timestamp 1644511149
transform 1 0 7544 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1298_
timestamp 1644511149
transform 1 0 19780 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1299_
timestamp 1644511149
transform 1 0 6900 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1300_
timestamp 1644511149
transform 1 0 10120 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1301_
timestamp 1644511149
transform 1 0 7268 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1302_
timestamp 1644511149
transform 1 0 10028 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1303_
timestamp 1644511149
transform 1 0 6532 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1304_
timestamp 1644511149
transform 1 0 9752 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1305_
timestamp 1644511149
transform 1 0 6716 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1306_
timestamp 1644511149
transform 1 0 9844 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1307_
timestamp 1644511149
transform 1 0 7728 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1308_
timestamp 1644511149
transform 1 0 19780 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1309_
timestamp 1644511149
transform 1 0 18124 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1310_
timestamp 1644511149
transform 1 0 18216 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1311_
timestamp 1644511149
transform 1 0 19688 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1312_
timestamp 1644511149
transform 1 0 20608 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1313_
timestamp 1644511149
transform 1 0 20148 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1314_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21252 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1315_
timestamp 1644511149
transform 1 0 20976 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1316_
timestamp 1644511149
transform 1 0 21804 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1317_
timestamp 1644511149
transform 1 0 23644 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1318_
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1319_
timestamp 1644511149
transform 1 0 24472 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1320_
timestamp 1644511149
transform 1 0 25024 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1321_
timestamp 1644511149
transform 1 0 25024 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1322_
timestamp 1644511149
transform 1 0 16652 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1323_
timestamp 1644511149
transform 1 0 15824 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1324_
timestamp 1644511149
transform 1 0 17940 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1325_
timestamp 1644511149
transform 1 0 19780 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1326_
timestamp 1644511149
transform 1 0 19780 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1327_
timestamp 1644511149
transform 1 0 19412 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1328_
timestamp 1644511149
transform 1 0 20608 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1329_
timestamp 1644511149
transform 1 0 19964 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1330_
timestamp 1644511149
transform 1 0 21712 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1331_
timestamp 1644511149
transform 1 0 21804 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1332_
timestamp 1644511149
transform 1 0 22448 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1333_
timestamp 1644511149
transform 1 0 24380 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1334_
timestamp 1644511149
transform 1 0 24288 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1335_
timestamp 1644511149
transform 1 0 24472 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1336_
timestamp 1644511149
transform 1 0 25024 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1337_
timestamp 1644511149
transform 1 0 24472 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1338_
timestamp 1644511149
transform 1 0 19964 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1339_
timestamp 1644511149
transform 1 0 21712 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1340_
timestamp 1644511149
transform 1 0 21160 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1341_
timestamp 1644511149
transform 1 0 22724 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1342_
timestamp 1644511149
transform 1 0 23552 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1343_
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1344_
timestamp 1644511149
transform 1 0 25024 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1345_
timestamp 1644511149
transform 1 0 25024 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1346_
timestamp 1644511149
transform 1 0 25024 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1347_
timestamp 1644511149
transform 1 0 13524 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1348_
timestamp 1644511149
transform 1 0 19688 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1349_
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1350_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16008 0 1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1351_
timestamp 1644511149
transform 1 0 13340 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1352_
timestamp 1644511149
transform 1 0 14260 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1353_
timestamp 1644511149
transform 1 0 16284 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1354_
timestamp 1644511149
transform 1 0 18308 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1355_
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1356_
timestamp 1644511149
transform 1 0 18584 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1357_
timestamp 1644511149
transform 1 0 19320 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1358_
timestamp 1644511149
transform 1 0 14168 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1359_
timestamp 1644511149
transform 1 0 21804 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1360_
timestamp 1644511149
transform 1 0 21252 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1361_
timestamp 1644511149
transform 1 0 22448 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1362_
timestamp 1644511149
transform 1 0 23644 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1363_
timestamp 1644511149
transform 1 0 24380 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1364_
timestamp 1644511149
transform 1 0 25024 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1365_
timestamp 1644511149
transform 1 0 24472 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1366_
timestamp 1644511149
transform 1 0 25024 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1367_
timestamp 1644511149
transform 1 0 17388 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1368_
timestamp 1644511149
transform 1 0 18952 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1369_
timestamp 1644511149
transform 1 0 17112 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1370_
timestamp 1644511149
transform 1 0 18492 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1371_
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1372_
timestamp 1644511149
transform 1 0 16376 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1373_
timestamp 1644511149
transform 1 0 15732 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1374_
timestamp 1644511149
transform 1 0 16284 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1375_
timestamp 1644511149
transform 1 0 19872 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1376_
timestamp 1644511149
transform 1 0 19320 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1377_
timestamp 1644511149
transform 1 0 15640 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1378_
timestamp 1644511149
transform 1 0 15548 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1379_
timestamp 1644511149
transform 1 0 15640 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1380_
timestamp 1644511149
transform 1 0 16192 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1381_
timestamp 1644511149
transform 1 0 14720 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1382_
timestamp 1644511149
transform 1 0 13984 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1383_
timestamp 1644511149
transform 1 0 14720 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1384_
timestamp 1644511149
transform 1 0 16560 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1385_
timestamp 1644511149
transform 1 0 17112 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1386_
timestamp 1644511149
transform 1 0 11500 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1387_
timestamp 1644511149
transform 1 0 12144 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1388_
timestamp 1644511149
transform 1 0 12512 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1389_
timestamp 1644511149
transform 1 0 11224 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1390_
timestamp 1644511149
transform 1 0 11224 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1391_
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1392_
timestamp 1644511149
transform 1 0 11408 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1393_
timestamp 1644511149
transform 1 0 12144 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1394_
timestamp 1644511149
transform 1 0 14076 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1395_
timestamp 1644511149
transform 1 0 11776 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1396_
timestamp 1644511149
transform 1 0 11500 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1397_
timestamp 1644511149
transform 1 0 11684 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1398_
timestamp 1644511149
transform 1 0 10948 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1399_
timestamp 1644511149
transform 1 0 11500 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1400_
timestamp 1644511149
transform 1 0 13340 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1401_
timestamp 1644511149
transform 1 0 13432 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1402_
timestamp 1644511149
transform 1 0 14260 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1403_
timestamp 1644511149
transform 1 0 14076 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1404_
timestamp 1644511149
transform 1 0 11776 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1405_
timestamp 1644511149
transform 1 0 13616 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1406_
timestamp 1644511149
transform 1 0 14076 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1407_
timestamp 1644511149
transform 1 0 14536 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1408_
timestamp 1644511149
transform 1 0 16376 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1409_
timestamp 1644511149
transform 1 0 16652 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1410_
timestamp 1644511149
transform 1 0 18492 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1411_
timestamp 1644511149
transform 1 0 16744 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1412_
timestamp 1644511149
transform 1 0 17480 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1413_
timestamp 1644511149
transform 1 0 20700 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1414_
timestamp 1644511149
transform 1 0 17204 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1415_
timestamp 1644511149
transform 1 0 18308 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1416_
timestamp 1644511149
transform 1 0 19228 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1417_
timestamp 1644511149
transform 1 0 18216 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1418_
timestamp 1644511149
transform 1 0 17664 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1419_
timestamp 1644511149
transform 1 0 18952 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1420_
timestamp 1644511149
transform 1 0 19872 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1421_
timestamp 1644511149
transform 1 0 19780 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1422__9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6992 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1423__10
timestamp 1644511149
transform 1 0 1564 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1424__11
timestamp 1644511149
transform 1 0 14260 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1425__12
timestamp 1644511149
transform 1 0 4416 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1426__13
timestamp 1644511149
transform 1 0 25760 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1427__14
timestamp 1644511149
transform 1 0 4324 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1428__15
timestamp 1644511149
transform 1 0 27876 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1429__16
timestamp 1644511149
transform 1 0 4968 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1430__17
timestamp 1644511149
transform 1 0 7544 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1431__18
timestamp 1644511149
transform 1 0 10120 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1432__19
timestamp 1644511149
transform 1 0 27876 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1433__20
timestamp 1644511149
transform 1 0 15640 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1434__21
timestamp 1644511149
transform 1 0 9108 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1435__22
timestamp 1644511149
transform 1 0 1472 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1436__23
timestamp 1644511149
transform 1 0 9476 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1437__24
timestamp 1644511149
transform 1 0 6532 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1438__25
timestamp 1644511149
transform 1 0 24288 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1439__26
timestamp 1644511149
transform 1 0 6072 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1440__27
timestamp 1644511149
transform 1 0 6348 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1441__28
timestamp 1644511149
transform 1 0 10028 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1442__29
timestamp 1644511149
transform 1 0 3128 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1443__30
timestamp 1644511149
transform 1 0 7636 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1444__31
timestamp 1644511149
transform 1 0 8464 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1445__32
timestamp 1644511149
transform 1 0 9016 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1446__33
timestamp 1644511149
transform 1 0 27232 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1447__34
timestamp 1644511149
transform 1 0 6072 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1448__35
timestamp 1644511149
transform 1 0 27140 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1449__36
timestamp 1644511149
transform 1 0 3036 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1450__37
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1451__38
timestamp 1644511149
transform 1 0 4416 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1452__39
timestamp 1644511149
transform 1 0 26220 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1453__40
timestamp 1644511149
transform 1 0 7820 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1454__41
timestamp 1644511149
transform 1 0 6900 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1455__42
timestamp 1644511149
transform 1 0 8188 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1456__43
timestamp 1644511149
transform 1 0 5060 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1457__44
timestamp 1644511149
transform 1 0 2208 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1458__45
timestamp 1644511149
transform 1 0 9476 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1459__46
timestamp 1644511149
transform 1 0 8188 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1460__47
timestamp 1644511149
transform 1 0 7452 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1461__48
timestamp 1644511149
transform 1 0 2208 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1462__49
timestamp 1644511149
transform 1 0 12328 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1463__50
timestamp 1644511149
transform 1 0 3036 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1464__51
timestamp 1644511149
transform 1 0 9384 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1465__52
timestamp 1644511149
transform 1 0 5612 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1466__53
timestamp 1644511149
transform 1 0 5704 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1467__54
timestamp 1644511149
transform 1 0 23644 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1468__55
timestamp 1644511149
transform 1 0 7544 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1469__56
timestamp 1644511149
transform 1 0 27048 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1470__57
timestamp 1644511149
transform 1 0 2300 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1471__58
timestamp 1644511149
transform 1 0 7176 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1472__59
timestamp 1644511149
transform 1 0 1380 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1473__60
timestamp 1644511149
transform 1 0 21436 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1474__61
timestamp 1644511149
transform 1 0 25024 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1475__62
timestamp 1644511149
transform 1 0 18492 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1476__63
timestamp 1644511149
transform 1 0 7544 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1477__64
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1478__65
timestamp 1644511149
transform 1 0 6900 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1479__66
timestamp 1644511149
transform 1 0 11684 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1480__67
timestamp 1644511149
transform 1 0 27048 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1481__68
timestamp 1644511149
transform 1 0 6348 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1482__69
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1483__70
timestamp 1644511149
transform 1 0 3956 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1484__71
timestamp 1644511149
transform 1 0 27232 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1485__72
timestamp 1644511149
transform 1 0 7360 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1486__73
timestamp 1644511149
transform 1 0 7544 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1487__74
timestamp 1644511149
transform 1 0 5520 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1488__75
timestamp 1644511149
transform 1 0 7544 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1489__76
timestamp 1644511149
transform 1 0 20608 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1490__77
timestamp 1644511149
transform 1 0 25668 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1491__78
timestamp 1644511149
transform 1 0 6900 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1492__79
timestamp 1644511149
transform 1 0 17756 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1493__80
timestamp 1644511149
transform 1 0 27692 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1494__81
timestamp 1644511149
transform 1 0 1748 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1495__82
timestamp 1644511149
transform 1 0 23644 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1496__83
timestamp 1644511149
transform 1 0 4416 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1497__84
timestamp 1644511149
transform 1 0 6992 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1498__85
timestamp 1644511149
transform 1 0 7912 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1499__86
timestamp 1644511149
transform 1 0 2208 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1500__87
timestamp 1644511149
transform 1 0 8832 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1501__88
timestamp 1644511149
transform 1 0 22264 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1502__89
timestamp 1644511149
transform 1 0 25392 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1503__90
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1504__91
timestamp 1644511149
transform 1 0 5060 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1505__92
timestamp 1644511149
transform 1 0 27048 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1506__93
timestamp 1644511149
transform 1 0 10120 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1507__94
timestamp 1644511149
transform 1 0 6900 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1508__95
timestamp 1644511149
transform 1 0 6164 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1509__96
timestamp 1644511149
transform 1 0 11040 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1510__97
timestamp 1644511149
transform 1 0 3772 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1511__98
timestamp 1644511149
transform 1 0 4232 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1512__99
timestamp 1644511149
transform 1 0 6900 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1513__100
timestamp 1644511149
transform 1 0 6256 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1514__101
timestamp 1644511149
transform 1 0 25668 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1515__102
timestamp 1644511149
transform 1 0 6900 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1516__103
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1517__104
timestamp 1644511149
transform 1 0 23644 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1518__105
timestamp 1644511149
transform 1 0 7544 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1519__106
timestamp 1644511149
transform 1 0 4416 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1520__107
timestamp 1644511149
transform 1 0 22816 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1521__108
timestamp 1644511149
transform 1 0 1656 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1522__109
timestamp 1644511149
transform 1 0 25024 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1523__110
timestamp 1644511149
transform 1 0 5060 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1524__111
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1525__112
timestamp 1644511149
transform 1 0 2208 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1526__113
timestamp 1644511149
transform 1 0 2852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1527_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5336 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1528_
timestamp 1644511149
transform 1 0 1472 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1529_
timestamp 1644511149
transform 1 0 14168 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1530_
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1531_
timestamp 1644511149
transform 1 0 25116 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1532_
timestamp 1644511149
transform 1 0 2300 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1533_
timestamp 1644511149
transform 1 0 26312 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1534_
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1535_
timestamp 1644511149
transform 1 0 26312 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1536_
timestamp 1644511149
transform 1 0 26312 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1537_
timestamp 1644511149
transform 1 0 26312 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1538_
timestamp 1644511149
transform 1 0 15640 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1539_
timestamp 1644511149
transform 1 0 24564 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1540_
timestamp 1644511149
transform 1 0 1472 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1541_
timestamp 1644511149
transform 1 0 12972 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1542_
timestamp 1644511149
transform 1 0 6900 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1543_
timestamp 1644511149
transform 1 0 26312 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1544_
timestamp 1644511149
transform 1 0 26312 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1545_
timestamp 1644511149
transform 1 0 1380 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1546_
timestamp 1644511149
transform 1 0 26312 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1547_
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1548_
timestamp 1644511149
transform 1 0 26312 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1549_
timestamp 1644511149
transform 1 0 15548 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1550_
timestamp 1644511149
transform 1 0 9016 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1551_
timestamp 1644511149
transform 1 0 26312 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1552_
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1553_
timestamp 1644511149
transform 1 0 26312 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1554_
timestamp 1644511149
transform 1 0 1656 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1555_
timestamp 1644511149
transform 1 0 24564 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1556_
timestamp 1644511149
transform 1 0 3956 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1557_
timestamp 1644511149
transform 1 0 26312 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1558_
timestamp 1644511149
transform 1 0 26312 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1559_
timestamp 1644511149
transform 1 0 26312 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1560_
timestamp 1644511149
transform 1 0 17480 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1561_
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1562_
timestamp 1644511149
transform 1 0 1656 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1563_
timestamp 1644511149
transform 1 0 26312 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1564_
timestamp 1644511149
transform 1 0 10304 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1565_
timestamp 1644511149
transform 1 0 24564 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1566_
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1567_
timestamp 1644511149
transform 1 0 12972 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1568_
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1569_
timestamp 1644511149
transform 1 0 26312 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1570_
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1571_
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1572_
timestamp 1644511149
transform 1 0 23460 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1573_
timestamp 1644511149
transform 1 0 26312 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1574_
timestamp 1644511149
transform 1 0 20332 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1575_
timestamp 1644511149
transform 1 0 26312 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1576_
timestamp 1644511149
transform 1 0 24564 0 -1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1577_
timestamp 1644511149
transform 1 0 26312 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1578_
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1579_
timestamp 1644511149
transform 1 0 22264 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1580_
timestamp 1644511149
transform 1 0 1380 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1581_
timestamp 1644511149
transform 1 0 21896 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1582_
timestamp 1644511149
transform 1 0 26312 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1583_
timestamp 1644511149
transform 1 0 18860 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1584_
timestamp 1644511149
transform 1 0 20148 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1585_
timestamp 1644511149
transform 1 0 3680 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1586_
timestamp 1644511149
transform 1 0 21804 0 -1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1587_
timestamp 1644511149
transform 1 0 11684 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1588_
timestamp 1644511149
transform 1 0 26312 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1589_
timestamp 1644511149
transform 1 0 2024 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1590_
timestamp 1644511149
transform 1 0 1472 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1591_
timestamp 1644511149
transform 1 0 1380 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1592_
timestamp 1644511149
transform 1 0 26312 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1593_
timestamp 1644511149
transform 1 0 26312 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1594_
timestamp 1644511149
transform 1 0 26312 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1595_
timestamp 1644511149
transform 1 0 4692 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1596_
timestamp 1644511149
transform 1 0 24564 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1597_
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1598_
timestamp 1644511149
transform 1 0 26312 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1599_
timestamp 1644511149
transform 1 0 21988 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1600_
timestamp 1644511149
transform 1 0 17480 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1601_
timestamp 1644511149
transform 1 0 26312 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1602_
timestamp 1644511149
transform 1 0 1380 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1603_
timestamp 1644511149
transform 1 0 26312 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1604_
timestamp 1644511149
transform 1 0 3772 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1605_
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1606_
timestamp 1644511149
transform 1 0 7176 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1607_
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1608_
timestamp 1644511149
transform 1 0 26312 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1609_
timestamp 1644511149
transform 1 0 26312 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1610_
timestamp 1644511149
transform 1 0 24564 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1611_
timestamp 1644511149
transform 1 0 1932 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1612_
timestamp 1644511149
transform 1 0 3772 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1613_
timestamp 1644511149
transform 1 0 26312 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1614_
timestamp 1644511149
transform 1 0 9108 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1615_
timestamp 1644511149
transform 1 0 19412 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1616_
timestamp 1644511149
transform 1 0 3864 0 -1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1617_
timestamp 1644511149
transform 1 0 24564 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1618_
timestamp 1644511149
transform 1 0 1380 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1619_
timestamp 1644511149
transform 1 0 3404 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1620_
timestamp 1644511149
transform 1 0 11592 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1621_
timestamp 1644511149
transform 1 0 12328 0 -1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1622_
timestamp 1644511149
transform 1 0 24564 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1623_
timestamp 1644511149
transform 1 0 24564 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1624_
timestamp 1644511149
transform 1 0 14260 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1625_
timestamp 1644511149
transform 1 0 24564 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1626_
timestamp 1644511149
transform 1 0 26312 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1627_
timestamp 1644511149
transform 1 0 1564 0 -1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1628_
timestamp 1644511149
transform 1 0 21988 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1629_
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1630_
timestamp 1644511149
transform 1 0 24564 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1631_
timestamp 1644511149
transform 1 0 1472 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1632_
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1633_
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1634_
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19596 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_0_0_wb_clk_i
timestamp 1644511149
transform 1 0 12512 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 13248 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_2_0_wb_clk_i
timestamp 1644511149
transform 1 0 11500 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_3_0_wb_clk_i
timestamp 1644511149
transform 1 0 9844 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_0_0_wb_clk_i
timestamp 1644511149
transform 1 0 16192 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 13524 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_2_0_wb_clk_i
timestamp 1644511149
transform 1 0 23552 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_3_0_wb_clk_i
timestamp 1644511149
transform 1 0 13248 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_4_0_wb_clk_i
timestamp 1644511149
transform 1 0 10672 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_5_0_wb_clk_i
timestamp 1644511149
transform 1 0 12604 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_6_0_wb_clk_i
timestamp 1644511149
transform 1 0 9936 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_7_0_wb_clk_i
timestamp 1644511149
transform 1 0 11684 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input1
timestamp 1644511149
transform 1 0 1380 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1644511149
transform 1 0 6256 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1644511149
transform 1 0 4416 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1644511149
transform 1 0 5612 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1644511149
transform 1 0 17020 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1644511149
transform 1 0 6716 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1644511149
transform 1 0 27876 0 -1 11968
box -38 -48 406 592
<< labels >>
rlabel metal3 s 0 33268 800 33508 6 active
port 0 nsew signal input
rlabel metal2 s 10938 0 11050 800 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 14158 41200 14270 42000 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 0 35988 800 36228 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 29200 35988 30000 36228 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 16734 0 16846 800 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 7718 41200 7830 42000 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 29200 37348 30000 37588 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 29200 8788 30000 9028 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 1278 41200 1390 42000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 2566 41200 2678 42000 6 io_in[18]
port 10 nsew signal input
rlabel metal3 s 29200 628 30000 868 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 0 11508 800 11748 6 io_in[1]
port 12 nsew signal input
rlabel metal3 s 0 20348 800 20588 6 io_in[20]
port 13 nsew signal input
rlabel metal3 s 0 13548 800 13788 6 io_in[21]
port 14 nsew signal input
rlabel metal3 s 29200 17628 30000 17868 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 634 41200 746 42000 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s 0 40748 800 40988 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 27038 0 27150 800 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 26394 0 26506 800 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 29200 13548 30000 13788 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 23818 0 23930 800 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 29614 41200 29726 42000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 11582 0 11694 800 6 io_in[2]
port 23 nsew signal input
rlabel metal3 s 29200 20348 30000 20588 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 0 31908 800 32148 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 21886 0 21998 800 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 0 18308 800 18548 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 21242 41200 21354 42000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 25106 41200 25218 42000 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 29200 28508 30000 28748 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 25750 41200 25862 42000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 14802 41200 14914 42000 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 29200 27828 30000 28068 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 29200 40068 30000 40308 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 0 21708 800 21948 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 0 14908 800 15148 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 29200 29868 30000 30108 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s -10 41200 102 42000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 18666 0 18778 800 6 io_oeb[0]
port 39 nsew signal tristate
rlabel metal3 s 0 12188 800 12428 6 io_oeb[10]
port 40 nsew signal tristate
rlabel metal3 s 29200 26468 30000 26708 6 io_oeb[11]
port 41 nsew signal tristate
rlabel metal3 s 29200 16268 30000 16508 6 io_oeb[12]
port 42 nsew signal tristate
rlabel metal3 s 29200 15588 30000 15828 6 io_oeb[13]
port 43 nsew signal tristate
rlabel metal3 s 0 3348 800 3588 6 io_oeb[14]
port 44 nsew signal tristate
rlabel metal2 s 3854 41200 3966 42000 6 io_oeb[15]
port 45 nsew signal tristate
rlabel metal3 s 29200 7428 30000 7668 6 io_oeb[16]
port 46 nsew signal tristate
rlabel metal2 s 9650 0 9762 800 6 io_oeb[17]
port 47 nsew signal tristate
rlabel metal2 s 19954 41200 20066 42000 6 io_oeb[18]
port 48 nsew signal tristate
rlabel metal2 s 4498 41200 4610 42000 6 io_oeb[19]
port 49 nsew signal tristate
rlabel metal2 s 28326 0 28438 800 6 io_oeb[1]
port 50 nsew signal tristate
rlabel metal3 s 29200 21708 30000 21948 6 io_oeb[20]
port 51 nsew signal tristate
rlabel metal3 s 0 37348 800 37588 6 io_oeb[21]
port 52 nsew signal tristate
rlabel metal2 s 3854 0 3966 800 6 io_oeb[22]
port 53 nsew signal tristate
rlabel metal2 s 12226 41200 12338 42000 6 io_oeb[23]
port 54 nsew signal tristate
rlabel metal2 s 12870 41200 12982 42000 6 io_oeb[24]
port 55 nsew signal tristate
rlabel metal3 s 29200 4028 30000 4268 6 io_oeb[25]
port 56 nsew signal tristate
rlabel metal3 s 29200 33948 30000 34188 6 io_oeb[26]
port 57 nsew signal tristate
rlabel metal2 s 15446 41200 15558 42000 6 io_oeb[27]
port 58 nsew signal tristate
rlabel metal3 s 29200 -52 30000 188 6 io_oeb[28]
port 59 nsew signal tristate
rlabel metal3 s 29200 29188 30000 29428 6 io_oeb[29]
port 60 nsew signal tristate
rlabel metal2 s 23818 41200 23930 42000 6 io_oeb[2]
port 61 nsew signal tristate
rlabel metal3 s 0 38028 800 38268 6 io_oeb[30]
port 62 nsew signal tristate
rlabel metal2 s 29614 0 29726 800 6 io_oeb[31]
port 63 nsew signal tristate
rlabel metal3 s 0 17628 800 17868 6 io_oeb[32]
port 64 nsew signal tristate
rlabel metal3 s 29200 4708 30000 4948 6 io_oeb[33]
port 65 nsew signal tristate
rlabel metal2 s 1922 41200 2034 42000 6 io_oeb[34]
port 66 nsew signal tristate
rlabel metal3 s 0 15588 800 15828 6 io_oeb[35]
port 67 nsew signal tristate
rlabel metal3 s 0 8108 800 8348 6 io_oeb[36]
port 68 nsew signal tristate
rlabel metal3 s 0 12868 800 13108 6 io_oeb[37]
port 69 nsew signal tristate
rlabel metal2 s 18022 0 18134 800 6 io_oeb[3]
port 70 nsew signal tristate
rlabel metal3 s 29200 6068 30000 6308 6 io_oeb[4]
port 71 nsew signal tristate
rlabel metal3 s 0 23068 800 23308 6 io_oeb[5]
port 72 nsew signal tristate
rlabel metal3 s 29200 18988 30000 19228 6 io_oeb[6]
port 73 nsew signal tristate
rlabel metal2 s 3210 41200 3322 42000 6 io_oeb[7]
port 74 nsew signal tristate
rlabel metal2 s 3210 0 3322 800 6 io_oeb[8]
port 75 nsew signal tristate
rlabel metal2 s 7718 0 7830 800 6 io_oeb[9]
port 76 nsew signal tristate
rlabel metal3 s 29200 39388 30000 39628 6 io_out[0]
port 77 nsew signal tristate
rlabel metal3 s 29200 25788 30000 26028 6 io_out[10]
port 78 nsew signal tristate
rlabel metal3 s 0 1988 800 2228 6 io_out[11]
port 79 nsew signal tristate
rlabel metal3 s 0 5388 800 5628 6 io_out[12]
port 80 nsew signal tristate
rlabel metal2 s 28970 0 29082 800 6 io_out[13]
port 81 nsew signal tristate
rlabel metal3 s 29200 34628 30000 34868 6 io_out[14]
port 82 nsew signal tristate
rlabel metal3 s 0 29868 800 30108 6 io_out[15]
port 83 nsew signal tristate
rlabel metal3 s 29200 25108 30000 25348 6 io_out[16]
port 84 nsew signal tristate
rlabel metal2 s 27038 41200 27150 42000 6 io_out[17]
port 85 nsew signal tristate
rlabel metal3 s 29200 3348 30000 3588 6 io_out[18]
port 86 nsew signal tristate
rlabel metal3 s 0 16948 800 17188 6 io_out[19]
port 87 nsew signal tristate
rlabel metal2 s 18022 41200 18134 42000 6 io_out[1]
port 88 nsew signal tristate
rlabel metal2 s 23174 41200 23286 42000 6 io_out[20]
port 89 nsew signal tristate
rlabel metal3 s 0 29188 800 29428 6 io_out[21]
port 90 nsew signal tristate
rlabel metal2 s 22530 0 22642 800 6 io_out[22]
port 91 nsew signal tristate
rlabel metal3 s 29200 22388 30000 22628 6 io_out[23]
port 92 nsew signal tristate
rlabel metal2 s 19310 0 19422 800 6 io_out[24]
port 93 nsew signal tristate
rlabel metal2 s 20598 41200 20710 42000 6 io_out[25]
port 94 nsew signal tristate
rlabel metal3 s 0 4028 800 4268 6 io_out[26]
port 95 nsew signal tristate
rlabel metal2 s 21886 41200 21998 42000 6 io_out[27]
port 96 nsew signal tristate
rlabel metal2 s 12226 0 12338 800 6 io_out[28]
port 97 nsew signal tristate
rlabel metal3 s 29200 6748 30000 6988 6 io_out[29]
port 98 nsew signal tristate
rlabel metal2 s 5142 0 5254 800 6 io_out[2]
port 99 nsew signal tristate
rlabel metal3 s 0 4708 800 4948 6 io_out[30]
port 100 nsew signal tristate
rlabel metal3 s 0 10148 800 10388 6 io_out[31]
port 101 nsew signal tristate
rlabel metal3 s 0 33948 800 34188 6 io_out[32]
port 102 nsew signal tristate
rlabel metal3 s 29200 10828 30000 11068 6 io_out[33]
port 103 nsew signal tristate
rlabel metal3 s 29200 35308 30000 35548 6 io_out[34]
port 104 nsew signal tristate
rlabel metal3 s 29200 33268 30000 33508 6 io_out[35]
port 105 nsew signal tristate
rlabel metal2 s 5142 41200 5254 42000 6 io_out[36]
port 106 nsew signal tristate
rlabel metal3 s 29200 38028 30000 38268 6 io_out[37]
port 107 nsew signal tristate
rlabel metal3 s 0 31228 800 31468 6 io_out[3]
port 108 nsew signal tristate
rlabel metal3 s 29200 27148 30000 27388 6 io_out[4]
port 109 nsew signal tristate
rlabel metal2 s 10938 41200 11050 42000 6 io_out[5]
port 110 nsew signal tristate
rlabel metal2 s 28326 41200 28438 42000 6 io_out[6]
port 111 nsew signal tristate
rlabel metal3 s 0 14228 800 14468 6 io_out[7]
port 112 nsew signal tristate
rlabel metal2 s 13514 0 13626 800 6 io_out[8]
port 113 nsew signal tristate
rlabel metal3 s 0 10828 800 11068 6 io_out[9]
port 114 nsew signal tristate
rlabel metal3 s 29200 11508 30000 11748 6 la1_data_in[0]
port 115 nsew signal input
rlabel metal2 s 15446 0 15558 800 6 la1_data_in[10]
port 116 nsew signal input
rlabel metal3 s 29200 10148 30000 10388 6 la1_data_in[11]
port 117 nsew signal input
rlabel metal3 s 0 27148 800 27388 6 la1_data_in[12]
port 118 nsew signal input
rlabel metal2 s 24462 0 24574 800 6 la1_data_in[13]
port 119 nsew signal input
rlabel metal3 s 0 9468 800 9708 6 la1_data_in[14]
port 120 nsew signal input
rlabel metal2 s 5786 41200 5898 42000 6 la1_data_in[15]
port 121 nsew signal input
rlabel metal2 s 16734 41200 16846 42000 6 la1_data_in[16]
port 122 nsew signal input
rlabel metal2 s 11582 41200 11694 42000 6 la1_data_in[17]
port 123 nsew signal input
rlabel metal3 s 29200 1308 30000 1548 6 la1_data_in[18]
port 124 nsew signal input
rlabel metal2 s 7074 41200 7186 42000 6 la1_data_in[19]
port 125 nsew signal input
rlabel metal2 s 14158 0 14270 800 6 la1_data_in[1]
port 126 nsew signal input
rlabel metal3 s 0 26468 800 26708 6 la1_data_in[20]
port 127 nsew signal input
rlabel metal2 s 28970 41200 29082 42000 6 la1_data_in[21]
port 128 nsew signal input
rlabel metal3 s 29200 12188 30000 12428 6 la1_data_in[22]
port 129 nsew signal input
rlabel metal3 s 0 628 800 868 6 la1_data_in[23]
port 130 nsew signal input
rlabel metal2 s 10294 0 10406 800 6 la1_data_in[24]
port 131 nsew signal input
rlabel metal3 s 0 27828 800 28068 6 la1_data_in[25]
port 132 nsew signal input
rlabel metal3 s 29200 8108 30000 8348 6 la1_data_in[26]
port 133 nsew signal input
rlabel metal2 s 20598 0 20710 800 6 la1_data_in[27]
port 134 nsew signal input
rlabel metal3 s 0 23748 800 23988 6 la1_data_in[28]
port 135 nsew signal input
rlabel metal3 s 0 36668 800 36908 6 la1_data_in[29]
port 136 nsew signal input
rlabel metal2 s 8362 0 8474 800 6 la1_data_in[2]
port 137 nsew signal input
rlabel metal2 s 1278 0 1390 800 6 la1_data_in[30]
port 138 nsew signal input
rlabel metal2 s 27682 0 27794 800 6 la1_data_in[31]
port 139 nsew signal input
rlabel metal3 s 0 22388 800 22628 6 la1_data_in[3]
port 140 nsew signal input
rlabel metal2 s 24462 41200 24574 42000 6 la1_data_in[4]
port 141 nsew signal input
rlabel metal3 s 29200 23748 30000 23988 6 la1_data_in[5]
port 142 nsew signal input
rlabel metal2 s 8362 41200 8474 42000 6 la1_data_in[6]
port 143 nsew signal input
rlabel metal3 s 0 16268 800 16508 6 la1_data_in[7]
port 144 nsew signal input
rlabel metal2 s 9006 41200 9118 42000 6 la1_data_in[8]
port 145 nsew signal input
rlabel metal3 s 0 25108 800 25348 6 la1_data_in[9]
port 146 nsew signal input
rlabel metal2 s 5786 0 5898 800 6 la1_data_out[0]
port 147 nsew signal tristate
rlabel metal3 s 29200 14228 30000 14468 6 la1_data_out[10]
port 148 nsew signal tristate
rlabel metal2 s 16090 0 16202 800 6 la1_data_out[11]
port 149 nsew signal tristate
rlabel metal3 s 29200 38708 30000 38948 6 la1_data_out[12]
port 150 nsew signal tristate
rlabel metal3 s 0 39388 800 39628 6 la1_data_out[13]
port 151 nsew signal tristate
rlabel metal2 s 13514 41200 13626 42000 6 la1_data_out[14]
port 152 nsew signal tristate
rlabel metal3 s 0 1308 800 1548 6 la1_data_out[15]
port 153 nsew signal tristate
rlabel metal3 s 29200 18308 30000 18548 6 la1_data_out[16]
port 154 nsew signal tristate
rlabel metal3 s 29200 31908 30000 32148 6 la1_data_out[17]
port 155 nsew signal tristate
rlabel metal3 s 0 40068 800 40308 6 la1_data_out[18]
port 156 nsew signal tristate
rlabel metal3 s 29200 24428 30000 24668 6 la1_data_out[19]
port 157 nsew signal tristate
rlabel metal3 s 0 32588 800 32828 6 la1_data_out[1]
port 158 nsew signal tristate
rlabel metal3 s 0 7428 800 7668 6 la1_data_out[20]
port 159 nsew signal tristate
rlabel metal3 s 29200 36668 30000 36908 6 la1_data_out[21]
port 160 nsew signal tristate
rlabel metal2 s 16090 41200 16202 42000 6 la1_data_out[22]
port 161 nsew signal tristate
rlabel metal2 s 9006 0 9118 800 6 la1_data_out[23]
port 162 nsew signal tristate
rlabel metal3 s 29200 19668 30000 19908 6 la1_data_out[24]
port 163 nsew signal tristate
rlabel metal3 s 0 2668 800 2908 6 la1_data_out[25]
port 164 nsew signal tristate
rlabel metal3 s 29200 9468 30000 9708 6 la1_data_out[26]
port 165 nsew signal tristate
rlabel metal3 s 0 34628 800 34868 6 la1_data_out[27]
port 166 nsew signal tristate
rlabel metal3 s 29200 1988 30000 2228 6 la1_data_out[28]
port 167 nsew signal tristate
rlabel metal2 s 4498 0 4610 800 6 la1_data_out[29]
port 168 nsew signal tristate
rlabel metal2 s 14802 0 14914 800 6 la1_data_out[2]
port 169 nsew signal tristate
rlabel metal3 s 29200 14908 30000 15148 6 la1_data_out[30]
port 170 nsew signal tristate
rlabel metal3 s 29200 40748 30000 40988 6 la1_data_out[31]
port 171 nsew signal tristate
rlabel metal3 s 0 6748 800 6988 6 la1_data_out[3]
port 172 nsew signal tristate
rlabel metal3 s 29200 2668 30000 2908 6 la1_data_out[4]
port 173 nsew signal tristate
rlabel metal2 s 2566 0 2678 800 6 la1_data_out[5]
port 174 nsew signal tristate
rlabel metal3 s 29200 21028 30000 21268 6 la1_data_out[6]
port 175 nsew signal tristate
rlabel metal2 s 634 0 746 800 6 la1_data_out[7]
port 176 nsew signal tristate
rlabel metal3 s 29200 32588 30000 32828 6 la1_data_out[8]
port 177 nsew signal tristate
rlabel metal2 s 27682 41200 27794 42000 6 la1_data_out[9]
port 178 nsew signal tristate
rlabel metal3 s 29200 5388 30000 5628 6 la1_oenb[0]
port 179 nsew signal input
rlabel metal2 s 26394 41200 26506 42000 6 la1_oenb[10]
port 180 nsew signal input
rlabel metal3 s 0 19668 800 19908 6 la1_oenb[11]
port 181 nsew signal input
rlabel metal3 s 0 21028 800 21268 6 la1_oenb[12]
port 182 nsew signal input
rlabel metal2 s 21242 0 21354 800 6 la1_oenb[13]
port 183 nsew signal input
rlabel metal2 s -10 0 102 800 6 la1_oenb[14]
port 184 nsew signal input
rlabel metal2 s 25750 0 25862 800 6 la1_oenb[15]
port 185 nsew signal input
rlabel metal3 s 0 25788 800 26028 6 la1_oenb[16]
port 186 nsew signal input
rlabel metal3 s 0 38708 800 38948 6 la1_oenb[17]
port 187 nsew signal input
rlabel metal2 s 10294 41200 10406 42000 6 la1_oenb[18]
port 188 nsew signal input
rlabel metal3 s 0 18988 800 19228 6 la1_oenb[19]
port 189 nsew signal input
rlabel metal2 s 6430 0 6542 800 6 la1_oenb[1]
port 190 nsew signal input
rlabel metal2 s 1922 0 2034 800 6 la1_oenb[20]
port 191 nsew signal input
rlabel metal2 s 17378 41200 17490 42000 6 la1_oenb[21]
port 192 nsew signal input
rlabel metal2 s 9650 41200 9762 42000 6 la1_oenb[22]
port 193 nsew signal input
rlabel metal2 s 17378 0 17490 800 6 la1_oenb[23]
port 194 nsew signal input
rlabel metal2 s 22530 41200 22642 42000 6 la1_oenb[24]
port 195 nsew signal input
rlabel metal3 s 29200 12868 30000 13108 6 la1_oenb[25]
port 196 nsew signal input
rlabel metal3 s 0 28508 800 28748 6 la1_oenb[26]
port 197 nsew signal input
rlabel metal3 s 29200 31228 30000 31468 6 la1_oenb[27]
port 198 nsew signal input
rlabel metal2 s 7074 0 7186 800 6 la1_oenb[28]
port 199 nsew signal input
rlabel metal2 s 12870 0 12982 800 6 la1_oenb[29]
port 200 nsew signal input
rlabel metal3 s 0 6068 800 6308 6 la1_oenb[2]
port 201 nsew signal input
rlabel metal3 s 29200 30548 30000 30788 6 la1_oenb[30]
port 202 nsew signal input
rlabel metal2 s 19954 0 20066 800 6 la1_oenb[31]
port 203 nsew signal input
rlabel metal2 s 19310 41200 19422 42000 6 la1_oenb[3]
port 204 nsew signal input
rlabel metal2 s 18666 41200 18778 42000 6 la1_oenb[4]
port 205 nsew signal input
rlabel metal3 s 0 35308 800 35548 6 la1_oenb[5]
port 206 nsew signal input
rlabel metal3 s 0 41428 800 41668 6 la1_oenb[6]
port 207 nsew signal input
rlabel metal2 s 25106 0 25218 800 6 la1_oenb[7]
port 208 nsew signal input
rlabel metal3 s 0 8788 800 9028 6 la1_oenb[8]
port 209 nsew signal input
rlabel metal3 s 0 30548 800 30788 6 la1_oenb[9]
port 210 nsew signal input
rlabel metal4 s 5576 2128 5896 39760 6 vccd1
port 211 nsew power input
rlabel metal4 s 14840 2128 15160 39760 6 vccd1
port 211 nsew power input
rlabel metal4 s 24104 2128 24424 39760 6 vccd1
port 211 nsew power input
rlabel metal4 s 10208 2128 10528 39760 6 vssd1
port 212 nsew ground input
rlabel metal4 s 19472 2128 19792 39760 6 vssd1
port 212 nsew ground input
rlabel metal3 s 29200 23068 30000 23308 6 wb_clk_i
port 213 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 30000 42000
<< end >>
