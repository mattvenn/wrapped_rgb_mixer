VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_rgb_mixer
  CLASS BLOCK ;
  FOREIGN wrapped_rgb_mixer ;
  ORIGIN 0.000 0.000 ;
  SIZE 180.000 BY 210.000 ;
  PIN active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 179.940 4.000 181.140 ;
    END
  END active
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.910 1.000 58.470 4.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.330 206.000 93.890 209.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 193.540 4.000 194.740 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 179.940 179.000 181.140 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.110 1.000 90.670 4.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.910 206.000 58.470 209.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 186.740 179.000 187.940 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 30.340 179.000 31.540 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.710 206.000 26.270 209.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.150 206.000 32.710 209.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.390 1.000 167.950 4.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 60.940 4.000 62.140 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 111.940 4.000 113.140 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 74.540 4.000 75.740 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 77.940 179.000 79.140 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.490 206.000 23.050 209.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.610 206.000 10.170 209.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.850 1.000 145.410 4.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.630 1.000 142.190 4.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 57.540 179.000 58.740 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.750 1.000 129.310 4.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.050 206.000 177.610 209.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.350 1.000 64.910 4.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 91.540 179.000 92.740 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 173.140 4.000 174.340 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.090 1.000 119.650 4.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 101.740 4.000 102.940 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.970 206.000 132.530 209.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.510 206.000 155.070 209.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 135.740 179.000 136.940 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.730 206.000 158.290 209.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.550 206.000 97.110 209.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 132.340 179.000 133.540 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 200.340 179.000 201.540 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 118.740 4.000 119.940 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 81.340 4.000 82.540 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 145.940 179.000 147.140 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.050 206.000 16.610 209.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.990 1.000 103.550 4.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 67.740 4.000 68.940 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 125.540 179.000 126.740 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 71.140 179.000 72.340 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 67.740 179.000 68.940 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 16.740 4.000 17.940 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.590 206.000 39.150 209.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 23.540 179.000 24.740 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.470 1.000 52.030 4.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.530 206.000 126.090 209.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.810 206.000 42.370 209.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.290 1.000 151.850 4.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 98.340 179.000 99.540 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 203.740 4.000 204.940 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.270 1.000 19.830 4.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.450 206.000 81.010 209.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.890 206.000 87.450 209.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 3.140 179.000 4.340 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 166.340 179.000 167.540 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.770 206.000 100.330 209.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.170 1.000 164.730 4.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 139.140 179.000 140.340 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.850 206.000 145.410 209.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 207.140 4.000 208.340 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.950 1.000 161.510 4.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 94.940 4.000 96.140 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 9.940 179.000 11.140 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.930 206.000 29.490 209.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 84.740 4.000 85.940 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 43.940 4.000 45.140 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 71.140 4.000 72.340 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.770 1.000 100.330 4.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 16.740 179.000 17.940 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 125.540 4.000 126.740 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 84.740 179.000 85.940 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.370 206.000 35.930 209.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.050 1.000 16.610 4.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.810 1.000 42.370 4.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 196.940 179.000 198.140 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 122.140 179.000 123.340 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 9.940 4.000 11.140 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 26.940 4.000 28.140 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.510 1.000 155.070 4.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 169.740 179.000 170.940 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 159.540 4.000 160.740 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 118.740 179.000 119.940 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.170 206.000 164.730 209.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 -0.260 179.000 0.940 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 91.540 4.000 92.740 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.650 206.000 113.210 209.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.630 206.000 142.190 209.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 156.140 4.000 157.340 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.310 1.000 122.870 4.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 101.740 179.000 102.940 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.210 1.000 106.770 4.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.750 206.000 129.310 209.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 20.140 4.000 21.340 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.190 206.000 135.750 209.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.570 1.000 68.130 4.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 20.140 179.000 21.340 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.710 1.000 26.270 4.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 23.540 4.000 24.740 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 54.140 4.000 55.340 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 183.340 4.000 184.540 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 43.940 179.000 45.140 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 173.140 179.000 174.340 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 162.940 179.000 164.140 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.030 206.000 45.590 209.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 190.140 179.000 191.340 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 169.740 4.000 170.940 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 128.940 179.000 130.140 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.010 206.000 74.570 209.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.610 206.000 171.170 209.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 77.940 4.000 79.140 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.010 1.000 74.570 4.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 57.540 4.000 58.740 ;
    END
  END io_out[9]
  PIN la1_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 47.340 179.000 48.540 ;
    END
  END la1_data_in[0]
  PIN la1_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.670 1.000 84.230 4.000 ;
    END
  END la1_data_in[10]
  PIN la1_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 37.140 179.000 38.340 ;
    END
  END la1_data_in[11]
  PIN la1_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 145.940 4.000 147.140 ;
    END
  END la1_data_in[12]
  PIN la1_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.970 1.000 132.530 4.000 ;
    END
  END la1_data_in[13]
  PIN la1_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 50.740 4.000 51.940 ;
    END
  END la1_data_in[14]
  PIN la1_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.250 206.000 48.810 209.000 ;
    END
  END la1_data_in[15]
  PIN la1_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.210 206.000 106.770 209.000 ;
    END
  END la1_data_in[16]
  PIN la1_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.230 206.000 77.790 209.000 ;
    END
  END la1_data_in[17]
  PIN la1_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.610 1.000 171.170 4.000 ;
    END
  END la1_data_in[18]
  PIN la1_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.690 206.000 55.250 209.000 ;
    END
  END la1_data_in[19]
  PIN la1_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.230 1.000 77.790 4.000 ;
    END
  END la1_data_in[1]
  PIN la1_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 142.540 4.000 143.740 ;
    END
  END la1_data_in[20]
  PIN la1_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.830 206.000 174.390 209.000 ;
    END
  END la1_data_in[21]
  PIN la1_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 50.740 179.000 51.940 ;
    END
  END la1_data_in[22]
  PIN la1_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 3.140 4.000 4.340 ;
    END
  END la1_data_in[23]
  PIN la1_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.690 1.000 55.250 4.000 ;
    END
  END la1_data_in[24]
  PIN la1_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 149.340 4.000 150.540 ;
    END
  END la1_data_in[25]
  PIN la1_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 26.940 179.000 28.140 ;
    END
  END la1_data_in[26]
  PIN la1_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.650 1.000 113.210 4.000 ;
    END
  END la1_data_in[27]
  PIN la1_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 128.940 4.000 130.140 ;
    END
  END la1_data_in[28]
  PIN la1_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 196.940 4.000 198.140 ;
    END
  END la1_data_in[29]
  PIN la1_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.030 1.000 45.590 4.000 ;
    END
  END la1_data_in[2]
  PIN la1_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.390 1.000 6.950 4.000 ;
    END
  END la1_data_in[30]
  PIN la1_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.070 1.000 148.630 4.000 ;
    END
  END la1_data_in[31]
  PIN la1_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 122.140 4.000 123.340 ;
    END
  END la1_data_in[3]
  PIN la1_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.290 206.000 151.850 209.000 ;
    END
  END la1_data_in[4]
  PIN la1_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 111.940 179.000 113.140 ;
    END
  END la1_data_in[5]
  PIN la1_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.130 206.000 61.690 209.000 ;
    END
  END la1_data_in[6]
  PIN la1_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 88.140 4.000 89.340 ;
    END
  END la1_data_in[7]
  PIN la1_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.350 206.000 64.910 209.000 ;
    END
  END la1_data_in[8]
  PIN la1_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 135.740 4.000 136.940 ;
    END
  END la1_data_in[9]
  PIN la1_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.150 1.000 32.710 4.000 ;
    END
  END la1_data_out[0]
  PIN la1_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 60.940 179.000 62.140 ;
    END
  END la1_data_out[10]
  PIN la1_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.890 1.000 87.450 4.000 ;
    END
  END la1_data_out[11]
  PIN la1_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 193.540 179.000 194.740 ;
    END
  END la1_data_out[12]
  PIN la1_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.170 206.000 3.730 209.000 ;
    END
  END la1_data_out[13]
  PIN la1_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.110 206.000 90.670 209.000 ;
    END
  END la1_data_out[14]
  PIN la1_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 6.540 4.000 7.740 ;
    END
  END la1_data_out[15]
  PIN la1_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 81.340 179.000 82.540 ;
    END
  END la1_data_out[16]
  PIN la1_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 156.140 179.000 157.340 ;
    END
  END la1_data_out[17]
  PIN la1_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.390 206.000 6.950 209.000 ;
    END
  END la1_data_out[18]
  PIN la1_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 115.340 179.000 116.540 ;
    END
  END la1_data_out[19]
  PIN la1_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 176.540 4.000 177.740 ;
    END
  END la1_data_out[1]
  PIN la1_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 40.540 4.000 41.740 ;
    END
  END la1_data_out[20]
  PIN la1_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 183.340 179.000 184.540 ;
    END
  END la1_data_out[21]
  PIN la1_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.990 206.000 103.550 209.000 ;
    END
  END la1_data_out[22]
  PIN la1_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.250 1.000 48.810 4.000 ;
    END
  END la1_data_out[23]
  PIN la1_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 88.140 179.000 89.340 ;
    END
  END la1_data_out[24]
  PIN la1_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 13.340 4.000 14.540 ;
    END
  END la1_data_out[25]
  PIN la1_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 33.740 179.000 34.940 ;
    END
  END la1_data_out[26]
  PIN la1_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 186.740 4.000 187.940 ;
    END
  END la1_data_out[27]
  PIN la1_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.830 1.000 174.390 4.000 ;
    END
  END la1_data_out[28]
  PIN la1_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.490 1.000 23.050 4.000 ;
    END
  END la1_data_out[29]
  PIN la1_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.450 1.000 81.010 4.000 ;
    END
  END la1_data_out[2]
  PIN la1_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 64.340 179.000 65.540 ;
    END
  END la1_data_out[30]
  PIN la1_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 203.740 179.000 204.940 ;
    END
  END la1_data_out[31]
  PIN la1_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 37.140 4.000 38.340 ;
    END
  END la1_data_out[3]
  PIN la1_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.050 1.000 177.610 4.000 ;
    END
  END la1_data_out[4]
  PIN la1_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.830 1.000 13.390 4.000 ;
    END
  END la1_data_out[5]
  PIN la1_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 94.940 179.000 96.140 ;
    END
  END la1_data_out[6]
  PIN la1_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.170 1.000 3.730 4.000 ;
    END
  END la1_data_out[7]
  PIN la1_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 159.540 179.000 160.740 ;
    END
  END la1_data_out[8]
  PIN la1_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.390 206.000 167.950 209.000 ;
    END
  END la1_data_out[9]
  PIN la1_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 13.340 179.000 14.540 ;
    END
  END la1_oenb[0]
  PIN la1_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.950 206.000 161.510 209.000 ;
    END
  END la1_oenb[10]
  PIN la1_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 108.540 4.000 109.740 ;
    END
  END la1_oenb[11]
  PIN la1_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 115.340 4.000 116.540 ;
    END
  END la1_oenb[12]
  PIN la1_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.870 1.000 116.430 4.000 ;
    END
  END la1_oenb[13]
  PIN la1_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT -0.050 1.000 0.510 4.000 ;
    END
  END la1_oenb[14]
  PIN la1_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.410 1.000 138.970 4.000 ;
    END
  END la1_oenb[15]
  PIN la1_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 139.140 4.000 140.340 ;
    END
  END la1_oenb[16]
  PIN la1_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT -0.050 206.000 0.510 209.000 ;
    END
  END la1_oenb[17]
  PIN la1_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.790 206.000 71.350 209.000 ;
    END
  END la1_oenb[18]
  PIN la1_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 105.140 4.000 106.340 ;
    END
  END la1_oenb[19]
  PIN la1_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.370 1.000 35.930 4.000 ;
    END
  END la1_oenb[1]
  PIN la1_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.610 1.000 10.170 4.000 ;
    END
  END la1_oenb[20]
  PIN la1_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.430 206.000 109.990 209.000 ;
    END
  END la1_oenb[21]
  PIN la1_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.570 206.000 68.130 209.000 ;
    END
  END la1_oenb[22]
  PIN la1_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.550 1.000 97.110 4.000 ;
    END
  END la1_oenb[23]
  PIN la1_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.410 206.000 138.970 209.000 ;
    END
  END la1_oenb[24]
  PIN la1_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 54.140 179.000 55.340 ;
    END
  END la1_oenb[25]
  PIN la1_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 152.740 4.000 153.940 ;
    END
  END la1_oenb[26]
  PIN la1_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 152.740 179.000 153.940 ;
    END
  END la1_oenb[27]
  PIN la1_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.590 1.000 39.150 4.000 ;
    END
  END la1_oenb[28]
  PIN la1_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.790 1.000 71.350 4.000 ;
    END
  END la1_oenb[29]
  PIN la1_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 33.740 4.000 34.940 ;
    END
  END la1_oenb[2]
  PIN la1_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 149.340 179.000 150.540 ;
    END
  END la1_oenb[30]
  PIN la1_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.430 1.000 109.990 4.000 ;
    END
  END la1_oenb[31]
  PIN la1_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.310 206.000 122.870 209.000 ;
    END
  END la1_oenb[3]
  PIN la1_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.090 206.000 119.650 209.000 ;
    END
  END la1_oenb[4]
  PIN la1_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 190.140 4.000 191.340 ;
    END
  END la1_oenb[5]
  PIN la1_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.830 206.000 13.390 209.000 ;
    END
  END la1_oenb[6]
  PIN la1_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.190 1.000 135.750 4.000 ;
    END
  END la1_oenb[7]
  PIN la1_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 47.340 4.000 48.540 ;
    END
  END la1_oenb[8]
  PIN la1_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 162.940 4.000 164.140 ;
    END
  END la1_oenb[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 25.820 10.640 27.420 198.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 68.025 10.640 69.625 198.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 110.230 10.640 111.830 198.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 152.435 10.640 154.035 198.800 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 46.920 10.640 48.520 198.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 89.125 10.640 90.725 198.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 131.330 10.640 132.930 198.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 173.535 10.640 175.135 198.800 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 105.140 179.000 106.340 ;
    END
  END wb_clk_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 174.340 198.645 ;
      LAYER met1 ;
        RECT 3.290 5.480 179.790 200.220 ;
      LAYER met2 ;
        RECT 4.010 205.720 6.110 207.925 ;
        RECT 7.230 205.720 9.330 207.925 ;
        RECT 10.450 205.720 12.550 207.925 ;
        RECT 13.670 205.720 15.770 207.925 ;
        RECT 16.890 205.720 22.210 207.925 ;
        RECT 23.330 205.720 25.430 207.925 ;
        RECT 26.550 205.720 28.650 207.925 ;
        RECT 29.770 205.720 31.870 207.925 ;
        RECT 32.990 205.720 35.090 207.925 ;
        RECT 36.210 205.720 38.310 207.925 ;
        RECT 39.430 205.720 41.530 207.925 ;
        RECT 42.650 205.720 44.750 207.925 ;
        RECT 45.870 205.720 47.970 207.925 ;
        RECT 49.090 205.720 54.410 207.925 ;
        RECT 55.530 205.720 57.630 207.925 ;
        RECT 58.750 205.720 60.850 207.925 ;
        RECT 61.970 205.720 64.070 207.925 ;
        RECT 65.190 205.720 67.290 207.925 ;
        RECT 68.410 205.720 70.510 207.925 ;
        RECT 71.630 205.720 73.730 207.925 ;
        RECT 74.850 205.720 76.950 207.925 ;
        RECT 78.070 205.720 80.170 207.925 ;
        RECT 81.290 205.720 86.610 207.925 ;
        RECT 87.730 205.720 89.830 207.925 ;
        RECT 90.950 205.720 93.050 207.925 ;
        RECT 94.170 205.720 96.270 207.925 ;
        RECT 97.390 205.720 99.490 207.925 ;
        RECT 100.610 205.720 102.710 207.925 ;
        RECT 103.830 205.720 105.930 207.925 ;
        RECT 107.050 205.720 109.150 207.925 ;
        RECT 110.270 205.720 112.370 207.925 ;
        RECT 113.490 205.720 118.810 207.925 ;
        RECT 119.930 205.720 122.030 207.925 ;
        RECT 123.150 205.720 125.250 207.925 ;
        RECT 126.370 205.720 128.470 207.925 ;
        RECT 129.590 205.720 131.690 207.925 ;
        RECT 132.810 205.720 134.910 207.925 ;
        RECT 136.030 205.720 138.130 207.925 ;
        RECT 139.250 205.720 141.350 207.925 ;
        RECT 142.470 205.720 144.570 207.925 ;
        RECT 145.690 205.720 151.010 207.925 ;
        RECT 152.130 205.720 154.230 207.925 ;
        RECT 155.350 205.720 157.450 207.925 ;
        RECT 158.570 205.720 160.670 207.925 ;
        RECT 161.790 205.720 163.890 207.925 ;
        RECT 165.010 205.720 167.110 207.925 ;
        RECT 168.230 205.720 170.330 207.925 ;
        RECT 171.450 205.720 173.550 207.925 ;
        RECT 174.670 205.720 176.770 207.925 ;
        RECT 177.890 205.720 179.770 207.925 ;
        RECT 3.320 4.280 179.770 205.720 ;
        RECT 4.010 0.720 6.110 4.280 ;
        RECT 7.230 0.720 9.330 4.280 ;
        RECT 10.450 0.720 12.550 4.280 ;
        RECT 13.670 0.720 15.770 4.280 ;
        RECT 16.890 0.720 18.990 4.280 ;
        RECT 20.110 0.720 22.210 4.280 ;
        RECT 23.330 0.720 25.430 4.280 ;
        RECT 26.550 0.720 31.870 4.280 ;
        RECT 32.990 0.720 35.090 4.280 ;
        RECT 36.210 0.720 38.310 4.280 ;
        RECT 39.430 0.720 41.530 4.280 ;
        RECT 42.650 0.720 44.750 4.280 ;
        RECT 45.870 0.720 47.970 4.280 ;
        RECT 49.090 0.720 51.190 4.280 ;
        RECT 52.310 0.720 54.410 4.280 ;
        RECT 55.530 0.720 57.630 4.280 ;
        RECT 58.750 0.720 64.070 4.280 ;
        RECT 65.190 0.720 67.290 4.280 ;
        RECT 68.410 0.720 70.510 4.280 ;
        RECT 71.630 0.720 73.730 4.280 ;
        RECT 74.850 0.720 76.950 4.280 ;
        RECT 78.070 0.720 80.170 4.280 ;
        RECT 81.290 0.720 83.390 4.280 ;
        RECT 84.510 0.720 86.610 4.280 ;
        RECT 87.730 0.720 89.830 4.280 ;
        RECT 90.950 0.720 96.270 4.280 ;
        RECT 97.390 0.720 99.490 4.280 ;
        RECT 100.610 0.720 102.710 4.280 ;
        RECT 103.830 0.720 105.930 4.280 ;
        RECT 107.050 0.720 109.150 4.280 ;
        RECT 110.270 0.720 112.370 4.280 ;
        RECT 113.490 0.720 115.590 4.280 ;
        RECT 116.710 0.720 118.810 4.280 ;
        RECT 119.930 0.720 122.030 4.280 ;
        RECT 123.150 0.720 128.470 4.280 ;
        RECT 129.590 0.720 131.690 4.280 ;
        RECT 132.810 0.720 134.910 4.280 ;
        RECT 136.030 0.720 138.130 4.280 ;
        RECT 139.250 0.720 141.350 4.280 ;
        RECT 142.470 0.720 144.570 4.280 ;
        RECT 145.690 0.720 147.790 4.280 ;
        RECT 148.910 0.720 151.010 4.280 ;
        RECT 152.130 0.720 154.230 4.280 ;
        RECT 155.350 0.720 160.670 4.280 ;
        RECT 161.790 0.720 163.890 4.280 ;
        RECT 165.010 0.720 167.110 4.280 ;
        RECT 168.230 0.720 170.330 4.280 ;
        RECT 171.450 0.720 173.550 4.280 ;
        RECT 174.670 0.720 176.770 4.280 ;
        RECT 177.890 0.720 179.770 4.280 ;
        RECT 3.320 0.155 179.770 0.720 ;
      LAYER met3 ;
        RECT 4.400 206.740 179.795 207.905 ;
        RECT 4.000 205.340 179.795 206.740 ;
        RECT 4.400 203.340 175.600 205.340 ;
        RECT 179.400 203.340 179.795 205.340 ;
        RECT 4.000 201.940 179.795 203.340 ;
        RECT 4.000 199.940 175.600 201.940 ;
        RECT 179.400 199.940 179.795 201.940 ;
        RECT 4.000 198.540 179.795 199.940 ;
        RECT 4.400 196.540 175.600 198.540 ;
        RECT 179.400 196.540 179.795 198.540 ;
        RECT 4.000 195.140 179.795 196.540 ;
        RECT 4.400 193.140 175.600 195.140 ;
        RECT 179.400 193.140 179.795 195.140 ;
        RECT 4.000 191.740 179.795 193.140 ;
        RECT 4.400 189.740 175.600 191.740 ;
        RECT 179.400 189.740 179.795 191.740 ;
        RECT 4.000 188.340 179.795 189.740 ;
        RECT 4.400 186.340 175.600 188.340 ;
        RECT 179.400 186.340 179.795 188.340 ;
        RECT 4.000 184.940 179.795 186.340 ;
        RECT 4.400 182.940 175.600 184.940 ;
        RECT 179.400 182.940 179.795 184.940 ;
        RECT 4.000 181.540 179.795 182.940 ;
        RECT 4.400 179.540 175.600 181.540 ;
        RECT 179.400 179.540 179.795 181.540 ;
        RECT 4.000 178.140 179.795 179.540 ;
        RECT 4.400 176.140 179.795 178.140 ;
        RECT 4.000 174.740 179.795 176.140 ;
        RECT 4.400 172.740 175.600 174.740 ;
        RECT 179.400 172.740 179.795 174.740 ;
        RECT 4.000 171.340 179.795 172.740 ;
        RECT 4.400 169.340 175.600 171.340 ;
        RECT 179.400 169.340 179.795 171.340 ;
        RECT 4.000 167.940 179.795 169.340 ;
        RECT 4.000 165.940 175.600 167.940 ;
        RECT 179.400 165.940 179.795 167.940 ;
        RECT 4.000 164.540 179.795 165.940 ;
        RECT 4.400 162.540 175.600 164.540 ;
        RECT 179.400 162.540 179.795 164.540 ;
        RECT 4.000 161.140 179.795 162.540 ;
        RECT 4.400 159.140 175.600 161.140 ;
        RECT 179.400 159.140 179.795 161.140 ;
        RECT 4.000 157.740 179.795 159.140 ;
        RECT 4.400 155.740 175.600 157.740 ;
        RECT 179.400 155.740 179.795 157.740 ;
        RECT 4.000 154.340 179.795 155.740 ;
        RECT 4.400 152.340 175.600 154.340 ;
        RECT 179.400 152.340 179.795 154.340 ;
        RECT 4.000 150.940 179.795 152.340 ;
        RECT 4.400 148.940 175.600 150.940 ;
        RECT 179.400 148.940 179.795 150.940 ;
        RECT 4.000 147.540 179.795 148.940 ;
        RECT 4.400 145.540 175.600 147.540 ;
        RECT 179.400 145.540 179.795 147.540 ;
        RECT 4.000 144.140 179.795 145.540 ;
        RECT 4.400 142.140 179.795 144.140 ;
        RECT 4.000 140.740 179.795 142.140 ;
        RECT 4.400 138.740 175.600 140.740 ;
        RECT 179.400 138.740 179.795 140.740 ;
        RECT 4.000 137.340 179.795 138.740 ;
        RECT 4.400 135.340 175.600 137.340 ;
        RECT 179.400 135.340 179.795 137.340 ;
        RECT 4.000 133.940 179.795 135.340 ;
        RECT 4.000 131.940 175.600 133.940 ;
        RECT 179.400 131.940 179.795 133.940 ;
        RECT 4.000 130.540 179.795 131.940 ;
        RECT 4.400 128.540 175.600 130.540 ;
        RECT 179.400 128.540 179.795 130.540 ;
        RECT 4.000 127.140 179.795 128.540 ;
        RECT 4.400 125.140 175.600 127.140 ;
        RECT 179.400 125.140 179.795 127.140 ;
        RECT 4.000 123.740 179.795 125.140 ;
        RECT 4.400 121.740 175.600 123.740 ;
        RECT 179.400 121.740 179.795 123.740 ;
        RECT 4.000 120.340 179.795 121.740 ;
        RECT 4.400 118.340 175.600 120.340 ;
        RECT 179.400 118.340 179.795 120.340 ;
        RECT 4.000 116.940 179.795 118.340 ;
        RECT 4.400 114.940 175.600 116.940 ;
        RECT 179.400 114.940 179.795 116.940 ;
        RECT 4.000 113.540 179.795 114.940 ;
        RECT 4.400 111.540 175.600 113.540 ;
        RECT 179.400 111.540 179.795 113.540 ;
        RECT 4.000 110.140 179.795 111.540 ;
        RECT 4.400 108.140 179.795 110.140 ;
        RECT 4.000 106.740 179.795 108.140 ;
        RECT 4.400 104.740 175.600 106.740 ;
        RECT 179.400 104.740 179.795 106.740 ;
        RECT 4.000 103.340 179.795 104.740 ;
        RECT 4.400 101.340 175.600 103.340 ;
        RECT 179.400 101.340 179.795 103.340 ;
        RECT 4.000 99.940 179.795 101.340 ;
        RECT 4.000 97.940 175.600 99.940 ;
        RECT 179.400 97.940 179.795 99.940 ;
        RECT 4.000 96.540 179.795 97.940 ;
        RECT 4.400 94.540 175.600 96.540 ;
        RECT 179.400 94.540 179.795 96.540 ;
        RECT 4.000 93.140 179.795 94.540 ;
        RECT 4.400 91.140 175.600 93.140 ;
        RECT 179.400 91.140 179.795 93.140 ;
        RECT 4.000 89.740 179.795 91.140 ;
        RECT 4.400 87.740 175.600 89.740 ;
        RECT 179.400 87.740 179.795 89.740 ;
        RECT 4.000 86.340 179.795 87.740 ;
        RECT 4.400 84.340 175.600 86.340 ;
        RECT 179.400 84.340 179.795 86.340 ;
        RECT 4.000 82.940 179.795 84.340 ;
        RECT 4.400 80.940 175.600 82.940 ;
        RECT 179.400 80.940 179.795 82.940 ;
        RECT 4.000 79.540 179.795 80.940 ;
        RECT 4.400 77.540 175.600 79.540 ;
        RECT 179.400 77.540 179.795 79.540 ;
        RECT 4.000 76.140 179.795 77.540 ;
        RECT 4.400 74.140 179.795 76.140 ;
        RECT 4.000 72.740 179.795 74.140 ;
        RECT 4.400 70.740 175.600 72.740 ;
        RECT 179.400 70.740 179.795 72.740 ;
        RECT 4.000 69.340 179.795 70.740 ;
        RECT 4.400 67.340 175.600 69.340 ;
        RECT 179.400 67.340 179.795 69.340 ;
        RECT 4.000 65.940 179.795 67.340 ;
        RECT 4.000 63.940 175.600 65.940 ;
        RECT 179.400 63.940 179.795 65.940 ;
        RECT 4.000 62.540 179.795 63.940 ;
        RECT 4.400 60.540 175.600 62.540 ;
        RECT 179.400 60.540 179.795 62.540 ;
        RECT 4.000 59.140 179.795 60.540 ;
        RECT 4.400 57.140 175.600 59.140 ;
        RECT 179.400 57.140 179.795 59.140 ;
        RECT 4.000 55.740 179.795 57.140 ;
        RECT 4.400 53.740 175.600 55.740 ;
        RECT 179.400 53.740 179.795 55.740 ;
        RECT 4.000 52.340 179.795 53.740 ;
        RECT 4.400 50.340 175.600 52.340 ;
        RECT 179.400 50.340 179.795 52.340 ;
        RECT 4.000 48.940 179.795 50.340 ;
        RECT 4.400 46.940 175.600 48.940 ;
        RECT 179.400 46.940 179.795 48.940 ;
        RECT 4.000 45.540 179.795 46.940 ;
        RECT 4.400 43.540 175.600 45.540 ;
        RECT 179.400 43.540 179.795 45.540 ;
        RECT 4.000 42.140 179.795 43.540 ;
        RECT 4.400 40.140 179.795 42.140 ;
        RECT 4.000 38.740 179.795 40.140 ;
        RECT 4.400 36.740 175.600 38.740 ;
        RECT 179.400 36.740 179.795 38.740 ;
        RECT 4.000 35.340 179.795 36.740 ;
        RECT 4.400 33.340 175.600 35.340 ;
        RECT 179.400 33.340 179.795 35.340 ;
        RECT 4.000 31.940 179.795 33.340 ;
        RECT 4.000 29.940 175.600 31.940 ;
        RECT 179.400 29.940 179.795 31.940 ;
        RECT 4.000 28.540 179.795 29.940 ;
        RECT 4.400 26.540 175.600 28.540 ;
        RECT 179.400 26.540 179.795 28.540 ;
        RECT 4.000 25.140 179.795 26.540 ;
        RECT 4.400 23.140 175.600 25.140 ;
        RECT 179.400 23.140 179.795 25.140 ;
        RECT 4.000 21.740 179.795 23.140 ;
        RECT 4.400 19.740 175.600 21.740 ;
        RECT 179.400 19.740 179.795 21.740 ;
        RECT 4.000 18.340 179.795 19.740 ;
        RECT 4.400 16.340 175.600 18.340 ;
        RECT 179.400 16.340 179.795 18.340 ;
        RECT 4.000 14.940 179.795 16.340 ;
        RECT 4.400 12.940 175.600 14.940 ;
        RECT 179.400 12.940 179.795 14.940 ;
        RECT 4.000 11.540 179.795 12.940 ;
        RECT 4.400 9.540 175.600 11.540 ;
        RECT 179.400 9.540 179.795 11.540 ;
        RECT 4.000 8.140 179.795 9.540 ;
        RECT 4.400 6.140 179.795 8.140 ;
        RECT 4.000 4.740 179.795 6.140 ;
        RECT 4.400 2.740 175.600 4.740 ;
        RECT 179.400 2.740 179.795 4.740 ;
        RECT 4.000 1.340 179.795 2.740 ;
        RECT 4.000 0.175 175.600 1.340 ;
        RECT 179.400 0.175 179.795 1.340 ;
      LAYER met4 ;
        RECT 117.135 58.655 130.930 197.025 ;
        RECT 133.330 58.655 152.035 197.025 ;
        RECT 154.435 58.655 170.825 197.025 ;
  END
END wrapped_rgb_mixer
END LIBRARY

