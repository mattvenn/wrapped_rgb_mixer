magic
tech sky130A
magscale 1 2
timestamp 1647517088
<< viali >>
rect 10333 39593 10367 39627
rect 23765 39593 23799 39627
rect 26433 39593 26467 39627
rect 8401 39525 8435 39559
rect 12265 39525 12299 39559
rect 25329 39525 25363 39559
rect 1685 39457 1719 39491
rect 13553 39457 13587 39491
rect 16681 39457 16715 39491
rect 17417 39457 17451 39491
rect 19441 39457 19475 39491
rect 19993 39457 20027 39491
rect 27445 39457 27479 39491
rect 30757 39457 30791 39491
rect 32505 39457 32539 39491
rect 34161 39457 34195 39491
rect 1409 39389 1443 39423
rect 3065 39389 3099 39423
rect 3801 39389 3835 39423
rect 4629 39389 4663 39423
rect 5273 39389 5307 39423
rect 6561 39389 6595 39423
rect 7389 39389 7423 39423
rect 9137 39389 9171 39423
rect 10977 39389 11011 39423
rect 12909 39389 12943 39423
rect 14473 39389 14507 39423
rect 15117 39389 15151 39423
rect 15761 39389 15795 39423
rect 15945 39389 15979 39423
rect 21925 39389 21959 39423
rect 22017 39389 22051 39423
rect 22661 39389 22695 39423
rect 23673 39389 23707 39423
rect 24593 39389 24627 39423
rect 25605 39399 25639 39433
rect 26157 39389 26191 39423
rect 26249 39389 26283 39423
rect 26985 39389 27019 39423
rect 30665 39389 30699 39423
rect 31401 39389 31435 39423
rect 32321 39389 32355 39423
rect 14565 39321 14599 39355
rect 16129 39321 16163 39355
rect 16865 39321 16899 39355
rect 19625 39321 19659 39355
rect 22753 39321 22787 39355
rect 25329 39321 25363 39355
rect 25513 39321 25547 39355
rect 27169 39321 27203 39355
rect 30021 39321 30055 39355
rect 3157 39253 3191 39287
rect 3893 39253 3927 39287
rect 15209 39253 15243 39287
rect 22201 39253 22235 39287
rect 24777 39253 24811 39287
rect 30113 39253 30147 39287
rect 31493 39253 31527 39287
rect 12909 39049 12943 39083
rect 13645 39049 13679 39083
rect 30389 39049 30423 39083
rect 3985 38981 4019 39015
rect 8033 38981 8067 39015
rect 8769 38981 8803 39015
rect 24685 38981 24719 39015
rect 27077 38981 27111 39015
rect 27261 38981 27295 39015
rect 27905 38981 27939 39015
rect 30941 38981 30975 39015
rect 32505 38981 32539 39015
rect 1501 38913 1535 38947
rect 7297 38913 7331 38947
rect 7941 38913 7975 38947
rect 8585 38913 8619 38947
rect 11805 38913 11839 38947
rect 12449 38913 12483 38947
rect 13093 38913 13127 38947
rect 13553 38913 13587 38947
rect 16681 38913 16715 38947
rect 16865 38913 16899 38947
rect 20157 38913 20191 38947
rect 22201 38913 22235 38947
rect 24501 38913 24535 38947
rect 30205 38913 30239 38947
rect 32321 38913 32355 38947
rect 1685 38845 1719 38879
rect 1961 38845 1995 38879
rect 3801 38845 3835 38879
rect 5457 38845 5491 38879
rect 9321 38845 9355 38879
rect 14197 38845 14231 38879
rect 14381 38845 14415 38879
rect 14841 38845 14875 38879
rect 17509 38845 17543 38879
rect 17693 38845 17727 38879
rect 18245 38845 18279 38879
rect 19901 38845 19935 38879
rect 22385 38845 22419 38879
rect 22661 38845 22695 38879
rect 25145 38845 25179 38879
rect 27721 38845 27755 38879
rect 28365 38845 28399 38879
rect 30021 38845 30055 38879
rect 33517 38845 33551 38879
rect 31125 38777 31159 38811
rect 6745 38709 6779 38743
rect 7389 38709 7423 38743
rect 17049 38709 17083 38743
rect 21281 38709 21315 38743
rect 11621 38505 11655 38539
rect 14473 38505 14507 38539
rect 18153 38505 18187 38539
rect 19349 38505 19383 38539
rect 12265 38437 12299 38471
rect 23765 38437 23799 38471
rect 1961 38369 1995 38403
rect 4261 38369 4295 38403
rect 5825 38369 5859 38403
rect 6561 38369 6595 38403
rect 7113 38369 7147 38403
rect 9137 38369 9171 38403
rect 9413 38369 9447 38403
rect 15669 38369 15703 38403
rect 16129 38369 16163 38403
rect 20269 38369 20303 38403
rect 20729 38369 20763 38403
rect 25329 38369 25363 38403
rect 25789 38369 25823 38403
rect 28641 38369 28675 38403
rect 30021 38369 30055 38403
rect 32321 38369 32355 38403
rect 34161 38369 34195 38403
rect 1409 38301 1443 38335
rect 8953 38301 8987 38335
rect 12909 38301 12943 38335
rect 13553 38301 13587 38335
rect 14381 38301 14415 38335
rect 15485 38301 15519 38335
rect 17785 38301 17819 38335
rect 17969 38301 18003 38335
rect 19257 38301 19291 38335
rect 20085 38301 20119 38335
rect 22385 38301 22419 38335
rect 24501 38301 24535 38335
rect 25145 38301 25179 38335
rect 27445 38301 27479 38335
rect 27629 38301 27663 38335
rect 28365 38301 28399 38335
rect 29561 38301 29595 38335
rect 1593 38233 1627 38267
rect 4445 38233 4479 38267
rect 6745 38233 6779 38267
rect 22641 38233 22675 38267
rect 29745 38233 29779 38267
rect 32505 38233 32539 38267
rect 12725 38165 12759 38199
rect 13369 38165 13403 38199
rect 24593 38165 24627 38199
rect 27813 38165 27847 38199
rect 1961 37961 1995 37995
rect 5365 37961 5399 37995
rect 6653 37961 6687 37995
rect 11621 37961 11655 37995
rect 12265 37961 12299 37995
rect 12909 37961 12943 37995
rect 23213 37961 23247 37995
rect 23949 37961 23983 37995
rect 24041 37961 24075 37995
rect 2789 37893 2823 37927
rect 14657 37893 14691 37927
rect 22078 37893 22112 37927
rect 25053 37893 25087 37927
rect 29929 37893 29963 37927
rect 31585 37893 31619 37927
rect 34161 37893 34195 37927
rect 1869 37825 1903 37859
rect 5273 37825 5307 37859
rect 6561 37825 6595 37859
rect 7205 37825 7239 37859
rect 10333 37825 10367 37859
rect 10977 37825 11011 37859
rect 11805 37825 11839 37859
rect 12449 37825 12483 37859
rect 13093 37825 13127 37859
rect 13737 37825 13771 37859
rect 14289 37825 14323 37859
rect 15945 37825 15979 37859
rect 16037 37825 16071 37859
rect 16948 37825 16982 37859
rect 18788 37825 18822 37859
rect 20545 37825 20579 37859
rect 21833 37825 21867 37859
rect 23857 37825 23891 37859
rect 24869 37825 24903 37859
rect 25697 37825 25731 37859
rect 27169 37825 27203 37859
rect 28457 37825 28491 37859
rect 32321 37825 32355 37859
rect 2605 37757 2639 37791
rect 3065 37757 3099 37791
rect 7389 37757 7423 37791
rect 7757 37757 7791 37791
rect 16681 37757 16715 37791
rect 18521 37757 18555 37791
rect 20361 37757 20395 37791
rect 24685 37757 24719 37791
rect 25513 37757 25547 37791
rect 26985 37757 27019 37791
rect 28641 37757 28675 37791
rect 29745 37757 29779 37791
rect 32505 37757 32539 37791
rect 9689 37689 9723 37723
rect 19901 37689 19935 37723
rect 23673 37689 23707 37723
rect 13553 37621 13587 37655
rect 18061 37621 18095 37655
rect 20729 37621 20763 37655
rect 24225 37621 24259 37655
rect 25881 37621 25915 37655
rect 27353 37621 27387 37655
rect 1685 37417 1719 37451
rect 7389 37417 7423 37451
rect 8125 37417 8159 37451
rect 9597 37417 9631 37451
rect 10885 37417 10919 37451
rect 11345 37417 11379 37451
rect 17785 37417 17819 37451
rect 19349 37417 19383 37451
rect 21465 37417 21499 37451
rect 26157 37417 26191 37451
rect 31493 37417 31527 37451
rect 3065 37281 3099 37315
rect 10241 37281 10275 37315
rect 18337 37281 18371 37315
rect 19441 37281 19475 37315
rect 21097 37281 21131 37315
rect 22385 37281 22419 37315
rect 24777 37281 24811 37315
rect 32873 37281 32907 37315
rect 1593 37213 1627 37247
rect 2421 37213 2455 37247
rect 3801 37213 3835 37247
rect 5365 37213 5399 37247
rect 7297 37213 7331 37247
rect 11529 37213 11563 37247
rect 12173 37213 12207 37247
rect 12817 37213 12851 37247
rect 13277 37213 13311 37247
rect 14381 37213 14415 37247
rect 15761 37213 15795 37247
rect 17049 37213 17083 37247
rect 17693 37213 17727 37247
rect 18521 37213 18555 37247
rect 19625 37213 19659 37247
rect 20269 37213 20303 37247
rect 20637 37213 20671 37247
rect 21281 37213 21315 37247
rect 26617 37213 26651 37247
rect 28641 37213 28675 37247
rect 29929 37213 29963 37247
rect 30665 37213 30699 37247
rect 32137 37213 32171 37247
rect 4629 37145 4663 37179
rect 5917 37145 5951 37179
rect 15025 37145 15059 37179
rect 16221 37145 16255 37179
rect 17141 37145 17175 37179
rect 18705 37145 18739 37179
rect 19349 37145 19383 37179
rect 20453 37145 20487 37179
rect 22630 37145 22664 37179
rect 25022 37145 25056 37179
rect 26862 37145 26896 37179
rect 31309 37145 31343 37179
rect 31525 37145 31559 37179
rect 32321 37145 32355 37179
rect 11989 37077 12023 37111
rect 12633 37077 12667 37111
rect 13461 37077 13495 37111
rect 19809 37077 19843 37111
rect 23765 37077 23799 37111
rect 27997 37077 28031 37111
rect 28733 37077 28767 37111
rect 31677 37077 31711 37111
rect 13553 36873 13587 36907
rect 21925 36873 21959 36907
rect 31493 36873 31527 36907
rect 1593 36805 1627 36839
rect 2329 36805 2363 36839
rect 3985 36805 4019 36839
rect 5089 36805 5123 36839
rect 16937 36805 16971 36839
rect 25605 36805 25639 36839
rect 27414 36805 27448 36839
rect 1501 36737 1535 36771
rect 4537 36737 4571 36771
rect 5825 36737 5859 36771
rect 10333 36737 10367 36771
rect 10977 36737 11011 36771
rect 11805 36737 11839 36771
rect 12449 36737 12483 36771
rect 13093 36737 13127 36771
rect 13737 36737 13771 36771
rect 14381 36737 14415 36771
rect 15945 36737 15979 36771
rect 16037 36737 16071 36771
rect 18521 36737 18555 36771
rect 18777 36737 18811 36771
rect 20545 36737 20579 36771
rect 21833 36737 21867 36771
rect 22477 36737 22511 36771
rect 22753 36737 22787 36771
rect 23397 36737 23431 36771
rect 23581 36737 23615 36771
rect 24225 36737 24259 36771
rect 24409 36737 24443 36771
rect 25881 36737 25915 36771
rect 29101 36737 29135 36771
rect 30297 36737 30331 36771
rect 31401 36737 31435 36771
rect 34161 36737 34195 36771
rect 2145 36669 2179 36703
rect 14565 36669 14599 36703
rect 16681 36669 16715 36703
rect 20361 36669 20395 36703
rect 22661 36669 22695 36703
rect 24593 36669 24627 36703
rect 25789 36669 25823 36703
rect 27169 36669 27203 36703
rect 29653 36669 29687 36703
rect 30573 36669 30607 36703
rect 32321 36669 32355 36703
rect 32505 36669 32539 36703
rect 12909 36601 12943 36635
rect 11621 36533 11655 36567
rect 12265 36533 12299 36567
rect 18061 36533 18095 36567
rect 19901 36533 19935 36567
rect 20729 36533 20763 36567
rect 22753 36533 22787 36567
rect 22937 36533 22971 36567
rect 23765 36533 23799 36567
rect 25605 36533 25639 36567
rect 26065 36533 26099 36567
rect 28549 36533 28583 36567
rect 4997 36329 5031 36363
rect 10793 36329 10827 36363
rect 15945 36329 15979 36363
rect 16865 36329 16899 36363
rect 18705 36329 18739 36363
rect 25789 36329 25823 36363
rect 28549 36329 28583 36363
rect 11621 36261 11655 36295
rect 12081 36261 12115 36295
rect 23581 36261 23615 36295
rect 26249 36261 26283 36295
rect 1409 36193 1443 36227
rect 2789 36193 2823 36227
rect 16497 36193 16531 36227
rect 19533 36193 19567 36227
rect 24409 36193 24443 36227
rect 27537 36193 27571 36227
rect 28733 36193 28767 36227
rect 31125 36193 31159 36227
rect 32321 36193 32355 36227
rect 32505 36193 32539 36227
rect 32965 36193 32999 36227
rect 3893 36125 3927 36159
rect 4445 36125 4479 36159
rect 5181 36125 5215 36159
rect 10977 36125 11011 36159
rect 12265 36125 12299 36159
rect 12909 36125 12943 36159
rect 13553 36125 13587 36159
rect 14289 36125 14323 36159
rect 15853 36125 15887 36159
rect 16681 36125 16715 36159
rect 17325 36125 17359 36159
rect 21373 36125 21407 36159
rect 21629 36125 21663 36159
rect 23213 36125 23247 36159
rect 23383 36125 23417 36159
rect 27721 36125 27755 36159
rect 28089 36125 28123 36159
rect 28825 36125 28859 36159
rect 29653 36125 29687 36159
rect 30849 36125 30883 36159
rect 1593 36057 1627 36091
rect 14657 36057 14691 36091
rect 17592 36057 17626 36091
rect 19778 36057 19812 36091
rect 24654 36057 24688 36091
rect 26433 36057 26467 36091
rect 26617 36057 26651 36091
rect 28549 36057 28583 36091
rect 30205 36057 30239 36091
rect 12725 35989 12759 36023
rect 13369 35989 13403 36023
rect 20913 35989 20947 36023
rect 22753 35989 22787 36023
rect 26525 35989 26559 36023
rect 26801 35989 26835 36023
rect 27813 35989 27847 36023
rect 27905 35989 27939 36023
rect 29009 35989 29043 36023
rect 2237 35785 2271 35819
rect 3249 35785 3283 35819
rect 11897 35785 11931 35819
rect 13185 35785 13219 35819
rect 19533 35785 19567 35819
rect 23765 35785 23799 35819
rect 25697 35785 25731 35819
rect 30481 35785 30515 35819
rect 16129 35717 16163 35751
rect 16926 35717 16960 35751
rect 19717 35717 19751 35751
rect 22100 35717 22134 35751
rect 1409 35649 1443 35683
rect 2145 35649 2179 35683
rect 3065 35649 3099 35683
rect 3985 35649 4019 35683
rect 4629 35649 4663 35683
rect 12081 35649 12115 35683
rect 12725 35649 12759 35683
rect 13369 35649 13403 35683
rect 14013 35649 14047 35683
rect 14657 35649 14691 35683
rect 15117 35649 15151 35683
rect 15945 35649 15979 35683
rect 18521 35649 18555 35683
rect 18705 35649 18739 35683
rect 19625 35649 19659 35683
rect 20545 35649 20579 35683
rect 23673 35649 23707 35683
rect 24317 35649 24351 35683
rect 24573 35649 24607 35683
rect 26249 35649 26283 35683
rect 26433 35649 26467 35683
rect 27261 35649 27295 35683
rect 27517 35649 27551 35683
rect 29368 35649 29402 35683
rect 31401 35649 31435 35683
rect 32137 35649 32171 35683
rect 32321 35649 32355 35683
rect 33333 35649 33367 35683
rect 15209 35581 15243 35615
rect 15761 35581 15795 35615
rect 16681 35581 16715 35615
rect 19349 35581 19383 35615
rect 20361 35581 20395 35615
rect 21833 35581 21867 35615
rect 29101 35581 29135 35615
rect 31217 35581 31251 35615
rect 32505 35581 32539 35615
rect 33609 35581 33643 35615
rect 1593 35513 1627 35547
rect 12541 35513 12575 35547
rect 19901 35513 19935 35547
rect 20729 35513 20763 35547
rect 28641 35513 28675 35547
rect 13829 35445 13863 35479
rect 14473 35445 14507 35479
rect 18061 35445 18095 35479
rect 18889 35445 18923 35479
rect 23213 35445 23247 35479
rect 31585 35445 31619 35479
rect 12081 35241 12115 35275
rect 14289 35241 14323 35275
rect 16957 35241 16991 35275
rect 20729 35241 20763 35275
rect 23397 35241 23431 35275
rect 13185 35173 13219 35207
rect 14933 35173 14967 35207
rect 31861 35173 31895 35207
rect 2789 35105 2823 35139
rect 18705 35105 18739 35139
rect 21557 35105 21591 35139
rect 25053 35105 25087 35139
rect 25697 35105 25731 35139
rect 32321 35105 32355 35139
rect 1409 35037 1443 35071
rect 12725 35037 12759 35071
rect 13369 35037 13403 35071
rect 14473 35037 14507 35071
rect 15117 35037 15151 35071
rect 15577 35037 15611 35071
rect 17417 35037 17451 35071
rect 17693 35037 17727 35071
rect 18521 35037 18555 35071
rect 19441 35037 19475 35071
rect 19533 35037 19567 35071
rect 19901 35037 19935 35071
rect 20453 35037 20487 35071
rect 20545 35037 20579 35071
rect 23581 35037 23615 35071
rect 23673 35037 23707 35071
rect 24593 35037 24627 35071
rect 27721 35037 27755 35071
rect 27813 35037 27847 35071
rect 28023 35037 28057 35071
rect 28181 35037 28215 35071
rect 29561 35037 29595 35071
rect 30481 35037 30515 35071
rect 1593 34969 1627 35003
rect 15822 34969 15856 35003
rect 19625 34969 19659 35003
rect 19763 34969 19797 35003
rect 21802 34969 21836 35003
rect 23397 34969 23431 35003
rect 24685 34969 24719 35003
rect 24777 34969 24811 35003
rect 24915 34969 24949 35003
rect 25964 34969 25998 35003
rect 27537 34969 27571 35003
rect 27905 34969 27939 35003
rect 28641 34969 28675 35003
rect 28825 34969 28859 35003
rect 29837 34969 29871 35003
rect 30748 34969 30782 35003
rect 32505 34969 32539 35003
rect 34161 34969 34195 35003
rect 12541 34901 12575 34935
rect 17601 34901 17635 34935
rect 17785 34901 17819 34935
rect 17969 34901 18003 34935
rect 19257 34901 19291 34935
rect 22937 34901 22971 34935
rect 23857 34901 23891 34935
rect 24409 34901 24443 34935
rect 27077 34901 27111 34935
rect 29009 34901 29043 34935
rect 12725 34697 12759 34731
rect 13369 34697 13403 34731
rect 14841 34697 14875 34731
rect 15301 34697 15335 34731
rect 17049 34697 17083 34731
rect 23489 34697 23523 34731
rect 26157 34697 26191 34731
rect 32137 34697 32171 34731
rect 33609 34697 33643 34731
rect 18797 34629 18831 34663
rect 22354 34629 22388 34663
rect 24216 34629 24250 34663
rect 25789 34629 25823 34663
rect 29009 34629 29043 34663
rect 33241 34629 33275 34663
rect 1777 34561 1811 34595
rect 12909 34561 12943 34595
rect 13553 34561 13587 34595
rect 14197 34561 14231 34595
rect 14657 34561 14691 34595
rect 14841 34561 14875 34595
rect 15485 34561 15519 34595
rect 15945 34561 15979 34595
rect 16129 34561 16163 34595
rect 16865 34561 16899 34595
rect 17509 34561 17543 34595
rect 17785 34561 17819 34595
rect 18429 34561 18463 34595
rect 18613 34561 18647 34595
rect 19625 34561 19659 34595
rect 19892 34561 19926 34595
rect 22109 34561 22143 34595
rect 25973 34561 26007 34595
rect 27077 34561 27111 34595
rect 28825 34561 28859 34595
rect 29101 34561 29135 34595
rect 29653 34561 29687 34595
rect 29920 34561 29954 34595
rect 32367 34561 32401 34595
rect 32505 34561 32539 34595
rect 32597 34561 32631 34595
rect 32781 34561 32815 34595
rect 33425 34561 33459 34595
rect 33701 34561 33735 34595
rect 16037 34493 16071 34527
rect 16681 34493 16715 34527
rect 17693 34493 17727 34527
rect 23949 34493 23983 34527
rect 27721 34493 27755 34527
rect 28181 34493 28215 34527
rect 2421 34425 2455 34459
rect 12265 34425 12299 34459
rect 14013 34425 14047 34459
rect 21005 34425 21039 34459
rect 27261 34425 27295 34459
rect 27997 34425 28031 34459
rect 17509 34357 17543 34391
rect 17969 34357 18003 34391
rect 25329 34357 25363 34391
rect 28641 34357 28675 34391
rect 31033 34357 31067 34391
rect 12909 34153 12943 34187
rect 20637 34153 20671 34187
rect 23581 34153 23615 34187
rect 30757 34153 30791 34187
rect 13369 34085 13403 34119
rect 18061 34085 18095 34119
rect 18613 34085 18647 34119
rect 24869 34085 24903 34119
rect 2789 34017 2823 34051
rect 16681 34017 16715 34051
rect 25329 34017 25363 34051
rect 34161 34017 34195 34051
rect 1409 33949 1443 33983
rect 12265 33949 12299 33983
rect 13553 33949 13587 33983
rect 14105 33949 14139 33983
rect 14289 33949 14323 33983
rect 14933 33949 14967 33983
rect 15577 33949 15611 33983
rect 16037 33949 16071 33983
rect 18521 33949 18555 33983
rect 19257 33949 19291 33983
rect 21833 33949 21867 33983
rect 22109 33949 22143 33983
rect 23029 33949 23063 33983
rect 23305 33949 23339 33983
rect 24593 33949 24627 33983
rect 24685 33949 24719 33983
rect 25585 33949 25619 33983
rect 27169 33949 27203 33983
rect 29653 33949 29687 33983
rect 30113 33949 30147 33983
rect 31033 33949 31067 33983
rect 31125 33949 31159 33983
rect 31217 33949 31251 33983
rect 31401 33949 31435 33983
rect 32321 33949 32355 33983
rect 1593 33881 1627 33915
rect 16129 33881 16163 33915
rect 16926 33881 16960 33915
rect 19502 33881 19536 33915
rect 27414 33881 27448 33915
rect 32505 33881 32539 33915
rect 14289 33813 14323 33847
rect 14749 33813 14783 33847
rect 15393 33813 15427 33847
rect 21649 33813 21683 33847
rect 22017 33813 22051 33847
rect 23213 33813 23247 33847
rect 23397 33813 23431 33847
rect 26709 33813 26743 33847
rect 28549 33813 28583 33847
rect 2605 33609 2639 33643
rect 12081 33609 12115 33643
rect 13553 33609 13587 33643
rect 21833 33609 21867 33643
rect 23213 33609 23247 33643
rect 25513 33609 25547 33643
rect 27813 33609 27847 33643
rect 28089 33609 28123 33643
rect 30297 33609 30331 33643
rect 31585 33609 31619 33643
rect 14994 33541 15028 33575
rect 18613 33541 18647 33575
rect 18829 33541 18863 33575
rect 20545 33541 20579 33575
rect 27930 33541 27964 33575
rect 30941 33541 30975 33575
rect 32505 33541 32539 33575
rect 2053 33473 2087 33507
rect 2513 33473 2547 33507
rect 12265 33473 12299 33507
rect 12725 33473 12759 33507
rect 12909 33473 12943 33507
rect 13369 33473 13403 33507
rect 13553 33473 13587 33507
rect 14105 33473 14139 33507
rect 14289 33473 14323 33507
rect 16865 33473 16899 33507
rect 17969 33473 18003 33507
rect 18153 33473 18187 33507
rect 19809 33473 19843 33507
rect 19901 33473 19935 33507
rect 20085 33473 20119 33507
rect 22017 33473 22051 33507
rect 22109 33473 22143 33507
rect 22278 33473 22312 33507
rect 22385 33473 22419 33507
rect 23029 33473 23063 33507
rect 24133 33473 24167 33507
rect 24389 33473 24423 33507
rect 26065 33473 26099 33507
rect 26249 33473 26283 33507
rect 26433 33473 26467 33507
rect 28733 33473 28767 33507
rect 28825 33473 28859 33507
rect 29101 33473 29135 33507
rect 30113 33473 30147 33507
rect 31309 33473 31343 33507
rect 32321 33473 32355 33507
rect 14197 33405 14231 33439
rect 14749 33405 14783 33439
rect 16681 33405 16715 33439
rect 17785 33405 17819 33439
rect 22845 33405 22879 33439
rect 27445 33405 27479 33439
rect 27721 33405 27755 33439
rect 29009 33405 29043 33439
rect 29653 33405 29687 33439
rect 30021 33405 30055 33439
rect 31401 33405 31435 33439
rect 34161 33405 34195 33439
rect 17049 33337 17083 33371
rect 20821 33337 20855 33371
rect 21005 33337 21039 33371
rect 23765 33337 23799 33371
rect 12817 33269 12851 33303
rect 16129 33269 16163 33303
rect 18797 33269 18831 33303
rect 18981 33269 19015 33303
rect 28549 33269 28583 33303
rect 12081 33065 12115 33099
rect 18705 33065 18739 33099
rect 29653 33065 29687 33099
rect 30573 33065 30607 33099
rect 12725 32997 12759 33031
rect 13461 32997 13495 33031
rect 22109 32997 22143 33031
rect 22569 32997 22603 33031
rect 23857 32997 23891 33031
rect 24685 32997 24719 33031
rect 25605 32997 25639 33031
rect 27537 32997 27571 33031
rect 27721 32997 27755 33031
rect 14657 32929 14691 32963
rect 19257 32929 19291 32963
rect 26065 32929 26099 32963
rect 27261 32929 27295 32963
rect 28457 32929 28491 32963
rect 30481 32929 30515 32963
rect 31861 32929 31895 32963
rect 32689 32929 32723 32963
rect 12265 32861 12299 32895
rect 12909 32861 12943 32895
rect 13369 32861 13403 32895
rect 13553 32861 13587 32895
rect 14289 32861 14323 32895
rect 14473 32861 14507 32895
rect 15117 32861 15151 32895
rect 17325 32861 17359 32895
rect 21373 32861 21407 32895
rect 21557 32861 21591 32895
rect 21649 32861 21683 32895
rect 21787 32861 21821 32895
rect 21925 32861 21959 32895
rect 22799 32861 22833 32895
rect 23029 32861 23063 32895
rect 23489 32861 23523 32895
rect 23673 32861 23707 32895
rect 24501 32861 24535 32895
rect 25421 32861 25455 32895
rect 26249 32861 26283 32895
rect 28181 32861 28215 32895
rect 28365 32861 28399 32895
rect 28549 32861 28583 32895
rect 28716 32861 28750 32895
rect 29561 32861 29595 32895
rect 30205 32861 30239 32895
rect 31493 32861 31527 32895
rect 31677 32861 31711 32895
rect 31769 32861 31803 32895
rect 32045 32861 32079 32895
rect 15362 32793 15396 32827
rect 17570 32793 17604 32827
rect 19524 32793 19558 32827
rect 25237 32793 25271 32827
rect 26433 32793 26467 32827
rect 32229 32793 32263 32827
rect 32934 32793 32968 32827
rect 16497 32725 16531 32759
rect 20637 32725 20671 32759
rect 22937 32725 22971 32759
rect 28917 32725 28951 32759
rect 30757 32725 30791 32759
rect 34069 32725 34103 32759
rect 12265 32521 12299 32555
rect 16865 32521 16899 32555
rect 17877 32521 17911 32555
rect 17969 32521 18003 32555
rect 19901 32521 19935 32555
rect 20913 32521 20947 32555
rect 21005 32521 21039 32555
rect 21281 32521 21315 32555
rect 29837 32521 29871 32555
rect 13001 32453 13035 32487
rect 15669 32453 15703 32487
rect 16773 32453 16807 32487
rect 17417 32453 17451 32487
rect 21122 32453 21156 32487
rect 23734 32453 23768 32487
rect 25513 32453 25547 32487
rect 34161 32453 34195 32487
rect 12449 32385 12483 32419
rect 12909 32385 12943 32419
rect 13093 32385 13127 32419
rect 13553 32385 13587 32419
rect 14197 32385 14231 32419
rect 15025 32385 15059 32419
rect 15945 32385 15979 32419
rect 17605 32385 17639 32419
rect 18061 32385 18095 32419
rect 18521 32385 18555 32419
rect 18777 32385 18811 32419
rect 20637 32385 20671 32419
rect 22017 32385 22051 32419
rect 22109 32385 22143 32419
rect 22385 32385 22419 32419
rect 22845 32385 22879 32419
rect 23489 32385 23523 32419
rect 25329 32385 25363 32419
rect 25605 32385 25639 32419
rect 26249 32385 26283 32419
rect 27537 32385 27571 32419
rect 28457 32385 28491 32419
rect 28622 32385 28656 32419
rect 28733 32385 28767 32419
rect 28825 32385 28859 32419
rect 29469 32385 29503 32419
rect 31033 32385 31067 32419
rect 32321 32385 32355 32419
rect 11805 32317 11839 32351
rect 14841 32317 14875 32351
rect 15853 32317 15887 32351
rect 17693 32317 17727 32351
rect 26065 32317 26099 32351
rect 27813 32317 27847 32351
rect 29561 32317 29595 32351
rect 30757 32317 30791 32351
rect 32505 32317 32539 32351
rect 25329 32249 25363 32283
rect 26433 32249 26467 32283
rect 27353 32249 27387 32283
rect 13645 32181 13679 32215
rect 14289 32181 14323 32215
rect 15209 32181 15243 32215
rect 15945 32181 15979 32215
rect 16129 32181 16163 32215
rect 21833 32181 21867 32215
rect 22293 32181 22327 32215
rect 22937 32181 22971 32215
rect 24869 32181 24903 32215
rect 27721 32181 27755 32215
rect 28273 32181 28307 32215
rect 12817 31977 12851 32011
rect 16681 31977 16715 32011
rect 18521 31977 18555 32011
rect 21005 31977 21039 32011
rect 23213 31977 23247 32011
rect 25881 31977 25915 32011
rect 30665 31977 30699 32011
rect 12173 31909 12207 31943
rect 14841 31909 14875 31943
rect 17141 31909 17175 31943
rect 18705 31909 18739 31943
rect 20821 31909 20855 31943
rect 31861 31909 31895 31943
rect 15301 31841 15335 31875
rect 17693 31841 17727 31875
rect 18429 31841 18463 31875
rect 20545 31841 20579 31875
rect 22109 31841 22143 31875
rect 24409 31841 24443 31875
rect 25053 31841 25087 31875
rect 27813 31841 27847 31875
rect 30205 31841 30239 31875
rect 31401 31841 31435 31875
rect 32321 31841 32355 31875
rect 32505 31841 32539 31875
rect 34161 31841 34195 31875
rect 1685 31773 1719 31807
rect 11713 31773 11747 31807
rect 12357 31773 12391 31807
rect 12817 31773 12851 31807
rect 13001 31773 13035 31807
rect 14657 31773 14691 31807
rect 17325 31773 17359 31807
rect 17417 31773 17451 31807
rect 18521 31773 18555 31807
rect 22201 31773 22235 31807
rect 23489 31773 23523 31807
rect 23581 31773 23615 31807
rect 23673 31773 23707 31807
rect 23857 31773 23891 31807
rect 24777 31773 24811 31807
rect 24869 31773 24903 31807
rect 25513 31773 25547 31807
rect 25697 31773 25731 31807
rect 25973 31773 26007 31807
rect 26663 31773 26697 31807
rect 26801 31773 26835 31807
rect 26893 31773 26927 31807
rect 27077 31773 27111 31807
rect 27721 31773 27755 31807
rect 28549 31773 28583 31807
rect 28733 31773 28767 31807
rect 29009 31773 29043 31807
rect 30297 31773 30331 31807
rect 31493 31773 31527 31807
rect 15546 31705 15580 31739
rect 18245 31705 18279 31739
rect 19625 31705 19659 31739
rect 19809 31705 19843 31739
rect 11529 31637 11563 31671
rect 17509 31637 17543 31671
rect 22569 31637 22603 31671
rect 26433 31637 26467 31671
rect 28089 31637 28123 31671
rect 28917 31637 28951 31671
rect 12909 31433 12943 31467
rect 30205 31433 30239 31467
rect 14994 31365 15028 31399
rect 16773 31365 16807 31399
rect 16957 31365 16991 31399
rect 18245 31365 18279 31399
rect 19625 31365 19659 31399
rect 20361 31365 20395 31399
rect 24501 31365 24535 31399
rect 31401 31365 31435 31399
rect 1501 31297 1535 31331
rect 12265 31297 12299 31331
rect 12817 31297 12851 31331
rect 13001 31297 13035 31331
rect 13461 31297 13495 31331
rect 13645 31297 13679 31331
rect 14105 31297 14139 31331
rect 14749 31297 14783 31331
rect 17601 31297 17635 31331
rect 18429 31297 18463 31331
rect 18685 31297 18719 31331
rect 20545 31297 20579 31331
rect 21005 31297 21039 31331
rect 21833 31297 21867 31331
rect 22845 31297 22879 31331
rect 23751 31297 23785 31331
rect 24869 31297 24903 31331
rect 25789 31297 25823 31331
rect 30389 31297 30423 31331
rect 30573 31297 30607 31331
rect 30665 31297 30699 31331
rect 31217 31297 31251 31331
rect 34161 31297 34195 31331
rect 1685 31229 1719 31263
rect 1961 31229 1995 31263
rect 14197 31229 14231 31263
rect 17417 31229 17451 31263
rect 21281 31229 21315 31263
rect 22109 31229 22143 31263
rect 23673 31229 23707 31263
rect 24961 31229 24995 31263
rect 25145 31229 25179 31263
rect 25697 31229 25731 31263
rect 27537 31229 27571 31263
rect 27721 31229 27755 31263
rect 27997 31229 28031 31263
rect 30481 31229 30515 31263
rect 31585 31229 31619 31263
rect 32321 31229 32355 31263
rect 32505 31229 32539 31263
rect 12081 31161 12115 31195
rect 16129 31161 16163 31195
rect 18613 31161 18647 31195
rect 21189 31161 21223 31195
rect 22385 31161 22419 31195
rect 22937 31161 22971 31195
rect 13553 31093 13587 31127
rect 17785 31093 17819 31127
rect 19717 31093 19751 31127
rect 21097 31093 21131 31127
rect 22201 31093 22235 31127
rect 23949 31093 23983 31127
rect 26065 31093 26099 31127
rect 1869 30889 1903 30923
rect 12081 30889 12115 30923
rect 13369 30889 13403 30923
rect 18705 30889 18739 30923
rect 23029 30889 23063 30923
rect 27905 30889 27939 30923
rect 33885 30889 33919 30923
rect 15669 30821 15703 30855
rect 25145 30821 25179 30855
rect 29009 30821 29043 30855
rect 12817 30753 12851 30787
rect 16129 30753 16163 30787
rect 17325 30753 17359 30787
rect 21373 30753 21407 30787
rect 21557 30753 21591 30787
rect 22109 30753 22143 30787
rect 23489 30753 23523 30787
rect 24685 30753 24719 30787
rect 28549 30753 28583 30787
rect 32137 30753 32171 30787
rect 32229 30753 32263 30787
rect 33333 30753 33367 30787
rect 1777 30685 1811 30719
rect 11621 30685 11655 30719
rect 12265 30685 12299 30719
rect 12725 30685 12759 30719
rect 12909 30685 12943 30719
rect 13369 30685 13403 30719
rect 13553 30685 13587 30719
rect 14749 30685 14783 30719
rect 16313 30685 16347 30719
rect 19257 30685 19291 30719
rect 19441 30685 19475 30719
rect 21281 30685 21315 30719
rect 22201 30685 22235 30719
rect 23213 30685 23247 30719
rect 23305 30685 23339 30719
rect 23397 30685 23431 30719
rect 24777 30685 24811 30719
rect 25789 30685 25823 30719
rect 25973 30685 26007 30719
rect 26065 30685 26099 30719
rect 26525 30685 26559 30719
rect 26781 30685 26815 30719
rect 28719 30685 28753 30719
rect 30113 30685 30147 30719
rect 32321 30685 32355 30719
rect 32413 30685 32447 30719
rect 32965 30685 32999 30719
rect 33149 30685 33183 30719
rect 33425 30685 33459 30719
rect 33885 30685 33919 30719
rect 34161 30685 34195 30719
rect 14933 30617 14967 30651
rect 15485 30617 15519 30651
rect 17570 30617 17604 30651
rect 20269 30617 20303 30651
rect 20453 30617 20487 30651
rect 30358 30617 30392 30651
rect 16497 30549 16531 30583
rect 19625 30549 19659 30583
rect 20913 30549 20947 30583
rect 22569 30549 22603 30583
rect 25605 30549 25639 30583
rect 31493 30549 31527 30583
rect 31953 30549 31987 30583
rect 34069 30549 34103 30583
rect 17055 30345 17089 30379
rect 31375 30345 31409 30379
rect 15209 30277 15243 30311
rect 16129 30277 16163 30311
rect 19800 30277 19834 30311
rect 21833 30277 21867 30311
rect 26433 30277 26467 30311
rect 27445 30277 27479 30311
rect 29929 30277 29963 30311
rect 31585 30277 31619 30311
rect 11897 30209 11931 30243
rect 12081 30209 12115 30243
rect 12541 30209 12575 30243
rect 12725 30209 12759 30243
rect 13185 30209 13219 30243
rect 13369 30209 13403 30243
rect 13829 30209 13863 30243
rect 14473 30209 14507 30243
rect 15393 30209 15427 30243
rect 15945 30209 15979 30243
rect 16957 30209 16991 30243
rect 17141 30209 17175 30243
rect 17233 30209 17267 30243
rect 17693 30209 17727 30243
rect 17949 30209 17983 30243
rect 19533 30209 19567 30243
rect 22063 30209 22097 30243
rect 22198 30212 22232 30246
rect 22293 30209 22327 30243
rect 22477 30209 22511 30243
rect 23121 30209 23155 30243
rect 23949 30209 23983 30243
rect 24777 30209 24811 30243
rect 25053 30209 25087 30243
rect 26249 30209 26283 30243
rect 27261 30209 27295 30243
rect 27537 30209 27571 30243
rect 28264 30209 28298 30243
rect 30205 30209 30239 30243
rect 30294 30209 30328 30243
rect 30410 30212 30444 30246
rect 30573 30209 30607 30243
rect 32505 30209 32539 30243
rect 33517 30209 33551 30243
rect 33793 30209 33827 30243
rect 11989 30141 12023 30175
rect 23029 30141 23063 30175
rect 24869 30141 24903 30175
rect 24961 30141 24995 30175
rect 26065 30141 26099 30175
rect 27997 30141 28031 30175
rect 32413 30141 32447 30175
rect 12633 30073 12667 30107
rect 23489 30073 23523 30107
rect 24593 30073 24627 30107
rect 29377 30073 29411 30107
rect 31217 30073 31251 30107
rect 13277 30005 13311 30039
rect 13921 30005 13955 30039
rect 14565 30005 14599 30039
rect 19073 30005 19107 30039
rect 20913 30005 20947 30039
rect 24041 30005 24075 30039
rect 27077 30005 27111 30039
rect 30849 30005 30883 30039
rect 31401 30005 31435 30039
rect 32781 30005 32815 30039
rect 33333 30005 33367 30039
rect 33701 30005 33735 30039
rect 22845 29801 22879 29835
rect 23581 29801 23615 29835
rect 23765 29801 23799 29835
rect 24777 29801 24811 29835
rect 28365 29801 28399 29835
rect 32229 29801 32263 29835
rect 34161 29801 34195 29835
rect 20913 29733 20947 29767
rect 22477 29733 22511 29767
rect 26709 29733 26743 29767
rect 12817 29665 12851 29699
rect 19533 29665 19567 29699
rect 26249 29665 26283 29699
rect 27261 29665 27295 29699
rect 30021 29665 30055 29699
rect 31217 29665 31251 29699
rect 32781 29665 32815 29699
rect 12265 29597 12299 29631
rect 12725 29597 12759 29631
rect 12909 29597 12943 29631
rect 13369 29597 13403 29631
rect 13553 29597 13587 29631
rect 14105 29597 14139 29631
rect 14289 29597 14323 29631
rect 14749 29597 14783 29631
rect 15393 29597 15427 29631
rect 15485 29597 15519 29631
rect 16037 29597 16071 29631
rect 17877 29597 17911 29631
rect 18061 29597 18095 29631
rect 21649 29597 21683 29631
rect 21741 29597 21775 29631
rect 21833 29597 21867 29631
rect 22017 29597 22051 29631
rect 22661 29597 22695 29631
rect 22937 29597 22971 29631
rect 25421 29597 25455 29631
rect 25513 29597 25547 29631
rect 26341 29597 26375 29631
rect 27353 29597 27387 29631
rect 28595 29597 28629 29631
rect 28733 29597 28767 29631
rect 28825 29594 28859 29628
rect 29009 29597 29043 29631
rect 29745 29597 29779 29631
rect 29838 29597 29872 29631
rect 30113 29597 30147 29631
rect 31387 29597 31421 29631
rect 32137 29597 32171 29631
rect 16282 29529 16316 29563
rect 19800 29529 19834 29563
rect 21373 29529 21407 29563
rect 23397 29529 23431 29563
rect 24409 29529 24443 29563
rect 24593 29529 24627 29563
rect 25697 29529 25731 29563
rect 33026 29529 33060 29563
rect 12081 29461 12115 29495
rect 13461 29461 13495 29495
rect 14289 29461 14323 29495
rect 14841 29461 14875 29495
rect 17417 29461 17451 29495
rect 18245 29461 18279 29495
rect 23597 29461 23631 29495
rect 27721 29461 27755 29495
rect 29561 29461 29595 29495
rect 31677 29461 31711 29495
rect 13001 29257 13035 29291
rect 32873 29257 32907 29291
rect 34069 29257 34103 29291
rect 14657 29189 14691 29223
rect 19993 29189 20027 29223
rect 21833 29189 21867 29223
rect 22017 29189 22051 29223
rect 22753 29189 22787 29223
rect 32229 29189 32263 29223
rect 11989 29121 12023 29155
rect 13185 29121 13219 29155
rect 13277 29121 13311 29155
rect 13461 29121 13495 29155
rect 13921 29121 13955 29155
rect 14105 29121 14139 29155
rect 14565 29121 14599 29155
rect 14749 29121 14783 29155
rect 15209 29121 15243 29155
rect 15853 29121 15887 29155
rect 16037 29121 16071 29155
rect 16129 29121 16163 29155
rect 17213 29121 17247 29155
rect 18981 29121 19015 29155
rect 19809 29121 19843 29155
rect 21005 29121 21039 29155
rect 21281 29121 21315 29155
rect 23009 29121 23043 29155
rect 23134 29121 23168 29155
rect 23234 29121 23268 29155
rect 23397 29121 23431 29155
rect 24133 29121 24167 29155
rect 24400 29121 24434 29155
rect 25973 29121 26007 29155
rect 26157 29121 26191 29155
rect 26341 29121 26375 29155
rect 26985 29121 27019 29155
rect 27241 29121 27275 29155
rect 28825 29121 28859 29155
rect 29092 29121 29126 29155
rect 31217 29121 31251 29155
rect 33149 29121 33183 29155
rect 33241 29121 33275 29155
rect 33333 29121 33367 29155
rect 33517 29121 33551 29155
rect 33977 29121 34011 29155
rect 12541 29053 12575 29087
rect 12909 29053 12943 29087
rect 14013 29053 14047 29087
rect 16957 29053 16991 29087
rect 18797 29053 18831 29087
rect 19625 29053 19659 29087
rect 22201 29053 22235 29087
rect 26249 29053 26283 29087
rect 26433 29053 26467 29087
rect 31309 29053 31343 29087
rect 15301 28985 15335 29019
rect 18337 28985 18371 29019
rect 19165 28985 19199 29019
rect 21005 28985 21039 29019
rect 21097 28985 21131 29019
rect 28365 28985 28399 29019
rect 31585 28985 31619 29019
rect 32413 28985 32447 29019
rect 12173 28917 12207 28951
rect 13461 28917 13495 28951
rect 13737 28917 13771 28951
rect 15853 28917 15887 28951
rect 25513 28917 25547 28951
rect 30205 28917 30239 28951
rect 12725 28713 12759 28747
rect 20637 28713 20671 28747
rect 28549 28713 28583 28747
rect 13369 28645 13403 28679
rect 21097 28645 21131 28679
rect 21465 28645 21499 28679
rect 27077 28645 27111 28679
rect 28917 28645 28951 28679
rect 33149 28645 33183 28679
rect 18153 28577 18187 28611
rect 19257 28577 19291 28611
rect 22477 28577 22511 28611
rect 30113 28577 30147 28611
rect 12909 28509 12943 28543
rect 13553 28509 13587 28543
rect 14657 28509 14691 28543
rect 14749 28509 14783 28543
rect 15301 28509 15335 28543
rect 15393 28509 15427 28543
rect 16313 28509 16347 28543
rect 21281 28509 21315 28543
rect 21557 28509 21591 28543
rect 22744 28509 22778 28543
rect 26341 28509 26375 28543
rect 26985 28509 27019 28543
rect 27261 28509 27295 28543
rect 27445 28509 27479 28543
rect 27813 28509 27847 28543
rect 27997 28509 28031 28543
rect 28733 28509 28767 28543
rect 29009 28509 29043 28543
rect 31953 28509 31987 28543
rect 32046 28509 32080 28543
rect 32418 28509 32452 28543
rect 33057 28509 33091 28543
rect 33333 28509 33367 28543
rect 33609 28509 33643 28543
rect 33793 28509 33827 28543
rect 16569 28441 16603 28475
rect 18429 28441 18463 28475
rect 19524 28441 19558 28475
rect 24777 28441 24811 28475
rect 30358 28441 30392 28475
rect 32229 28441 32263 28475
rect 32321 28441 32355 28475
rect 17693 28373 17727 28407
rect 18337 28373 18371 28407
rect 18521 28373 18555 28407
rect 18705 28373 18739 28407
rect 23857 28373 23891 28407
rect 31493 28373 31527 28407
rect 32597 28373 32631 28407
rect 13277 28169 13311 28203
rect 17325 28169 17359 28203
rect 21281 28169 21315 28203
rect 23949 28169 23983 28203
rect 26341 28169 26375 28203
rect 26985 28169 27019 28203
rect 14657 28101 14691 28135
rect 16037 28101 16071 28135
rect 18306 28101 18340 28135
rect 20168 28101 20202 28135
rect 22017 28101 22051 28135
rect 24317 28101 24351 28135
rect 32505 28101 32539 28135
rect 13461 28033 13495 28067
rect 13921 28033 13955 28067
rect 14105 28033 14139 28067
rect 14565 28033 14599 28067
rect 14749 28033 14783 28067
rect 15209 28033 15243 28067
rect 15301 28033 15335 28067
rect 15853 28033 15887 28067
rect 16129 28033 16163 28067
rect 17141 28033 17175 28067
rect 18061 28033 18095 28067
rect 19901 28033 19935 28067
rect 22201 28033 22235 28067
rect 22293 28033 22327 28067
rect 22753 28033 22787 28067
rect 22846 28033 22880 28067
rect 23029 28033 23063 28067
rect 23121 28033 23155 28067
rect 23259 28033 23293 28067
rect 23857 28033 23891 28067
rect 24777 28033 24811 28067
rect 24961 28033 24995 28067
rect 25053 28033 25087 28067
rect 25329 28033 25363 28067
rect 26157 28033 26191 28067
rect 27169 28033 27203 28067
rect 27261 28033 27295 28067
rect 27537 28033 27571 28067
rect 28540 28033 28574 28067
rect 30297 28033 30331 28067
rect 30389 28033 30423 28067
rect 30573 28033 30607 28067
rect 30665 28033 30699 28067
rect 31125 28033 31159 28067
rect 32321 28033 32355 28067
rect 16957 27965 16991 27999
rect 24225 27965 24259 27999
rect 25145 27965 25179 27999
rect 25973 27965 26007 27999
rect 28273 27965 28307 27999
rect 34161 27965 34195 27999
rect 19441 27897 19475 27931
rect 22017 27897 22051 27931
rect 27445 27897 27479 27931
rect 29653 27897 29687 27931
rect 30113 27897 30147 27931
rect 13921 27829 13955 27863
rect 15853 27829 15887 27863
rect 23397 27829 23431 27863
rect 24133 27829 24167 27863
rect 25513 27829 25547 27863
rect 31309 27829 31343 27863
rect 31585 27829 31619 27863
rect 19257 27625 19291 27659
rect 26525 27625 26559 27659
rect 32321 27625 32355 27659
rect 34161 27625 34195 27659
rect 13369 27557 13403 27591
rect 19717 27557 19751 27591
rect 24961 27557 24995 27591
rect 28917 27557 28951 27591
rect 14749 27489 14783 27523
rect 16129 27489 16163 27523
rect 16681 27489 16715 27523
rect 17509 27489 17543 27523
rect 19441 27489 19475 27523
rect 21741 27489 21775 27523
rect 28825 27489 28859 27523
rect 29561 27489 29595 27523
rect 30941 27489 30975 27523
rect 31125 27489 31159 27523
rect 31861 27489 31895 27523
rect 31953 27489 31987 27523
rect 13553 27421 13587 27455
rect 14657 27421 14691 27455
rect 14841 27421 14875 27455
rect 15301 27421 15335 27455
rect 15485 27421 15519 27455
rect 16037 27421 16071 27455
rect 16865 27421 16899 27455
rect 17693 27421 17727 27455
rect 18337 27421 18371 27455
rect 19533 27421 19567 27455
rect 20913 27421 20947 27455
rect 21005 27421 21039 27455
rect 21189 27421 21223 27455
rect 21281 27421 21315 27455
rect 22017 27421 22051 27455
rect 23489 27421 23523 27455
rect 24409 27421 24443 27455
rect 24685 27421 24719 27455
rect 24777 27421 24811 27455
rect 25881 27421 25915 27455
rect 25974 27421 26008 27455
rect 26249 27421 26283 27455
rect 26346 27421 26380 27455
rect 27261 27421 27295 27455
rect 27721 27421 27755 27455
rect 28549 27421 28583 27455
rect 28917 27421 28951 27455
rect 29837 27421 29871 27455
rect 30849 27421 30883 27455
rect 31585 27421 31619 27455
rect 31769 27421 31803 27455
rect 32137 27421 32171 27455
rect 32781 27421 32815 27455
rect 17049 27353 17083 27387
rect 17877 27353 17911 27387
rect 18521 27353 18555 27387
rect 19257 27353 19291 27387
rect 23673 27353 23707 27387
rect 23857 27353 23891 27387
rect 24593 27353 24627 27387
rect 26157 27353 26191 27387
rect 27077 27353 27111 27387
rect 31125 27353 31159 27387
rect 33048 27353 33082 27387
rect 15393 27285 15427 27319
rect 18705 27285 18739 27319
rect 20729 27285 20763 27319
rect 27905 27285 27939 27319
rect 28641 27285 28675 27319
rect 15393 27081 15427 27115
rect 17601 27081 17635 27115
rect 17785 27081 17819 27115
rect 21281 27081 21315 27115
rect 22661 27081 22695 27115
rect 25237 27081 25271 27115
rect 28365 27081 28399 27115
rect 28825 27081 28859 27115
rect 31585 27081 31619 27115
rect 32229 27081 32263 27115
rect 33517 27081 33551 27115
rect 18981 27013 19015 27047
rect 19073 27013 19107 27047
rect 24102 27013 24136 27047
rect 30205 27013 30239 27047
rect 30297 27013 30331 27047
rect 31217 27013 31251 27047
rect 13553 26945 13587 26979
rect 14197 26945 14231 26979
rect 14841 26945 14875 26979
rect 15301 26945 15335 26979
rect 15485 26945 15519 26979
rect 15945 26945 15979 26979
rect 16037 26945 16071 26979
rect 16773 26945 16807 26979
rect 17693 26945 17727 26979
rect 17969 26945 18003 26979
rect 18889 26945 18923 26979
rect 19191 26945 19225 26979
rect 19349 26945 19383 26979
rect 20168 26945 20202 26979
rect 21925 26945 21959 26979
rect 22109 26945 22143 26979
rect 22477 26945 22511 26979
rect 23121 26945 23155 26979
rect 23305 26945 23339 26979
rect 23397 26945 23431 26979
rect 25789 26945 25823 26979
rect 25881 26945 25915 26979
rect 27241 26945 27275 26979
rect 29009 26945 29043 26979
rect 29929 26945 29963 26979
rect 30022 26945 30056 26979
rect 30435 26945 30469 26979
rect 31033 26945 31067 26979
rect 31309 26945 31343 26979
rect 31401 26945 31435 26979
rect 32137 26945 32171 26979
rect 32781 26945 32815 26979
rect 32969 26943 33003 26977
rect 33333 26945 33367 26979
rect 33977 26945 34011 26979
rect 17417 26877 17451 26911
rect 19901 26877 19935 26911
rect 22201 26877 22235 26911
rect 22293 26877 22327 26911
rect 23857 26877 23891 26911
rect 26985 26877 27019 26911
rect 29285 26877 29319 26911
rect 33057 26877 33091 26911
rect 33149 26877 33183 26911
rect 14013 26809 14047 26843
rect 30573 26809 30607 26843
rect 14657 26741 14691 26775
rect 16865 26741 16899 26775
rect 18705 26741 18739 26775
rect 23121 26741 23155 26775
rect 26065 26741 26099 26775
rect 29193 26741 29227 26775
rect 34069 26741 34103 26775
rect 14289 26537 14323 26571
rect 16957 26537 16991 26571
rect 17509 26537 17543 26571
rect 17877 26537 17911 26571
rect 21097 26537 21131 26571
rect 23489 26537 23523 26571
rect 23673 26537 23707 26571
rect 26249 26537 26283 26571
rect 28825 26537 28859 26571
rect 29009 26537 29043 26571
rect 31401 26537 31435 26571
rect 33701 26537 33735 26571
rect 31309 26469 31343 26503
rect 17601 26401 17635 26435
rect 22017 26401 22051 26435
rect 29653 26401 29687 26435
rect 29929 26401 29963 26435
rect 30941 26401 30975 26435
rect 14473 26333 14507 26367
rect 14933 26333 14967 26367
rect 15117 26333 15151 26367
rect 15577 26333 15611 26367
rect 15833 26333 15867 26367
rect 17693 26333 17727 26367
rect 18337 26333 18371 26367
rect 18521 26333 18555 26367
rect 19257 26333 19291 26367
rect 19524 26333 19558 26367
rect 21281 26333 21315 26367
rect 21465 26333 21499 26367
rect 21557 26333 21591 26367
rect 22293 26333 22327 26367
rect 24869 26333 24903 26367
rect 26709 26333 26743 26367
rect 32321 26333 32355 26367
rect 32577 26333 32611 26367
rect 23535 26299 23569 26333
rect 17417 26265 17451 26299
rect 23305 26265 23339 26299
rect 25136 26265 25170 26299
rect 26954 26265 26988 26299
rect 28641 26265 28675 26299
rect 15025 26197 15059 26231
rect 18705 26197 18739 26231
rect 20637 26197 20671 26231
rect 28089 26197 28123 26231
rect 28841 26197 28875 26231
rect 25605 25993 25639 26027
rect 26985 25993 27019 26027
rect 29745 25993 29779 26027
rect 15393 25925 15427 25959
rect 19708 25925 19742 25959
rect 24032 25925 24066 25959
rect 30205 25925 30239 25959
rect 30421 25925 30455 25959
rect 14013 25857 14047 25891
rect 14473 25857 14507 25891
rect 14657 25857 14691 25891
rect 15209 25857 15243 25891
rect 15945 25857 15979 25891
rect 17397 25857 17431 25891
rect 19441 25857 19475 25891
rect 21925 25857 21959 25891
rect 22181 25857 22215 25891
rect 23765 25857 23799 25891
rect 25789 25857 25823 25891
rect 26065 25857 26099 25891
rect 27169 25857 27203 25891
rect 27353 25857 27387 25891
rect 28632 25857 28666 25891
rect 31309 25857 31343 25891
rect 34161 25857 34195 25891
rect 17141 25789 17175 25823
rect 27445 25789 27479 25823
rect 28365 25789 28399 25823
rect 31493 25789 31527 25823
rect 31585 25789 31619 25823
rect 32321 25789 32355 25823
rect 32505 25789 32539 25823
rect 14473 25721 14507 25755
rect 18521 25721 18555 25755
rect 23305 25721 23339 25755
rect 25145 25721 25179 25755
rect 31125 25721 31159 25755
rect 13829 25653 13863 25687
rect 16037 25653 16071 25687
rect 20821 25653 20855 25687
rect 25973 25653 26007 25687
rect 30389 25653 30423 25687
rect 30573 25653 30607 25687
rect 14381 25449 14415 25483
rect 17141 25449 17175 25483
rect 23857 25449 23891 25483
rect 24593 25449 24627 25483
rect 25513 25449 25547 25483
rect 26249 25449 26283 25483
rect 26433 25449 26467 25483
rect 27997 25449 28031 25483
rect 29009 25449 29043 25483
rect 20085 25381 20119 25415
rect 22201 25381 22235 25415
rect 24777 25381 24811 25415
rect 27261 25381 27295 25415
rect 1869 25313 1903 25347
rect 15761 25313 15795 25347
rect 20821 25313 20855 25347
rect 23489 25313 23523 25347
rect 31769 25313 31803 25347
rect 31861 25313 31895 25347
rect 32321 25313 32355 25347
rect 1409 25245 1443 25279
rect 14565 25245 14599 25279
rect 16017 25245 16051 25279
rect 18429 25245 18463 25279
rect 18521 25245 18555 25279
rect 19809 25245 19843 25279
rect 19901 25245 19935 25279
rect 21077 25245 21111 25279
rect 23673 25245 23707 25279
rect 25421 25245 25455 25279
rect 27077 25245 27111 25279
rect 27813 25245 27847 25279
rect 28733 25245 28767 25279
rect 28825 25245 28859 25279
rect 29561 25245 29595 25279
rect 31585 25245 31619 25279
rect 34161 25245 34195 25279
rect 24639 25211 24673 25245
rect 26295 25211 26329 25245
rect 1593 25177 1627 25211
rect 15117 25177 15151 25211
rect 15301 25177 15335 25211
rect 17693 25177 17727 25211
rect 17877 25177 17911 25211
rect 22661 25177 22695 25211
rect 22845 25177 22879 25211
rect 24409 25177 24443 25211
rect 26065 25177 26099 25211
rect 29828 25177 29862 25211
rect 32505 25177 32539 25211
rect 18705 25109 18739 25143
rect 23029 25109 23063 25143
rect 30941 25109 30975 25143
rect 31401 25109 31435 25143
rect 2697 24905 2731 24939
rect 13737 24905 13771 24939
rect 16129 24905 16163 24939
rect 28825 24905 28859 24939
rect 27813 24837 27847 24871
rect 28029 24837 28063 24871
rect 29377 24837 29411 24871
rect 29577 24837 29611 24871
rect 32382 24837 32416 24871
rect 2053 24769 2087 24803
rect 2605 24769 2639 24803
rect 13921 24769 13955 24803
rect 14565 24769 14599 24803
rect 15117 24769 15151 24803
rect 15945 24769 15979 24803
rect 17233 24769 17267 24803
rect 17417 24769 17451 24803
rect 18061 24769 18095 24803
rect 18317 24769 18351 24803
rect 20453 24769 20487 24803
rect 20729 24769 20763 24803
rect 21833 24769 21867 24803
rect 22017 24769 22051 24803
rect 22845 24769 22879 24803
rect 23949 24769 23983 24803
rect 25513 24769 25547 24803
rect 25697 24769 25731 24803
rect 25789 24769 25823 24803
rect 26249 24769 26283 24803
rect 27077 24769 27111 24803
rect 28733 24769 28767 24803
rect 30472 24769 30506 24803
rect 33977 24769 34011 24803
rect 34069 24769 34103 24803
rect 15761 24701 15795 24735
rect 22661 24701 22695 24735
rect 23673 24701 23707 24735
rect 27353 24701 27387 24735
rect 30205 24701 30239 24735
rect 32137 24701 32171 24735
rect 15301 24633 15335 24667
rect 17601 24633 17635 24667
rect 19441 24633 19475 24667
rect 26341 24633 26375 24667
rect 28181 24633 28215 24667
rect 14381 24565 14415 24599
rect 22201 24565 22235 24599
rect 23029 24565 23063 24599
rect 25329 24565 25363 24599
rect 27169 24565 27203 24599
rect 27261 24565 27295 24599
rect 27997 24565 28031 24599
rect 29561 24565 29595 24599
rect 29745 24565 29779 24599
rect 31585 24565 31619 24599
rect 33517 24565 33551 24599
rect 17509 24361 17543 24395
rect 18245 24361 18279 24395
rect 31769 24361 31803 24395
rect 18429 24293 18463 24327
rect 21281 24293 21315 24327
rect 29561 24293 29595 24327
rect 32505 24225 32539 24259
rect 34161 24225 34195 24259
rect 14933 24157 14967 24191
rect 15485 24157 15519 24191
rect 15669 24157 15703 24191
rect 16129 24157 16163 24191
rect 17969 24157 18003 24191
rect 18153 24157 18187 24191
rect 18245 24157 18279 24191
rect 19717 24157 19751 24191
rect 19809 24157 19843 24191
rect 19901 24157 19935 24191
rect 20085 24157 20119 24191
rect 22201 24157 22235 24191
rect 22477 24157 22511 24191
rect 23213 24157 23247 24191
rect 23397 24157 23431 24191
rect 23489 24157 23523 24191
rect 24685 24157 24719 24191
rect 26709 24157 26743 24191
rect 27629 24157 27663 24191
rect 29837 24157 29871 24191
rect 30389 24157 30423 24191
rect 32321 24157 32355 24191
rect 16396 24089 16430 24123
rect 21005 24089 21039 24123
rect 24930 24089 24964 24123
rect 26525 24089 26559 24123
rect 27896 24089 27930 24123
rect 29561 24089 29595 24123
rect 30656 24089 30690 24123
rect 14749 24021 14783 24055
rect 19441 24021 19475 24055
rect 21465 24021 21499 24055
rect 22017 24021 22051 24055
rect 22385 24021 22419 24055
rect 23029 24021 23063 24055
rect 26065 24021 26099 24055
rect 26893 24021 26927 24055
rect 29009 24021 29043 24055
rect 29745 24021 29779 24055
rect 17325 23817 17359 23851
rect 22477 23817 22511 23851
rect 27445 23817 27479 23851
rect 31125 23817 31159 23851
rect 18306 23749 18340 23783
rect 20146 23749 20180 23783
rect 24317 23749 24351 23783
rect 34161 23749 34195 23783
rect 15025 23681 15059 23715
rect 15945 23681 15979 23715
rect 17049 23681 17083 23715
rect 17233 23681 17267 23715
rect 17417 23681 17451 23715
rect 17601 23681 17635 23715
rect 19901 23681 19935 23715
rect 21833 23681 21867 23715
rect 22201 23681 22235 23715
rect 22318 23681 22352 23715
rect 23113 23681 23147 23715
rect 23286 23681 23320 23715
rect 23397 23681 23431 23715
rect 23489 23681 23523 23715
rect 24133 23681 24167 23715
rect 24409 23681 24443 23715
rect 25237 23681 25271 23715
rect 25421 23681 25455 23715
rect 25789 23681 25823 23715
rect 27261 23681 27295 23715
rect 27537 23681 27571 23715
rect 28273 23681 28307 23715
rect 28549 23681 28583 23715
rect 30941 23681 30975 23715
rect 15761 23613 15795 23647
rect 18061 23613 18095 23647
rect 22109 23613 22143 23647
rect 22937 23613 22971 23647
rect 25513 23613 25547 23647
rect 25605 23613 25639 23647
rect 28457 23613 28491 23647
rect 29055 23613 29089 23647
rect 29285 23613 29319 23647
rect 30757 23613 30791 23647
rect 32321 23613 32355 23647
rect 32505 23613 32539 23647
rect 14841 23545 14875 23579
rect 28089 23545 28123 23579
rect 16129 23477 16163 23511
rect 19441 23477 19475 23511
rect 21281 23477 21315 23511
rect 23949 23477 23983 23511
rect 25973 23477 26007 23511
rect 27077 23477 27111 23511
rect 14473 23273 14507 23307
rect 17969 23273 18003 23307
rect 24869 23273 24903 23307
rect 28457 23273 28491 23307
rect 30941 23273 30975 23307
rect 31493 23273 31527 23307
rect 16037 23205 16071 23239
rect 16589 23137 16623 23171
rect 22109 23137 22143 23171
rect 22201 23137 22235 23171
rect 23029 23137 23063 23171
rect 23305 23137 23339 23171
rect 25145 23137 25179 23171
rect 25237 23137 25271 23171
rect 31677 23137 31711 23171
rect 34161 23137 34195 23171
rect 14657 23069 14691 23103
rect 15301 23069 15335 23103
rect 15945 23069 15979 23103
rect 16129 23069 16163 23103
rect 18429 23069 18463 23103
rect 19257 23069 19291 23103
rect 21833 23069 21867 23103
rect 22017 23069 22051 23103
rect 22396 23069 22430 23103
rect 25053 23069 25087 23103
rect 25329 23069 25363 23103
rect 26065 23069 26099 23103
rect 26332 23069 26366 23103
rect 27905 23069 27939 23103
rect 28273 23069 28307 23103
rect 29561 23069 29595 23103
rect 31401 23069 31435 23103
rect 32321 23069 32355 23103
rect 16856 23001 16890 23035
rect 19502 23001 19536 23035
rect 21189 23001 21223 23035
rect 21373 23001 21407 23035
rect 28089 23001 28123 23035
rect 28181 23001 28215 23035
rect 29806 23001 29840 23035
rect 32505 23001 32539 23035
rect 15117 22933 15151 22967
rect 18613 22933 18647 22967
rect 20637 22933 20671 22967
rect 22569 22933 22603 22967
rect 27445 22933 27479 22967
rect 31677 22933 31711 22967
rect 18061 22729 18095 22763
rect 19073 22729 19107 22763
rect 20269 22729 20303 22763
rect 23581 22729 23615 22763
rect 28641 22729 28675 22763
rect 31033 22729 31067 22763
rect 32321 22729 32355 22763
rect 16129 22661 16163 22695
rect 29460 22661 29494 22695
rect 33149 22661 33183 22695
rect 15301 22593 15335 22627
rect 15945 22593 15979 22627
rect 16681 22593 16715 22627
rect 16937 22593 16971 22627
rect 19349 22593 19383 22627
rect 19533 22593 19567 22627
rect 20085 22593 20119 22627
rect 20361 22593 20395 22627
rect 22201 22593 22235 22627
rect 22468 22593 22502 22627
rect 24041 22593 24075 22627
rect 24133 22593 24167 22627
rect 24915 22593 24949 22627
rect 25053 22593 25087 22627
rect 25145 22593 25179 22627
rect 25329 22593 25363 22627
rect 25973 22593 26007 22627
rect 26065 22593 26099 22627
rect 28549 22593 28583 22627
rect 31033 22593 31067 22627
rect 32137 22593 32171 22627
rect 32413 22593 32447 22627
rect 32873 22593 32907 22627
rect 32965 22593 32999 22627
rect 33793 22593 33827 22627
rect 15761 22525 15795 22559
rect 19257 22525 19291 22559
rect 19441 22525 19475 22559
rect 20821 22525 20855 22559
rect 26157 22525 26191 22559
rect 26249 22525 26283 22559
rect 27261 22525 27295 22559
rect 27537 22525 27571 22559
rect 29193 22525 29227 22559
rect 31309 22525 31343 22559
rect 33149 22525 33183 22559
rect 15117 22457 15151 22491
rect 21097 22457 21131 22491
rect 25789 22457 25823 22491
rect 31125 22457 31159 22491
rect 33609 22457 33643 22491
rect 20085 22389 20119 22423
rect 21281 22389 21315 22423
rect 24685 22389 24719 22423
rect 30573 22389 30607 22423
rect 32137 22389 32171 22423
rect 17785 22185 17819 22219
rect 19349 22185 19383 22219
rect 20361 22185 20395 22219
rect 21005 22185 21039 22219
rect 22201 22185 22235 22219
rect 22937 22185 22971 22219
rect 29745 22185 29779 22219
rect 20545 22117 20579 22151
rect 27445 22117 27479 22151
rect 31125 22117 31159 22151
rect 16405 22049 16439 22083
rect 18245 22049 18279 22083
rect 24501 22049 24535 22083
rect 24961 22049 24995 22083
rect 27905 22049 27939 22083
rect 28365 22049 28399 22083
rect 30461 22049 30495 22083
rect 32137 22049 32171 22083
rect 32873 22049 32907 22083
rect 33701 22049 33735 22083
rect 18429 21981 18463 22015
rect 19441 21981 19475 22015
rect 19533 21981 19567 22015
rect 21005 21981 21039 22015
rect 21281 21981 21315 22015
rect 21741 21981 21775 22015
rect 21925 21981 21959 22015
rect 22017 21981 22051 22015
rect 22293 21981 22327 22015
rect 23213 21981 23247 22015
rect 23305 21981 23339 22015
rect 23397 21981 23431 22015
rect 23581 21981 23615 22015
rect 24593 21981 24627 22015
rect 25421 21981 25455 22015
rect 26065 21981 26099 22015
rect 26332 21981 26366 22015
rect 28072 21981 28106 22015
rect 28181 21981 28215 22015
rect 28457 21981 28491 22015
rect 30573 21981 30607 22015
rect 30665 21981 30699 22015
rect 31401 21981 31435 22015
rect 31861 21981 31895 22015
rect 31953 21981 31987 22015
rect 32689 21981 32723 22015
rect 33609 21981 33643 22015
rect 16672 21913 16706 21947
rect 19257 21913 19291 21947
rect 20177 21913 20211 21947
rect 20377 21913 20411 21947
rect 21189 21913 21223 21947
rect 29561 21913 29595 21947
rect 30389 21913 30423 21947
rect 31125 21913 31159 21947
rect 18613 21845 18647 21879
rect 19717 21845 19751 21879
rect 25513 21845 25547 21879
rect 29761 21845 29795 21879
rect 29929 21845 29963 21879
rect 31309 21845 31343 21879
rect 32137 21845 32171 21879
rect 21281 21641 21315 21675
rect 23029 21641 23063 21675
rect 27905 21641 27939 21675
rect 32321 21641 32355 21675
rect 33425 21641 33459 21675
rect 34069 21641 34103 21675
rect 22661 21573 22695 21607
rect 27537 21573 27571 21607
rect 31125 21573 31159 21607
rect 17417 21505 17451 21539
rect 18328 21505 18362 21539
rect 20157 21505 20191 21539
rect 21833 21505 21867 21539
rect 22017 21505 22051 21539
rect 22845 21505 22879 21539
rect 23121 21505 23155 21539
rect 23581 21505 23615 21539
rect 23765 21505 23799 21539
rect 24041 21505 24075 21539
rect 24777 21505 24811 21539
rect 24869 21505 24903 21539
rect 24961 21505 24995 21539
rect 25145 21505 25179 21539
rect 25789 21505 25823 21539
rect 27353 21505 27387 21539
rect 27629 21505 27663 21539
rect 27745 21505 27779 21539
rect 28457 21505 28491 21539
rect 29469 21505 29503 21539
rect 30113 21505 30147 21539
rect 30205 21505 30239 21539
rect 30849 21505 30883 21539
rect 32229 21505 32263 21539
rect 33333 21505 33367 21539
rect 33977 21505 34011 21539
rect 17233 21437 17267 21471
rect 18061 21437 18095 21471
rect 19901 21437 19935 21471
rect 25697 21437 25731 21471
rect 26157 21437 26191 21471
rect 29285 21437 29319 21471
rect 30389 21437 30423 21471
rect 22201 21369 22235 21403
rect 30297 21369 30331 21403
rect 30849 21369 30883 21403
rect 30941 21369 30975 21403
rect 17601 21301 17635 21335
rect 19441 21301 19475 21335
rect 23949 21301 23983 21335
rect 24501 21301 24535 21335
rect 28549 21301 28583 21335
rect 29653 21301 29687 21335
rect 17049 21097 17083 21131
rect 17693 21097 17727 21131
rect 20545 21097 20579 21131
rect 22477 21097 22511 21131
rect 24501 21097 24535 21131
rect 28273 21097 28307 21131
rect 30941 21097 30975 21131
rect 31585 21097 31619 21131
rect 33885 21097 33919 21131
rect 26801 21029 26835 21063
rect 18705 20961 18739 20995
rect 21097 20961 21131 20995
rect 22937 20961 22971 20995
rect 27721 20961 27755 20995
rect 17233 20893 17267 20927
rect 17877 20893 17911 20927
rect 18337 20893 18371 20927
rect 18521 20893 18555 20927
rect 19809 20893 19843 20927
rect 19993 20893 20027 20927
rect 20453 20893 20487 20927
rect 21364 20893 21398 20927
rect 23213 20893 23247 20927
rect 23305 20893 23339 20927
rect 23397 20893 23431 20927
rect 23581 20893 23615 20927
rect 24685 20893 24719 20927
rect 24961 20893 24995 20927
rect 25421 20893 25455 20927
rect 27445 20893 27479 20927
rect 27537 20893 27571 20927
rect 27813 20893 27847 20927
rect 28457 20893 28491 20927
rect 28733 20893 28767 20927
rect 29561 20893 29595 20927
rect 31493 20893 31527 20927
rect 32137 20893 32171 20927
rect 32321 20893 32355 20927
rect 33241 20893 33275 20927
rect 34069 20893 34103 20927
rect 25688 20825 25722 20859
rect 29828 20825 29862 20859
rect 32229 20825 32263 20859
rect 19901 20757 19935 20791
rect 24869 20757 24903 20791
rect 27261 20757 27295 20791
rect 28641 20757 28675 20791
rect 33333 20757 33367 20791
rect 23581 20553 23615 20587
rect 28825 20553 28859 20587
rect 29485 20553 29519 20587
rect 31033 20553 31067 20587
rect 21189 20485 21223 20519
rect 28457 20485 28491 20519
rect 28549 20485 28583 20519
rect 29285 20485 29319 20519
rect 30941 20485 30975 20519
rect 32505 20485 32539 20519
rect 18521 20417 18555 20451
rect 20453 20417 20487 20451
rect 21097 20417 21131 20451
rect 21281 20417 21315 20451
rect 21925 20417 21959 20451
rect 22845 20417 22879 20451
rect 23029 20417 23063 20451
rect 24961 20417 24995 20451
rect 25973 20417 26007 20451
rect 26157 20417 26191 20451
rect 26341 20417 26375 20451
rect 26985 20417 27019 20451
rect 27169 20417 27203 20451
rect 27353 20417 27387 20451
rect 27537 20417 27571 20451
rect 27721 20417 27755 20451
rect 28181 20417 28215 20451
rect 28274 20417 28308 20451
rect 28646 20417 28680 20451
rect 30113 20417 30147 20451
rect 30389 20417 30423 20451
rect 34161 20417 34195 20451
rect 22109 20349 22143 20383
rect 22753 20349 22787 20383
rect 22937 20349 22971 20383
rect 23949 20349 23983 20383
rect 24041 20349 24075 20383
rect 24685 20349 24719 20383
rect 26433 20349 26467 20383
rect 27261 20349 27295 20383
rect 32321 20349 32355 20383
rect 18337 20281 18371 20315
rect 20545 20281 20579 20315
rect 29653 20281 29687 20315
rect 30205 20281 30239 20315
rect 22569 20213 22603 20247
rect 24225 20213 24259 20247
rect 29469 20213 29503 20247
rect 30113 20213 30147 20247
rect 20453 20009 20487 20043
rect 22569 20009 22603 20043
rect 26249 20009 26283 20043
rect 27353 20009 27387 20043
rect 27997 20009 28031 20043
rect 28273 20009 28307 20043
rect 30481 20009 30515 20043
rect 23765 19941 23799 19975
rect 28733 19941 28767 19975
rect 29929 19941 29963 19975
rect 22293 19873 22327 19907
rect 23305 19873 23339 19907
rect 24501 19873 24535 19907
rect 25697 19873 25731 19907
rect 1961 19805 1995 19839
rect 20453 19805 20487 19839
rect 20637 19805 20671 19839
rect 22201 19805 22235 19839
rect 23397 19805 23431 19839
rect 24593 19805 24627 19839
rect 26157 19805 26191 19839
rect 26801 19805 26835 19839
rect 27169 19805 27203 19839
rect 27813 19805 27847 19839
rect 28917 19805 28951 19839
rect 29009 19805 29043 19839
rect 29745 19805 29779 19839
rect 30021 19805 30055 19839
rect 30665 19805 30699 19839
rect 30757 19805 30791 19839
rect 31217 19805 31251 19839
rect 32321 19805 32355 19839
rect 21373 19737 21407 19771
rect 25513 19737 25547 19771
rect 26985 19737 27019 19771
rect 27077 19737 27111 19771
rect 28733 19737 28767 19771
rect 30481 19737 30515 19771
rect 32505 19737 32539 19771
rect 34161 19737 34195 19771
rect 21465 19669 21499 19703
rect 24961 19669 24995 19703
rect 29561 19669 29595 19703
rect 31309 19669 31343 19703
rect 22569 19465 22603 19499
rect 26341 19465 26375 19499
rect 30665 19465 30699 19499
rect 31217 19465 31251 19499
rect 32137 19465 32171 19499
rect 33241 19465 33275 19499
rect 33977 19465 34011 19499
rect 20729 19397 20763 19431
rect 24133 19397 24167 19431
rect 24317 19397 24351 19431
rect 28365 19397 28399 19431
rect 29530 19397 29564 19431
rect 1777 19329 1811 19363
rect 20637 19329 20671 19363
rect 20821 19329 20855 19363
rect 22385 19329 22419 19363
rect 22661 19329 22695 19363
rect 23305 19329 23339 19363
rect 24961 19329 24995 19363
rect 26249 19329 26283 19363
rect 27261 19329 27295 19363
rect 27445 19329 27479 19363
rect 28181 19329 28215 19363
rect 29285 19329 29319 19363
rect 31125 19329 31159 19363
rect 32321 19329 32355 19363
rect 33149 19329 33183 19363
rect 33885 19329 33919 19363
rect 1961 19261 1995 19295
rect 2237 19261 2271 19295
rect 23213 19261 23247 19295
rect 23673 19261 23707 19295
rect 24501 19261 24535 19295
rect 25237 19261 25271 19295
rect 27537 19261 27571 19295
rect 27997 19261 28031 19295
rect 22201 19125 22235 19159
rect 27077 19125 27111 19159
rect 2513 18921 2547 18955
rect 21741 18921 21775 18955
rect 22753 18921 22787 18955
rect 24593 18921 24627 18955
rect 28733 18921 28767 18955
rect 30941 18921 30975 18955
rect 31493 18921 31527 18955
rect 23305 18785 23339 18819
rect 23765 18785 23799 18819
rect 24777 18785 24811 18819
rect 34161 18785 34195 18819
rect 1685 18717 1719 18751
rect 2421 18717 2455 18751
rect 21741 18717 21775 18751
rect 21925 18717 21959 18751
rect 22385 18717 22419 18751
rect 22569 18717 22603 18751
rect 23397 18717 23431 18751
rect 24501 18717 24535 18751
rect 25237 18717 25271 18751
rect 27353 18717 27387 18751
rect 29561 18717 29595 18751
rect 29828 18717 29862 18751
rect 31401 18717 31435 18751
rect 32321 18717 32355 18751
rect 25504 18649 25538 18683
rect 27620 18649 27654 18683
rect 32505 18649 32539 18683
rect 24777 18581 24811 18615
rect 26617 18581 26651 18615
rect 22477 18377 22511 18411
rect 24593 18377 24627 18411
rect 26433 18377 26467 18411
rect 28365 18377 28399 18411
rect 29653 18377 29687 18411
rect 30297 18377 30331 18411
rect 31493 18377 31527 18411
rect 32597 18377 32631 18411
rect 33701 18377 33735 18411
rect 27230 18309 27264 18343
rect 1501 18241 1535 18275
rect 22385 18241 22419 18275
rect 22569 18241 22603 18275
rect 23581 18241 23615 18275
rect 24409 18241 24443 18275
rect 24593 18241 24627 18275
rect 25053 18241 25087 18275
rect 25309 18241 25343 18275
rect 26985 18241 27019 18275
rect 28825 18241 28859 18275
rect 29561 18241 29595 18275
rect 29745 18241 29779 18275
rect 30205 18241 30239 18275
rect 30389 18241 30423 18275
rect 31401 18241 31435 18275
rect 31585 18241 31619 18275
rect 32505 18241 32539 18275
rect 33609 18241 33643 18275
rect 1685 18173 1719 18207
rect 2881 18173 2915 18207
rect 23673 18173 23707 18207
rect 29101 18173 29135 18207
rect 23949 18105 23983 18139
rect 28917 18037 28951 18071
rect 29009 18037 29043 18071
rect 1869 17833 1903 17867
rect 24961 17833 24995 17867
rect 25789 17833 25823 17867
rect 26525 17833 26559 17867
rect 27353 17833 27387 17867
rect 28549 17833 28583 17867
rect 30113 17833 30147 17867
rect 31217 17833 31251 17867
rect 30573 17765 30607 17799
rect 25973 17697 26007 17731
rect 34161 17697 34195 17731
rect 1777 17629 1811 17663
rect 24961 17629 24995 17663
rect 25237 17629 25271 17663
rect 25697 17629 25731 17663
rect 26433 17629 26467 17663
rect 27537 17629 27571 17663
rect 27629 17629 27663 17663
rect 28549 17629 28583 17663
rect 28733 17629 28767 17663
rect 30573 17629 30607 17663
rect 30757 17629 30791 17663
rect 31217 17629 31251 17663
rect 31401 17629 31435 17663
rect 32321 17629 32355 17663
rect 25145 17561 25179 17595
rect 27353 17561 27387 17595
rect 32505 17561 32539 17595
rect 25973 17493 26007 17527
rect 24869 17289 24903 17323
rect 25513 17289 25547 17323
rect 27905 17289 27939 17323
rect 31493 17289 31527 17323
rect 24685 17221 24719 17255
rect 24961 17153 24995 17187
rect 25421 17153 25455 17187
rect 25605 17153 25639 17187
rect 27813 17153 27847 17187
rect 27997 17153 28031 17187
rect 30297 17153 30331 17187
rect 30941 17153 30975 17187
rect 31401 17153 31435 17187
rect 31585 17153 31619 17187
rect 1501 17085 1535 17119
rect 1685 17085 1719 17119
rect 1961 17085 1995 17119
rect 29653 17085 29687 17119
rect 32321 17085 32355 17119
rect 32505 17085 32539 17119
rect 34161 17085 34195 17119
rect 24685 17017 24719 17051
rect 1869 16745 1903 16779
rect 2605 16745 2639 16779
rect 31033 16745 31067 16779
rect 31677 16745 31711 16779
rect 30389 16677 30423 16711
rect 1777 16541 1811 16575
rect 32137 16541 32171 16575
rect 32321 16541 32355 16575
rect 33057 16541 33091 16575
rect 33149 16541 33183 16575
rect 33701 16541 33735 16575
rect 33793 16541 33827 16575
rect 32229 16405 32263 16439
rect 34161 16133 34195 16167
rect 31585 16065 31619 16099
rect 32321 16065 32355 16099
rect 30941 15997 30975 16031
rect 32505 15997 32539 16031
rect 1869 15861 1903 15895
rect 33701 15657 33735 15691
rect 33149 15589 33183 15623
rect 1409 15521 1443 15555
rect 2789 15521 2823 15555
rect 33609 15453 33643 15487
rect 1593 15385 1627 15419
rect 2053 15113 2087 15147
rect 1961 14977 1995 15011
rect 33057 14977 33091 15011
rect 33701 14977 33735 15011
rect 2789 14773 2823 14807
rect 32597 14773 32631 14807
rect 33149 14773 33183 14807
rect 33793 14773 33827 14807
rect 1409 14433 1443 14467
rect 1961 14433 1995 14467
rect 32321 14433 32355 14467
rect 32505 14433 32539 14467
rect 1593 14297 1627 14331
rect 34161 14297 34195 14331
rect 1869 14025 1903 14059
rect 32505 13957 32539 13991
rect 1777 13889 1811 13923
rect 2605 13889 2639 13923
rect 31585 13821 31619 13855
rect 32321 13821 32355 13855
rect 34161 13821 34195 13855
rect 2697 13685 2731 13719
rect 3433 13685 3467 13719
rect 1409 13345 1443 13379
rect 1593 13345 1627 13379
rect 2789 13345 2823 13379
rect 32505 13277 32539 13311
rect 33149 13277 33183 13311
rect 33609 13277 33643 13311
rect 33701 13141 33735 13175
rect 32505 12869 32539 12903
rect 34161 12869 34195 12903
rect 32321 12801 32355 12835
rect 1869 12597 1903 12631
rect 32321 12257 32355 12291
rect 34161 12257 34195 12291
rect 1961 12189 1995 12223
rect 32505 12121 32539 12155
rect 2053 12053 2087 12087
rect 1777 11781 1811 11815
rect 32505 11781 32539 11815
rect 1593 11713 1627 11747
rect 2789 11645 2823 11679
rect 32321 11645 32355 11679
rect 32781 11645 32815 11679
rect 33701 11305 33735 11339
rect 1869 11169 1903 11203
rect 1409 11101 1443 11135
rect 33609 11101 33643 11135
rect 1593 11033 1627 11067
rect 1961 10761 1995 10795
rect 1869 10625 1903 10659
rect 33977 10625 34011 10659
rect 2697 10557 2731 10591
rect 34069 10217 34103 10251
rect 1777 10013 1811 10047
rect 2605 10013 2639 10047
rect 33241 10013 33275 10047
rect 33977 9945 34011 9979
rect 1869 9877 1903 9911
rect 33333 9877 33367 9911
rect 1685 9605 1719 9639
rect 32505 9605 32539 9639
rect 1501 9469 1535 9503
rect 2881 9469 2915 9503
rect 32321 9469 32355 9503
rect 34161 9469 34195 9503
rect 33977 9129 34011 9163
rect 2789 8993 2823 9027
rect 1409 8925 1443 8959
rect 1593 8857 1627 8891
rect 1961 8585 1995 8619
rect 1869 8449 1903 8483
rect 2697 8449 2731 8483
rect 2053 8041 2087 8075
rect 1961 7837 1995 7871
rect 2789 7837 2823 7871
rect 33977 7837 34011 7871
rect 1593 7361 1627 7395
rect 1777 7293 1811 7327
rect 2789 7293 2823 7327
rect 4077 7157 4111 7191
rect 33333 7157 33367 7191
rect 33977 7157 34011 7191
rect 2053 6953 2087 6987
rect 32321 6817 32355 6851
rect 34161 6817 34195 6851
rect 1961 6749 1995 6783
rect 2789 6749 2823 6783
rect 3801 6749 3835 6783
rect 31861 6749 31895 6783
rect 32505 6681 32539 6715
rect 3893 6613 3927 6647
rect 33701 6409 33735 6443
rect 32965 6273 32999 6307
rect 33609 6273 33643 6307
rect 2053 6205 2087 6239
rect 2237 6205 2271 6239
rect 3249 6205 3283 6239
rect 1593 6069 1627 6103
rect 4537 6069 4571 6103
rect 5181 6069 5215 6103
rect 31585 6069 31619 6103
rect 32505 6069 32539 6103
rect 33057 6069 33091 6103
rect 31217 5865 31251 5899
rect 1409 5729 1443 5763
rect 1869 5729 1903 5763
rect 3801 5729 3835 5763
rect 3985 5729 4019 5763
rect 4261 5729 4295 5763
rect 31677 5729 31711 5763
rect 33149 5729 33183 5763
rect 6285 5661 6319 5695
rect 30573 5661 30607 5695
rect 33977 5661 34011 5695
rect 1593 5593 1627 5627
rect 31861 5593 31895 5627
rect 34069 5525 34103 5559
rect 1869 5321 1903 5355
rect 31493 5253 31527 5287
rect 32505 5253 32539 5287
rect 1777 5185 1811 5219
rect 2605 5185 2639 5219
rect 6561 5185 6595 5219
rect 29469 5185 29503 5219
rect 30757 5185 30791 5219
rect 31401 5185 31435 5219
rect 2789 5117 2823 5151
rect 3065 5117 3099 5151
rect 32321 5117 32355 5151
rect 34161 5117 34195 5151
rect 5089 4981 5123 5015
rect 5733 4981 5767 5015
rect 29561 4981 29595 5015
rect 30297 4981 30331 5015
rect 30849 4981 30883 5015
rect 3893 4777 3927 4811
rect 2789 4641 2823 4675
rect 5181 4641 5215 4675
rect 5641 4641 5675 4675
rect 29837 4641 29871 4675
rect 30021 4641 30055 4675
rect 30941 4641 30975 4675
rect 32321 4641 32355 4675
rect 32505 4641 32539 4675
rect 1869 4573 1903 4607
rect 2697 4573 2731 4607
rect 3801 4573 3835 4607
rect 4445 4573 4479 4607
rect 8033 4573 8067 4607
rect 9873 4573 9907 4607
rect 10517 4573 10551 4607
rect 5365 4505 5399 4539
rect 34161 4505 34195 4539
rect 1961 4437 1995 4471
rect 4537 4437 4571 4471
rect 29929 4165 29963 4199
rect 4077 4097 4111 4131
rect 4721 4097 4755 4131
rect 7757 4097 7791 4131
rect 10241 4097 10275 4131
rect 20545 4097 20579 4131
rect 29101 4097 29135 4131
rect 29193 4097 29227 4131
rect 29745 4097 29779 4131
rect 32137 4097 32171 4131
rect 1777 4029 1811 4063
rect 1961 4029 1995 4063
rect 2881 4029 2915 4063
rect 6561 4029 6595 4063
rect 7941 4029 7975 4063
rect 8401 4029 8435 4063
rect 31585 4029 31619 4063
rect 32321 4029 32355 4063
rect 33057 4029 33091 4063
rect 4169 3961 4203 3995
rect 20361 3961 20395 3995
rect 4813 3893 4847 3927
rect 5549 3893 5583 3927
rect 7205 3893 7239 3927
rect 10333 3893 10367 3927
rect 14565 3893 14599 3927
rect 15761 3893 15795 3927
rect 19717 3893 19751 3927
rect 21281 3893 21315 3927
rect 28641 3893 28675 3927
rect 8033 3689 8067 3723
rect 28917 3689 28951 3723
rect 27721 3621 27755 3655
rect 1409 3553 1443 3587
rect 1593 3553 1627 3587
rect 1869 3553 1903 3587
rect 4445 3553 4479 3587
rect 4629 3553 4663 3587
rect 5181 3553 5215 3587
rect 6929 3553 6963 3587
rect 9597 3553 9631 3587
rect 9781 3553 9815 3587
rect 10057 3553 10091 3587
rect 15485 3553 15519 3587
rect 16129 3553 16163 3587
rect 20821 3553 20855 3587
rect 22201 3553 22235 3587
rect 28365 3553 28399 3587
rect 30481 3553 30515 3587
rect 32321 3553 32355 3587
rect 3801 3485 3835 3519
rect 7941 3485 7975 3519
rect 8953 3485 8987 3519
rect 12081 3485 12115 3519
rect 13185 3485 13219 3519
rect 14289 3485 14323 3519
rect 17969 3485 18003 3519
rect 19441 3485 19475 3519
rect 20361 3485 20395 3519
rect 24593 3485 24627 3519
rect 28825 3485 28859 3519
rect 29561 3485 29595 3519
rect 32965 3485 32999 3519
rect 15669 3417 15703 3451
rect 21005 3417 21039 3451
rect 29837 3417 29871 3451
rect 30665 3417 30699 3451
rect 33793 3417 33827 3451
rect 3893 3349 3927 3383
rect 9045 3349 9079 3383
rect 14381 3349 14415 3383
rect 19533 3349 19567 3383
rect 21925 3145 21959 3179
rect 29101 3145 29135 3179
rect 2513 3077 2547 3111
rect 5733 3077 5767 3111
rect 6561 3077 6595 3111
rect 14473 3077 14507 3111
rect 23305 3077 23339 3111
rect 24041 3077 24075 3111
rect 32505 3077 32539 3111
rect 1685 3009 1719 3043
rect 2329 3009 2363 3043
rect 4629 3009 4663 3043
rect 5641 3009 5675 3043
rect 6377 3009 6411 3043
rect 9137 3009 9171 3043
rect 11989 3009 12023 3043
rect 14289 3009 14323 3043
rect 16865 3009 16899 3043
rect 19441 3009 19475 3043
rect 21833 3009 21867 3043
rect 23213 3009 23247 3043
rect 23857 3009 23891 3043
rect 27721 3009 27755 3043
rect 28365 3009 28399 3043
rect 29009 3009 29043 3043
rect 29653 3009 29687 3043
rect 2789 2941 2823 2975
rect 6837 2941 6871 2975
rect 9321 2941 9355 2975
rect 9689 2941 9723 2975
rect 12173 2941 12207 2975
rect 13553 2941 13587 2975
rect 14841 2941 14875 2975
rect 17049 2941 17083 2975
rect 17417 2941 17451 2975
rect 19625 2941 19659 2975
rect 20637 2941 20671 2975
rect 24501 2941 24535 2975
rect 28457 2941 28491 2975
rect 29837 2941 29871 2975
rect 30297 2941 30331 2975
rect 32321 2941 32355 2975
rect 34161 2941 34195 2975
rect 1777 2805 1811 2839
rect 4721 2805 4755 2839
rect 27813 2805 27847 2839
rect 13277 2601 13311 2635
rect 15853 2601 15887 2635
rect 16957 2601 16991 2635
rect 18337 2601 18371 2635
rect 21925 2601 21959 2635
rect 28917 2601 28951 2635
rect 1593 2465 1627 2499
rect 2789 2465 2823 2499
rect 3893 2465 3927 2499
rect 4077 2465 4111 2499
rect 4813 2465 4847 2499
rect 6377 2465 6411 2499
rect 7021 2465 7055 2499
rect 9137 2465 9171 2499
rect 9321 2465 9355 2499
rect 10333 2465 10367 2499
rect 14197 2465 14231 2499
rect 19441 2465 19475 2499
rect 19625 2465 19659 2499
rect 19993 2465 20027 2499
rect 29745 2465 29779 2499
rect 29929 2465 29963 2499
rect 31585 2465 31619 2499
rect 1409 2397 1443 2431
rect 13185 2397 13219 2431
rect 14105 2397 14139 2431
rect 15761 2397 15795 2431
rect 16865 2397 16899 2431
rect 21833 2397 21867 2431
rect 28825 2397 28859 2431
rect 32321 2397 32355 2431
rect 6561 2329 6595 2363
rect 18245 2329 18279 2363
rect 32505 2329 32539 2363
rect 34161 2329 34195 2363
<< metal1 >>
rect 13630 40876 13636 40928
rect 13688 40916 13694 40928
rect 20162 40916 20168 40928
rect 13688 40888 20168 40916
rect 13688 40876 13694 40888
rect 20162 40876 20168 40888
rect 20220 40876 20226 40928
rect 12066 40808 12072 40860
rect 12124 40848 12130 40860
rect 30374 40848 30380 40860
rect 12124 40820 30380 40848
rect 12124 40808 12130 40820
rect 30374 40808 30380 40820
rect 30432 40808 30438 40860
rect 4430 40740 4436 40792
rect 4488 40780 4494 40792
rect 18598 40780 18604 40792
rect 4488 40752 18604 40780
rect 4488 40740 4494 40752
rect 18598 40740 18604 40752
rect 18656 40740 18662 40792
rect 14734 40672 14740 40724
rect 14792 40712 14798 40724
rect 19886 40712 19892 40724
rect 14792 40684 19892 40712
rect 14792 40672 14798 40684
rect 19886 40672 19892 40684
rect 19944 40672 19950 40724
rect 11698 40604 11704 40656
rect 11756 40644 11762 40656
rect 11756 40616 12434 40644
rect 11756 40604 11762 40616
rect 12406 40304 12434 40616
rect 12986 40604 12992 40656
rect 13044 40644 13050 40656
rect 26418 40644 26424 40656
rect 13044 40616 26424 40644
rect 13044 40604 13050 40616
rect 26418 40604 26424 40616
rect 26476 40604 26482 40656
rect 12618 40536 12624 40588
rect 12676 40576 12682 40588
rect 31846 40576 31852 40588
rect 12676 40548 31852 40576
rect 12676 40536 12682 40548
rect 31846 40536 31852 40548
rect 31904 40536 31910 40588
rect 16022 40468 16028 40520
rect 16080 40508 16086 40520
rect 29914 40508 29920 40520
rect 16080 40480 29920 40508
rect 16080 40468 16086 40480
rect 29914 40468 29920 40480
rect 29972 40468 29978 40520
rect 15378 40400 15384 40452
rect 15436 40440 15442 40452
rect 30098 40440 30104 40452
rect 15436 40412 30104 40440
rect 15436 40400 15442 40412
rect 30098 40400 30104 40412
rect 30156 40400 30162 40452
rect 14458 40332 14464 40384
rect 14516 40372 14522 40384
rect 30282 40372 30288 40384
rect 14516 40344 30288 40372
rect 14516 40332 14522 40344
rect 30282 40332 30288 40344
rect 30340 40332 30346 40384
rect 30006 40304 30012 40316
rect 12406 40276 30012 40304
rect 30006 40264 30012 40276
rect 30064 40264 30070 40316
rect 15838 40196 15844 40248
rect 15896 40236 15902 40248
rect 19794 40236 19800 40248
rect 15896 40208 19800 40236
rect 15896 40196 15902 40208
rect 19794 40196 19800 40208
rect 19852 40196 19858 40248
rect 19886 40196 19892 40248
rect 19944 40236 19950 40248
rect 27246 40236 27252 40248
rect 19944 40208 27252 40236
rect 19944 40196 19950 40208
rect 27246 40196 27252 40208
rect 27304 40196 27310 40248
rect 13538 40128 13544 40180
rect 13596 40168 13602 40180
rect 31938 40168 31944 40180
rect 13596 40140 31944 40168
rect 13596 40128 13602 40140
rect 31938 40128 31944 40140
rect 31996 40128 32002 40180
rect 12710 40060 12716 40112
rect 12768 40100 12774 40112
rect 15930 40100 15936 40112
rect 12768 40072 15936 40100
rect 12768 40060 12774 40072
rect 15930 40060 15936 40072
rect 15988 40100 15994 40112
rect 19610 40100 19616 40112
rect 15988 40072 19616 40100
rect 15988 40060 15994 40072
rect 19610 40060 19616 40072
rect 19668 40060 19674 40112
rect 11790 39992 11796 40044
rect 11848 40032 11854 40044
rect 19242 40032 19248 40044
rect 11848 40004 19248 40032
rect 11848 39992 11854 40004
rect 19242 39992 19248 40004
rect 19300 39992 19306 40044
rect 22646 39992 22652 40044
rect 22704 40032 22710 40044
rect 29638 40032 29644 40044
rect 22704 40004 29644 40032
rect 22704 39992 22710 40004
rect 29638 39992 29644 40004
rect 29696 39992 29702 40044
rect 12250 39924 12256 39976
rect 12308 39964 12314 39976
rect 22186 39964 22192 39976
rect 12308 39936 22192 39964
rect 12308 39924 12314 39936
rect 22186 39924 22192 39936
rect 22244 39924 22250 39976
rect 23750 39924 23756 39976
rect 23808 39964 23814 39976
rect 32490 39964 32496 39976
rect 23808 39936 32496 39964
rect 23808 39924 23814 39936
rect 32490 39924 32496 39936
rect 32548 39924 32554 39976
rect 13906 39856 13912 39908
rect 13964 39896 13970 39908
rect 18874 39896 18880 39908
rect 13964 39868 18880 39896
rect 13964 39856 13970 39868
rect 18874 39856 18880 39868
rect 18932 39856 18938 39908
rect 18966 39856 18972 39908
rect 19024 39896 19030 39908
rect 26694 39896 26700 39908
rect 19024 39868 26700 39896
rect 19024 39856 19030 39868
rect 26694 39856 26700 39868
rect 26752 39856 26758 39908
rect 12894 39788 12900 39840
rect 12952 39828 12958 39840
rect 17770 39828 17776 39840
rect 12952 39800 17776 39828
rect 12952 39788 12958 39800
rect 17770 39788 17776 39800
rect 17828 39788 17834 39840
rect 20806 39788 20812 39840
rect 20864 39828 20870 39840
rect 27890 39828 27896 39840
rect 20864 39800 27896 39828
rect 20864 39788 20870 39800
rect 27890 39788 27896 39800
rect 27948 39788 27954 39840
rect 1104 39738 34868 39760
rect 1104 39686 6582 39738
rect 6634 39686 6646 39738
rect 6698 39686 6710 39738
rect 6762 39686 6774 39738
rect 6826 39686 6838 39738
rect 6890 39686 17846 39738
rect 17898 39686 17910 39738
rect 17962 39686 17974 39738
rect 18026 39686 18038 39738
rect 18090 39686 18102 39738
rect 18154 39686 29110 39738
rect 29162 39686 29174 39738
rect 29226 39686 29238 39738
rect 29290 39686 29302 39738
rect 29354 39686 29366 39738
rect 29418 39686 34868 39738
rect 1104 39664 34868 39686
rect 10318 39624 10324 39636
rect 10279 39596 10324 39624
rect 10318 39584 10324 39596
rect 10376 39584 10382 39636
rect 12820 39596 15976 39624
rect 8294 39556 8300 39568
rect 1688 39528 8300 39556
rect 1688 39497 1716 39528
rect 8294 39516 8300 39528
rect 8352 39516 8358 39568
rect 8389 39559 8447 39565
rect 8389 39525 8401 39559
rect 8435 39556 8447 39559
rect 9582 39556 9588 39568
rect 8435 39528 9588 39556
rect 8435 39525 8447 39528
rect 8389 39519 8447 39525
rect 9582 39516 9588 39528
rect 9640 39516 9646 39568
rect 12250 39556 12256 39568
rect 12211 39528 12256 39556
rect 12250 39516 12256 39528
rect 12308 39516 12314 39568
rect 1673 39491 1731 39497
rect 1673 39457 1685 39491
rect 1719 39457 1731 39491
rect 1673 39451 1731 39457
rect 4982 39448 4988 39500
rect 5040 39488 5046 39500
rect 12820 39488 12848 39596
rect 15948 39504 15976 39596
rect 16390 39584 16396 39636
rect 16448 39624 16454 39636
rect 17310 39624 17316 39636
rect 16448 39596 17316 39624
rect 16448 39584 16454 39596
rect 17310 39584 17316 39596
rect 17368 39584 17374 39636
rect 19058 39584 19064 39636
rect 19116 39624 19122 39636
rect 23750 39624 23756 39636
rect 19116 39596 23612 39624
rect 23711 39596 23756 39624
rect 19116 39584 19122 39596
rect 16298 39516 16304 39568
rect 16356 39556 16362 39568
rect 23584 39556 23612 39596
rect 23750 39584 23756 39596
rect 23808 39584 23814 39636
rect 25682 39624 25688 39636
rect 25148 39596 25688 39624
rect 25148 39556 25176 39596
rect 25682 39584 25688 39596
rect 25740 39624 25746 39636
rect 26234 39624 26240 39636
rect 25740 39596 26240 39624
rect 25740 39584 25746 39596
rect 26234 39584 26240 39596
rect 26292 39584 26298 39636
rect 26418 39624 26424 39636
rect 26379 39596 26424 39624
rect 26418 39584 26424 39596
rect 26476 39584 26482 39636
rect 26510 39584 26516 39636
rect 26568 39624 26574 39636
rect 31570 39624 31576 39636
rect 26568 39596 31576 39624
rect 26568 39584 26574 39596
rect 31570 39584 31576 39596
rect 31628 39584 31634 39636
rect 16356 39528 23244 39556
rect 23584 39528 25176 39556
rect 16356 39516 16362 39528
rect 5040 39460 12848 39488
rect 5040 39448 5046 39460
rect 13538 39448 13544 39500
rect 13596 39488 13602 39500
rect 13596 39460 13641 39488
rect 15948 39476 16068 39504
rect 16666 39488 16672 39500
rect 13596 39448 13602 39460
rect 1394 39420 1400 39432
rect 1355 39392 1400 39420
rect 1394 39380 1400 39392
rect 1452 39380 1458 39432
rect 3053 39423 3111 39429
rect 3053 39389 3065 39423
rect 3099 39389 3111 39423
rect 3053 39383 3111 39389
rect 3068 39352 3096 39383
rect 3602 39380 3608 39432
rect 3660 39420 3666 39432
rect 3789 39423 3847 39429
rect 3789 39420 3801 39423
rect 3660 39392 3801 39420
rect 3660 39380 3666 39392
rect 3789 39389 3801 39392
rect 3835 39420 3847 39423
rect 4062 39420 4068 39432
rect 3835 39392 4068 39420
rect 3835 39389 3847 39392
rect 3789 39383 3847 39389
rect 4062 39380 4068 39392
rect 4120 39380 4126 39432
rect 4614 39420 4620 39432
rect 4575 39392 4620 39420
rect 4614 39380 4620 39392
rect 4672 39380 4678 39432
rect 5258 39420 5264 39432
rect 5219 39392 5264 39420
rect 5258 39380 5264 39392
rect 5316 39380 5322 39432
rect 5350 39380 5356 39432
rect 5408 39420 5414 39432
rect 6549 39423 6607 39429
rect 6549 39420 6561 39423
rect 5408 39392 6561 39420
rect 5408 39380 5414 39392
rect 6549 39389 6561 39392
rect 6595 39389 6607 39423
rect 6549 39383 6607 39389
rect 7190 39380 7196 39432
rect 7248 39420 7254 39432
rect 7377 39423 7435 39429
rect 7377 39420 7389 39423
rect 7248 39392 7389 39420
rect 7248 39380 7254 39392
rect 7377 39389 7389 39392
rect 7423 39389 7435 39423
rect 7377 39383 7435 39389
rect 8570 39380 8576 39432
rect 8628 39420 8634 39432
rect 9125 39423 9183 39429
rect 9125 39420 9137 39423
rect 8628 39392 9137 39420
rect 8628 39380 8634 39392
rect 9125 39389 9137 39392
rect 9171 39389 9183 39423
rect 10962 39420 10968 39432
rect 10923 39392 10968 39420
rect 9125 39383 9183 39389
rect 10962 39380 10968 39392
rect 11020 39380 11026 39432
rect 12897 39423 12955 39429
rect 12897 39389 12909 39423
rect 12943 39420 12955 39423
rect 13446 39420 13452 39432
rect 12943 39392 13452 39420
rect 12943 39389 12955 39392
rect 12897 39383 12955 39389
rect 13446 39380 13452 39392
rect 13504 39380 13510 39432
rect 13814 39380 13820 39432
rect 13872 39420 13878 39432
rect 14458 39420 14464 39432
rect 13872 39392 14464 39420
rect 13872 39380 13878 39392
rect 14458 39380 14464 39392
rect 14516 39380 14522 39432
rect 14918 39380 14924 39432
rect 14976 39420 14982 39432
rect 15105 39423 15163 39429
rect 15105 39420 15117 39423
rect 14976 39392 15117 39420
rect 14976 39380 14982 39392
rect 15105 39389 15117 39392
rect 15151 39389 15163 39423
rect 15105 39383 15163 39389
rect 15194 39380 15200 39432
rect 15252 39420 15258 39432
rect 15749 39423 15807 39429
rect 15749 39420 15761 39423
rect 15252 39392 15761 39420
rect 15252 39380 15258 39392
rect 15749 39389 15761 39392
rect 15795 39389 15807 39423
rect 15749 39383 15807 39389
rect 15933 39423 15991 39429
rect 15933 39389 15945 39423
rect 15979 39414 15991 39423
rect 16040 39414 16068 39476
rect 16627 39460 16672 39488
rect 16666 39448 16672 39460
rect 16724 39448 16730 39500
rect 17402 39488 17408 39500
rect 17363 39460 17408 39488
rect 17402 39448 17408 39460
rect 17460 39448 17466 39500
rect 17494 39448 17500 39500
rect 17552 39488 17558 39500
rect 19429 39491 19487 39497
rect 19429 39488 19441 39491
rect 17552 39460 19441 39488
rect 17552 39448 17558 39460
rect 19429 39457 19441 39460
rect 19475 39457 19487 39491
rect 19978 39488 19984 39500
rect 19939 39460 19984 39488
rect 19429 39451 19487 39457
rect 19978 39448 19984 39460
rect 20036 39448 20042 39500
rect 23216 39488 23244 39528
rect 25222 39516 25228 39568
rect 25280 39556 25286 39568
rect 25317 39559 25375 39565
rect 25317 39556 25329 39559
rect 25280 39528 25329 39556
rect 25280 39516 25286 39528
rect 25317 39525 25329 39528
rect 25363 39525 25375 39559
rect 25317 39519 25375 39525
rect 26786 39516 26792 39568
rect 26844 39556 26850 39568
rect 30190 39556 30196 39568
rect 26844 39528 30196 39556
rect 26844 39516 26850 39528
rect 30190 39516 30196 39528
rect 30248 39516 30254 39568
rect 25516 39488 25728 39504
rect 23216 39476 26464 39488
rect 23216 39460 25544 39476
rect 25700 39460 26464 39476
rect 25593 39433 25651 39439
rect 15979 39389 16068 39414
rect 15933 39386 16068 39389
rect 15933 39383 15991 39386
rect 18046 39380 18052 39432
rect 18104 39420 18110 39432
rect 19334 39420 19340 39432
rect 18104 39392 19340 39420
rect 18104 39380 18110 39392
rect 19334 39380 19340 39392
rect 19392 39380 19398 39432
rect 21910 39420 21916 39432
rect 21871 39392 21916 39420
rect 21910 39380 21916 39392
rect 21968 39380 21974 39432
rect 22002 39380 22008 39432
rect 22060 39420 22066 39432
rect 22646 39420 22652 39432
rect 22060 39392 22105 39420
rect 22607 39392 22652 39420
rect 22060 39380 22066 39392
rect 22646 39380 22652 39392
rect 22704 39380 22710 39432
rect 23658 39420 23664 39432
rect 23619 39392 23664 39420
rect 23658 39380 23664 39392
rect 23716 39380 23722 39432
rect 24578 39420 24584 39432
rect 24539 39392 24584 39420
rect 24578 39380 24584 39392
rect 24636 39380 24642 39432
rect 24688 39392 25452 39420
rect 25593 39399 25605 39433
rect 25639 39430 25651 39433
rect 25639 39420 25728 39430
rect 26142 39420 26148 39432
rect 25639 39402 26004 39420
rect 25639 39399 25651 39402
rect 25593 39393 25651 39399
rect 25700 39392 26004 39402
rect 26103 39392 26148 39420
rect 7006 39352 7012 39364
rect 3068 39324 7012 39352
rect 7006 39312 7012 39324
rect 7064 39312 7070 39364
rect 7926 39312 7932 39364
rect 7984 39352 7990 39364
rect 12710 39352 12716 39364
rect 7984 39324 12716 39352
rect 7984 39312 7990 39324
rect 12710 39312 12716 39324
rect 12768 39312 12774 39364
rect 14553 39355 14611 39361
rect 14553 39321 14565 39355
rect 14599 39352 14611 39355
rect 15654 39352 15660 39364
rect 14599 39324 15660 39352
rect 14599 39321 14611 39324
rect 14553 39315 14611 39321
rect 15654 39312 15660 39324
rect 15712 39312 15718 39364
rect 16114 39352 16120 39364
rect 16075 39324 16120 39352
rect 16114 39312 16120 39324
rect 16172 39312 16178 39364
rect 16574 39312 16580 39364
rect 16632 39352 16638 39364
rect 16853 39355 16911 39361
rect 16853 39352 16865 39355
rect 16632 39324 16865 39352
rect 16632 39312 16638 39324
rect 16853 39321 16865 39324
rect 16899 39321 16911 39355
rect 16853 39315 16911 39321
rect 17310 39312 17316 39364
rect 17368 39352 17374 39364
rect 18782 39352 18788 39364
rect 17368 39324 18788 39352
rect 17368 39312 17374 39324
rect 18782 39312 18788 39324
rect 18840 39312 18846 39364
rect 19426 39312 19432 39364
rect 19484 39352 19490 39364
rect 19613 39355 19671 39361
rect 19613 39352 19625 39355
rect 19484 39324 19625 39352
rect 19484 39312 19490 39324
rect 19613 39321 19625 39324
rect 19659 39321 19671 39355
rect 19613 39315 19671 39321
rect 20438 39312 20444 39364
rect 20496 39352 20502 39364
rect 22741 39355 22799 39361
rect 22741 39352 22753 39355
rect 20496 39324 22753 39352
rect 20496 39312 20502 39324
rect 22741 39321 22753 39324
rect 22787 39321 22799 39355
rect 22741 39315 22799 39321
rect 22830 39312 22836 39364
rect 22888 39352 22894 39364
rect 24688 39352 24716 39392
rect 22888 39324 24716 39352
rect 25317 39355 25375 39361
rect 22888 39312 22894 39324
rect 25317 39321 25329 39355
rect 25363 39321 25375 39355
rect 25424 39352 25452 39392
rect 25501 39355 25559 39361
rect 25501 39352 25513 39355
rect 25424 39324 25513 39352
rect 25317 39315 25375 39321
rect 25501 39321 25513 39324
rect 25547 39321 25559 39355
rect 25976 39352 26004 39392
rect 26142 39380 26148 39392
rect 26200 39380 26206 39432
rect 26234 39380 26240 39432
rect 26292 39420 26298 39432
rect 26292 39392 26337 39420
rect 26292 39380 26298 39392
rect 26050 39352 26056 39364
rect 25976 39324 26056 39352
rect 25501 39315 25559 39321
rect 3142 39284 3148 39296
rect 3103 39256 3148 39284
rect 3142 39244 3148 39256
rect 3200 39244 3206 39296
rect 3234 39244 3240 39296
rect 3292 39284 3298 39296
rect 3881 39287 3939 39293
rect 3881 39284 3893 39287
rect 3292 39256 3893 39284
rect 3292 39244 3298 39256
rect 3881 39253 3893 39256
rect 3927 39253 3939 39287
rect 15194 39284 15200 39296
rect 15155 39256 15200 39284
rect 3881 39247 3939 39253
rect 15194 39244 15200 39256
rect 15252 39244 15258 39296
rect 15562 39244 15568 39296
rect 15620 39284 15626 39296
rect 16390 39284 16396 39296
rect 15620 39256 16396 39284
rect 15620 39244 15626 39256
rect 16390 39244 16396 39256
rect 16448 39244 16454 39296
rect 16482 39244 16488 39296
rect 16540 39284 16546 39296
rect 18966 39284 18972 39296
rect 16540 39256 18972 39284
rect 16540 39244 16546 39256
rect 18966 39244 18972 39256
rect 19024 39244 19030 39296
rect 20714 39244 20720 39296
rect 20772 39284 20778 39296
rect 22189 39287 22247 39293
rect 22189 39284 22201 39287
rect 20772 39256 22201 39284
rect 20772 39244 20778 39256
rect 22189 39253 22201 39256
rect 22235 39253 22247 39287
rect 22189 39247 22247 39253
rect 23842 39244 23848 39296
rect 23900 39284 23906 39296
rect 24765 39287 24823 39293
rect 24765 39284 24777 39287
rect 23900 39256 24777 39284
rect 23900 39244 23906 39256
rect 24765 39253 24777 39256
rect 24811 39253 24823 39287
rect 25332 39284 25360 39315
rect 26050 39312 26056 39324
rect 26108 39312 26114 39364
rect 26436 39352 26464 39460
rect 27154 39448 27160 39500
rect 27212 39488 27218 39500
rect 27433 39491 27491 39497
rect 27433 39488 27445 39491
rect 27212 39460 27445 39488
rect 27212 39448 27218 39460
rect 27433 39457 27445 39460
rect 27479 39457 27491 39491
rect 27433 39451 27491 39457
rect 30466 39448 30472 39500
rect 30524 39488 30530 39500
rect 30745 39491 30803 39497
rect 30524 39460 30696 39488
rect 30524 39448 30530 39460
rect 26970 39420 26976 39432
rect 26931 39392 26976 39420
rect 26970 39380 26976 39392
rect 27028 39380 27034 39432
rect 30668 39429 30696 39460
rect 30745 39457 30757 39491
rect 30791 39488 30803 39491
rect 32493 39491 32551 39497
rect 32493 39488 32505 39491
rect 30791 39460 32505 39488
rect 30791 39457 30803 39460
rect 30745 39451 30803 39457
rect 32493 39457 32505 39460
rect 32539 39457 32551 39491
rect 34146 39488 34152 39500
rect 34107 39460 34152 39488
rect 32493 39451 32551 39457
rect 34146 39448 34152 39460
rect 34204 39448 34210 39500
rect 30653 39423 30711 39429
rect 28828 39392 30604 39420
rect 27157 39355 27215 39361
rect 27157 39352 27169 39355
rect 26436 39324 27169 39352
rect 27157 39321 27169 39324
rect 27203 39321 27215 39355
rect 27157 39315 27215 39321
rect 28828 39284 28856 39392
rect 29454 39312 29460 39364
rect 29512 39352 29518 39364
rect 30009 39355 30067 39361
rect 30009 39352 30021 39355
rect 29512 39324 30021 39352
rect 29512 39312 29518 39324
rect 30009 39321 30021 39324
rect 30055 39321 30067 39355
rect 30576 39352 30604 39392
rect 30653 39389 30665 39423
rect 30699 39389 30711 39423
rect 30653 39383 30711 39389
rect 30834 39380 30840 39432
rect 30892 39420 30898 39432
rect 31389 39423 31447 39429
rect 31389 39420 31401 39423
rect 30892 39392 31401 39420
rect 30892 39380 30898 39392
rect 31389 39389 31401 39392
rect 31435 39389 31447 39423
rect 32306 39420 32312 39432
rect 32267 39392 32312 39420
rect 31389 39383 31447 39389
rect 32306 39380 32312 39392
rect 32364 39380 32370 39432
rect 30926 39352 30932 39364
rect 30576 39324 30932 39352
rect 30009 39315 30067 39321
rect 30926 39312 30932 39324
rect 30984 39312 30990 39364
rect 25332 39256 28856 39284
rect 24765 39247 24823 39253
rect 28902 39244 28908 39296
rect 28960 39284 28966 39296
rect 30101 39287 30159 39293
rect 30101 39284 30113 39287
rect 28960 39256 30113 39284
rect 28960 39244 28966 39256
rect 30101 39253 30113 39256
rect 30147 39253 30159 39287
rect 30101 39247 30159 39253
rect 30834 39244 30840 39296
rect 30892 39284 30898 39296
rect 31481 39287 31539 39293
rect 31481 39284 31493 39287
rect 30892 39256 31493 39284
rect 30892 39244 30898 39256
rect 31481 39253 31493 39256
rect 31527 39253 31539 39287
rect 31481 39247 31539 39253
rect 1104 39194 34868 39216
rect 1104 39142 12214 39194
rect 12266 39142 12278 39194
rect 12330 39142 12342 39194
rect 12394 39142 12406 39194
rect 12458 39142 12470 39194
rect 12522 39142 23478 39194
rect 23530 39142 23542 39194
rect 23594 39142 23606 39194
rect 23658 39142 23670 39194
rect 23722 39142 23734 39194
rect 23786 39142 34868 39194
rect 1104 39120 34868 39142
rect 4614 39080 4620 39092
rect 1504 39052 4620 39080
rect 1504 38953 1532 39052
rect 4614 39040 4620 39052
rect 4672 39040 4678 39092
rect 12894 39080 12900 39092
rect 6886 39052 12756 39080
rect 12855 39052 12900 39080
rect 3142 38972 3148 39024
rect 3200 39012 3206 39024
rect 3973 39015 4031 39021
rect 3973 39012 3985 39015
rect 3200 38984 3985 39012
rect 3200 38972 3206 38984
rect 3973 38981 3985 38984
rect 4019 38981 4031 39015
rect 3973 38975 4031 38981
rect 4062 38972 4068 39024
rect 4120 39012 4126 39024
rect 6886 39012 6914 39052
rect 4120 38984 6914 39012
rect 8021 39015 8079 39021
rect 4120 38972 4126 38984
rect 8021 38981 8033 39015
rect 8067 39012 8079 39015
rect 8757 39015 8815 39021
rect 8757 39012 8769 39015
rect 8067 38984 8769 39012
rect 8067 38981 8079 38984
rect 8021 38975 8079 38981
rect 8757 38981 8769 38984
rect 8803 38981 8815 39015
rect 8757 38975 8815 38981
rect 1489 38947 1547 38953
rect 1489 38913 1501 38947
rect 1535 38913 1547 38947
rect 1489 38907 1547 38913
rect 7285 38947 7343 38953
rect 7285 38913 7297 38947
rect 7331 38913 7343 38947
rect 7926 38944 7932 38956
rect 7887 38916 7932 38944
rect 7285 38907 7343 38913
rect 1670 38876 1676 38888
rect 1631 38848 1676 38876
rect 1670 38836 1676 38848
rect 1728 38836 1734 38888
rect 1949 38879 2007 38885
rect 1949 38845 1961 38879
rect 1995 38845 2007 38879
rect 1949 38839 2007 38845
rect 3789 38879 3847 38885
rect 3789 38845 3801 38879
rect 3835 38876 3847 38879
rect 5350 38876 5356 38888
rect 3835 38848 5356 38876
rect 3835 38845 3847 38848
rect 3789 38839 3847 38845
rect 658 38768 664 38820
rect 716 38808 722 38820
rect 1964 38808 1992 38839
rect 5350 38836 5356 38848
rect 5408 38836 5414 38888
rect 5445 38879 5503 38885
rect 5445 38845 5457 38879
rect 5491 38845 5503 38879
rect 5445 38839 5503 38845
rect 716 38780 1992 38808
rect 716 38768 722 38780
rect 4154 38768 4160 38820
rect 4212 38808 4218 38820
rect 5460 38808 5488 38839
rect 7006 38836 7012 38888
rect 7064 38876 7070 38888
rect 7300 38876 7328 38907
rect 7926 38904 7932 38916
rect 7984 38904 7990 38956
rect 8570 38944 8576 38956
rect 8531 38916 8576 38944
rect 8570 38904 8576 38916
rect 8628 38904 8634 38956
rect 11790 38944 11796 38956
rect 11751 38916 11796 38944
rect 11790 38904 11796 38916
rect 11848 38904 11854 38956
rect 12437 38947 12495 38953
rect 12437 38913 12449 38947
rect 12483 38944 12495 38947
rect 12618 38944 12624 38956
rect 12483 38916 12624 38944
rect 12483 38913 12495 38916
rect 12437 38907 12495 38913
rect 12618 38904 12624 38916
rect 12676 38904 12682 38956
rect 9214 38876 9220 38888
rect 7064 38848 9220 38876
rect 7064 38836 7070 38848
rect 9214 38836 9220 38848
rect 9272 38836 9278 38888
rect 9306 38836 9312 38888
rect 9364 38876 9370 38888
rect 12728 38876 12756 39052
rect 12894 39040 12900 39052
rect 12952 39040 12958 39092
rect 13446 39040 13452 39092
rect 13504 39080 13510 39092
rect 13633 39083 13691 39089
rect 13633 39080 13645 39083
rect 13504 39052 13645 39080
rect 13504 39040 13510 39052
rect 13633 39049 13645 39052
rect 13679 39049 13691 39083
rect 13633 39043 13691 39049
rect 13722 39040 13728 39092
rect 13780 39080 13786 39092
rect 14918 39080 14924 39092
rect 13780 39052 14924 39080
rect 13780 39040 13786 39052
rect 14918 39040 14924 39052
rect 14976 39040 14982 39092
rect 15194 39040 15200 39092
rect 15252 39080 15258 39092
rect 15252 39052 18644 39080
rect 15252 39040 15258 39052
rect 16114 39012 16120 39024
rect 13096 38984 16120 39012
rect 13096 38953 13124 38984
rect 16114 38972 16120 38984
rect 16172 38972 16178 39024
rect 18046 39012 18052 39024
rect 16684 38984 17172 39012
rect 13081 38947 13139 38953
rect 13081 38913 13093 38947
rect 13127 38913 13139 38947
rect 13081 38907 13139 38913
rect 13541 38947 13599 38953
rect 13541 38913 13553 38947
rect 13587 38944 13599 38947
rect 13814 38944 13820 38956
rect 13587 38916 13820 38944
rect 13587 38913 13599 38916
rect 13541 38907 13599 38913
rect 13556 38876 13584 38907
rect 13814 38904 13820 38916
rect 13872 38904 13878 38956
rect 16684 38953 16712 38984
rect 17144 38956 17172 38984
rect 17236 38984 18052 39012
rect 16669 38947 16727 38953
rect 16669 38944 16681 38947
rect 15580 38916 16681 38944
rect 14182 38876 14188 38888
rect 9364 38848 9409 38876
rect 12728 38848 13584 38876
rect 14143 38848 14188 38876
rect 9364 38836 9370 38848
rect 14182 38836 14188 38848
rect 14240 38836 14246 38888
rect 14366 38876 14372 38888
rect 14327 38848 14372 38876
rect 14366 38836 14372 38848
rect 14424 38836 14430 38888
rect 14826 38876 14832 38888
rect 14787 38848 14832 38876
rect 14826 38836 14832 38848
rect 14884 38836 14890 38888
rect 15102 38836 15108 38888
rect 15160 38876 15166 38888
rect 15580 38876 15608 38916
rect 16669 38913 16681 38916
rect 16715 38913 16727 38947
rect 16853 38947 16911 38953
rect 16853 38942 16865 38947
rect 16669 38907 16727 38913
rect 16776 38914 16865 38942
rect 15160 38848 15608 38876
rect 15160 38836 15166 38848
rect 15746 38836 15752 38888
rect 15804 38876 15810 38888
rect 16482 38876 16488 38888
rect 15804 38848 16488 38876
rect 15804 38836 15810 38848
rect 16482 38836 16488 38848
rect 16540 38836 16546 38888
rect 4212 38780 5488 38808
rect 4212 38768 4218 38780
rect 8294 38768 8300 38820
rect 8352 38808 8358 38820
rect 16776 38808 16804 38914
rect 16853 38913 16865 38914
rect 16899 38913 16911 38947
rect 16853 38907 16911 38913
rect 17126 38904 17132 38956
rect 17184 38904 17190 38956
rect 16942 38836 16948 38888
rect 17000 38876 17006 38888
rect 17236 38876 17264 38984
rect 18046 38972 18052 38984
rect 18104 38972 18110 39024
rect 18616 39012 18644 39052
rect 18782 39040 18788 39092
rect 18840 39080 18846 39092
rect 20990 39080 20996 39092
rect 18840 39052 20996 39080
rect 18840 39040 18846 39052
rect 20990 39040 20996 39052
rect 21048 39040 21054 39092
rect 22094 39040 22100 39092
rect 22152 39080 22158 39092
rect 26786 39080 26792 39092
rect 22152 39052 26792 39080
rect 22152 39040 22158 39052
rect 26786 39040 26792 39052
rect 26844 39040 26850 39092
rect 30374 39080 30380 39092
rect 27080 39052 29592 39080
rect 30335 39052 30380 39080
rect 27080 39021 27108 39052
rect 24673 39015 24731 39021
rect 24673 39012 24685 39015
rect 18616 38984 24685 39012
rect 24673 38981 24685 38984
rect 24719 38981 24731 39015
rect 24673 38975 24731 38981
rect 27065 39015 27123 39021
rect 27065 38981 27077 39015
rect 27111 38981 27123 39015
rect 27246 39012 27252 39024
rect 27207 38984 27252 39012
rect 27065 38975 27123 38981
rect 27246 38972 27252 38984
rect 27304 38972 27310 39024
rect 27890 39012 27896 39024
rect 27851 38984 27896 39012
rect 27890 38972 27896 38984
rect 27948 38972 27954 39024
rect 29564 39012 29592 39052
rect 30374 39040 30380 39052
rect 30432 39040 30438 39092
rect 29822 39012 29828 39024
rect 29564 38984 29828 39012
rect 29822 38972 29828 38984
rect 29880 39012 29886 39024
rect 30929 39015 30987 39021
rect 30929 39012 30941 39015
rect 29880 38984 30941 39012
rect 29880 38972 29886 38984
rect 30929 38981 30941 38984
rect 30975 38981 30987 39015
rect 32490 39012 32496 39024
rect 32451 38984 32496 39012
rect 30929 38975 30987 38981
rect 32490 38972 32496 38984
rect 32548 38972 32554 39024
rect 18874 38904 18880 38956
rect 18932 38944 18938 38956
rect 20145 38947 20203 38953
rect 20145 38944 20157 38947
rect 18932 38916 20157 38944
rect 18932 38904 18938 38916
rect 20145 38913 20157 38916
rect 20191 38913 20203 38947
rect 22186 38944 22192 38956
rect 20145 38907 20203 38913
rect 20916 38916 22094 38944
rect 22147 38916 22192 38944
rect 17000 38848 17264 38876
rect 17497 38879 17555 38885
rect 17000 38836 17006 38848
rect 17497 38845 17509 38879
rect 17543 38845 17555 38879
rect 17497 38839 17555 38845
rect 17681 38879 17739 38885
rect 17681 38845 17693 38879
rect 17727 38860 17739 38879
rect 18230 38876 18236 38888
rect 17727 38845 17816 38860
rect 18191 38848 18236 38876
rect 17681 38839 17816 38845
rect 8352 38780 16804 38808
rect 8352 38768 8358 38780
rect 17218 38768 17224 38820
rect 17276 38808 17282 38820
rect 17512 38808 17540 38839
rect 17696 38832 17816 38839
rect 18230 38836 18236 38848
rect 18288 38836 18294 38888
rect 18322 38836 18328 38888
rect 18380 38876 18386 38888
rect 19702 38876 19708 38888
rect 18380 38848 19708 38876
rect 18380 38836 18386 38848
rect 19702 38836 19708 38848
rect 19760 38836 19766 38888
rect 19886 38876 19892 38888
rect 19847 38848 19892 38876
rect 19886 38836 19892 38848
rect 19944 38836 19950 38888
rect 17276 38780 17540 38808
rect 17788 38808 17816 38832
rect 19334 38808 19340 38820
rect 17788 38780 19340 38808
rect 17276 38768 17282 38780
rect 19334 38768 19340 38780
rect 19392 38768 19398 38820
rect 6454 38700 6460 38752
rect 6512 38740 6518 38752
rect 6733 38743 6791 38749
rect 6733 38740 6745 38743
rect 6512 38712 6745 38740
rect 6512 38700 6518 38712
rect 6733 38709 6745 38712
rect 6779 38709 6791 38743
rect 6733 38703 6791 38709
rect 7377 38743 7435 38749
rect 7377 38709 7389 38743
rect 7423 38740 7435 38743
rect 9122 38740 9128 38752
rect 7423 38712 9128 38740
rect 7423 38709 7435 38712
rect 7377 38703 7435 38709
rect 9122 38700 9128 38712
rect 9180 38700 9186 38752
rect 9214 38700 9220 38752
rect 9272 38740 9278 38752
rect 13722 38740 13728 38752
rect 9272 38712 13728 38740
rect 9272 38700 9278 38712
rect 13722 38700 13728 38712
rect 13780 38700 13786 38752
rect 13814 38700 13820 38752
rect 13872 38740 13878 38752
rect 17037 38743 17095 38749
rect 17037 38740 17049 38743
rect 13872 38712 17049 38740
rect 13872 38700 13878 38712
rect 17037 38709 17049 38712
rect 17083 38709 17095 38743
rect 17037 38703 17095 38709
rect 17310 38700 17316 38752
rect 17368 38740 17374 38752
rect 20916 38740 20944 38916
rect 22066 38876 22094 38916
rect 22186 38904 22192 38916
rect 22244 38904 22250 38956
rect 24486 38944 24492 38956
rect 24447 38916 24492 38944
rect 24486 38904 24492 38916
rect 24544 38904 24550 38956
rect 30193 38947 30251 38953
rect 30193 38913 30205 38947
rect 30239 38913 30251 38947
rect 30193 38907 30251 38913
rect 22373 38879 22431 38885
rect 22066 38848 22324 38876
rect 20990 38768 20996 38820
rect 21048 38808 21054 38820
rect 22094 38808 22100 38820
rect 21048 38780 22100 38808
rect 21048 38768 21054 38780
rect 22094 38768 22100 38780
rect 22152 38768 22158 38820
rect 22296 38808 22324 38848
rect 22373 38845 22385 38879
rect 22419 38876 22431 38879
rect 22462 38876 22468 38888
rect 22419 38848 22468 38876
rect 22419 38845 22431 38848
rect 22373 38839 22431 38845
rect 22462 38836 22468 38848
rect 22520 38836 22526 38888
rect 22554 38836 22560 38888
rect 22612 38876 22618 38888
rect 22649 38879 22707 38885
rect 22649 38876 22661 38879
rect 22612 38848 22661 38876
rect 22612 38836 22618 38848
rect 22649 38845 22661 38848
rect 22695 38845 22707 38879
rect 25130 38876 25136 38888
rect 25091 38848 25136 38876
rect 22649 38839 22707 38845
rect 25130 38836 25136 38848
rect 25188 38836 25194 38888
rect 27706 38876 27712 38888
rect 27667 38848 27712 38876
rect 27706 38836 27712 38848
rect 27764 38836 27770 38888
rect 28350 38876 28356 38888
rect 28311 38848 28356 38876
rect 28350 38836 28356 38848
rect 28408 38836 28414 38888
rect 28442 38836 28448 38888
rect 28500 38876 28506 38888
rect 30009 38879 30067 38885
rect 30009 38876 30021 38879
rect 28500 38848 30021 38876
rect 28500 38836 28506 38848
rect 30009 38845 30021 38848
rect 30055 38845 30067 38879
rect 30009 38839 30067 38845
rect 22296 38780 27476 38808
rect 17368 38712 20944 38740
rect 17368 38700 17374 38712
rect 21082 38700 21088 38752
rect 21140 38740 21146 38752
rect 21269 38743 21327 38749
rect 21269 38740 21281 38743
rect 21140 38712 21281 38740
rect 21140 38700 21146 38712
rect 21269 38709 21281 38712
rect 21315 38709 21327 38743
rect 21269 38703 21327 38709
rect 21910 38700 21916 38752
rect 21968 38740 21974 38752
rect 22554 38740 22560 38752
rect 21968 38712 22560 38740
rect 21968 38700 21974 38712
rect 22554 38700 22560 38712
rect 22612 38740 22618 38752
rect 23750 38740 23756 38752
rect 22612 38712 23756 38740
rect 22612 38700 22618 38712
rect 23750 38700 23756 38712
rect 23808 38700 23814 38752
rect 27448 38740 27476 38780
rect 27522 38768 27528 38820
rect 27580 38808 27586 38820
rect 30208 38808 30236 38907
rect 31938 38904 31944 38956
rect 31996 38944 32002 38956
rect 32309 38947 32367 38953
rect 32309 38944 32321 38947
rect 31996 38916 32321 38944
rect 31996 38904 32002 38916
rect 32309 38913 32321 38916
rect 32355 38913 32367 38947
rect 32309 38907 32367 38913
rect 33502 38876 33508 38888
rect 33463 38848 33508 38876
rect 33502 38836 33508 38848
rect 33560 38836 33566 38888
rect 27580 38780 30236 38808
rect 31113 38811 31171 38817
rect 27580 38768 27586 38780
rect 31113 38777 31125 38811
rect 31159 38808 31171 38811
rect 31478 38808 31484 38820
rect 31159 38780 31484 38808
rect 31159 38777 31171 38780
rect 31113 38771 31171 38777
rect 31478 38768 31484 38780
rect 31536 38768 31542 38820
rect 30650 38740 30656 38752
rect 27448 38712 30656 38740
rect 30650 38700 30656 38712
rect 30708 38700 30714 38752
rect 1104 38650 34868 38672
rect 1104 38598 6582 38650
rect 6634 38598 6646 38650
rect 6698 38598 6710 38650
rect 6762 38598 6774 38650
rect 6826 38598 6838 38650
rect 6890 38598 17846 38650
rect 17898 38598 17910 38650
rect 17962 38598 17974 38650
rect 18026 38598 18038 38650
rect 18090 38598 18102 38650
rect 18154 38598 29110 38650
rect 29162 38598 29174 38650
rect 29226 38598 29238 38650
rect 29290 38598 29302 38650
rect 29354 38598 29366 38650
rect 29418 38598 34868 38650
rect 1104 38576 34868 38598
rect 11609 38539 11667 38545
rect 11609 38505 11621 38539
rect 11655 38536 11667 38539
rect 14182 38536 14188 38548
rect 11655 38508 14188 38536
rect 11655 38505 11667 38508
rect 11609 38499 11667 38505
rect 14182 38496 14188 38508
rect 14240 38496 14246 38548
rect 14366 38496 14372 38548
rect 14424 38536 14430 38548
rect 14461 38539 14519 38545
rect 14461 38536 14473 38539
rect 14424 38508 14473 38536
rect 14424 38496 14430 38508
rect 14461 38505 14473 38508
rect 14507 38505 14519 38539
rect 14461 38499 14519 38505
rect 14642 38496 14648 38548
rect 14700 38536 14706 38548
rect 18141 38539 18199 38545
rect 18141 38536 18153 38539
rect 14700 38508 18153 38536
rect 14700 38496 14706 38508
rect 18141 38505 18153 38508
rect 18187 38505 18199 38539
rect 18141 38499 18199 38505
rect 18414 38496 18420 38548
rect 18472 38536 18478 38548
rect 18782 38536 18788 38548
rect 18472 38508 18788 38536
rect 18472 38496 18478 38508
rect 18782 38496 18788 38508
rect 18840 38496 18846 38548
rect 19334 38536 19340 38548
rect 19295 38508 19340 38536
rect 19334 38496 19340 38508
rect 19392 38496 19398 38548
rect 19430 38508 25360 38536
rect 1854 38428 1860 38480
rect 1912 38468 1918 38480
rect 1912 38440 8064 38468
rect 1912 38428 1918 38440
rect 1302 38360 1308 38412
rect 1360 38400 1366 38412
rect 1949 38403 2007 38409
rect 1949 38400 1961 38403
rect 1360 38372 1961 38400
rect 1360 38360 1366 38372
rect 1949 38369 1961 38372
rect 1995 38369 2007 38403
rect 1949 38363 2007 38369
rect 4249 38403 4307 38409
rect 4249 38369 4261 38403
rect 4295 38400 4307 38403
rect 5626 38400 5632 38412
rect 4295 38372 5632 38400
rect 4295 38369 4307 38372
rect 4249 38363 4307 38369
rect 5626 38360 5632 38372
rect 5684 38360 5690 38412
rect 5810 38400 5816 38412
rect 5771 38372 5816 38400
rect 5810 38360 5816 38372
rect 5868 38360 5874 38412
rect 6454 38360 6460 38412
rect 6512 38400 6518 38412
rect 6549 38403 6607 38409
rect 6549 38400 6561 38403
rect 6512 38372 6561 38400
rect 6512 38360 6518 38372
rect 6549 38369 6561 38372
rect 6595 38369 6607 38403
rect 7098 38400 7104 38412
rect 7059 38372 7104 38400
rect 6549 38363 6607 38369
rect 7098 38360 7104 38372
rect 7156 38360 7162 38412
rect 1397 38335 1455 38341
rect 1397 38301 1409 38335
rect 1443 38301 1455 38335
rect 1397 38295 1455 38301
rect 1412 38196 1440 38295
rect 1578 38264 1584 38276
rect 1539 38236 1584 38264
rect 1578 38224 1584 38236
rect 1636 38224 1642 38276
rect 4433 38267 4491 38273
rect 4433 38233 4445 38267
rect 4479 38264 4491 38267
rect 5350 38264 5356 38276
rect 4479 38236 5356 38264
rect 4479 38233 4491 38236
rect 4433 38227 4491 38233
rect 5350 38224 5356 38236
rect 5408 38224 5414 38276
rect 6730 38264 6736 38276
rect 6691 38236 6736 38264
rect 6730 38224 6736 38236
rect 6788 38224 6794 38276
rect 8036 38264 8064 38440
rect 8386 38428 8392 38480
rect 8444 38468 8450 38480
rect 12250 38468 12256 38480
rect 8444 38440 9444 38468
rect 12211 38440 12256 38468
rect 8444 38428 8450 38440
rect 9122 38400 9128 38412
rect 9083 38372 9128 38400
rect 9122 38360 9128 38372
rect 9180 38360 9186 38412
rect 9416 38409 9444 38440
rect 12250 38428 12256 38440
rect 12308 38428 12314 38480
rect 13446 38428 13452 38480
rect 13504 38468 13510 38480
rect 17678 38468 17684 38480
rect 13504 38440 17684 38468
rect 13504 38428 13510 38440
rect 17678 38428 17684 38440
rect 17736 38428 17742 38480
rect 19430 38468 19458 38508
rect 17880 38440 19458 38468
rect 9401 38403 9459 38409
rect 9401 38369 9413 38403
rect 9447 38369 9459 38403
rect 9401 38363 9459 38369
rect 11330 38360 11336 38412
rect 11388 38400 11394 38412
rect 13078 38400 13084 38412
rect 11388 38372 13084 38400
rect 11388 38360 11394 38372
rect 13078 38360 13084 38372
rect 13136 38360 13142 38412
rect 14642 38400 14648 38412
rect 13556 38372 14648 38400
rect 8110 38292 8116 38344
rect 8168 38332 8174 38344
rect 8941 38335 8999 38341
rect 8941 38332 8953 38335
rect 8168 38304 8953 38332
rect 8168 38292 8174 38304
rect 8941 38301 8953 38304
rect 8987 38301 8999 38335
rect 12894 38332 12900 38344
rect 12855 38304 12900 38332
rect 8941 38295 8999 38301
rect 12894 38292 12900 38304
rect 12952 38292 12958 38344
rect 13556 38341 13584 38372
rect 14642 38360 14648 38372
rect 14700 38360 14706 38412
rect 15654 38400 15660 38412
rect 15615 38372 15660 38400
rect 15654 38360 15660 38372
rect 15712 38360 15718 38412
rect 16110 38400 16116 38412
rect 16168 38409 16174 38412
rect 16075 38372 16116 38400
rect 16110 38360 16116 38372
rect 16168 38363 16175 38409
rect 16168 38360 16174 38363
rect 17402 38360 17408 38412
rect 17460 38400 17466 38412
rect 17880 38400 17908 38440
rect 19702 38428 19708 38480
rect 19760 38468 19766 38480
rect 21910 38468 21916 38480
rect 19760 38440 21916 38468
rect 19760 38428 19766 38440
rect 21910 38428 21916 38440
rect 21968 38428 21974 38480
rect 23750 38468 23756 38480
rect 23711 38440 23756 38468
rect 23750 38428 23756 38440
rect 23808 38468 23814 38480
rect 24026 38468 24032 38480
rect 23808 38440 24032 38468
rect 23808 38428 23814 38440
rect 24026 38428 24032 38440
rect 24084 38428 24090 38480
rect 17460 38372 17908 38400
rect 17460 38360 17466 38372
rect 18138 38360 18144 38412
rect 18196 38400 18202 38412
rect 19978 38400 19984 38412
rect 18196 38372 19984 38400
rect 18196 38360 18202 38372
rect 19978 38360 19984 38372
rect 20036 38360 20042 38412
rect 20254 38360 20260 38412
rect 20312 38400 20318 38412
rect 20312 38372 20357 38400
rect 20312 38360 20318 38372
rect 20622 38360 20628 38412
rect 20680 38400 20686 38412
rect 20717 38403 20775 38409
rect 20717 38400 20729 38403
rect 20680 38372 20729 38400
rect 20680 38360 20686 38372
rect 20717 38369 20729 38372
rect 20763 38369 20775 38403
rect 20717 38363 20775 38369
rect 21726 38360 21732 38412
rect 21784 38400 21790 38412
rect 22278 38400 22284 38412
rect 21784 38372 22284 38400
rect 21784 38360 21790 38372
rect 22278 38360 22284 38372
rect 22336 38360 22342 38412
rect 25332 38409 25360 38508
rect 25317 38403 25375 38409
rect 25317 38369 25329 38403
rect 25363 38369 25375 38403
rect 25774 38400 25780 38412
rect 25735 38372 25780 38400
rect 25317 38363 25375 38369
rect 25774 38360 25780 38372
rect 25832 38360 25838 38412
rect 28626 38400 28632 38412
rect 28587 38372 28632 38400
rect 28626 38360 28632 38372
rect 28684 38360 28690 38412
rect 28994 38360 29000 38412
rect 29052 38400 29058 38412
rect 30009 38403 30067 38409
rect 30009 38400 30021 38403
rect 29052 38372 30021 38400
rect 29052 38360 29058 38372
rect 30009 38369 30021 38372
rect 30055 38369 30067 38403
rect 30009 38363 30067 38369
rect 31846 38360 31852 38412
rect 31904 38400 31910 38412
rect 32309 38403 32367 38409
rect 32309 38400 32321 38403
rect 31904 38372 32321 38400
rect 31904 38360 31910 38372
rect 32309 38369 32321 38372
rect 32355 38369 32367 38403
rect 34146 38400 34152 38412
rect 34107 38372 34152 38400
rect 32309 38363 32367 38369
rect 34146 38360 34152 38372
rect 34204 38360 34210 38412
rect 13541 38335 13599 38341
rect 13541 38301 13553 38335
rect 13587 38301 13599 38335
rect 14366 38332 14372 38344
rect 14327 38304 14372 38332
rect 13541 38295 13599 38301
rect 14366 38292 14372 38304
rect 14424 38292 14430 38344
rect 14458 38292 14464 38344
rect 14516 38332 14522 38344
rect 15473 38335 15531 38341
rect 15473 38332 15485 38335
rect 14516 38304 15485 38332
rect 14516 38292 14522 38304
rect 15473 38301 15485 38304
rect 15519 38301 15531 38335
rect 15473 38295 15531 38301
rect 16850 38292 16856 38344
rect 16908 38332 16914 38344
rect 16908 38304 17080 38332
rect 16908 38292 16914 38304
rect 13262 38264 13268 38276
rect 8036 38236 13268 38264
rect 13262 38224 13268 38236
rect 13320 38224 13326 38276
rect 16942 38264 16948 38276
rect 13372 38236 16948 38264
rect 5258 38196 5264 38208
rect 1412 38168 5264 38196
rect 5258 38156 5264 38168
rect 5316 38156 5322 38208
rect 11606 38156 11612 38208
rect 11664 38196 11670 38208
rect 12618 38196 12624 38208
rect 11664 38168 12624 38196
rect 11664 38156 11670 38168
rect 12618 38156 12624 38168
rect 12676 38156 12682 38208
rect 12713 38199 12771 38205
rect 12713 38165 12725 38199
rect 12759 38196 12771 38199
rect 13078 38196 13084 38208
rect 12759 38168 13084 38196
rect 12759 38165 12771 38168
rect 12713 38159 12771 38165
rect 13078 38156 13084 38168
rect 13136 38156 13142 38208
rect 13372 38205 13400 38236
rect 16942 38224 16948 38236
rect 17000 38224 17006 38276
rect 17052 38264 17080 38304
rect 17126 38292 17132 38344
rect 17184 38332 17190 38344
rect 17773 38335 17831 38341
rect 17773 38332 17785 38335
rect 17184 38304 17785 38332
rect 17184 38292 17190 38304
rect 17773 38301 17785 38304
rect 17819 38301 17831 38335
rect 17773 38295 17831 38301
rect 17862 38292 17868 38344
rect 17920 38332 17926 38344
rect 17957 38335 18015 38341
rect 17957 38332 17969 38335
rect 17920 38304 17969 38332
rect 17920 38292 17926 38304
rect 17957 38301 17969 38304
rect 18003 38301 18015 38335
rect 19058 38332 19064 38344
rect 17957 38295 18015 38301
rect 18708 38304 19064 38332
rect 18708 38264 18736 38304
rect 19058 38292 19064 38304
rect 19116 38292 19122 38344
rect 19150 38292 19156 38344
rect 19208 38332 19214 38344
rect 19245 38335 19303 38341
rect 19245 38332 19257 38335
rect 19208 38304 19257 38332
rect 19208 38292 19214 38304
rect 19245 38301 19257 38304
rect 19291 38301 19303 38335
rect 19245 38295 19303 38301
rect 19334 38292 19340 38344
rect 19392 38332 19398 38344
rect 20073 38335 20131 38341
rect 20073 38332 20085 38335
rect 19392 38304 20085 38332
rect 19392 38292 19398 38304
rect 20073 38301 20085 38304
rect 20119 38301 20131 38335
rect 22370 38332 22376 38344
rect 22331 38304 22376 38332
rect 20073 38295 20131 38301
rect 22370 38292 22376 38304
rect 22428 38292 22434 38344
rect 24489 38335 24547 38341
rect 24489 38332 24501 38335
rect 22480 38304 24501 38332
rect 22480 38264 22508 38304
rect 24489 38301 24501 38304
rect 24535 38301 24547 38335
rect 25130 38332 25136 38344
rect 25091 38304 25136 38332
rect 24489 38295 24547 38301
rect 25130 38292 25136 38304
rect 25188 38292 25194 38344
rect 26510 38292 26516 38344
rect 26568 38332 26574 38344
rect 27433 38335 27491 38341
rect 27433 38332 27445 38335
rect 26568 38304 27445 38332
rect 26568 38292 26574 38304
rect 27433 38301 27445 38304
rect 27479 38301 27491 38335
rect 27433 38295 27491 38301
rect 27522 38292 27528 38344
rect 27580 38332 27586 38344
rect 27617 38335 27675 38341
rect 27617 38332 27629 38335
rect 27580 38304 27629 38332
rect 27580 38292 27586 38304
rect 27617 38301 27629 38304
rect 27663 38301 27675 38335
rect 27617 38295 27675 38301
rect 28353 38335 28411 38341
rect 28353 38301 28365 38335
rect 28399 38332 28411 38335
rect 28810 38332 28816 38344
rect 28399 38304 28816 38332
rect 28399 38301 28411 38304
rect 28353 38295 28411 38301
rect 28810 38292 28816 38304
rect 28868 38292 28874 38344
rect 29546 38332 29552 38344
rect 29507 38304 29552 38332
rect 29546 38292 29552 38304
rect 29604 38292 29610 38344
rect 17052 38236 18736 38264
rect 22066 38236 22508 38264
rect 22629 38267 22687 38273
rect 13357 38199 13415 38205
rect 13357 38165 13369 38199
rect 13403 38165 13415 38199
rect 13357 38159 13415 38165
rect 13722 38156 13728 38208
rect 13780 38196 13786 38208
rect 15010 38196 15016 38208
rect 13780 38168 15016 38196
rect 13780 38156 13786 38168
rect 15010 38156 15016 38168
rect 15068 38156 15074 38208
rect 15102 38156 15108 38208
rect 15160 38196 15166 38208
rect 22066 38196 22094 38236
rect 22629 38233 22641 38267
rect 22675 38233 22687 38267
rect 22629 38227 22687 38233
rect 15160 38168 22094 38196
rect 15160 38156 15166 38168
rect 22186 38156 22192 38208
rect 22244 38196 22250 38208
rect 22633 38196 22661 38227
rect 22738 38224 22744 38276
rect 22796 38264 22802 38276
rect 24762 38264 24768 38276
rect 22796 38236 24768 38264
rect 22796 38224 22802 38236
rect 24762 38224 24768 38236
rect 24820 38224 24826 38276
rect 25038 38224 25044 38276
rect 25096 38264 25102 38276
rect 29733 38267 29791 38273
rect 29733 38264 29745 38267
rect 25096 38236 29745 38264
rect 25096 38224 25102 38236
rect 29733 38233 29745 38236
rect 29779 38233 29791 38267
rect 32490 38264 32496 38276
rect 32451 38236 32496 38264
rect 29733 38227 29791 38233
rect 32490 38224 32496 38236
rect 32548 38224 32554 38276
rect 22244 38168 22661 38196
rect 24581 38199 24639 38205
rect 22244 38156 22250 38168
rect 24581 38165 24593 38199
rect 24627 38196 24639 38199
rect 24670 38196 24676 38208
rect 24627 38168 24676 38196
rect 24627 38165 24639 38168
rect 24581 38159 24639 38165
rect 24670 38156 24676 38168
rect 24728 38156 24734 38208
rect 27798 38196 27804 38208
rect 27759 38168 27804 38196
rect 27798 38156 27804 38168
rect 27856 38156 27862 38208
rect 1104 38106 34868 38128
rect 1104 38054 12214 38106
rect 12266 38054 12278 38106
rect 12330 38054 12342 38106
rect 12394 38054 12406 38106
rect 12458 38054 12470 38106
rect 12522 38054 23478 38106
rect 23530 38054 23542 38106
rect 23594 38054 23606 38106
rect 23658 38054 23670 38106
rect 23722 38054 23734 38106
rect 23786 38054 34868 38106
rect 1104 38032 34868 38054
rect 1670 37952 1676 38004
rect 1728 37992 1734 38004
rect 1949 37995 2007 38001
rect 1949 37992 1961 37995
rect 1728 37964 1961 37992
rect 1728 37952 1734 37964
rect 1949 37961 1961 37964
rect 1995 37961 2007 37995
rect 5350 37992 5356 38004
rect 5311 37964 5356 37992
rect 1949 37955 2007 37961
rect 5350 37952 5356 37964
rect 5408 37952 5414 38004
rect 6641 37995 6699 38001
rect 6641 37961 6653 37995
rect 6687 37992 6699 37995
rect 6730 37992 6736 38004
rect 6687 37964 6736 37992
rect 6687 37961 6699 37964
rect 6641 37955 6699 37961
rect 6730 37952 6736 37964
rect 6788 37952 6794 38004
rect 11606 37992 11612 38004
rect 11567 37964 11612 37992
rect 11606 37952 11612 37964
rect 11664 37952 11670 38004
rect 12253 37995 12311 38001
rect 12253 37961 12265 37995
rect 12299 37992 12311 37995
rect 12710 37992 12716 38004
rect 12299 37964 12716 37992
rect 12299 37961 12311 37964
rect 12253 37955 12311 37961
rect 12710 37952 12716 37964
rect 12768 37952 12774 38004
rect 12897 37995 12955 38001
rect 12897 37961 12909 37995
rect 12943 37992 12955 37995
rect 13906 37992 13912 38004
rect 12943 37964 13912 37992
rect 12943 37961 12955 37964
rect 12897 37955 12955 37961
rect 13906 37952 13912 37964
rect 13964 37952 13970 38004
rect 14182 37952 14188 38004
rect 14240 37992 14246 38004
rect 14240 37964 14688 37992
rect 14240 37952 14246 37964
rect 2777 37927 2835 37933
rect 2777 37893 2789 37927
rect 2823 37924 2835 37927
rect 3234 37924 3240 37936
rect 2823 37896 3240 37924
rect 2823 37893 2835 37896
rect 2777 37887 2835 37893
rect 3234 37884 3240 37896
rect 3292 37884 3298 37936
rect 10410 37884 10416 37936
rect 10468 37924 10474 37936
rect 14458 37924 14464 37936
rect 10468 37896 14464 37924
rect 10468 37884 10474 37896
rect 14458 37884 14464 37896
rect 14516 37884 14522 37936
rect 14660 37933 14688 37964
rect 14936 37964 20944 37992
rect 14645 37927 14703 37933
rect 14645 37893 14657 37927
rect 14691 37893 14703 37927
rect 14645 37887 14703 37893
rect 1854 37856 1860 37868
rect 1815 37828 1860 37856
rect 1854 37816 1860 37828
rect 1912 37816 1918 37868
rect 4798 37816 4804 37868
rect 4856 37856 4862 37868
rect 5261 37859 5319 37865
rect 5261 37856 5273 37859
rect 4856 37828 5273 37856
rect 4856 37816 4862 37828
rect 5261 37825 5273 37828
rect 5307 37825 5319 37859
rect 5261 37819 5319 37825
rect 5534 37816 5540 37868
rect 5592 37856 5598 37868
rect 6549 37859 6607 37865
rect 6549 37856 6561 37859
rect 5592 37828 6561 37856
rect 5592 37816 5598 37828
rect 6549 37825 6561 37828
rect 6595 37825 6607 37859
rect 7190 37856 7196 37868
rect 7151 37828 7196 37856
rect 6549 37819 6607 37825
rect 7190 37816 7196 37828
rect 7248 37816 7254 37868
rect 10318 37856 10324 37868
rect 10279 37828 10324 37856
rect 10318 37816 10324 37828
rect 10376 37816 10382 37868
rect 10962 37856 10968 37868
rect 10923 37828 10968 37856
rect 10962 37816 10968 37828
rect 11020 37816 11026 37868
rect 11793 37859 11851 37865
rect 11793 37825 11805 37859
rect 11839 37856 11851 37859
rect 12066 37856 12072 37868
rect 11839 37828 12072 37856
rect 11839 37825 11851 37828
rect 11793 37819 11851 37825
rect 12066 37816 12072 37828
rect 12124 37816 12130 37868
rect 12434 37816 12440 37868
rect 12492 37856 12498 37868
rect 13081 37859 13139 37865
rect 12492 37828 12537 37856
rect 12492 37816 12498 37828
rect 13081 37825 13093 37859
rect 13127 37825 13139 37859
rect 13081 37819 13139 37825
rect 13725 37859 13783 37865
rect 13725 37825 13737 37859
rect 13771 37856 13783 37859
rect 13814 37856 13820 37868
rect 13771 37828 13820 37856
rect 13771 37825 13783 37828
rect 13725 37819 13783 37825
rect 2593 37791 2651 37797
rect 2593 37757 2605 37791
rect 2639 37757 2651 37791
rect 2593 37751 2651 37757
rect 2608 37720 2636 37751
rect 2958 37748 2964 37800
rect 3016 37788 3022 37800
rect 3053 37791 3111 37797
rect 3053 37788 3065 37791
rect 3016 37760 3065 37788
rect 3016 37748 3022 37760
rect 3053 37757 3065 37760
rect 3099 37757 3111 37791
rect 7374 37788 7380 37800
rect 7335 37760 7380 37788
rect 3053 37751 3111 37757
rect 7374 37748 7380 37760
rect 7432 37748 7438 37800
rect 7742 37788 7748 37800
rect 7703 37760 7748 37788
rect 7742 37748 7748 37760
rect 7800 37748 7806 37800
rect 13096 37788 13124 37819
rect 13814 37816 13820 37828
rect 13872 37816 13878 37868
rect 14277 37859 14335 37865
rect 14277 37825 14289 37859
rect 14323 37856 14335 37859
rect 14366 37856 14372 37868
rect 14323 37828 14372 37856
rect 14323 37825 14335 37828
rect 14277 37819 14335 37825
rect 14366 37816 14372 37828
rect 14424 37816 14430 37868
rect 14936 37856 14964 37964
rect 15010 37884 15016 37936
rect 15068 37924 15074 37936
rect 18138 37924 18144 37936
rect 15068 37896 18144 37924
rect 15068 37884 15074 37896
rect 18138 37884 18144 37896
rect 18196 37884 18202 37936
rect 18230 37884 18236 37936
rect 18288 37924 18294 37936
rect 18288 37896 19012 37924
rect 18288 37884 18294 37896
rect 15930 37856 15936 37868
rect 14844 37828 14964 37856
rect 15891 37828 15936 37856
rect 13096 37760 13860 37788
rect 4614 37720 4620 37732
rect 2608 37692 4620 37720
rect 4614 37680 4620 37692
rect 4672 37680 4678 37732
rect 9674 37720 9680 37732
rect 9635 37692 9680 37720
rect 9674 37680 9680 37692
rect 9732 37680 9738 37732
rect 12710 37680 12716 37732
rect 12768 37720 12774 37732
rect 13722 37720 13728 37732
rect 12768 37692 13728 37720
rect 12768 37680 12774 37692
rect 13722 37680 13728 37692
rect 13780 37680 13786 37732
rect 13832 37720 13860 37760
rect 13906 37748 13912 37800
rect 13964 37788 13970 37800
rect 14844 37788 14872 37828
rect 15930 37816 15936 37828
rect 15988 37816 15994 37868
rect 16022 37816 16028 37868
rect 16080 37856 16086 37868
rect 16758 37856 16764 37868
rect 16080 37828 16125 37856
rect 16224 37828 16764 37856
rect 16080 37816 16086 37828
rect 13964 37760 14872 37788
rect 13964 37748 13970 37760
rect 14918 37748 14924 37800
rect 14976 37788 14982 37800
rect 16224 37788 16252 37828
rect 16758 37816 16764 37828
rect 16816 37816 16822 37868
rect 16942 37865 16948 37868
rect 16936 37856 16948 37865
rect 16903 37828 16948 37856
rect 16936 37819 16948 37828
rect 16942 37816 16948 37819
rect 17000 37816 17006 37868
rect 17218 37816 17224 37868
rect 17276 37856 17282 37868
rect 18322 37856 18328 37868
rect 17276 37828 18328 37856
rect 17276 37816 17282 37828
rect 18322 37816 18328 37828
rect 18380 37816 18386 37868
rect 18782 37865 18788 37868
rect 18776 37819 18788 37865
rect 18840 37856 18846 37868
rect 18984 37856 19012 37896
rect 19886 37884 19892 37936
rect 19944 37924 19950 37936
rect 20916 37924 20944 37964
rect 20990 37952 20996 38004
rect 21048 37992 21054 38004
rect 23014 37992 23020 38004
rect 21048 37964 23020 37992
rect 21048 37952 21054 37964
rect 23014 37952 23020 37964
rect 23072 37952 23078 38004
rect 23201 37995 23259 38001
rect 23201 37961 23213 37995
rect 23247 37992 23259 37995
rect 23382 37992 23388 38004
rect 23247 37964 23388 37992
rect 23247 37961 23259 37964
rect 23201 37955 23259 37961
rect 23382 37952 23388 37964
rect 23440 37992 23446 38004
rect 23937 37995 23995 38001
rect 23937 37992 23949 37995
rect 23440 37964 23949 37992
rect 23440 37952 23446 37964
rect 23937 37961 23949 37964
rect 23983 37961 23995 37995
rect 23937 37955 23995 37961
rect 24026 37952 24032 38004
rect 24084 37992 24090 38004
rect 24084 37964 24129 37992
rect 24084 37952 24090 37964
rect 22066 37927 22124 37933
rect 22066 37924 22078 37927
rect 19944 37896 20852 37924
rect 20916 37896 22078 37924
rect 19944 37884 19950 37896
rect 20254 37856 20260 37868
rect 18840 37828 18876 37856
rect 18984 37828 20260 37856
rect 18782 37816 18788 37819
rect 18840 37816 18846 37828
rect 20254 37816 20260 37828
rect 20312 37816 20318 37868
rect 20530 37856 20536 37868
rect 20491 37828 20536 37856
rect 20530 37816 20536 37828
rect 20588 37816 20594 37868
rect 20824 37856 20852 37896
rect 22066 37893 22078 37896
rect 22112 37893 22124 37927
rect 22066 37887 22124 37893
rect 22186 37884 22192 37936
rect 22244 37924 22250 37936
rect 25041 37927 25099 37933
rect 25041 37924 25053 37927
rect 22244 37896 25053 37924
rect 22244 37884 22250 37896
rect 25041 37893 25053 37896
rect 25087 37893 25099 37927
rect 29914 37924 29920 37936
rect 29875 37896 29920 37924
rect 25041 37887 25099 37893
rect 29914 37884 29920 37896
rect 29972 37884 29978 37936
rect 31573 37927 31631 37933
rect 31573 37893 31585 37927
rect 31619 37924 31631 37927
rect 33042 37924 33048 37936
rect 31619 37896 33048 37924
rect 31619 37893 31631 37896
rect 31573 37887 31631 37893
rect 33042 37884 33048 37896
rect 33100 37884 33106 37936
rect 34054 37884 34060 37936
rect 34112 37924 34118 37936
rect 34149 37927 34207 37933
rect 34149 37924 34161 37927
rect 34112 37896 34161 37924
rect 34112 37884 34118 37896
rect 34149 37893 34161 37896
rect 34195 37893 34207 37927
rect 34149 37887 34207 37893
rect 21821 37859 21879 37865
rect 21821 37856 21833 37859
rect 20824 37828 21833 37856
rect 21821 37825 21833 37828
rect 21867 37856 21879 37859
rect 22370 37856 22376 37868
rect 21867 37828 22376 37856
rect 21867 37825 21879 37828
rect 21821 37819 21879 37825
rect 22370 37816 22376 37828
rect 22428 37816 22434 37868
rect 23014 37816 23020 37868
rect 23072 37856 23078 37868
rect 23845 37859 23903 37865
rect 23845 37856 23857 37859
rect 23072 37828 23857 37856
rect 23072 37816 23078 37828
rect 23845 37825 23857 37828
rect 23891 37825 23903 37859
rect 23845 37819 23903 37825
rect 24394 37816 24400 37868
rect 24452 37856 24458 37868
rect 24857 37859 24915 37865
rect 24857 37856 24869 37859
rect 24452 37828 24869 37856
rect 24452 37816 24458 37828
rect 24857 37825 24869 37828
rect 24903 37825 24915 37859
rect 25682 37856 25688 37868
rect 25643 37828 25688 37856
rect 24857 37819 24915 37825
rect 25682 37816 25688 37828
rect 25740 37856 25746 37868
rect 27157 37859 27215 37865
rect 27157 37856 27169 37859
rect 25740 37828 27169 37856
rect 25740 37816 25746 37828
rect 27157 37825 27169 37828
rect 27203 37856 27215 37859
rect 27522 37856 27528 37868
rect 27203 37828 27528 37856
rect 27203 37825 27215 37828
rect 27157 37819 27215 37825
rect 27522 37816 27528 37828
rect 27580 37816 27586 37868
rect 28445 37859 28503 37865
rect 28445 37825 28457 37859
rect 28491 37856 28503 37859
rect 28902 37856 28908 37868
rect 28491 37828 28908 37856
rect 28491 37825 28503 37828
rect 28445 37819 28503 37825
rect 28902 37816 28908 37828
rect 28960 37816 28966 37868
rect 32030 37816 32036 37868
rect 32088 37856 32094 37868
rect 32309 37859 32367 37865
rect 32309 37856 32321 37859
rect 32088 37828 32321 37856
rect 32088 37816 32094 37828
rect 32309 37825 32321 37828
rect 32355 37825 32367 37859
rect 32309 37819 32367 37825
rect 14976 37760 16252 37788
rect 14976 37748 14982 37760
rect 16574 37748 16580 37800
rect 16632 37788 16638 37800
rect 16669 37791 16727 37797
rect 16669 37788 16681 37791
rect 16632 37760 16681 37788
rect 16632 37748 16638 37760
rect 16669 37757 16681 37760
rect 16715 37757 16727 37791
rect 16669 37751 16727 37757
rect 17678 37748 17684 37800
rect 17736 37788 17742 37800
rect 18230 37788 18236 37800
rect 17736 37760 18236 37788
rect 17736 37748 17742 37760
rect 18230 37748 18236 37760
rect 18288 37748 18294 37800
rect 18506 37788 18512 37800
rect 18467 37760 18512 37788
rect 18506 37748 18512 37760
rect 18564 37748 18570 37800
rect 20349 37791 20407 37797
rect 20349 37788 20361 37791
rect 19904 37760 20361 37788
rect 19904 37729 19932 37760
rect 20349 37757 20361 37760
rect 20395 37788 20407 37791
rect 20990 37788 20996 37800
rect 20395 37760 20996 37788
rect 20395 37757 20407 37760
rect 20349 37751 20407 37757
rect 20990 37748 20996 37760
rect 21048 37748 21054 37800
rect 24673 37791 24731 37797
rect 24673 37757 24685 37791
rect 24719 37788 24731 37791
rect 25406 37788 25412 37800
rect 24719 37760 25412 37788
rect 24719 37757 24731 37760
rect 24673 37751 24731 37757
rect 25406 37748 25412 37760
rect 25464 37748 25470 37800
rect 25501 37791 25559 37797
rect 25501 37757 25513 37791
rect 25547 37788 25559 37791
rect 25866 37788 25872 37800
rect 25547 37760 25872 37788
rect 25547 37757 25559 37760
rect 25501 37751 25559 37757
rect 25866 37748 25872 37760
rect 25924 37748 25930 37800
rect 26602 37748 26608 37800
rect 26660 37788 26666 37800
rect 26973 37791 27031 37797
rect 26973 37788 26985 37791
rect 26660 37760 26985 37788
rect 26660 37748 26666 37760
rect 26973 37757 26985 37760
rect 27019 37757 27031 37791
rect 26973 37751 27031 37757
rect 28534 37748 28540 37800
rect 28592 37788 28598 37800
rect 28629 37791 28687 37797
rect 28629 37788 28641 37791
rect 28592 37760 28641 37788
rect 28592 37748 28598 37760
rect 28629 37757 28641 37760
rect 28675 37757 28687 37791
rect 29730 37788 29736 37800
rect 29691 37760 29736 37788
rect 28629 37751 28687 37757
rect 29730 37748 29736 37760
rect 29788 37748 29794 37800
rect 32493 37791 32551 37797
rect 32493 37757 32505 37791
rect 32539 37757 32551 37791
rect 32493 37751 32551 37757
rect 19889 37723 19947 37729
rect 13832 37692 16574 37720
rect 13541 37655 13599 37661
rect 13541 37621 13553 37655
rect 13587 37652 13599 37655
rect 15562 37652 15568 37664
rect 13587 37624 15568 37652
rect 13587 37621 13599 37624
rect 13541 37615 13599 37621
rect 15562 37612 15568 37624
rect 15620 37612 15626 37664
rect 16546 37652 16574 37692
rect 17696 37692 18184 37720
rect 17696 37652 17724 37692
rect 16546 37624 17724 37652
rect 17770 37612 17776 37664
rect 17828 37652 17834 37664
rect 18049 37655 18107 37661
rect 18049 37652 18061 37655
rect 17828 37624 18061 37652
rect 17828 37612 17834 37624
rect 18049 37621 18061 37624
rect 18095 37621 18107 37655
rect 18156 37652 18184 37692
rect 19889 37689 19901 37723
rect 19935 37689 19947 37723
rect 19889 37683 19947 37689
rect 22830 37680 22836 37732
rect 22888 37720 22894 37732
rect 23661 37723 23719 37729
rect 23661 37720 23673 37723
rect 22888 37692 23673 37720
rect 22888 37680 22894 37692
rect 23661 37689 23673 37692
rect 23707 37689 23719 37723
rect 32508 37720 32536 37751
rect 23661 37683 23719 37689
rect 23748 37692 32536 37720
rect 20717 37655 20775 37661
rect 20717 37652 20729 37655
rect 18156 37624 20729 37652
rect 18049 37615 18107 37621
rect 20717 37621 20729 37624
rect 20763 37621 20775 37655
rect 20717 37615 20775 37621
rect 22002 37612 22008 37664
rect 22060 37652 22066 37664
rect 23748 37652 23776 37692
rect 22060 37624 23776 37652
rect 24213 37655 24271 37661
rect 22060 37612 22066 37624
rect 24213 37621 24225 37655
rect 24259 37652 24271 37655
rect 24578 37652 24584 37664
rect 24259 37624 24584 37652
rect 24259 37621 24271 37624
rect 24213 37615 24271 37621
rect 24578 37612 24584 37624
rect 24636 37612 24642 37664
rect 24762 37612 24768 37664
rect 24820 37652 24826 37664
rect 25869 37655 25927 37661
rect 25869 37652 25881 37655
rect 24820 37624 25881 37652
rect 24820 37612 24826 37624
rect 25869 37621 25881 37624
rect 25915 37621 25927 37655
rect 25869 37615 25927 37621
rect 26234 37612 26240 37664
rect 26292 37652 26298 37664
rect 27341 37655 27399 37661
rect 27341 37652 27353 37655
rect 26292 37624 27353 37652
rect 26292 37612 26298 37624
rect 27341 37621 27353 37624
rect 27387 37621 27399 37655
rect 27341 37615 27399 37621
rect 1104 37562 34868 37584
rect 1104 37510 6582 37562
rect 6634 37510 6646 37562
rect 6698 37510 6710 37562
rect 6762 37510 6774 37562
rect 6826 37510 6838 37562
rect 6890 37510 17846 37562
rect 17898 37510 17910 37562
rect 17962 37510 17974 37562
rect 18026 37510 18038 37562
rect 18090 37510 18102 37562
rect 18154 37510 29110 37562
rect 29162 37510 29174 37562
rect 29226 37510 29238 37562
rect 29290 37510 29302 37562
rect 29354 37510 29366 37562
rect 29418 37510 34868 37562
rect 1104 37488 34868 37510
rect 1578 37408 1584 37460
rect 1636 37448 1642 37460
rect 1673 37451 1731 37457
rect 1673 37448 1685 37451
rect 1636 37420 1685 37448
rect 1636 37408 1642 37420
rect 1673 37417 1685 37420
rect 1719 37417 1731 37451
rect 7374 37448 7380 37460
rect 7335 37420 7380 37448
rect 1673 37411 1731 37417
rect 7374 37408 7380 37420
rect 7432 37408 7438 37460
rect 8110 37448 8116 37460
rect 8071 37420 8116 37448
rect 8110 37408 8116 37420
rect 8168 37408 8174 37460
rect 9585 37451 9643 37457
rect 9585 37417 9597 37451
rect 9631 37448 9643 37451
rect 9766 37448 9772 37460
rect 9631 37420 9772 37448
rect 9631 37417 9643 37420
rect 9585 37411 9643 37417
rect 9766 37408 9772 37420
rect 9824 37408 9830 37460
rect 10870 37448 10876 37460
rect 10831 37420 10876 37448
rect 10870 37408 10876 37420
rect 10928 37408 10934 37460
rect 11333 37451 11391 37457
rect 11333 37417 11345 37451
rect 11379 37448 11391 37451
rect 12342 37448 12348 37460
rect 11379 37420 12348 37448
rect 11379 37417 11391 37420
rect 11333 37411 11391 37417
rect 12342 37408 12348 37420
rect 12400 37408 12406 37460
rect 12434 37408 12440 37460
rect 12492 37448 12498 37460
rect 16482 37448 16488 37460
rect 12492 37420 16488 37448
rect 12492 37408 12498 37420
rect 16482 37408 16488 37420
rect 16540 37408 16546 37460
rect 16850 37408 16856 37460
rect 16908 37448 16914 37460
rect 17494 37448 17500 37460
rect 16908 37420 17500 37448
rect 16908 37408 16914 37420
rect 17494 37408 17500 37420
rect 17552 37408 17558 37460
rect 17773 37451 17831 37457
rect 17773 37417 17785 37451
rect 17819 37448 17831 37451
rect 18230 37448 18236 37460
rect 17819 37420 18236 37448
rect 17819 37417 17831 37420
rect 17773 37411 17831 37417
rect 18230 37408 18236 37420
rect 18288 37408 18294 37460
rect 18322 37408 18328 37460
rect 18380 37448 18386 37460
rect 18690 37448 18696 37460
rect 18380 37420 18696 37448
rect 18380 37408 18386 37420
rect 18690 37408 18696 37420
rect 18748 37448 18754 37460
rect 19334 37448 19340 37460
rect 18748 37420 19340 37448
rect 18748 37408 18754 37420
rect 19334 37408 19340 37420
rect 19392 37408 19398 37460
rect 21450 37448 21456 37460
rect 21411 37420 21456 37448
rect 21450 37408 21456 37420
rect 21508 37408 21514 37460
rect 26145 37451 26203 37457
rect 22066 37420 25728 37448
rect 2976 37352 3188 37380
rect 1581 37247 1639 37253
rect 1581 37213 1593 37247
rect 1627 37244 1639 37247
rect 2314 37244 2320 37256
rect 1627 37216 2320 37244
rect 1627 37213 1639 37216
rect 1581 37207 1639 37213
rect 2314 37204 2320 37216
rect 2372 37204 2378 37256
rect 2409 37247 2467 37253
rect 2409 37213 2421 37247
rect 2455 37244 2467 37247
rect 2976 37244 3004 37352
rect 3053 37315 3111 37321
rect 3053 37281 3065 37315
rect 3099 37281 3111 37315
rect 3053 37275 3111 37281
rect 2455 37216 3004 37244
rect 2455 37213 2467 37216
rect 2409 37207 2467 37213
rect 3068 37188 3096 37275
rect 3160 37244 3188 37352
rect 12618 37340 12624 37392
rect 12676 37380 12682 37392
rect 15654 37380 15660 37392
rect 12676 37352 15660 37380
rect 12676 37340 12682 37352
rect 15654 37340 15660 37352
rect 15712 37340 15718 37392
rect 15746 37340 15752 37392
rect 15804 37380 15810 37392
rect 16206 37380 16212 37392
rect 15804 37352 16212 37380
rect 15804 37340 15810 37352
rect 16206 37340 16212 37352
rect 16264 37340 16270 37392
rect 17218 37380 17224 37392
rect 16868 37352 17224 37380
rect 3326 37272 3332 37324
rect 3384 37312 3390 37324
rect 5166 37312 5172 37324
rect 3384 37284 5172 37312
rect 3384 37272 3390 37284
rect 5166 37272 5172 37284
rect 5224 37272 5230 37324
rect 10226 37312 10232 37324
rect 10187 37284 10232 37312
rect 10226 37272 10232 37284
rect 10284 37272 10290 37324
rect 11532 37284 12756 37312
rect 3786 37244 3792 37256
rect 3160 37216 3792 37244
rect 3786 37204 3792 37216
rect 3844 37244 3850 37256
rect 11532 37253 11560 37284
rect 5353 37247 5411 37253
rect 5353 37244 5365 37247
rect 3844 37216 5365 37244
rect 3844 37204 3850 37216
rect 5353 37213 5365 37216
rect 5399 37213 5411 37247
rect 5353 37207 5411 37213
rect 7285 37247 7343 37253
rect 7285 37213 7297 37247
rect 7331 37213 7343 37247
rect 7285 37207 7343 37213
rect 11517 37247 11575 37253
rect 11517 37213 11529 37247
rect 11563 37213 11575 37247
rect 11517 37207 11575 37213
rect 12161 37247 12219 37253
rect 12161 37213 12173 37247
rect 12207 37213 12219 37247
rect 12161 37207 12219 37213
rect 3050 37176 3056 37188
rect 2963 37148 3056 37176
rect 3050 37136 3056 37148
rect 3108 37176 3114 37188
rect 4617 37179 4675 37185
rect 3108 37148 4384 37176
rect 3108 37136 3114 37148
rect 4356 37108 4384 37148
rect 4617 37145 4629 37179
rect 4663 37176 4675 37179
rect 4706 37176 4712 37188
rect 4663 37148 4712 37176
rect 4663 37145 4675 37148
rect 4617 37139 4675 37145
rect 4706 37136 4712 37148
rect 4764 37136 4770 37188
rect 5905 37179 5963 37185
rect 5905 37145 5917 37179
rect 5951 37176 5963 37179
rect 7006 37176 7012 37188
rect 5951 37148 7012 37176
rect 5951 37145 5963 37148
rect 5905 37139 5963 37145
rect 7006 37136 7012 37148
rect 7064 37136 7070 37188
rect 7300 37108 7328 37207
rect 12176 37176 12204 37207
rect 12434 37176 12440 37188
rect 12176 37148 12440 37176
rect 12434 37136 12440 37148
rect 12492 37136 12498 37188
rect 12728 37176 12756 37284
rect 12894 37272 12900 37324
rect 12952 37312 12958 37324
rect 16868 37312 16896 37352
rect 17218 37340 17224 37352
rect 17276 37340 17282 37392
rect 17678 37340 17684 37392
rect 17736 37380 17742 37392
rect 22066 37380 22094 37420
rect 17736 37352 22094 37380
rect 25700 37380 25728 37420
rect 26145 37417 26157 37451
rect 26191 37448 26203 37451
rect 26510 37448 26516 37460
rect 26191 37420 26516 37448
rect 26191 37417 26203 37420
rect 26145 37411 26203 37417
rect 26510 37408 26516 37420
rect 26568 37408 26574 37460
rect 31202 37408 31208 37460
rect 31260 37448 31266 37460
rect 31481 37451 31539 37457
rect 31481 37448 31493 37451
rect 31260 37420 31493 37448
rect 31260 37408 31266 37420
rect 31481 37417 31493 37420
rect 31527 37417 31539 37451
rect 31481 37411 31539 37417
rect 26326 37380 26332 37392
rect 25700 37352 26332 37380
rect 17736 37340 17742 37352
rect 26326 37340 26332 37352
rect 26384 37340 26390 37392
rect 18322 37312 18328 37324
rect 12952 37284 16896 37312
rect 16960 37284 18184 37312
rect 18283 37284 18328 37312
rect 12952 37272 12958 37284
rect 12805 37247 12863 37253
rect 12805 37213 12817 37247
rect 12851 37244 12863 37247
rect 13170 37244 13176 37256
rect 12851 37216 13176 37244
rect 12851 37213 12863 37216
rect 12805 37207 12863 37213
rect 13170 37204 13176 37216
rect 13228 37204 13234 37256
rect 13262 37204 13268 37256
rect 13320 37244 13326 37256
rect 14366 37244 14372 37256
rect 13320 37216 13365 37244
rect 14279 37216 14372 37244
rect 13320 37204 13326 37216
rect 14366 37204 14372 37216
rect 14424 37244 14430 37256
rect 15749 37247 15807 37253
rect 15749 37244 15761 37247
rect 14424 37216 15761 37244
rect 14424 37204 14430 37216
rect 15749 37213 15761 37216
rect 15795 37213 15807 37247
rect 15749 37207 15807 37213
rect 15838 37204 15844 37256
rect 15896 37244 15902 37256
rect 16960 37244 16988 37284
rect 15896 37216 16988 37244
rect 15896 37204 15902 37216
rect 17034 37204 17040 37256
rect 17092 37244 17098 37256
rect 17092 37216 17137 37244
rect 17092 37204 17098 37216
rect 17494 37204 17500 37256
rect 17552 37244 17558 37256
rect 17681 37247 17739 37253
rect 17681 37246 17693 37247
rect 17604 37244 17693 37246
rect 17552 37218 17693 37244
rect 17552 37216 17632 37218
rect 17552 37204 17558 37216
rect 17681 37213 17693 37218
rect 17727 37213 17739 37247
rect 18156 37244 18184 37284
rect 18322 37272 18328 37284
rect 18380 37272 18386 37324
rect 19150 37312 19156 37324
rect 18432 37284 19156 37312
rect 18432 37244 18460 37284
rect 19150 37272 19156 37284
rect 19208 37272 19214 37324
rect 19429 37315 19487 37321
rect 19429 37281 19441 37315
rect 19475 37312 19487 37315
rect 19794 37312 19800 37324
rect 19475 37284 19800 37312
rect 19475 37281 19487 37284
rect 19429 37275 19487 37281
rect 19794 37272 19800 37284
rect 19852 37272 19858 37324
rect 21082 37312 21088 37324
rect 21043 37284 21088 37312
rect 21082 37272 21088 37284
rect 21140 37312 21146 37324
rect 21726 37312 21732 37324
rect 21140 37284 21732 37312
rect 21140 37272 21146 37284
rect 21726 37272 21732 37284
rect 21784 37272 21790 37324
rect 22370 37312 22376 37324
rect 22331 37284 22376 37312
rect 22370 37272 22376 37284
rect 22428 37272 22434 37324
rect 24118 37272 24124 37324
rect 24176 37312 24182 37324
rect 24670 37312 24676 37324
rect 24176 37284 24676 37312
rect 24176 37272 24182 37284
rect 24670 37272 24676 37284
rect 24728 37312 24734 37324
rect 24765 37315 24823 37321
rect 24765 37312 24777 37315
rect 24728 37284 24777 37312
rect 24728 37272 24734 37284
rect 24765 37281 24777 37284
rect 24811 37281 24823 37315
rect 32858 37312 32864 37324
rect 32819 37284 32864 37312
rect 24765 37275 24823 37281
rect 18156 37216 18460 37244
rect 18509 37247 18567 37253
rect 17681 37207 17739 37213
rect 18509 37213 18521 37247
rect 18555 37244 18567 37247
rect 18598 37244 18604 37256
rect 18555 37216 18604 37244
rect 18555 37213 18567 37216
rect 18509 37207 18567 37213
rect 18598 37204 18604 37216
rect 18656 37204 18662 37256
rect 19242 37204 19248 37256
rect 19300 37244 19306 37256
rect 19613 37247 19671 37253
rect 19300 37216 19458 37244
rect 19300 37204 19306 37216
rect 15010 37176 15016 37188
rect 12728 37148 14872 37176
rect 14971 37148 15016 37176
rect 11974 37108 11980 37120
rect 4356 37080 7328 37108
rect 11935 37080 11980 37108
rect 11974 37068 11980 37080
rect 12032 37068 12038 37120
rect 12618 37108 12624 37120
rect 12579 37080 12624 37108
rect 12618 37068 12624 37080
rect 12676 37068 12682 37120
rect 13449 37111 13507 37117
rect 13449 37077 13461 37111
rect 13495 37108 13507 37111
rect 14366 37108 14372 37120
rect 13495 37080 14372 37108
rect 13495 37077 13507 37080
rect 13449 37071 13507 37077
rect 14366 37068 14372 37080
rect 14424 37068 14430 37120
rect 14844 37108 14872 37148
rect 15010 37136 15016 37148
rect 15068 37136 15074 37188
rect 16206 37136 16212 37188
rect 16264 37176 16270 37188
rect 16264 37148 16309 37176
rect 16264 37136 16270 37148
rect 16390 37136 16396 37188
rect 16448 37176 16454 37188
rect 17129 37179 17187 37185
rect 16448 37148 17080 37176
rect 16448 37136 16454 37148
rect 16666 37108 16672 37120
rect 14844 37080 16672 37108
rect 16666 37068 16672 37080
rect 16724 37068 16730 37120
rect 17052 37108 17080 37148
rect 17129 37145 17141 37179
rect 17175 37176 17187 37179
rect 17310 37176 17316 37188
rect 17175 37148 17316 37176
rect 17175 37145 17187 37148
rect 17129 37139 17187 37145
rect 17310 37136 17316 37148
rect 17368 37136 17374 37188
rect 18693 37179 18751 37185
rect 18693 37176 18705 37179
rect 17420 37148 18705 37176
rect 17420 37108 17448 37148
rect 18693 37145 18705 37148
rect 18739 37145 18751 37179
rect 18693 37139 18751 37145
rect 19337 37179 19395 37185
rect 19337 37145 19349 37179
rect 19383 37145 19395 37179
rect 19430 37176 19458 37216
rect 19613 37213 19625 37247
rect 19659 37244 19671 37247
rect 19886 37244 19892 37256
rect 19659 37216 19892 37244
rect 19659 37213 19671 37216
rect 19613 37207 19671 37213
rect 19886 37204 19892 37216
rect 19944 37204 19950 37256
rect 20254 37244 20260 37256
rect 20215 37216 20260 37244
rect 20254 37204 20260 37216
rect 20312 37204 20318 37256
rect 20346 37204 20352 37256
rect 20404 37244 20410 37256
rect 20625 37247 20683 37253
rect 20625 37244 20637 37247
rect 20404 37216 20637 37244
rect 20404 37204 20410 37216
rect 20625 37213 20637 37216
rect 20671 37213 20683 37247
rect 20625 37207 20683 37213
rect 20806 37204 20812 37256
rect 20864 37244 20870 37256
rect 21269 37247 21327 37253
rect 21269 37244 21281 37247
rect 20864 37216 21281 37244
rect 20864 37204 20870 37216
rect 21269 37213 21281 37216
rect 21315 37213 21327 37247
rect 21269 37207 21327 37213
rect 21358 37204 21364 37256
rect 21416 37244 21422 37256
rect 24302 37244 24308 37256
rect 21416 37216 24308 37244
rect 21416 37204 21422 37216
rect 24302 37204 24308 37216
rect 24360 37204 24366 37256
rect 24780 37244 24808 37275
rect 32858 37272 32864 37284
rect 32916 37272 32922 37324
rect 26605 37247 26663 37253
rect 26605 37244 26617 37247
rect 24780 37216 26617 37244
rect 26605 37213 26617 37216
rect 26651 37244 26663 37247
rect 27154 37244 27160 37256
rect 26651 37216 27160 37244
rect 26651 37213 26663 37216
rect 26605 37207 26663 37213
rect 27154 37204 27160 37216
rect 27212 37204 27218 37256
rect 28629 37247 28687 37253
rect 28629 37213 28641 37247
rect 28675 37244 28687 37247
rect 28902 37244 28908 37256
rect 28675 37216 28908 37244
rect 28675 37213 28687 37216
rect 28629 37207 28687 37213
rect 28902 37204 28908 37216
rect 28960 37244 28966 37256
rect 29917 37247 29975 37253
rect 29917 37244 29929 37247
rect 28960 37216 29929 37244
rect 28960 37204 28966 37216
rect 29917 37213 29929 37216
rect 29963 37213 29975 37247
rect 30650 37244 30656 37256
rect 30611 37216 30656 37244
rect 29917 37207 29975 37213
rect 30650 37204 30656 37216
rect 30708 37204 30714 37256
rect 32122 37244 32128 37256
rect 32083 37216 32128 37244
rect 32122 37204 32128 37216
rect 32180 37204 32186 37256
rect 20441 37179 20499 37185
rect 20441 37176 20453 37179
rect 19430 37148 20453 37176
rect 19337 37139 19395 37145
rect 20441 37145 20453 37148
rect 20487 37145 20499 37179
rect 20441 37139 20499 37145
rect 17052 37080 17448 37108
rect 17586 37068 17592 37120
rect 17644 37108 17650 37120
rect 18322 37108 18328 37120
rect 17644 37080 18328 37108
rect 17644 37068 17650 37080
rect 18322 37068 18328 37080
rect 18380 37068 18386 37120
rect 19352 37108 19380 37139
rect 20714 37136 20720 37188
rect 20772 37176 20778 37188
rect 22618 37179 22676 37185
rect 22618 37176 22630 37179
rect 20772 37148 22630 37176
rect 20772 37136 20778 37148
rect 22618 37145 22630 37148
rect 22664 37145 22676 37179
rect 22618 37139 22676 37145
rect 23216 37148 23888 37176
rect 19702 37108 19708 37120
rect 19352 37080 19708 37108
rect 19702 37068 19708 37080
rect 19760 37068 19766 37120
rect 19797 37111 19855 37117
rect 19797 37077 19809 37111
rect 19843 37108 19855 37111
rect 20254 37108 20260 37120
rect 19843 37080 20260 37108
rect 19843 37077 19855 37080
rect 19797 37071 19855 37077
rect 20254 37068 20260 37080
rect 20312 37068 20318 37120
rect 21542 37068 21548 37120
rect 21600 37108 21606 37120
rect 23216 37108 23244 37148
rect 21600 37080 23244 37108
rect 21600 37068 21606 37080
rect 23290 37068 23296 37120
rect 23348 37108 23354 37120
rect 23753 37111 23811 37117
rect 23753 37108 23765 37111
rect 23348 37080 23765 37108
rect 23348 37068 23354 37080
rect 23753 37077 23765 37080
rect 23799 37077 23811 37111
rect 23860 37108 23888 37148
rect 24854 37136 24860 37188
rect 24912 37176 24918 37188
rect 25010 37179 25068 37185
rect 25010 37176 25022 37179
rect 24912 37148 25022 37176
rect 24912 37136 24918 37148
rect 25010 37145 25022 37148
rect 25056 37145 25068 37179
rect 26234 37176 26240 37188
rect 25010 37139 25068 37145
rect 25148 37148 26240 37176
rect 25148 37108 25176 37148
rect 26234 37136 26240 37148
rect 26292 37136 26298 37188
rect 26326 37136 26332 37188
rect 26384 37176 26390 37188
rect 26850 37179 26908 37185
rect 26850 37176 26862 37179
rect 26384 37148 26862 37176
rect 26384 37136 26390 37148
rect 26850 37145 26862 37148
rect 26896 37145 26908 37179
rect 30558 37176 30564 37188
rect 26850 37139 26908 37145
rect 27908 37148 30564 37176
rect 23860 37080 25176 37108
rect 23753 37071 23811 37077
rect 25314 37068 25320 37120
rect 25372 37108 25378 37120
rect 27908 37108 27936 37148
rect 30558 37136 30564 37148
rect 30616 37136 30622 37188
rect 31294 37176 31300 37188
rect 31255 37148 31300 37176
rect 31294 37136 31300 37148
rect 31352 37136 31358 37188
rect 31513 37179 31571 37185
rect 31513 37145 31525 37179
rect 31559 37176 31571 37179
rect 32306 37176 32312 37188
rect 31559 37148 32168 37176
rect 32267 37148 32312 37176
rect 31559 37145 31571 37148
rect 31513 37139 31571 37145
rect 25372 37080 27936 37108
rect 27985 37111 28043 37117
rect 25372 37068 25378 37080
rect 27985 37077 27997 37111
rect 28031 37108 28043 37111
rect 28442 37108 28448 37120
rect 28031 37080 28448 37108
rect 28031 37077 28043 37080
rect 27985 37071 28043 37077
rect 28442 37068 28448 37080
rect 28500 37068 28506 37120
rect 28718 37108 28724 37120
rect 28679 37080 28724 37108
rect 28718 37068 28724 37080
rect 28776 37068 28782 37120
rect 31662 37108 31668 37120
rect 31623 37080 31668 37108
rect 31662 37068 31668 37080
rect 31720 37068 31726 37120
rect 32140 37108 32168 37148
rect 32306 37136 32312 37148
rect 32364 37136 32370 37188
rect 33410 37108 33416 37120
rect 32140 37080 33416 37108
rect 33410 37068 33416 37080
rect 33468 37068 33474 37120
rect 1104 37018 34868 37040
rect 1104 36966 12214 37018
rect 12266 36966 12278 37018
rect 12330 36966 12342 37018
rect 12394 36966 12406 37018
rect 12458 36966 12470 37018
rect 12522 36966 23478 37018
rect 23530 36966 23542 37018
rect 23594 36966 23606 37018
rect 23658 36966 23670 37018
rect 23722 36966 23734 37018
rect 23786 36966 34868 37018
rect 1104 36944 34868 36966
rect 4706 36864 4712 36916
rect 4764 36904 4770 36916
rect 7926 36904 7932 36916
rect 4764 36876 7932 36904
rect 4764 36864 4770 36876
rect 7926 36864 7932 36876
rect 7984 36864 7990 36916
rect 10870 36864 10876 36916
rect 10928 36904 10934 36916
rect 13446 36904 13452 36916
rect 10928 36876 13452 36904
rect 10928 36864 10934 36876
rect 13446 36864 13452 36876
rect 13504 36864 13510 36916
rect 13541 36907 13599 36913
rect 13541 36873 13553 36907
rect 13587 36904 13599 36907
rect 13587 36876 16528 36904
rect 13587 36873 13599 36876
rect 13541 36867 13599 36873
rect 1581 36839 1639 36845
rect 1581 36805 1593 36839
rect 1627 36836 1639 36839
rect 2317 36839 2375 36845
rect 2317 36836 2329 36839
rect 1627 36808 2329 36836
rect 1627 36805 1639 36808
rect 1581 36799 1639 36805
rect 2317 36805 2329 36808
rect 2363 36805 2375 36839
rect 3970 36836 3976 36848
rect 3931 36808 3976 36836
rect 2317 36799 2375 36805
rect 3970 36796 3976 36808
rect 4028 36796 4034 36848
rect 5074 36836 5080 36848
rect 4987 36808 5080 36836
rect 5074 36796 5080 36808
rect 5132 36836 5138 36848
rect 5534 36836 5540 36848
rect 5132 36808 5540 36836
rect 5132 36796 5138 36808
rect 5534 36796 5540 36808
rect 5592 36796 5598 36848
rect 12894 36836 12900 36848
rect 11808 36808 12900 36836
rect 1489 36771 1547 36777
rect 1489 36737 1501 36771
rect 1535 36737 1547 36771
rect 1489 36731 1547 36737
rect 1504 36632 1532 36731
rect 3786 36728 3792 36780
rect 3844 36768 3850 36780
rect 4525 36771 4583 36777
rect 4525 36768 4537 36771
rect 3844 36740 4537 36768
rect 3844 36728 3850 36740
rect 4525 36737 4537 36740
rect 4571 36737 4583 36771
rect 4525 36731 4583 36737
rect 5626 36728 5632 36780
rect 5684 36768 5690 36780
rect 5813 36771 5871 36777
rect 5813 36768 5825 36771
rect 5684 36740 5825 36768
rect 5684 36728 5690 36740
rect 5813 36737 5825 36740
rect 5859 36737 5871 36771
rect 5813 36731 5871 36737
rect 10321 36771 10379 36777
rect 10321 36737 10333 36771
rect 10367 36768 10379 36771
rect 10410 36768 10416 36780
rect 10367 36740 10416 36768
rect 10367 36737 10379 36740
rect 10321 36731 10379 36737
rect 10410 36728 10416 36740
rect 10468 36728 10474 36780
rect 10778 36728 10784 36780
rect 10836 36768 10842 36780
rect 11808 36777 11836 36808
rect 12894 36796 12900 36808
rect 12952 36796 12958 36848
rect 16390 36836 16396 36848
rect 13096 36808 16396 36836
rect 10965 36771 11023 36777
rect 10965 36768 10977 36771
rect 10836 36740 10977 36768
rect 10836 36728 10842 36740
rect 10965 36737 10977 36740
rect 11011 36737 11023 36771
rect 10965 36731 11023 36737
rect 11793 36771 11851 36777
rect 11793 36737 11805 36771
rect 11839 36737 11851 36771
rect 12434 36768 12440 36780
rect 12395 36740 12440 36768
rect 11793 36731 11851 36737
rect 12434 36728 12440 36740
rect 12492 36728 12498 36780
rect 13096 36777 13124 36808
rect 16390 36796 16396 36808
rect 16448 36796 16454 36848
rect 16500 36836 16528 36876
rect 16666 36864 16672 36916
rect 16724 36904 16730 36916
rect 21358 36904 21364 36916
rect 16724 36876 21364 36904
rect 16724 36864 16730 36876
rect 21358 36864 21364 36876
rect 21416 36864 21422 36916
rect 21913 36907 21971 36913
rect 21913 36873 21925 36907
rect 21959 36904 21971 36907
rect 22002 36904 22008 36916
rect 21959 36876 22008 36904
rect 21959 36873 21971 36876
rect 21913 36867 21971 36873
rect 22002 36864 22008 36876
rect 22060 36864 22066 36916
rect 22922 36864 22928 36916
rect 22980 36904 22986 36916
rect 31110 36904 31116 36916
rect 22980 36876 31116 36904
rect 22980 36864 22986 36876
rect 31110 36864 31116 36876
rect 31168 36864 31174 36916
rect 31481 36907 31539 36913
rect 31481 36873 31493 36907
rect 31527 36904 31539 36907
rect 32490 36904 32496 36916
rect 31527 36876 32496 36904
rect 31527 36873 31539 36876
rect 31481 36867 31539 36873
rect 32490 36864 32496 36876
rect 32548 36864 32554 36916
rect 16925 36839 16983 36845
rect 16925 36836 16937 36839
rect 16500 36808 16937 36836
rect 16925 36805 16937 36808
rect 16971 36805 16983 36839
rect 16925 36799 16983 36805
rect 17034 36796 17040 36848
rect 17092 36836 17098 36848
rect 17218 36836 17224 36848
rect 17092 36808 17224 36836
rect 17092 36796 17098 36808
rect 17218 36796 17224 36808
rect 17276 36836 17282 36848
rect 21542 36836 21548 36848
rect 17276 36808 18460 36836
rect 17276 36796 17282 36808
rect 13081 36771 13139 36777
rect 13081 36737 13093 36771
rect 13127 36737 13139 36771
rect 13081 36731 13139 36737
rect 13725 36771 13783 36777
rect 13725 36737 13737 36771
rect 13771 36768 13783 36771
rect 13906 36768 13912 36780
rect 13771 36740 13912 36768
rect 13771 36737 13783 36740
rect 13725 36731 13783 36737
rect 13906 36728 13912 36740
rect 13964 36728 13970 36780
rect 14366 36768 14372 36780
rect 14327 36740 14372 36768
rect 14366 36728 14372 36740
rect 14424 36728 14430 36780
rect 14462 36740 14780 36768
rect 2133 36703 2191 36709
rect 2133 36669 2145 36703
rect 2179 36700 2191 36703
rect 3878 36700 3884 36712
rect 2179 36672 3884 36700
rect 2179 36669 2191 36672
rect 2133 36663 2191 36669
rect 3878 36660 3884 36672
rect 3936 36660 3942 36712
rect 14462 36700 14490 36740
rect 12406 36672 14490 36700
rect 2682 36632 2688 36644
rect 1504 36604 2688 36632
rect 2682 36592 2688 36604
rect 2740 36592 2746 36644
rect 4798 36592 4804 36644
rect 4856 36632 4862 36644
rect 12066 36632 12072 36644
rect 4856 36604 12072 36632
rect 4856 36592 4862 36604
rect 12066 36592 12072 36604
rect 12124 36592 12130 36644
rect 11609 36567 11667 36573
rect 11609 36533 11621 36567
rect 11655 36564 11667 36567
rect 12158 36564 12164 36576
rect 11655 36536 12164 36564
rect 11655 36533 11667 36536
rect 11609 36527 11667 36533
rect 12158 36524 12164 36536
rect 12216 36524 12222 36576
rect 12253 36567 12311 36573
rect 12253 36533 12265 36567
rect 12299 36564 12311 36567
rect 12406 36564 12434 36672
rect 14550 36660 14556 36712
rect 14608 36700 14614 36712
rect 14752 36700 14780 36740
rect 15194 36728 15200 36780
rect 15252 36768 15258 36780
rect 15930 36768 15936 36780
rect 15252 36740 15936 36768
rect 15252 36728 15258 36740
rect 15930 36728 15936 36740
rect 15988 36728 15994 36780
rect 16022 36728 16028 36780
rect 16080 36768 16086 36780
rect 16080 36740 16125 36768
rect 16080 36728 16086 36740
rect 16298 36728 16304 36780
rect 16356 36768 16362 36780
rect 18230 36768 18236 36780
rect 16356 36740 18236 36768
rect 16356 36728 16362 36740
rect 18230 36728 18236 36740
rect 18288 36728 18294 36780
rect 18432 36768 18460 36808
rect 18616 36808 21548 36836
rect 18506 36768 18512 36780
rect 18419 36740 18512 36768
rect 18506 36728 18512 36740
rect 18564 36728 18570 36780
rect 16390 36700 16396 36712
rect 14608 36672 14653 36700
rect 14752 36672 16396 36700
rect 14608 36660 14614 36672
rect 16390 36660 16396 36672
rect 16448 36660 16454 36712
rect 16666 36700 16672 36712
rect 16627 36672 16672 36700
rect 16666 36660 16672 36672
rect 16724 36660 16730 36712
rect 18616 36700 18644 36808
rect 21542 36796 21548 36808
rect 21600 36796 21606 36848
rect 21726 36796 21732 36848
rect 21784 36836 21790 36848
rect 22830 36836 22836 36848
rect 21784 36808 22836 36836
rect 21784 36796 21790 36808
rect 18782 36777 18788 36780
rect 18765 36771 18788 36777
rect 18765 36737 18777 36771
rect 18765 36731 18788 36737
rect 18782 36728 18788 36731
rect 18840 36728 18846 36780
rect 19150 36728 19156 36780
rect 19208 36768 19214 36780
rect 20533 36771 20591 36777
rect 19208 36740 20484 36768
rect 19208 36728 19214 36740
rect 17696 36672 18644 36700
rect 12897 36635 12955 36641
rect 12897 36601 12909 36635
rect 12943 36632 12955 36635
rect 16482 36632 16488 36644
rect 12943 36604 16488 36632
rect 12943 36601 12955 36604
rect 12897 36595 12955 36601
rect 16482 36592 16488 36604
rect 16540 36592 16546 36644
rect 12299 36536 12434 36564
rect 12299 36533 12311 36536
rect 12253 36527 12311 36533
rect 12710 36524 12716 36576
rect 12768 36564 12774 36576
rect 17696 36564 17724 36672
rect 19518 36660 19524 36712
rect 19576 36700 19582 36712
rect 19886 36700 19892 36712
rect 19576 36672 19892 36700
rect 19576 36660 19582 36672
rect 19886 36660 19892 36672
rect 19944 36700 19950 36712
rect 20349 36703 20407 36709
rect 20349 36700 20361 36703
rect 19944 36672 20361 36700
rect 19944 36660 19950 36672
rect 20349 36669 20361 36672
rect 20395 36669 20407 36703
rect 20456 36700 20484 36740
rect 20533 36737 20545 36771
rect 20579 36768 20591 36771
rect 20622 36768 20628 36780
rect 20579 36740 20628 36768
rect 20579 36737 20591 36740
rect 20533 36731 20591 36737
rect 20622 36728 20628 36740
rect 20680 36728 20686 36780
rect 21174 36728 21180 36780
rect 21232 36768 21238 36780
rect 21818 36768 21824 36780
rect 21232 36740 21824 36768
rect 21232 36728 21238 36740
rect 21818 36728 21824 36740
rect 21876 36728 21882 36780
rect 22465 36771 22523 36777
rect 22465 36737 22477 36771
rect 22511 36768 22523 36771
rect 22554 36768 22560 36780
rect 22511 36740 22560 36768
rect 22511 36737 22523 36740
rect 22465 36731 22523 36737
rect 22554 36728 22560 36740
rect 22612 36728 22618 36780
rect 22756 36777 22784 36808
rect 22830 36796 22836 36808
rect 22888 36796 22894 36848
rect 23198 36796 23204 36848
rect 23256 36836 23262 36848
rect 25593 36839 25651 36845
rect 23256 36808 24256 36836
rect 23256 36796 23262 36808
rect 22741 36771 22799 36777
rect 22741 36737 22753 36771
rect 22787 36737 22799 36771
rect 23382 36768 23388 36780
rect 23343 36740 23388 36768
rect 22741 36731 22799 36737
rect 23382 36728 23388 36740
rect 23440 36728 23446 36780
rect 23474 36728 23480 36780
rect 23532 36768 23538 36780
rect 24228 36777 24256 36808
rect 25593 36805 25605 36839
rect 25639 36836 25651 36839
rect 25774 36836 25780 36848
rect 25639 36808 25780 36836
rect 25639 36805 25651 36808
rect 25593 36799 25651 36805
rect 25774 36796 25780 36808
rect 25832 36836 25838 36848
rect 26602 36836 26608 36848
rect 25832 36808 26608 36836
rect 25832 36796 25838 36808
rect 26602 36796 26608 36808
rect 26660 36796 26666 36848
rect 26694 36796 26700 36848
rect 26752 36836 26758 36848
rect 27402 36839 27460 36845
rect 27402 36836 27414 36839
rect 26752 36808 27414 36836
rect 26752 36796 26758 36808
rect 27402 36805 27414 36808
rect 27448 36805 27460 36839
rect 32306 36836 32312 36848
rect 27402 36799 27460 36805
rect 27540 36808 32312 36836
rect 23569 36771 23627 36777
rect 23569 36768 23581 36771
rect 23532 36740 23581 36768
rect 23532 36728 23538 36740
rect 23569 36737 23581 36740
rect 23615 36737 23627 36771
rect 23569 36731 23627 36737
rect 24213 36771 24271 36777
rect 24213 36737 24225 36771
rect 24259 36737 24271 36771
rect 24213 36731 24271 36737
rect 22649 36703 22707 36709
rect 20456 36672 22600 36700
rect 20349 36663 20407 36669
rect 17770 36592 17776 36644
rect 17828 36632 17834 36644
rect 21542 36632 21548 36644
rect 17828 36604 18552 36632
rect 17828 36592 17834 36604
rect 12768 36536 17724 36564
rect 18049 36567 18107 36573
rect 12768 36524 12774 36536
rect 18049 36533 18061 36567
rect 18095 36564 18107 36567
rect 18414 36564 18420 36576
rect 18095 36536 18420 36564
rect 18095 36533 18107 36536
rect 18049 36527 18107 36533
rect 18414 36524 18420 36536
rect 18472 36524 18478 36576
rect 18524 36564 18552 36604
rect 19781 36604 21548 36632
rect 19781 36564 19809 36604
rect 21542 36592 21548 36604
rect 21600 36592 21606 36644
rect 22572 36632 22600 36672
rect 22649 36669 22661 36703
rect 22695 36700 22707 36703
rect 23400 36700 23428 36728
rect 22695 36672 23428 36700
rect 23584 36700 23612 36731
rect 24394 36728 24400 36780
rect 24452 36768 24458 36780
rect 25866 36768 25872 36780
rect 24452 36740 24545 36768
rect 25827 36740 25872 36768
rect 24452 36728 24458 36740
rect 25866 36728 25872 36740
rect 25924 36728 25930 36780
rect 25958 36728 25964 36780
rect 26016 36768 26022 36780
rect 27540 36768 27568 36808
rect 32306 36796 32312 36808
rect 32364 36796 32370 36848
rect 26016 36740 27568 36768
rect 26016 36728 26022 36740
rect 28902 36728 28908 36780
rect 28960 36768 28966 36780
rect 29089 36771 29147 36777
rect 29089 36768 29101 36771
rect 28960 36740 29101 36768
rect 28960 36728 28966 36740
rect 29089 36737 29101 36740
rect 29135 36737 29147 36771
rect 30282 36768 30288 36780
rect 30243 36740 30288 36768
rect 29089 36731 29147 36737
rect 30282 36728 30288 36740
rect 30340 36728 30346 36780
rect 31386 36768 31392 36780
rect 31347 36740 31392 36768
rect 31386 36728 31392 36740
rect 31444 36768 31450 36780
rect 31846 36768 31852 36780
rect 31444 36740 31852 36768
rect 31444 36728 31450 36740
rect 31846 36728 31852 36740
rect 31904 36728 31910 36780
rect 34146 36768 34152 36780
rect 34107 36740 34152 36768
rect 34146 36728 34152 36740
rect 34204 36728 34210 36780
rect 24412 36700 24440 36728
rect 23584 36672 24440 36700
rect 24581 36703 24639 36709
rect 22695 36669 22707 36672
rect 22649 36663 22707 36669
rect 24581 36669 24593 36703
rect 24627 36700 24639 36703
rect 24670 36700 24676 36712
rect 24627 36672 24676 36700
rect 24627 36669 24639 36672
rect 24581 36663 24639 36669
rect 24670 36660 24676 36672
rect 24728 36660 24734 36712
rect 25777 36703 25835 36709
rect 25777 36669 25789 36703
rect 25823 36700 25835 36703
rect 26510 36700 26516 36712
rect 25823 36672 26516 36700
rect 25823 36669 25835 36672
rect 25777 36663 25835 36669
rect 26510 36660 26516 36672
rect 26568 36660 26574 36712
rect 27154 36700 27160 36712
rect 27115 36672 27160 36700
rect 27154 36660 27160 36672
rect 27212 36660 27218 36712
rect 28166 36660 28172 36712
rect 28224 36700 28230 36712
rect 29641 36703 29699 36709
rect 29641 36700 29653 36703
rect 28224 36672 29653 36700
rect 28224 36660 28230 36672
rect 29641 36669 29653 36672
rect 29687 36669 29699 36703
rect 30558 36700 30564 36712
rect 30519 36672 30564 36700
rect 29641 36663 29699 36669
rect 23566 36632 23572 36644
rect 22572 36604 23572 36632
rect 23566 36592 23572 36604
rect 23624 36592 23630 36644
rect 23658 36592 23664 36644
rect 23716 36632 23722 36644
rect 23716 36604 24256 36632
rect 23716 36592 23722 36604
rect 18524 36536 19809 36564
rect 19886 36524 19892 36576
rect 19944 36564 19950 36576
rect 20714 36564 20720 36576
rect 19944 36536 19989 36564
rect 20675 36536 20720 36564
rect 19944 36524 19950 36536
rect 20714 36524 20720 36536
rect 20772 36524 20778 36576
rect 22738 36564 22744 36576
rect 22699 36536 22744 36564
rect 22738 36524 22744 36536
rect 22796 36524 22802 36576
rect 22922 36564 22928 36576
rect 22883 36536 22928 36564
rect 22922 36524 22928 36536
rect 22980 36524 22986 36576
rect 23106 36524 23112 36576
rect 23164 36564 23170 36576
rect 23474 36564 23480 36576
rect 23164 36536 23480 36564
rect 23164 36524 23170 36536
rect 23474 36524 23480 36536
rect 23532 36524 23538 36576
rect 23750 36564 23756 36576
rect 23711 36536 23756 36564
rect 23750 36524 23756 36536
rect 23808 36524 23814 36576
rect 24228 36564 24256 36604
rect 24302 36592 24308 36644
rect 24360 36632 24366 36644
rect 24360 36604 26188 36632
rect 24360 36592 24366 36604
rect 25314 36564 25320 36576
rect 24228 36536 25320 36564
rect 25314 36524 25320 36536
rect 25372 36524 25378 36576
rect 25406 36524 25412 36576
rect 25464 36564 25470 36576
rect 25593 36567 25651 36573
rect 25593 36564 25605 36567
rect 25464 36536 25605 36564
rect 25464 36524 25470 36536
rect 25593 36533 25605 36536
rect 25639 36533 25651 36567
rect 25593 36527 25651 36533
rect 25682 36524 25688 36576
rect 25740 36564 25746 36576
rect 26053 36567 26111 36573
rect 26053 36564 26065 36567
rect 25740 36536 26065 36564
rect 25740 36524 25746 36536
rect 26053 36533 26065 36536
rect 26099 36533 26111 36567
rect 26160 36564 26188 36604
rect 27798 36564 27804 36576
rect 26160 36536 27804 36564
rect 26053 36527 26111 36533
rect 27798 36524 27804 36536
rect 27856 36524 27862 36576
rect 28350 36524 28356 36576
rect 28408 36564 28414 36576
rect 28537 36567 28595 36573
rect 28537 36564 28549 36567
rect 28408 36536 28549 36564
rect 28408 36524 28414 36536
rect 28537 36533 28549 36536
rect 28583 36533 28595 36567
rect 29656 36564 29684 36663
rect 30558 36660 30564 36672
rect 30616 36700 30622 36712
rect 31018 36700 31024 36712
rect 30616 36672 31024 36700
rect 30616 36660 30622 36672
rect 31018 36660 31024 36672
rect 31076 36660 31082 36712
rect 31938 36660 31944 36712
rect 31996 36700 32002 36712
rect 32309 36703 32367 36709
rect 32309 36700 32321 36703
rect 31996 36672 32321 36700
rect 31996 36660 32002 36672
rect 32309 36669 32321 36672
rect 32355 36669 32367 36703
rect 32309 36663 32367 36669
rect 32493 36703 32551 36709
rect 32493 36669 32505 36703
rect 32539 36669 32551 36703
rect 32493 36663 32551 36669
rect 29730 36592 29736 36644
rect 29788 36632 29794 36644
rect 32508 36632 32536 36663
rect 29788 36604 32536 36632
rect 29788 36592 29794 36604
rect 30558 36564 30564 36576
rect 29656 36536 30564 36564
rect 28537 36527 28595 36533
rect 30558 36524 30564 36536
rect 30616 36524 30622 36576
rect 30650 36524 30656 36576
rect 30708 36564 30714 36576
rect 34330 36564 34336 36576
rect 30708 36536 34336 36564
rect 30708 36524 30714 36536
rect 34330 36524 34336 36536
rect 34388 36524 34394 36576
rect 1104 36474 34868 36496
rect 1104 36422 6582 36474
rect 6634 36422 6646 36474
rect 6698 36422 6710 36474
rect 6762 36422 6774 36474
rect 6826 36422 6838 36474
rect 6890 36422 17846 36474
rect 17898 36422 17910 36474
rect 17962 36422 17974 36474
rect 18026 36422 18038 36474
rect 18090 36422 18102 36474
rect 18154 36422 29110 36474
rect 29162 36422 29174 36474
rect 29226 36422 29238 36474
rect 29290 36422 29302 36474
rect 29354 36422 29366 36474
rect 29418 36422 34868 36474
rect 1104 36400 34868 36422
rect 2314 36320 2320 36372
rect 2372 36360 2378 36372
rect 4982 36360 4988 36372
rect 2372 36332 3648 36360
rect 4943 36332 4988 36360
rect 2372 36320 2378 36332
rect 2682 36252 2688 36304
rect 2740 36292 2746 36304
rect 3620 36292 3648 36332
rect 4982 36320 4988 36332
rect 5040 36320 5046 36372
rect 10781 36363 10839 36369
rect 10781 36329 10793 36363
rect 10827 36360 10839 36363
rect 10870 36360 10876 36372
rect 10827 36332 10876 36360
rect 10827 36329 10839 36332
rect 10781 36323 10839 36329
rect 10870 36320 10876 36332
rect 10928 36320 10934 36372
rect 13630 36360 13636 36372
rect 12636 36332 13636 36360
rect 11422 36292 11428 36304
rect 2740 36264 3556 36292
rect 3620 36264 11428 36292
rect 2740 36252 2746 36264
rect 1397 36227 1455 36233
rect 1397 36193 1409 36227
rect 1443 36224 1455 36227
rect 2406 36224 2412 36236
rect 1443 36196 2412 36224
rect 1443 36193 1455 36196
rect 1397 36187 1455 36193
rect 2406 36184 2412 36196
rect 2464 36184 2470 36236
rect 2774 36224 2780 36236
rect 2735 36196 2780 36224
rect 2774 36184 2780 36196
rect 2832 36184 2838 36236
rect 3528 36224 3556 36264
rect 11422 36252 11428 36264
rect 11480 36252 11486 36304
rect 11606 36292 11612 36304
rect 11567 36264 11612 36292
rect 11606 36252 11612 36264
rect 11664 36252 11670 36304
rect 12069 36295 12127 36301
rect 12069 36261 12081 36295
rect 12115 36292 12127 36295
rect 12636 36292 12664 36332
rect 13630 36320 13636 36332
rect 13688 36320 13694 36372
rect 13906 36320 13912 36372
rect 13964 36360 13970 36372
rect 15838 36360 15844 36372
rect 13964 36332 15844 36360
rect 13964 36320 13970 36332
rect 15838 36320 15844 36332
rect 15896 36320 15902 36372
rect 15933 36363 15991 36369
rect 15933 36329 15945 36363
rect 15979 36360 15991 36363
rect 16114 36360 16120 36372
rect 15979 36332 16120 36360
rect 15979 36329 15991 36332
rect 15933 36323 15991 36329
rect 16114 36320 16120 36332
rect 16172 36320 16178 36372
rect 16206 36320 16212 36372
rect 16264 36360 16270 36372
rect 16853 36363 16911 36369
rect 16853 36360 16865 36363
rect 16264 36332 16865 36360
rect 16264 36320 16270 36332
rect 16853 36329 16865 36332
rect 16899 36329 16911 36363
rect 16853 36323 16911 36329
rect 16942 36320 16948 36372
rect 17000 36360 17006 36372
rect 18690 36360 18696 36372
rect 17000 36332 18552 36360
rect 18651 36332 18696 36360
rect 17000 36320 17006 36332
rect 12115 36264 12664 36292
rect 12115 36261 12127 36264
rect 12069 36255 12127 36261
rect 12894 36252 12900 36304
rect 12952 36292 12958 36304
rect 16390 36292 16396 36304
rect 12952 36264 16396 36292
rect 12952 36252 12958 36264
rect 16390 36252 16396 36264
rect 16448 36252 16454 36304
rect 17310 36292 17316 36304
rect 16500 36264 17316 36292
rect 12342 36224 12348 36236
rect 3528 36196 12348 36224
rect 12342 36184 12348 36196
rect 12400 36184 12406 36236
rect 12434 36184 12440 36236
rect 12492 36224 12498 36236
rect 16500 36233 16528 36264
rect 17310 36252 17316 36264
rect 17368 36252 17374 36304
rect 18524 36292 18552 36332
rect 18690 36320 18696 36332
rect 18748 36320 18754 36372
rect 20714 36360 20720 36372
rect 18791 36332 20720 36360
rect 18791 36292 18819 36332
rect 20714 36320 20720 36332
rect 20772 36320 20778 36372
rect 21542 36320 21548 36372
rect 21600 36360 21606 36372
rect 23750 36360 23756 36372
rect 21600 36332 23756 36360
rect 21600 36320 21606 36332
rect 23750 36320 23756 36332
rect 23808 36320 23814 36372
rect 24026 36320 24032 36372
rect 24084 36360 24090 36372
rect 25777 36363 25835 36369
rect 24084 36332 25452 36360
rect 24084 36320 24090 36332
rect 18524 36264 18819 36292
rect 23290 36252 23296 36304
rect 23348 36252 23354 36304
rect 23566 36292 23572 36304
rect 23527 36264 23572 36292
rect 23566 36252 23572 36264
rect 23624 36252 23630 36304
rect 16485 36227 16543 36233
rect 12492 36196 15976 36224
rect 12492 36184 12498 36196
rect 3510 36116 3516 36168
rect 3568 36156 3574 36168
rect 3786 36156 3792 36168
rect 3568 36128 3792 36156
rect 3568 36116 3574 36128
rect 3786 36116 3792 36128
rect 3844 36156 3850 36168
rect 3881 36159 3939 36165
rect 3881 36156 3893 36159
rect 3844 36128 3893 36156
rect 3844 36116 3850 36128
rect 3881 36125 3893 36128
rect 3927 36125 3939 36159
rect 4430 36156 4436 36168
rect 4391 36128 4436 36156
rect 3881 36119 3939 36125
rect 4430 36116 4436 36128
rect 4488 36116 4494 36168
rect 5166 36156 5172 36168
rect 5127 36128 5172 36156
rect 5166 36116 5172 36128
rect 5224 36116 5230 36168
rect 10965 36159 11023 36165
rect 10965 36125 10977 36159
rect 11011 36156 11023 36159
rect 11330 36156 11336 36168
rect 11011 36128 11336 36156
rect 11011 36125 11023 36128
rect 10965 36119 11023 36125
rect 11330 36116 11336 36128
rect 11388 36116 11394 36168
rect 12253 36159 12311 36165
rect 12253 36125 12265 36159
rect 12299 36156 12311 36159
rect 12802 36156 12808 36168
rect 12299 36128 12808 36156
rect 12299 36125 12311 36128
rect 12253 36119 12311 36125
rect 12802 36116 12808 36128
rect 12860 36116 12866 36168
rect 12894 36116 12900 36168
rect 12952 36156 12958 36168
rect 13538 36156 13544 36168
rect 12952 36128 12997 36156
rect 13499 36128 13544 36156
rect 12952 36116 12958 36128
rect 13538 36116 13544 36128
rect 13596 36116 13602 36168
rect 14277 36159 14335 36165
rect 14277 36125 14289 36159
rect 14323 36156 14335 36159
rect 14366 36156 14372 36168
rect 14323 36128 14372 36156
rect 14323 36125 14335 36128
rect 14277 36119 14335 36125
rect 14366 36116 14372 36128
rect 14424 36116 14430 36168
rect 14458 36116 14464 36168
rect 14516 36156 14522 36168
rect 14918 36156 14924 36168
rect 14516 36128 14924 36156
rect 14516 36116 14522 36128
rect 14918 36116 14924 36128
rect 14976 36116 14982 36168
rect 15286 36116 15292 36168
rect 15344 36156 15350 36168
rect 15470 36156 15476 36168
rect 15344 36128 15476 36156
rect 15344 36116 15350 36128
rect 15470 36116 15476 36128
rect 15528 36116 15534 36168
rect 15841 36159 15899 36165
rect 15841 36125 15853 36159
rect 15887 36125 15899 36159
rect 15948 36156 15976 36196
rect 16485 36193 16497 36227
rect 16531 36193 16543 36227
rect 16942 36224 16948 36236
rect 16485 36187 16543 36193
rect 16592 36196 16948 36224
rect 16592 36156 16620 36196
rect 16942 36184 16948 36196
rect 17000 36184 17006 36236
rect 17236 36196 17428 36224
rect 15948 36128 16620 36156
rect 16669 36159 16727 36165
rect 15841 36119 15899 36125
rect 16669 36125 16681 36159
rect 16715 36156 16727 36159
rect 16758 36156 16764 36168
rect 16715 36128 16764 36156
rect 16715 36125 16727 36128
rect 16669 36119 16727 36125
rect 1578 36088 1584 36100
rect 1539 36060 1584 36088
rect 1578 36048 1584 36060
rect 1636 36048 1642 36100
rect 13722 36048 13728 36100
rect 13780 36088 13786 36100
rect 14645 36091 14703 36097
rect 14645 36088 14657 36091
rect 13780 36060 14657 36088
rect 13780 36048 13786 36060
rect 14645 36057 14657 36060
rect 14691 36088 14703 36091
rect 15194 36088 15200 36100
rect 14691 36060 15200 36088
rect 14691 36057 14703 36060
rect 14645 36051 14703 36057
rect 15194 36048 15200 36060
rect 15252 36048 15258 36100
rect 15562 36048 15568 36100
rect 15620 36088 15626 36100
rect 15856 36088 15884 36119
rect 16758 36116 16764 36128
rect 16816 36116 16822 36168
rect 17236 36156 17264 36196
rect 16868 36128 17264 36156
rect 17313 36159 17371 36165
rect 16868 36088 16896 36128
rect 17313 36125 17325 36159
rect 17359 36125 17371 36159
rect 17400 36156 17428 36196
rect 18506 36184 18512 36236
rect 18564 36224 18570 36236
rect 18690 36224 18696 36236
rect 18564 36196 18696 36224
rect 18564 36184 18570 36196
rect 18690 36184 18696 36196
rect 18748 36224 18754 36236
rect 19521 36227 19579 36233
rect 19521 36224 19533 36227
rect 18748 36196 19533 36224
rect 18748 36184 18754 36196
rect 19521 36193 19533 36196
rect 19567 36193 19579 36227
rect 19521 36187 19579 36193
rect 18966 36156 18972 36168
rect 17400 36128 18972 36156
rect 17313 36119 17371 36125
rect 15620 36060 16896 36088
rect 15620 36048 15626 36060
rect 16942 36048 16948 36100
rect 17000 36088 17006 36100
rect 17126 36088 17132 36100
rect 17000 36060 17132 36088
rect 17000 36048 17006 36060
rect 17126 36048 17132 36060
rect 17184 36048 17190 36100
rect 17218 36048 17224 36100
rect 17276 36088 17282 36100
rect 17328 36088 17356 36119
rect 18966 36116 18972 36128
rect 19024 36116 19030 36168
rect 19536 36156 19564 36187
rect 20530 36184 20536 36236
rect 20588 36224 20594 36236
rect 20588 36196 21496 36224
rect 20588 36184 20594 36196
rect 21266 36156 21272 36168
rect 19536 36128 21272 36156
rect 21266 36116 21272 36128
rect 21324 36156 21330 36168
rect 21361 36159 21419 36165
rect 21361 36156 21373 36159
rect 21324 36128 21373 36156
rect 21324 36116 21330 36128
rect 21361 36125 21373 36128
rect 21407 36125 21419 36159
rect 21468 36156 21496 36196
rect 21617 36159 21675 36165
rect 21617 36156 21629 36159
rect 21468 36128 21629 36156
rect 21361 36119 21419 36125
rect 21617 36125 21629 36128
rect 21663 36125 21675 36159
rect 22370 36156 22376 36168
rect 21617 36119 21675 36125
rect 21744 36128 22376 36156
rect 17276 36060 17356 36088
rect 17580 36091 17638 36097
rect 17276 36048 17282 36060
rect 17580 36057 17592 36091
rect 17626 36057 17638 36091
rect 17580 36051 17638 36057
rect 12710 36020 12716 36032
rect 12671 35992 12716 36020
rect 12710 35980 12716 35992
rect 12768 35980 12774 36032
rect 13354 36020 13360 36032
rect 13315 35992 13360 36020
rect 13354 35980 13360 35992
rect 13412 35980 13418 36032
rect 13538 35980 13544 36032
rect 13596 36020 13602 36032
rect 14366 36020 14372 36032
rect 13596 35992 14372 36020
rect 13596 35980 13602 35992
rect 14366 35980 14372 35992
rect 14424 35980 14430 36032
rect 15010 35980 15016 36032
rect 15068 36020 15074 36032
rect 17590 36020 17618 36051
rect 17770 36048 17776 36100
rect 17828 36088 17834 36100
rect 19766 36091 19824 36097
rect 19766 36088 19778 36091
rect 17828 36060 19778 36088
rect 17828 36048 17834 36060
rect 19766 36057 19778 36060
rect 19812 36057 19824 36091
rect 21376 36088 21404 36119
rect 21744 36088 21772 36128
rect 22370 36116 22376 36128
rect 22428 36116 22434 36168
rect 22738 36116 22744 36168
rect 22796 36156 22802 36168
rect 23201 36159 23259 36165
rect 23201 36156 23213 36159
rect 22796 36128 23213 36156
rect 22796 36116 22802 36128
rect 23201 36125 23213 36128
rect 23247 36156 23259 36159
rect 23308 36156 23336 36252
rect 24118 36184 24124 36236
rect 24176 36224 24182 36236
rect 24397 36227 24455 36233
rect 24397 36224 24409 36227
rect 24176 36196 24409 36224
rect 24176 36184 24182 36196
rect 24397 36193 24409 36196
rect 24443 36193 24455 36227
rect 25424 36224 25452 36332
rect 25777 36329 25789 36363
rect 25823 36360 25835 36363
rect 25866 36360 25872 36372
rect 25823 36332 25872 36360
rect 25823 36329 25835 36332
rect 25777 36323 25835 36329
rect 25866 36320 25872 36332
rect 25924 36320 25930 36372
rect 28350 36360 28356 36372
rect 27540 36332 28356 36360
rect 25498 36252 25504 36304
rect 25556 36292 25562 36304
rect 25682 36292 25688 36304
rect 25556 36264 25688 36292
rect 25556 36252 25562 36264
rect 25682 36252 25688 36264
rect 25740 36252 25746 36304
rect 25884 36292 25912 36320
rect 26237 36295 26295 36301
rect 26237 36292 26249 36295
rect 25884 36264 26249 36292
rect 26237 36261 26249 36264
rect 26283 36261 26295 36295
rect 26237 36255 26295 36261
rect 25958 36224 25964 36236
rect 25424 36196 25964 36224
rect 24397 36187 24455 36193
rect 25958 36184 25964 36196
rect 26016 36184 26022 36236
rect 26142 36184 26148 36236
rect 26200 36224 26206 36236
rect 27540 36233 27568 36332
rect 28350 36320 28356 36332
rect 28408 36320 28414 36372
rect 28442 36320 28448 36372
rect 28500 36360 28506 36372
rect 28537 36363 28595 36369
rect 28537 36360 28549 36363
rect 28500 36332 28549 36360
rect 28500 36320 28506 36332
rect 28537 36329 28549 36332
rect 28583 36329 28595 36363
rect 28537 36323 28595 36329
rect 29638 36320 29644 36372
rect 29696 36360 29702 36372
rect 30006 36360 30012 36372
rect 29696 36332 30012 36360
rect 29696 36320 29702 36332
rect 30006 36320 30012 36332
rect 30064 36320 30070 36372
rect 27890 36252 27896 36304
rect 27948 36292 27954 36304
rect 27948 36264 32536 36292
rect 27948 36252 27954 36264
rect 27525 36227 27583 36233
rect 27525 36224 27537 36227
rect 26200 36196 27537 36224
rect 26200 36184 26206 36196
rect 27525 36193 27537 36196
rect 27571 36193 27583 36227
rect 28442 36224 28448 36236
rect 27525 36187 27583 36193
rect 27724 36196 28448 36224
rect 23247 36128 23336 36156
rect 23371 36159 23429 36165
rect 23247 36125 23259 36128
rect 23201 36119 23259 36125
rect 23371 36125 23383 36159
rect 23417 36156 23429 36159
rect 23474 36156 23480 36168
rect 23417 36128 23480 36156
rect 23417 36125 23429 36128
rect 23371 36119 23429 36125
rect 23474 36116 23480 36128
rect 23532 36116 23538 36168
rect 27724 36165 27752 36196
rect 28442 36184 28448 36196
rect 28500 36184 28506 36236
rect 28721 36227 28779 36233
rect 28721 36193 28733 36227
rect 28767 36224 28779 36227
rect 28994 36224 29000 36236
rect 28767 36196 29000 36224
rect 28767 36193 28779 36196
rect 28721 36187 28779 36193
rect 27709 36159 27767 36165
rect 27709 36125 27721 36159
rect 27755 36125 27767 36159
rect 27709 36119 27767 36125
rect 27798 36116 27804 36168
rect 27856 36156 27862 36168
rect 28077 36159 28135 36165
rect 28077 36156 28089 36159
rect 27856 36128 28089 36156
rect 27856 36116 27862 36128
rect 28077 36125 28089 36128
rect 28123 36125 28135 36159
rect 28736 36156 28764 36187
rect 28994 36184 29000 36196
rect 29052 36184 29058 36236
rect 31110 36224 31116 36236
rect 31071 36196 31116 36224
rect 31110 36184 31116 36196
rect 31168 36184 31174 36236
rect 32306 36224 32312 36236
rect 32267 36196 32312 36224
rect 32306 36184 32312 36196
rect 32364 36184 32370 36236
rect 32508 36233 32536 36264
rect 32493 36227 32551 36233
rect 32493 36193 32505 36227
rect 32539 36193 32551 36227
rect 32950 36224 32956 36236
rect 32911 36196 32956 36224
rect 32493 36187 32551 36193
rect 32950 36184 32956 36196
rect 33008 36184 33014 36236
rect 28077 36119 28135 36125
rect 28460 36128 28764 36156
rect 28813 36159 28871 36165
rect 24642 36091 24700 36097
rect 24642 36088 24654 36091
rect 19766 36051 19824 36057
rect 19904 36060 21036 36088
rect 21376 36060 21772 36088
rect 22066 36060 24654 36088
rect 15068 35992 17618 36020
rect 15068 35980 15074 35992
rect 17678 35980 17684 36032
rect 17736 36020 17742 36032
rect 18506 36020 18512 36032
rect 17736 35992 18512 36020
rect 17736 35980 17742 35992
rect 18506 35980 18512 35992
rect 18564 35980 18570 36032
rect 18782 35980 18788 36032
rect 18840 36020 18846 36032
rect 19904 36020 19932 36060
rect 18840 35992 19932 36020
rect 18840 35980 18846 35992
rect 19978 35980 19984 36032
rect 20036 36020 20042 36032
rect 20901 36023 20959 36029
rect 20901 36020 20913 36023
rect 20036 35992 20913 36020
rect 20036 35980 20042 35992
rect 20901 35989 20913 35992
rect 20947 35989 20959 36023
rect 21008 36020 21036 36060
rect 22066 36020 22094 36060
rect 24642 36057 24654 36060
rect 24688 36057 24700 36091
rect 24642 36051 24700 36057
rect 25406 36048 25412 36100
rect 25464 36088 25470 36100
rect 26421 36091 26479 36097
rect 26421 36088 26433 36091
rect 25464 36060 26433 36088
rect 25464 36048 25470 36060
rect 26421 36057 26433 36060
rect 26467 36057 26479 36091
rect 26602 36088 26608 36100
rect 26563 36060 26608 36088
rect 26421 36051 26479 36057
rect 26602 36048 26608 36060
rect 26660 36048 26666 36100
rect 28460 36088 28488 36128
rect 28813 36125 28825 36159
rect 28859 36125 28871 36159
rect 29638 36156 29644 36168
rect 29599 36128 29644 36156
rect 28813 36119 28871 36125
rect 27816 36060 28488 36088
rect 21008 35992 22094 36020
rect 20901 35983 20959 35989
rect 22370 35980 22376 36032
rect 22428 36020 22434 36032
rect 22741 36023 22799 36029
rect 22741 36020 22753 36023
rect 22428 35992 22753 36020
rect 22428 35980 22434 35992
rect 22741 35989 22753 35992
rect 22787 35989 22799 36023
rect 22741 35983 22799 35989
rect 22922 35980 22928 36032
rect 22980 36020 22986 36032
rect 25958 36020 25964 36032
rect 22980 35992 25964 36020
rect 22980 35980 22986 35992
rect 25958 35980 25964 35992
rect 26016 35980 26022 36032
rect 26510 35980 26516 36032
rect 26568 36020 26574 36032
rect 26789 36023 26847 36029
rect 26568 35992 26613 36020
rect 26568 35980 26574 35992
rect 26789 35989 26801 36023
rect 26835 36020 26847 36023
rect 27614 36020 27620 36032
rect 26835 35992 27620 36020
rect 26835 35989 26847 35992
rect 26789 35983 26847 35989
rect 27614 35980 27620 35992
rect 27672 35980 27678 36032
rect 27816 36029 27844 36060
rect 28534 36048 28540 36100
rect 28592 36088 28598 36100
rect 28592 36060 28637 36088
rect 28592 36048 28598 36060
rect 27801 36023 27859 36029
rect 27801 35989 27813 36023
rect 27847 35989 27859 36023
rect 27801 35983 27859 35989
rect 27890 35980 27896 36032
rect 27948 36020 27954 36032
rect 27948 35992 27993 36020
rect 27948 35980 27954 35992
rect 28350 35980 28356 36032
rect 28408 36020 28414 36032
rect 28828 36020 28856 36119
rect 29638 36116 29644 36128
rect 29696 36156 29702 36168
rect 30282 36156 30288 36168
rect 29696 36128 30288 36156
rect 29696 36116 29702 36128
rect 30282 36116 30288 36128
rect 30340 36156 30346 36168
rect 30837 36159 30895 36165
rect 30837 36156 30849 36159
rect 30340 36128 30849 36156
rect 30340 36116 30346 36128
rect 30837 36125 30849 36128
rect 30883 36125 30895 36159
rect 30837 36119 30895 36125
rect 30193 36091 30251 36097
rect 30193 36057 30205 36091
rect 30239 36088 30251 36091
rect 30374 36088 30380 36100
rect 30239 36060 30380 36088
rect 30239 36057 30251 36060
rect 30193 36051 30251 36057
rect 30374 36048 30380 36060
rect 30432 36048 30438 36100
rect 28408 35992 28856 36020
rect 28997 36023 29055 36029
rect 28408 35980 28414 35992
rect 28997 35989 29009 36023
rect 29043 36020 29055 36023
rect 29546 36020 29552 36032
rect 29043 35992 29552 36020
rect 29043 35989 29055 35992
rect 28997 35983 29055 35989
rect 29546 35980 29552 35992
rect 29604 35980 29610 36032
rect 1104 35930 34868 35952
rect 1104 35878 12214 35930
rect 12266 35878 12278 35930
rect 12330 35878 12342 35930
rect 12394 35878 12406 35930
rect 12458 35878 12470 35930
rect 12522 35878 23478 35930
rect 23530 35878 23542 35930
rect 23594 35878 23606 35930
rect 23658 35878 23670 35930
rect 23722 35878 23734 35930
rect 23786 35878 34868 35930
rect 1104 35856 34868 35878
rect 1578 35776 1584 35828
rect 1636 35816 1642 35828
rect 2225 35819 2283 35825
rect 2225 35816 2237 35819
rect 1636 35788 2237 35816
rect 1636 35776 1642 35788
rect 2225 35785 2237 35788
rect 2271 35785 2283 35819
rect 2225 35779 2283 35785
rect 3237 35819 3295 35825
rect 3237 35785 3249 35819
rect 3283 35816 3295 35819
rect 3510 35816 3516 35828
rect 3283 35788 3516 35816
rect 3283 35785 3295 35788
rect 3237 35779 3295 35785
rect 3510 35776 3516 35788
rect 3568 35776 3574 35828
rect 11698 35776 11704 35828
rect 11756 35816 11762 35828
rect 11885 35819 11943 35825
rect 11885 35816 11897 35819
rect 11756 35788 11897 35816
rect 11756 35776 11762 35788
rect 11885 35785 11897 35788
rect 11931 35785 11943 35819
rect 11885 35779 11943 35785
rect 13173 35819 13231 35825
rect 13173 35785 13185 35819
rect 13219 35816 13231 35819
rect 13219 35788 16252 35816
rect 13219 35785 13231 35788
rect 13173 35779 13231 35785
rect 13262 35748 13268 35760
rect 3068 35720 13268 35748
rect 1394 35680 1400 35692
rect 1355 35652 1400 35680
rect 1394 35640 1400 35652
rect 1452 35640 1458 35692
rect 2130 35680 2136 35692
rect 2091 35652 2136 35680
rect 2130 35640 2136 35652
rect 2188 35640 2194 35692
rect 3068 35689 3096 35720
rect 13262 35708 13268 35720
rect 13320 35708 13326 35760
rect 16117 35751 16175 35757
rect 16117 35748 16129 35751
rect 13372 35720 16129 35748
rect 3053 35683 3111 35689
rect 3053 35649 3065 35683
rect 3099 35649 3111 35683
rect 3053 35643 3111 35649
rect 1581 35547 1639 35553
rect 1581 35513 1593 35547
rect 1627 35544 1639 35547
rect 3068 35544 3096 35643
rect 3878 35640 3884 35692
rect 3936 35680 3942 35692
rect 3973 35683 4031 35689
rect 3973 35680 3985 35683
rect 3936 35652 3985 35680
rect 3936 35640 3942 35652
rect 3973 35649 3985 35652
rect 4019 35649 4031 35683
rect 4614 35680 4620 35692
rect 4575 35652 4620 35680
rect 3973 35643 4031 35649
rect 4614 35640 4620 35652
rect 4672 35640 4678 35692
rect 12069 35683 12127 35689
rect 12069 35649 12081 35683
rect 12115 35649 12127 35683
rect 12069 35643 12127 35649
rect 12713 35683 12771 35689
rect 12713 35649 12725 35683
rect 12759 35680 12771 35683
rect 13170 35680 13176 35692
rect 12759 35652 13176 35680
rect 12759 35649 12771 35652
rect 12713 35643 12771 35649
rect 12084 35612 12112 35643
rect 13170 35640 13176 35652
rect 13228 35640 13234 35692
rect 13372 35689 13400 35720
rect 16117 35717 16129 35720
rect 16163 35717 16175 35751
rect 16224 35748 16252 35788
rect 16758 35776 16764 35828
rect 16816 35816 16822 35828
rect 18690 35816 18696 35828
rect 16816 35788 18696 35816
rect 16816 35776 16822 35788
rect 18690 35776 18696 35788
rect 18748 35776 18754 35828
rect 19334 35776 19340 35828
rect 19392 35816 19398 35828
rect 19521 35819 19579 35825
rect 19521 35816 19533 35819
rect 19392 35788 19533 35816
rect 19392 35776 19398 35788
rect 19521 35785 19533 35788
rect 19567 35785 19579 35819
rect 19521 35779 19579 35785
rect 19628 35788 20024 35816
rect 16914 35751 16972 35757
rect 16914 35748 16926 35751
rect 16224 35720 16926 35748
rect 16117 35711 16175 35717
rect 16914 35717 16926 35720
rect 16960 35717 16972 35751
rect 16914 35711 16972 35717
rect 17126 35708 17132 35760
rect 17184 35748 17190 35760
rect 19628 35748 19656 35788
rect 17184 35720 19656 35748
rect 17184 35708 17190 35720
rect 19702 35708 19708 35760
rect 19760 35748 19766 35760
rect 19886 35748 19892 35760
rect 19760 35720 19892 35748
rect 19760 35708 19766 35720
rect 19886 35708 19892 35720
rect 19944 35708 19950 35760
rect 19996 35748 20024 35788
rect 20070 35776 20076 35828
rect 20128 35816 20134 35828
rect 20530 35816 20536 35828
rect 20128 35788 20536 35816
rect 20128 35776 20134 35788
rect 20530 35776 20536 35788
rect 20588 35776 20594 35828
rect 21358 35776 21364 35828
rect 21416 35816 21422 35828
rect 21416 35788 22416 35816
rect 21416 35776 21422 35788
rect 20990 35748 20996 35760
rect 19996 35720 20996 35748
rect 20990 35708 20996 35720
rect 21048 35708 21054 35760
rect 22094 35757 22100 35760
rect 22088 35711 22100 35757
rect 22152 35748 22158 35760
rect 22388 35748 22416 35788
rect 22462 35776 22468 35828
rect 22520 35816 22526 35828
rect 23753 35819 23811 35825
rect 23753 35816 23765 35819
rect 22520 35788 23765 35816
rect 22520 35776 22526 35788
rect 23753 35785 23765 35788
rect 23799 35785 23811 35819
rect 23753 35779 23811 35785
rect 25685 35819 25743 35825
rect 25685 35785 25697 35819
rect 25731 35816 25743 35819
rect 25774 35816 25780 35828
rect 25731 35788 25780 35816
rect 25731 35785 25743 35788
rect 25685 35779 25743 35785
rect 25774 35776 25780 35788
rect 25832 35776 25838 35828
rect 28994 35776 29000 35828
rect 29052 35816 29058 35828
rect 30469 35819 30527 35825
rect 30469 35816 30481 35819
rect 29052 35788 30481 35816
rect 29052 35776 29058 35788
rect 30469 35785 30481 35788
rect 30515 35785 30527 35819
rect 30469 35779 30527 35785
rect 24210 35748 24216 35760
rect 22152 35720 22188 35748
rect 22388 35720 24216 35748
rect 22094 35708 22100 35711
rect 22152 35708 22158 35720
rect 13357 35683 13415 35689
rect 13357 35649 13369 35683
rect 13403 35649 13415 35683
rect 13357 35643 13415 35649
rect 14001 35683 14059 35689
rect 14001 35649 14013 35683
rect 14047 35649 14059 35683
rect 14001 35643 14059 35649
rect 13906 35612 13912 35624
rect 12084 35584 13912 35612
rect 13906 35572 13912 35584
rect 13964 35572 13970 35624
rect 14016 35612 14044 35643
rect 14366 35640 14372 35692
rect 14424 35680 14430 35692
rect 14645 35683 14703 35689
rect 14645 35680 14657 35683
rect 14424 35652 14657 35680
rect 14424 35640 14430 35652
rect 14645 35649 14657 35652
rect 14691 35649 14703 35683
rect 14645 35643 14703 35649
rect 15105 35683 15163 35689
rect 15105 35649 15117 35683
rect 15151 35680 15163 35683
rect 15286 35680 15292 35692
rect 15151 35652 15292 35680
rect 15151 35649 15163 35652
rect 15105 35643 15163 35649
rect 15286 35640 15292 35652
rect 15344 35640 15350 35692
rect 15580 35652 15884 35680
rect 14918 35612 14924 35624
rect 14016 35584 14924 35612
rect 14918 35572 14924 35584
rect 14976 35572 14982 35624
rect 15197 35615 15255 35621
rect 15197 35581 15209 35615
rect 15243 35612 15255 35615
rect 15580 35612 15608 35652
rect 15746 35612 15752 35624
rect 15243 35584 15608 35612
rect 15707 35584 15752 35612
rect 15243 35581 15255 35584
rect 15197 35575 15255 35581
rect 15746 35572 15752 35584
rect 15804 35572 15810 35624
rect 15856 35612 15884 35652
rect 15930 35640 15936 35692
rect 15988 35680 15994 35692
rect 15988 35652 16033 35680
rect 15988 35640 15994 35652
rect 16206 35640 16212 35692
rect 16264 35640 16270 35692
rect 16390 35640 16396 35692
rect 16448 35680 16454 35692
rect 16448 35678 16804 35680
rect 16951 35678 17724 35680
rect 16448 35652 17724 35678
rect 16448 35640 16454 35652
rect 16776 35650 16979 35652
rect 16224 35612 16252 35640
rect 15856 35584 16252 35612
rect 16482 35572 16488 35624
rect 16540 35572 16546 35624
rect 16666 35612 16672 35624
rect 16627 35584 16672 35612
rect 16666 35572 16672 35584
rect 16724 35572 16730 35624
rect 17696 35612 17724 35652
rect 17770 35640 17776 35692
rect 17828 35680 17834 35692
rect 18414 35680 18420 35692
rect 17828 35652 18420 35680
rect 17828 35640 17834 35652
rect 18414 35640 18420 35652
rect 18472 35680 18478 35692
rect 18509 35683 18567 35689
rect 18509 35680 18521 35683
rect 18472 35652 18521 35680
rect 18472 35640 18478 35652
rect 18509 35649 18521 35652
rect 18555 35649 18567 35683
rect 18690 35680 18696 35692
rect 18651 35652 18696 35680
rect 18509 35643 18567 35649
rect 18690 35640 18696 35652
rect 18748 35640 18754 35692
rect 19613 35683 19671 35689
rect 19613 35649 19625 35683
rect 19659 35680 19671 35683
rect 19794 35680 19800 35692
rect 19659 35652 19800 35680
rect 19659 35649 19671 35652
rect 19613 35643 19671 35649
rect 19794 35640 19800 35652
rect 19852 35680 19858 35692
rect 20533 35683 20591 35689
rect 19852 35652 20484 35680
rect 19852 35640 19858 35652
rect 19337 35615 19395 35621
rect 17696 35584 18276 35612
rect 12526 35544 12532 35556
rect 1627 35516 3096 35544
rect 12487 35516 12532 35544
rect 1627 35513 1639 35516
rect 1581 35507 1639 35513
rect 12526 35504 12532 35516
rect 12584 35504 12590 35556
rect 13170 35504 13176 35556
rect 13228 35544 13234 35556
rect 16500 35544 16528 35572
rect 18248 35544 18276 35584
rect 19337 35581 19349 35615
rect 19383 35612 19395 35615
rect 19426 35612 19432 35624
rect 19383 35584 19432 35612
rect 19383 35581 19395 35584
rect 19337 35575 19395 35581
rect 19426 35572 19432 35584
rect 19484 35572 19490 35624
rect 19527 35584 20024 35612
rect 19527 35544 19555 35584
rect 13228 35516 16528 35544
rect 17590 35516 18184 35544
rect 18248 35516 19555 35544
rect 19889 35547 19947 35553
rect 13228 35504 13234 35516
rect 2130 35436 2136 35488
rect 2188 35476 2194 35488
rect 13446 35476 13452 35488
rect 2188 35448 13452 35476
rect 2188 35436 2194 35448
rect 13446 35436 13452 35448
rect 13504 35436 13510 35488
rect 13814 35436 13820 35488
rect 13872 35476 13878 35488
rect 14458 35476 14464 35488
rect 13872 35448 13917 35476
rect 14419 35448 14464 35476
rect 13872 35436 13878 35448
rect 14458 35436 14464 35448
rect 14516 35436 14522 35488
rect 14918 35436 14924 35488
rect 14976 35476 14982 35488
rect 17590 35476 17618 35516
rect 14976 35448 17618 35476
rect 14976 35436 14982 35448
rect 17770 35436 17776 35488
rect 17828 35476 17834 35488
rect 18049 35479 18107 35485
rect 18049 35476 18061 35479
rect 17828 35448 18061 35476
rect 17828 35436 17834 35448
rect 18049 35445 18061 35448
rect 18095 35445 18107 35479
rect 18156 35476 18184 35516
rect 19889 35513 19901 35547
rect 19935 35513 19947 35547
rect 19996 35544 20024 35584
rect 20070 35572 20076 35624
rect 20128 35612 20134 35624
rect 20349 35615 20407 35621
rect 20349 35612 20361 35615
rect 20128 35584 20361 35612
rect 20128 35572 20134 35584
rect 20349 35581 20361 35584
rect 20395 35581 20407 35615
rect 20456 35612 20484 35652
rect 20533 35649 20545 35683
rect 20579 35680 20591 35683
rect 20622 35680 20628 35692
rect 20579 35652 20628 35680
rect 20579 35649 20591 35652
rect 20533 35643 20591 35649
rect 20622 35640 20628 35652
rect 20680 35640 20686 35692
rect 22370 35680 22376 35692
rect 20732 35652 22376 35680
rect 20732 35612 20760 35652
rect 22370 35640 22376 35652
rect 22428 35640 22434 35692
rect 22554 35640 22560 35692
rect 22612 35680 22618 35692
rect 23566 35680 23572 35692
rect 22612 35652 23572 35680
rect 22612 35640 22618 35652
rect 23566 35640 23572 35652
rect 23624 35640 23630 35692
rect 23676 35689 23704 35720
rect 24210 35708 24216 35720
rect 24268 35708 24274 35760
rect 27264 35720 28994 35748
rect 23661 35683 23719 35689
rect 23661 35649 23673 35683
rect 23707 35649 23719 35683
rect 23661 35643 23719 35649
rect 24118 35640 24124 35692
rect 24176 35680 24182 35692
rect 24305 35683 24363 35689
rect 24305 35680 24317 35683
rect 24176 35652 24317 35680
rect 24176 35640 24182 35652
rect 24305 35649 24317 35652
rect 24351 35649 24363 35683
rect 24561 35683 24619 35689
rect 24561 35680 24573 35683
rect 24305 35643 24363 35649
rect 24392 35652 24573 35680
rect 20456 35584 20760 35612
rect 20349 35575 20407 35581
rect 21266 35572 21272 35624
rect 21324 35612 21330 35624
rect 21821 35615 21879 35621
rect 21821 35612 21833 35615
rect 21324 35584 21833 35612
rect 21324 35572 21330 35584
rect 21821 35581 21833 35584
rect 21867 35581 21879 35615
rect 24392 35612 24420 35652
rect 24561 35649 24573 35652
rect 24607 35649 24619 35683
rect 26234 35680 26240 35692
rect 26195 35652 26240 35680
rect 24561 35643 24619 35649
rect 26234 35640 26240 35652
rect 26292 35640 26298 35692
rect 26421 35683 26479 35689
rect 26421 35649 26433 35683
rect 26467 35680 26479 35683
rect 27062 35680 27068 35692
rect 26467 35652 27068 35680
rect 26467 35649 26479 35652
rect 26421 35643 26479 35649
rect 27062 35640 27068 35652
rect 27120 35640 27126 35692
rect 27154 35640 27160 35692
rect 27212 35680 27218 35692
rect 27264 35689 27292 35720
rect 27249 35683 27307 35689
rect 27249 35680 27261 35683
rect 27212 35652 27261 35680
rect 27212 35640 27218 35652
rect 27249 35649 27261 35652
rect 27295 35649 27307 35683
rect 27505 35683 27563 35689
rect 27505 35680 27517 35683
rect 27249 35643 27307 35649
rect 27356 35652 27517 35680
rect 21821 35575 21879 35581
rect 23446 35584 24420 35612
rect 20717 35547 20775 35553
rect 20717 35544 20729 35547
rect 19996 35516 20729 35544
rect 19889 35507 19947 35513
rect 20717 35513 20729 35516
rect 20763 35513 20775 35547
rect 23446 35544 23474 35584
rect 25314 35572 25320 35624
rect 25372 35612 25378 35624
rect 27356 35612 27384 35652
rect 27505 35649 27517 35652
rect 27551 35649 27563 35683
rect 27505 35643 27563 35649
rect 27890 35640 27896 35692
rect 27948 35680 27954 35692
rect 28534 35680 28540 35692
rect 27948 35652 28540 35680
rect 27948 35640 27954 35652
rect 28534 35640 28540 35652
rect 28592 35680 28598 35692
rect 28592 35652 28672 35680
rect 28592 35640 28598 35652
rect 25372 35584 27384 35612
rect 25372 35572 25378 35584
rect 26694 35544 26700 35556
rect 20717 35507 20775 35513
rect 22756 35516 23474 35544
rect 25240 35516 26700 35544
rect 18877 35479 18935 35485
rect 18877 35476 18889 35479
rect 18156 35448 18889 35476
rect 18049 35439 18107 35445
rect 18877 35445 18889 35448
rect 18923 35445 18935 35479
rect 18877 35439 18935 35445
rect 19518 35436 19524 35488
rect 19576 35476 19582 35488
rect 19904 35476 19932 35507
rect 19576 35448 19932 35476
rect 19576 35436 19582 35448
rect 20346 35436 20352 35488
rect 20404 35476 20410 35488
rect 22756 35476 22784 35516
rect 20404 35448 22784 35476
rect 20404 35436 20410 35448
rect 22922 35436 22928 35488
rect 22980 35476 22986 35488
rect 23201 35479 23259 35485
rect 23201 35476 23213 35479
rect 22980 35448 23213 35476
rect 22980 35436 22986 35448
rect 23201 35445 23213 35448
rect 23247 35445 23259 35479
rect 23201 35439 23259 35445
rect 23290 35436 23296 35488
rect 23348 35476 23354 35488
rect 25240 35476 25268 35516
rect 26694 35504 26700 35516
rect 26752 35504 26758 35556
rect 28644 35553 28672 35652
rect 28966 35612 28994 35720
rect 29178 35708 29184 35760
rect 29236 35748 29242 35760
rect 29236 35720 30144 35748
rect 29236 35708 29242 35720
rect 29356 35683 29414 35689
rect 29356 35649 29368 35683
rect 29402 35680 29414 35683
rect 29914 35680 29920 35692
rect 29402 35652 29920 35680
rect 29402 35649 29414 35652
rect 29356 35643 29414 35649
rect 29914 35640 29920 35652
rect 29972 35640 29978 35692
rect 29089 35615 29147 35621
rect 29089 35612 29101 35615
rect 28966 35584 29101 35612
rect 29089 35581 29101 35584
rect 29135 35581 29147 35615
rect 29089 35575 29147 35581
rect 28629 35547 28687 35553
rect 28629 35513 28641 35547
rect 28675 35513 28687 35547
rect 28629 35507 28687 35513
rect 23348 35448 25268 35476
rect 23348 35436 23354 35448
rect 25774 35436 25780 35488
rect 25832 35476 25838 35488
rect 27982 35476 27988 35488
rect 25832 35448 27988 35476
rect 25832 35436 25838 35448
rect 27982 35436 27988 35448
rect 28040 35436 28046 35488
rect 29104 35476 29132 35575
rect 30116 35544 30144 35720
rect 31294 35708 31300 35760
rect 31352 35748 31358 35760
rect 32490 35748 32496 35760
rect 31352 35720 32496 35748
rect 31352 35708 31358 35720
rect 31404 35689 31432 35720
rect 32490 35708 32496 35720
rect 32548 35708 32554 35760
rect 31389 35683 31447 35689
rect 31389 35649 31401 35683
rect 31435 35649 31447 35683
rect 31389 35643 31447 35649
rect 32030 35640 32036 35692
rect 32088 35680 32094 35692
rect 32125 35683 32183 35689
rect 32125 35680 32137 35683
rect 32088 35652 32137 35680
rect 32088 35640 32094 35652
rect 32125 35649 32137 35652
rect 32171 35649 32183 35683
rect 32125 35643 32183 35649
rect 32309 35683 32367 35689
rect 32309 35649 32321 35683
rect 32355 35680 32367 35683
rect 32398 35680 32404 35692
rect 32355 35652 32404 35680
rect 32355 35649 32367 35652
rect 32309 35643 32367 35649
rect 32398 35640 32404 35652
rect 32456 35640 32462 35692
rect 33318 35680 33324 35692
rect 33279 35652 33324 35680
rect 33318 35640 33324 35652
rect 33376 35640 33382 35692
rect 31205 35615 31263 35621
rect 31205 35581 31217 35615
rect 31251 35612 31263 35615
rect 32493 35615 32551 35621
rect 32493 35612 32505 35615
rect 31251 35584 32505 35612
rect 31251 35581 31263 35584
rect 31205 35575 31263 35581
rect 32493 35581 32505 35584
rect 32539 35581 32551 35615
rect 32493 35575 32551 35581
rect 33597 35615 33655 35621
rect 33597 35581 33609 35615
rect 33643 35581 33655 35615
rect 33597 35575 33655 35581
rect 33612 35544 33640 35575
rect 30116 35516 33640 35544
rect 29454 35476 29460 35488
rect 29104 35448 29460 35476
rect 29454 35436 29460 35448
rect 29512 35436 29518 35488
rect 30466 35436 30472 35488
rect 30524 35476 30530 35488
rect 31573 35479 31631 35485
rect 31573 35476 31585 35479
rect 30524 35448 31585 35476
rect 30524 35436 30530 35448
rect 31573 35445 31585 35448
rect 31619 35476 31631 35479
rect 32214 35476 32220 35488
rect 31619 35448 32220 35476
rect 31619 35445 31631 35448
rect 31573 35439 31631 35445
rect 32214 35436 32220 35448
rect 32272 35436 32278 35488
rect 1104 35386 34868 35408
rect 1104 35334 6582 35386
rect 6634 35334 6646 35386
rect 6698 35334 6710 35386
rect 6762 35334 6774 35386
rect 6826 35334 6838 35386
rect 6890 35334 17846 35386
rect 17898 35334 17910 35386
rect 17962 35334 17974 35386
rect 18026 35334 18038 35386
rect 18090 35334 18102 35386
rect 18154 35334 29110 35386
rect 29162 35334 29174 35386
rect 29226 35334 29238 35386
rect 29290 35334 29302 35386
rect 29354 35334 29366 35386
rect 29418 35334 34868 35386
rect 1104 35312 34868 35334
rect 1762 35232 1768 35284
rect 1820 35272 1826 35284
rect 12069 35275 12127 35281
rect 1820 35244 6914 35272
rect 1820 35232 1826 35244
rect 2774 35136 2780 35148
rect 2735 35108 2780 35136
rect 2774 35096 2780 35108
rect 2832 35096 2838 35148
rect 6886 35136 6914 35244
rect 12069 35241 12081 35275
rect 12115 35272 12127 35275
rect 14090 35272 14096 35284
rect 12115 35244 14096 35272
rect 12115 35241 12127 35244
rect 12069 35235 12127 35241
rect 14090 35232 14096 35244
rect 14148 35232 14154 35284
rect 14277 35275 14335 35281
rect 14277 35241 14289 35275
rect 14323 35272 14335 35275
rect 15010 35272 15016 35284
rect 14323 35244 15016 35272
rect 14323 35241 14335 35244
rect 14277 35235 14335 35241
rect 15010 35232 15016 35244
rect 15068 35232 15074 35284
rect 15746 35232 15752 35284
rect 15804 35272 15810 35284
rect 16942 35272 16948 35284
rect 15804 35244 16948 35272
rect 15804 35232 15810 35244
rect 16942 35232 16948 35244
rect 17000 35232 17006 35284
rect 17126 35232 17132 35284
rect 17184 35272 17190 35284
rect 18322 35272 18328 35284
rect 17184 35244 18328 35272
rect 17184 35232 17190 35244
rect 18322 35232 18328 35244
rect 18380 35232 18386 35284
rect 20717 35275 20775 35281
rect 20717 35272 20729 35275
rect 18524 35244 20729 35272
rect 13170 35204 13176 35216
rect 13131 35176 13176 35204
rect 13170 35164 13176 35176
rect 13228 35164 13234 35216
rect 14918 35204 14924 35216
rect 14879 35176 14924 35204
rect 14918 35164 14924 35176
rect 14976 35164 14982 35216
rect 15194 35164 15200 35216
rect 15252 35204 15258 35216
rect 15252 35176 15608 35204
rect 15252 35164 15258 35176
rect 14274 35136 14280 35148
rect 6886 35108 14280 35136
rect 14274 35096 14280 35108
rect 14332 35096 14338 35148
rect 15470 35136 15476 35148
rect 14476 35108 15476 35136
rect 1394 35068 1400 35080
rect 1355 35040 1400 35068
rect 1394 35028 1400 35040
rect 1452 35028 1458 35080
rect 12713 35071 12771 35077
rect 12713 35037 12725 35071
rect 12759 35037 12771 35071
rect 12713 35031 12771 35037
rect 1581 35003 1639 35009
rect 1581 34969 1593 35003
rect 1627 35000 1639 35003
rect 2038 35000 2044 35012
rect 1627 34972 2044 35000
rect 1627 34969 1639 34972
rect 1581 34963 1639 34969
rect 2038 34960 2044 34972
rect 2096 34960 2102 35012
rect 12728 35000 12756 35031
rect 12802 35028 12808 35080
rect 12860 35068 12866 35080
rect 13357 35071 13415 35077
rect 13357 35068 13369 35071
rect 12860 35040 13369 35068
rect 12860 35028 12866 35040
rect 13357 35037 13369 35040
rect 13403 35068 13415 35071
rect 13538 35068 13544 35080
rect 13403 35040 13544 35068
rect 13403 35037 13415 35040
rect 13357 35031 13415 35037
rect 13538 35028 13544 35040
rect 13596 35028 13602 35080
rect 13906 35068 13912 35080
rect 13740 35040 13912 35068
rect 13740 35000 13768 35040
rect 13906 35028 13912 35040
rect 13964 35028 13970 35080
rect 14476 35077 14504 35108
rect 15470 35096 15476 35108
rect 15528 35096 15534 35148
rect 15580 35136 15608 35176
rect 16574 35164 16580 35216
rect 16632 35204 16638 35216
rect 18524 35204 18552 35244
rect 20717 35241 20729 35244
rect 20763 35241 20775 35275
rect 20717 35235 20775 35241
rect 20898 35232 20904 35284
rect 20956 35272 20962 35284
rect 20956 35244 22508 35272
rect 20956 35232 20962 35244
rect 19334 35204 19340 35216
rect 16632 35176 18552 35204
rect 18616 35176 19340 35204
rect 16632 35164 16638 35176
rect 15580 35108 15700 35136
rect 14461 35071 14519 35077
rect 14461 35037 14473 35071
rect 14507 35037 14519 35071
rect 14461 35031 14519 35037
rect 14642 35028 14648 35080
rect 14700 35068 14706 35080
rect 15105 35071 15163 35077
rect 15105 35068 15117 35071
rect 14700 35040 15117 35068
rect 14700 35028 14706 35040
rect 15105 35037 15117 35040
rect 15151 35037 15163 35071
rect 15105 35031 15163 35037
rect 15286 35028 15292 35080
rect 15344 35068 15350 35080
rect 15565 35071 15623 35077
rect 15565 35068 15577 35071
rect 15344 35040 15577 35068
rect 15344 35028 15350 35040
rect 15565 35037 15577 35040
rect 15611 35037 15623 35071
rect 15672 35068 15700 35108
rect 16666 35096 16672 35148
rect 16724 35136 16730 35148
rect 17218 35136 17224 35148
rect 16724 35108 17224 35136
rect 16724 35096 16730 35108
rect 17218 35096 17224 35108
rect 17276 35096 17282 35148
rect 17310 35096 17316 35148
rect 17368 35136 17374 35148
rect 18616 35136 18644 35176
rect 19334 35164 19340 35176
rect 19392 35164 19398 35216
rect 19610 35164 19616 35216
rect 19668 35204 19674 35216
rect 20806 35204 20812 35216
rect 19668 35176 20812 35204
rect 19668 35164 19674 35176
rect 20806 35164 20812 35176
rect 20864 35164 20870 35216
rect 22480 35204 22508 35244
rect 23382 35232 23388 35284
rect 23440 35272 23446 35284
rect 23440 35244 23485 35272
rect 23440 35232 23446 35244
rect 23566 35232 23572 35284
rect 23624 35272 23630 35284
rect 23624 35244 31754 35272
rect 23624 35232 23630 35244
rect 25314 35204 25320 35216
rect 22480 35176 25320 35204
rect 25314 35164 25320 35176
rect 25372 35164 25378 35216
rect 27062 35164 27068 35216
rect 27120 35204 27126 35216
rect 29638 35204 29644 35216
rect 27120 35176 29644 35204
rect 27120 35164 27126 35176
rect 29638 35164 29644 35176
rect 29696 35164 29702 35216
rect 30466 35204 30472 35216
rect 29748 35176 30472 35204
rect 17368 35108 18644 35136
rect 18693 35139 18751 35145
rect 17368 35096 17374 35108
rect 18693 35105 18705 35139
rect 18739 35136 18751 35139
rect 18782 35136 18788 35148
rect 18739 35108 18788 35136
rect 18739 35105 18751 35108
rect 18693 35099 18751 35105
rect 18782 35096 18788 35108
rect 18840 35136 18846 35148
rect 19150 35136 19156 35148
rect 18840 35108 19156 35136
rect 18840 35096 18846 35108
rect 19150 35096 19156 35108
rect 19208 35096 19214 35148
rect 21082 35136 21088 35148
rect 19260 35108 21088 35136
rect 17034 35068 17040 35080
rect 15672 35040 17040 35068
rect 15565 35031 15623 35037
rect 17034 35028 17040 35040
rect 17092 35028 17098 35080
rect 17405 35071 17463 35077
rect 17405 35037 17417 35071
rect 17451 35068 17463 35071
rect 17494 35068 17500 35080
rect 17451 35040 17500 35068
rect 17451 35037 17463 35040
rect 17405 35031 17463 35037
rect 17494 35028 17500 35040
rect 17552 35028 17558 35080
rect 17681 35071 17739 35077
rect 17681 35037 17693 35071
rect 17727 35068 17739 35071
rect 17770 35068 17776 35080
rect 17727 35040 17776 35068
rect 17727 35037 17739 35040
rect 17681 35031 17739 35037
rect 17770 35028 17776 35040
rect 17828 35028 17834 35080
rect 18414 35028 18420 35080
rect 18472 35068 18478 35080
rect 18509 35071 18567 35077
rect 18509 35068 18521 35071
rect 18472 35040 18521 35068
rect 18472 35028 18478 35040
rect 18509 35037 18521 35040
rect 18555 35037 18567 35071
rect 18509 35031 18567 35037
rect 18598 35028 18604 35080
rect 18656 35068 18662 35080
rect 19260 35068 19288 35108
rect 21082 35096 21088 35108
rect 21140 35096 21146 35148
rect 21266 35096 21272 35148
rect 21324 35136 21330 35148
rect 21545 35139 21603 35145
rect 21545 35136 21557 35139
rect 21324 35108 21557 35136
rect 21324 35096 21330 35108
rect 21545 35105 21557 35108
rect 21591 35105 21603 35139
rect 21545 35099 21603 35105
rect 22572 35108 24716 35136
rect 18656 35040 19288 35068
rect 19429 35071 19487 35077
rect 18656 35028 18662 35040
rect 19429 35037 19441 35071
rect 19475 35037 19487 35071
rect 19429 35031 19487 35037
rect 12728 34972 13768 35000
rect 13814 34960 13820 35012
rect 13872 35000 13878 35012
rect 15810 35003 15868 35009
rect 15810 35000 15822 35003
rect 13872 34972 15822 35000
rect 13872 34960 13878 34972
rect 15810 34969 15822 34972
rect 15856 34969 15868 35003
rect 15810 34963 15868 34969
rect 15930 34960 15936 35012
rect 15988 35000 15994 35012
rect 16574 35000 16580 35012
rect 15988 34972 16580 35000
rect 15988 34960 15994 34972
rect 16574 34960 16580 34972
rect 16632 34960 16638 35012
rect 17218 34960 17224 35012
rect 17276 35000 17282 35012
rect 18966 35000 18972 35012
rect 17276 34972 18972 35000
rect 17276 34960 17282 34972
rect 18966 34960 18972 34972
rect 19024 34960 19030 35012
rect 19444 35000 19472 35031
rect 19518 35028 19524 35080
rect 19576 35068 19582 35080
rect 19886 35068 19892 35080
rect 19576 35040 19621 35068
rect 19847 35040 19892 35068
rect 19576 35028 19582 35040
rect 19886 35028 19892 35040
rect 19944 35028 19950 35080
rect 20254 35068 20260 35080
rect 19996 35040 20260 35068
rect 19610 35000 19616 35012
rect 19076 34972 19472 35000
rect 19571 34972 19616 35000
rect 12529 34935 12587 34941
rect 12529 34901 12541 34935
rect 12575 34932 12587 34935
rect 14366 34932 14372 34944
rect 12575 34904 14372 34932
rect 12575 34901 12587 34904
rect 12529 34895 12587 34901
rect 14366 34892 14372 34904
rect 14424 34892 14430 34944
rect 14550 34892 14556 34944
rect 14608 34932 14614 34944
rect 17034 34932 17040 34944
rect 14608 34904 17040 34932
rect 14608 34892 14614 34904
rect 17034 34892 17040 34904
rect 17092 34892 17098 34944
rect 17402 34892 17408 34944
rect 17460 34932 17466 34944
rect 17589 34935 17647 34941
rect 17589 34932 17601 34935
rect 17460 34904 17601 34932
rect 17460 34892 17466 34904
rect 17589 34901 17601 34904
rect 17635 34901 17647 34935
rect 17589 34895 17647 34901
rect 17770 34892 17776 34944
rect 17828 34932 17834 34944
rect 17957 34935 18015 34941
rect 17828 34904 17873 34932
rect 17828 34892 17834 34904
rect 17957 34901 17969 34935
rect 18003 34932 18015 34935
rect 19076 34932 19104 34972
rect 19610 34960 19616 34972
rect 19668 34960 19674 35012
rect 19751 35003 19809 35009
rect 19751 34969 19763 35003
rect 19797 35000 19809 35003
rect 19996 35000 20024 35040
rect 20254 35028 20260 35040
rect 20312 35028 20318 35080
rect 20438 35068 20444 35080
rect 20399 35040 20444 35068
rect 20438 35028 20444 35040
rect 20496 35028 20502 35080
rect 20533 35071 20591 35077
rect 20533 35037 20545 35071
rect 20579 35068 20591 35071
rect 20622 35068 20628 35080
rect 20579 35040 20628 35068
rect 20579 35037 20591 35040
rect 20533 35031 20591 35037
rect 20622 35028 20628 35040
rect 20680 35028 20686 35080
rect 20806 35028 20812 35080
rect 20864 35068 20870 35080
rect 22572 35068 22600 35108
rect 23290 35068 23296 35080
rect 20864 35040 22600 35068
rect 22848 35040 23296 35068
rect 20864 35028 20870 35040
rect 19797 34972 20024 35000
rect 19797 34969 19809 34972
rect 19751 34963 19809 34969
rect 20070 34960 20076 35012
rect 20128 35000 20134 35012
rect 21790 35003 21848 35009
rect 21790 35000 21802 35003
rect 20128 34972 21802 35000
rect 20128 34960 20134 34972
rect 21790 34969 21802 34972
rect 21836 34969 21848 35003
rect 21790 34963 21848 34969
rect 18003 34904 19104 34932
rect 18003 34901 18015 34904
rect 17957 34895 18015 34901
rect 19150 34892 19156 34944
rect 19208 34932 19214 34944
rect 19245 34935 19303 34941
rect 19245 34932 19257 34935
rect 19208 34904 19257 34932
rect 19208 34892 19214 34904
rect 19245 34901 19257 34904
rect 19291 34901 19303 34935
rect 19245 34895 19303 34901
rect 19334 34892 19340 34944
rect 19392 34932 19398 34944
rect 22848 34932 22876 35040
rect 23290 35028 23296 35040
rect 23348 35028 23354 35080
rect 23474 35028 23480 35080
rect 23532 35068 23538 35080
rect 23569 35071 23627 35077
rect 23569 35068 23581 35071
rect 23532 35040 23581 35068
rect 23532 35028 23538 35040
rect 23569 35037 23581 35040
rect 23615 35037 23627 35071
rect 23569 35031 23627 35037
rect 23661 35071 23719 35077
rect 23661 35037 23673 35071
rect 23707 35037 23719 35071
rect 24578 35068 24584 35080
rect 24539 35040 24584 35068
rect 23661 35031 23719 35037
rect 23198 35000 23204 35012
rect 22940 34972 23204 35000
rect 22940 34941 22968 34972
rect 23198 34960 23204 34972
rect 23256 35000 23262 35012
rect 23385 35003 23443 35009
rect 23385 35000 23397 35003
rect 23256 34972 23397 35000
rect 23256 34960 23262 34972
rect 23385 34969 23397 34972
rect 23431 34969 23443 35003
rect 23385 34963 23443 34969
rect 19392 34904 22876 34932
rect 22925 34935 22983 34941
rect 19392 34892 19398 34904
rect 22925 34901 22937 34935
rect 22971 34901 22983 34935
rect 22925 34895 22983 34901
rect 23014 34892 23020 34944
rect 23072 34932 23078 34944
rect 23676 34932 23704 35031
rect 24578 35028 24584 35040
rect 24636 35028 24642 35080
rect 24688 35068 24716 35108
rect 24854 35096 24860 35148
rect 24912 35136 24918 35148
rect 25041 35139 25099 35145
rect 25041 35136 25053 35139
rect 24912 35108 25053 35136
rect 24912 35096 24918 35108
rect 25041 35105 25053 35108
rect 25087 35105 25099 35139
rect 25041 35099 25099 35105
rect 25130 35096 25136 35148
rect 25188 35136 25194 35148
rect 25685 35139 25743 35145
rect 25685 35136 25697 35139
rect 25188 35108 25697 35136
rect 25188 35096 25194 35108
rect 25685 35105 25697 35108
rect 25731 35105 25743 35139
rect 25685 35099 25743 35105
rect 26694 35096 26700 35148
rect 26752 35136 26758 35148
rect 29362 35136 29368 35148
rect 26752 35108 29368 35136
rect 26752 35096 26758 35108
rect 29362 35096 29368 35108
rect 29420 35096 29426 35148
rect 26418 35068 26424 35080
rect 24688 35040 26424 35068
rect 26418 35028 26424 35040
rect 26476 35028 26482 35080
rect 27614 35028 27620 35080
rect 27672 35068 27678 35080
rect 27709 35071 27767 35077
rect 27709 35068 27721 35071
rect 27672 35040 27721 35068
rect 27672 35028 27678 35040
rect 27709 35037 27721 35040
rect 27755 35037 27767 35071
rect 27709 35031 27767 35037
rect 27798 35028 27804 35080
rect 27856 35068 27862 35080
rect 27856 35040 27901 35068
rect 27856 35028 27862 35040
rect 27982 35028 27988 35080
rect 28040 35077 28046 35080
rect 28040 35071 28069 35077
rect 28057 35037 28069 35071
rect 28040 35031 28069 35037
rect 28040 35028 28046 35031
rect 28166 35028 28172 35080
rect 28224 35068 28230 35080
rect 29549 35071 29607 35077
rect 28224 35040 28269 35068
rect 28644 35040 29500 35068
rect 28224 35028 28230 35040
rect 28644 35012 28672 35040
rect 23750 34960 23756 35012
rect 23808 35000 23814 35012
rect 24670 35000 24676 35012
rect 23808 34972 24532 35000
rect 24631 34972 24676 35000
rect 23808 34960 23814 34972
rect 23842 34932 23848 34944
rect 23072 34904 23704 34932
rect 23803 34904 23848 34932
rect 23072 34892 23078 34904
rect 23842 34892 23848 34904
rect 23900 34892 23906 34944
rect 24394 34932 24400 34944
rect 24355 34904 24400 34932
rect 24394 34892 24400 34904
rect 24452 34892 24458 34944
rect 24504 34932 24532 34972
rect 24670 34960 24676 34972
rect 24728 34960 24734 35012
rect 24762 34960 24768 35012
rect 24820 35000 24826 35012
rect 24903 35003 24961 35009
rect 24820 34972 24865 35000
rect 24820 34960 24854 34972
rect 24903 34969 24915 35003
rect 24949 35000 24961 35003
rect 25952 35003 26010 35009
rect 24949 34972 25912 35000
rect 24949 34969 24961 34972
rect 24903 34963 24961 34969
rect 24826 34932 24854 34960
rect 24504 34904 24854 34932
rect 25884 34932 25912 34972
rect 25952 34969 25964 35003
rect 25998 35000 26010 35003
rect 27525 35003 27583 35009
rect 27525 35000 27537 35003
rect 25998 34972 27537 35000
rect 25998 34969 26010 34972
rect 25952 34963 26010 34969
rect 27525 34969 27537 34972
rect 27571 34969 27583 35003
rect 27525 34963 27583 34969
rect 27893 35003 27951 35009
rect 27893 34969 27905 35003
rect 27939 35000 27951 35003
rect 28350 35000 28356 35012
rect 27939 34972 28356 35000
rect 27939 34969 27951 34972
rect 27893 34963 27951 34969
rect 28350 34960 28356 34972
rect 28408 34960 28414 35012
rect 28626 35000 28632 35012
rect 28587 34972 28632 35000
rect 28626 34960 28632 34972
rect 28684 34960 28690 35012
rect 28813 35003 28871 35009
rect 28813 34969 28825 35003
rect 28859 34969 28871 35003
rect 29472 35000 29500 35040
rect 29549 35037 29561 35071
rect 29595 35068 29607 35071
rect 29638 35068 29644 35080
rect 29595 35040 29644 35068
rect 29595 35037 29607 35040
rect 29549 35031 29607 35037
rect 29638 35028 29644 35040
rect 29696 35028 29702 35080
rect 29748 35000 29776 35176
rect 30466 35164 30472 35176
rect 30524 35164 30530 35216
rect 31726 35136 31754 35244
rect 31849 35207 31907 35213
rect 31849 35173 31861 35207
rect 31895 35204 31907 35207
rect 32398 35204 32404 35216
rect 31895 35176 32404 35204
rect 31895 35173 31907 35176
rect 31849 35167 31907 35173
rect 32398 35164 32404 35176
rect 32456 35204 32462 35216
rect 33502 35204 33508 35216
rect 32456 35176 33508 35204
rect 32456 35164 32462 35176
rect 33502 35164 33508 35176
rect 33560 35164 33566 35216
rect 32309 35139 32367 35145
rect 32309 35136 32321 35139
rect 31726 35108 32321 35136
rect 32309 35105 32321 35108
rect 32355 35105 32367 35139
rect 32309 35099 32367 35105
rect 30466 35068 30472 35080
rect 30379 35040 30472 35068
rect 30466 35028 30472 35040
rect 30524 35068 30530 35080
rect 31938 35068 31944 35080
rect 30524 35040 31944 35068
rect 30524 35028 30530 35040
rect 31938 35028 31944 35040
rect 31996 35028 32002 35080
rect 29472 34972 29776 35000
rect 29825 35003 29883 35009
rect 28813 34963 28871 34969
rect 29825 34969 29837 35003
rect 29871 35000 29883 35003
rect 30190 35000 30196 35012
rect 29871 34972 30196 35000
rect 29871 34969 29883 34972
rect 29825 34963 29883 34969
rect 26142 34932 26148 34944
rect 25884 34904 26148 34932
rect 26142 34892 26148 34904
rect 26200 34892 26206 34944
rect 27065 34935 27123 34941
rect 27065 34901 27077 34935
rect 27111 34932 27123 34935
rect 27430 34932 27436 34944
rect 27111 34904 27436 34932
rect 27111 34901 27123 34904
rect 27065 34895 27123 34901
rect 27430 34892 27436 34904
rect 27488 34892 27494 34944
rect 28534 34892 28540 34944
rect 28592 34932 28598 34944
rect 28828 34932 28856 34963
rect 30190 34960 30196 34972
rect 30248 34960 30254 35012
rect 30736 35003 30794 35009
rect 30736 34969 30748 35003
rect 30782 35000 30794 35003
rect 32122 35000 32128 35012
rect 30782 34972 32128 35000
rect 30782 34969 30794 34972
rect 30736 34963 30794 34969
rect 32122 34960 32128 34972
rect 32180 34960 32186 35012
rect 32493 35003 32551 35009
rect 32493 35000 32505 35003
rect 32416 34972 32505 35000
rect 32416 34944 32444 34972
rect 32493 34969 32505 34972
rect 32539 34969 32551 35003
rect 34146 35000 34152 35012
rect 34107 34972 34152 35000
rect 32493 34963 32551 34969
rect 34146 34960 34152 34972
rect 34204 34960 34210 35012
rect 28592 34904 28856 34932
rect 28997 34935 29055 34941
rect 28592 34892 28598 34904
rect 28997 34901 29009 34935
rect 29043 34932 29055 34935
rect 31294 34932 31300 34944
rect 29043 34904 31300 34932
rect 29043 34901 29055 34904
rect 28997 34895 29055 34901
rect 31294 34892 31300 34904
rect 31352 34892 31358 34944
rect 32398 34892 32404 34944
rect 32456 34892 32462 34944
rect 1104 34842 34868 34864
rect 1104 34790 12214 34842
rect 12266 34790 12278 34842
rect 12330 34790 12342 34842
rect 12394 34790 12406 34842
rect 12458 34790 12470 34842
rect 12522 34790 23478 34842
rect 23530 34790 23542 34842
rect 23594 34790 23606 34842
rect 23658 34790 23670 34842
rect 23722 34790 23734 34842
rect 23786 34790 34868 34842
rect 1104 34768 34868 34790
rect 12710 34728 12716 34740
rect 12671 34700 12716 34728
rect 12710 34688 12716 34700
rect 12768 34688 12774 34740
rect 13354 34728 13360 34740
rect 13315 34700 13360 34728
rect 13354 34688 13360 34700
rect 13412 34688 13418 34740
rect 14829 34731 14887 34737
rect 14829 34697 14841 34731
rect 14875 34728 14887 34731
rect 15010 34728 15016 34740
rect 14875 34700 15016 34728
rect 14875 34697 14887 34700
rect 14829 34691 14887 34697
rect 15010 34688 15016 34700
rect 15068 34688 15074 34740
rect 15289 34731 15347 34737
rect 15289 34697 15301 34731
rect 15335 34728 15347 34731
rect 15470 34728 15476 34740
rect 15335 34700 15476 34728
rect 15335 34697 15347 34700
rect 15289 34691 15347 34697
rect 15470 34688 15476 34700
rect 15528 34688 15534 34740
rect 17037 34731 17095 34737
rect 17037 34728 17049 34731
rect 15856 34700 17049 34728
rect 13630 34620 13636 34672
rect 13688 34660 13694 34672
rect 15194 34660 15200 34672
rect 13688 34632 15200 34660
rect 13688 34620 13694 34632
rect 15194 34620 15200 34632
rect 15252 34620 15258 34672
rect 1394 34552 1400 34604
rect 1452 34592 1458 34604
rect 1765 34595 1823 34601
rect 1765 34592 1777 34595
rect 1452 34564 1777 34592
rect 1452 34552 1458 34564
rect 1765 34561 1777 34564
rect 1811 34561 1823 34595
rect 1765 34555 1823 34561
rect 12897 34595 12955 34601
rect 12897 34561 12909 34595
rect 12943 34592 12955 34595
rect 12986 34592 12992 34604
rect 12943 34564 12992 34592
rect 12943 34561 12955 34564
rect 12897 34555 12955 34561
rect 12986 34552 12992 34564
rect 13044 34552 13050 34604
rect 13541 34595 13599 34601
rect 13541 34561 13553 34595
rect 13587 34561 13599 34595
rect 14182 34592 14188 34604
rect 14143 34564 14188 34592
rect 13541 34555 13599 34561
rect 13556 34524 13584 34555
rect 14182 34552 14188 34564
rect 14240 34552 14246 34604
rect 14550 34552 14556 34604
rect 14608 34592 14614 34604
rect 14645 34595 14703 34601
rect 14645 34592 14657 34595
rect 14608 34564 14657 34592
rect 14608 34552 14614 34564
rect 14645 34561 14657 34564
rect 14691 34561 14703 34595
rect 14645 34555 14703 34561
rect 14734 34552 14740 34604
rect 14792 34592 14798 34604
rect 14829 34595 14887 34601
rect 14829 34592 14841 34595
rect 14792 34564 14841 34592
rect 14792 34552 14798 34564
rect 14829 34561 14841 34564
rect 14875 34592 14887 34595
rect 15010 34592 15016 34604
rect 14875 34564 15016 34592
rect 14875 34561 14887 34564
rect 14829 34555 14887 34561
rect 15010 34552 15016 34564
rect 15068 34552 15074 34604
rect 15473 34595 15531 34601
rect 15473 34561 15485 34595
rect 15519 34592 15531 34595
rect 15746 34592 15752 34604
rect 15519 34564 15752 34592
rect 15519 34561 15531 34564
rect 15473 34555 15531 34561
rect 15746 34552 15752 34564
rect 15804 34552 15810 34604
rect 14458 34524 14464 34536
rect 13556 34496 14464 34524
rect 14458 34484 14464 34496
rect 14516 34484 14522 34536
rect 15856 34524 15884 34700
rect 17037 34697 17049 34700
rect 17083 34697 17095 34731
rect 20990 34728 20996 34740
rect 17037 34691 17095 34697
rect 17328 34700 20996 34728
rect 16482 34660 16488 34672
rect 15948 34632 16488 34660
rect 15948 34601 15976 34632
rect 16482 34620 16488 34632
rect 16540 34620 16546 34672
rect 16574 34620 16580 34672
rect 16632 34660 16638 34672
rect 16758 34660 16764 34672
rect 16632 34632 16764 34660
rect 16632 34620 16638 34632
rect 16758 34620 16764 34632
rect 16816 34620 16822 34672
rect 17328 34660 17356 34700
rect 20990 34688 20996 34700
rect 21048 34688 21054 34740
rect 23382 34688 23388 34740
rect 23440 34728 23446 34740
rect 23477 34731 23535 34737
rect 23477 34728 23489 34731
rect 23440 34700 23489 34728
rect 23440 34688 23446 34700
rect 23477 34697 23489 34700
rect 23523 34697 23535 34731
rect 23477 34691 23535 34697
rect 23842 34688 23848 34740
rect 23900 34728 23906 34740
rect 26142 34728 26148 34740
rect 23900 34700 25820 34728
rect 26103 34700 26148 34728
rect 23900 34688 23906 34700
rect 18046 34660 18052 34672
rect 16951 34632 17356 34660
rect 17512 34632 18052 34660
rect 15933 34595 15991 34601
rect 15933 34561 15945 34595
rect 15979 34561 15991 34595
rect 15933 34555 15991 34561
rect 16117 34595 16175 34601
rect 16117 34561 16129 34595
rect 16163 34592 16175 34595
rect 16390 34592 16396 34604
rect 16163 34564 16396 34592
rect 16163 34561 16175 34564
rect 16117 34555 16175 34561
rect 16390 34552 16396 34564
rect 16448 34552 16454 34604
rect 16853 34595 16911 34601
rect 16500 34564 16804 34592
rect 14568 34496 15884 34524
rect 16025 34527 16083 34533
rect 2406 34456 2412 34468
rect 2367 34428 2412 34456
rect 2406 34416 2412 34428
rect 2464 34416 2470 34468
rect 12250 34456 12256 34468
rect 12211 34428 12256 34456
rect 12250 34416 12256 34428
rect 12308 34416 12314 34468
rect 13998 34456 14004 34468
rect 13959 34428 14004 34456
rect 13998 34416 14004 34428
rect 14056 34416 14062 34468
rect 14568 34456 14596 34496
rect 16025 34493 16037 34527
rect 16071 34524 16083 34527
rect 16500 34524 16528 34564
rect 16071 34496 16528 34524
rect 16071 34493 16083 34496
rect 16025 34487 16083 34493
rect 16574 34484 16580 34536
rect 16632 34524 16638 34536
rect 16669 34527 16727 34533
rect 16669 34524 16681 34527
rect 16632 34496 16681 34524
rect 16632 34484 16638 34496
rect 16669 34493 16681 34496
rect 16715 34493 16727 34527
rect 16776 34524 16804 34564
rect 16853 34561 16865 34595
rect 16899 34590 16911 34595
rect 16951 34590 16979 34632
rect 16899 34562 16979 34590
rect 16899 34561 16911 34562
rect 16853 34555 16911 34561
rect 17034 34552 17040 34604
rect 17092 34592 17098 34604
rect 17512 34601 17540 34632
rect 18046 34620 18052 34632
rect 18104 34620 18110 34672
rect 18230 34620 18236 34672
rect 18288 34660 18294 34672
rect 18785 34663 18843 34669
rect 18785 34660 18797 34663
rect 18288 34632 18797 34660
rect 18288 34620 18294 34632
rect 18785 34629 18797 34632
rect 18831 34629 18843 34663
rect 18785 34623 18843 34629
rect 18966 34620 18972 34672
rect 19024 34660 19030 34672
rect 19024 34632 21036 34660
rect 19024 34620 19030 34632
rect 17497 34595 17555 34601
rect 17497 34592 17509 34595
rect 17092 34564 17509 34592
rect 17092 34552 17098 34564
rect 17497 34561 17509 34564
rect 17543 34561 17555 34595
rect 17497 34555 17555 34561
rect 17586 34552 17592 34604
rect 17644 34592 17650 34604
rect 17773 34595 17831 34601
rect 17773 34592 17785 34595
rect 17644 34564 17785 34592
rect 17644 34552 17650 34564
rect 17773 34561 17785 34564
rect 17819 34561 17831 34595
rect 18417 34595 18475 34601
rect 18417 34592 18429 34595
rect 17773 34555 17831 34561
rect 17952 34564 18429 34592
rect 17678 34524 17684 34536
rect 16776 34496 17540 34524
rect 17639 34496 17684 34524
rect 16669 34487 16727 34493
rect 14108 34428 14596 34456
rect 11882 34348 11888 34400
rect 11940 34388 11946 34400
rect 14108 34388 14136 34428
rect 14918 34416 14924 34468
rect 14976 34456 14982 34468
rect 15194 34456 15200 34468
rect 14976 34428 15200 34456
rect 14976 34416 14982 34428
rect 15194 34416 15200 34428
rect 15252 34416 15258 34468
rect 15286 34416 15292 34468
rect 15344 34456 15350 34468
rect 16298 34456 16304 34468
rect 15344 34428 16304 34456
rect 15344 34416 15350 34428
rect 16298 34416 16304 34428
rect 16356 34416 16362 34468
rect 16482 34416 16488 34468
rect 16540 34456 16546 34468
rect 17218 34456 17224 34468
rect 16540 34428 17224 34456
rect 16540 34416 16546 34428
rect 17218 34416 17224 34428
rect 17276 34416 17282 34468
rect 17512 34456 17540 34496
rect 17678 34484 17684 34496
rect 17736 34524 17742 34536
rect 17952 34524 17980 34564
rect 18417 34561 18429 34564
rect 18463 34561 18475 34595
rect 18417 34555 18475 34561
rect 18601 34595 18659 34601
rect 18601 34561 18613 34595
rect 18647 34592 18659 34595
rect 18690 34592 18696 34604
rect 18647 34564 18696 34592
rect 18647 34561 18659 34564
rect 18601 34555 18659 34561
rect 18690 34552 18696 34564
rect 18748 34552 18754 34604
rect 19242 34552 19248 34604
rect 19300 34592 19306 34604
rect 19613 34595 19671 34601
rect 19613 34592 19625 34595
rect 19300 34564 19625 34592
rect 19300 34552 19306 34564
rect 19613 34561 19625 34564
rect 19659 34561 19671 34595
rect 19613 34555 19671 34561
rect 19702 34552 19708 34604
rect 19760 34592 19766 34604
rect 19886 34601 19892 34604
rect 19880 34592 19892 34601
rect 19760 34564 19892 34592
rect 19760 34552 19766 34564
rect 19880 34555 19892 34564
rect 19944 34592 19950 34604
rect 19944 34564 20028 34592
rect 19886 34552 19892 34555
rect 19944 34552 19950 34564
rect 18782 34524 18788 34536
rect 17736 34496 17980 34524
rect 18156 34496 18788 34524
rect 17736 34484 17742 34496
rect 18156 34456 18184 34496
rect 18782 34484 18788 34496
rect 18840 34484 18846 34536
rect 18874 34484 18880 34536
rect 18932 34524 18938 34536
rect 19518 34524 19524 34536
rect 18932 34496 19524 34524
rect 18932 34484 18938 34496
rect 19518 34484 19524 34496
rect 19576 34484 19582 34536
rect 21008 34468 21036 34632
rect 21082 34620 21088 34672
rect 21140 34660 21146 34672
rect 22342 34663 22400 34669
rect 22342 34660 22354 34663
rect 21140 34632 22354 34660
rect 21140 34620 21146 34632
rect 22342 34629 22354 34632
rect 22388 34629 22400 34663
rect 22342 34623 22400 34629
rect 24204 34663 24262 34669
rect 24204 34629 24216 34663
rect 24250 34660 24262 34663
rect 24394 34660 24400 34672
rect 24250 34632 24400 34660
rect 24250 34629 24262 34632
rect 24204 34623 24262 34629
rect 24394 34620 24400 34632
rect 24452 34620 24458 34672
rect 25792 34669 25820 34700
rect 26142 34688 26148 34700
rect 26200 34688 26206 34740
rect 31570 34728 31576 34740
rect 26252 34700 31576 34728
rect 25777 34663 25835 34669
rect 25777 34629 25789 34663
rect 25823 34629 25835 34663
rect 26252 34660 26280 34700
rect 31570 34688 31576 34700
rect 31628 34688 31634 34740
rect 32122 34728 32128 34740
rect 32083 34700 32128 34728
rect 32122 34688 32128 34700
rect 32180 34688 32186 34740
rect 32490 34688 32496 34740
rect 32548 34728 32554 34740
rect 33597 34731 33655 34737
rect 33597 34728 33609 34731
rect 32548 34700 33609 34728
rect 32548 34688 32554 34700
rect 33597 34697 33609 34700
rect 33643 34697 33655 34731
rect 33597 34691 33655 34697
rect 25777 34623 25835 34629
rect 25884 34632 26280 34660
rect 21266 34552 21272 34604
rect 21324 34592 21330 34604
rect 22097 34595 22155 34601
rect 22097 34592 22109 34595
rect 21324 34564 22109 34592
rect 21324 34552 21330 34564
rect 22097 34561 22109 34564
rect 22143 34561 22155 34595
rect 22097 34555 22155 34561
rect 22646 34552 22652 34604
rect 22704 34592 22710 34604
rect 22704 34564 24992 34592
rect 22704 34552 22710 34564
rect 23750 34484 23756 34536
rect 23808 34524 23814 34536
rect 23937 34527 23995 34533
rect 23937 34524 23949 34527
rect 23808 34496 23949 34524
rect 23808 34484 23814 34496
rect 23937 34493 23949 34496
rect 23983 34493 23995 34527
rect 24964 34524 24992 34564
rect 25314 34552 25320 34604
rect 25372 34592 25378 34604
rect 25884 34592 25912 34632
rect 27338 34620 27344 34672
rect 27396 34660 27402 34672
rect 28166 34660 28172 34672
rect 27396 34632 28172 34660
rect 27396 34620 27402 34632
rect 28166 34620 28172 34632
rect 28224 34620 28230 34672
rect 28997 34663 29055 34669
rect 28997 34629 29009 34663
rect 29043 34660 29055 34663
rect 29362 34660 29368 34672
rect 29043 34632 29368 34660
rect 29043 34629 29055 34632
rect 28997 34623 29055 34629
rect 29362 34620 29368 34632
rect 29420 34620 29426 34672
rect 29454 34620 29460 34672
rect 29512 34660 29518 34672
rect 30466 34660 30472 34672
rect 29512 34632 30472 34660
rect 29512 34620 29518 34632
rect 25372 34564 25912 34592
rect 25372 34552 25378 34564
rect 25958 34552 25964 34604
rect 26016 34592 26022 34604
rect 27065 34595 27123 34601
rect 26016 34564 26061 34592
rect 26016 34552 26022 34564
rect 27065 34561 27077 34595
rect 27111 34561 27123 34595
rect 27065 34555 27123 34561
rect 27080 34524 27108 34555
rect 27614 34552 27620 34604
rect 27672 34592 27678 34604
rect 27890 34592 27896 34604
rect 27672 34564 27896 34592
rect 27672 34552 27678 34564
rect 27890 34552 27896 34564
rect 27948 34552 27954 34604
rect 28810 34592 28816 34604
rect 28771 34564 28816 34592
rect 28810 34552 28816 34564
rect 28868 34552 28874 34604
rect 28902 34552 28908 34604
rect 28960 34592 28966 34604
rect 29656 34601 29684 34632
rect 30466 34620 30472 34632
rect 30524 34620 30530 34672
rect 32674 34660 32680 34672
rect 32600 34632 32680 34660
rect 29089 34595 29147 34601
rect 29089 34592 29101 34595
rect 28960 34564 29101 34592
rect 28960 34552 28966 34564
rect 29089 34561 29101 34564
rect 29135 34561 29147 34595
rect 29089 34555 29147 34561
rect 29641 34595 29699 34601
rect 29641 34561 29653 34595
rect 29687 34561 29699 34595
rect 29641 34555 29699 34561
rect 29908 34595 29966 34601
rect 29908 34561 29920 34595
rect 29954 34592 29966 34595
rect 30742 34592 30748 34604
rect 29954 34564 30748 34592
rect 29954 34561 29966 34564
rect 29908 34555 29966 34561
rect 30742 34552 30748 34564
rect 30800 34552 30806 34604
rect 31570 34552 31576 34604
rect 31628 34592 31634 34604
rect 32306 34592 32312 34604
rect 31628 34564 32312 34592
rect 31628 34552 31634 34564
rect 32306 34552 32312 34564
rect 32364 34601 32370 34604
rect 32364 34595 32413 34601
rect 32364 34561 32367 34595
rect 32401 34561 32413 34595
rect 32490 34592 32496 34604
rect 32451 34564 32496 34592
rect 32364 34555 32413 34561
rect 32364 34552 32370 34555
rect 32490 34552 32496 34564
rect 32548 34552 32554 34604
rect 32600 34601 32628 34632
rect 32674 34620 32680 34632
rect 32732 34620 32738 34672
rect 33226 34660 33232 34672
rect 33187 34632 33232 34660
rect 33226 34620 33232 34632
rect 33284 34620 33290 34672
rect 32585 34595 32643 34601
rect 32585 34561 32597 34595
rect 32631 34561 32643 34595
rect 32585 34555 32643 34561
rect 32766 34552 32772 34604
rect 32824 34592 32830 34604
rect 33410 34592 33416 34604
rect 32824 34564 32869 34592
rect 33371 34564 33416 34592
rect 32824 34552 32830 34564
rect 33410 34552 33416 34564
rect 33468 34552 33474 34604
rect 33686 34592 33692 34604
rect 33647 34564 33692 34592
rect 33686 34552 33692 34564
rect 33744 34552 33750 34604
rect 24964 34496 27108 34524
rect 23937 34487 23995 34493
rect 27430 34484 27436 34536
rect 27488 34524 27494 34536
rect 27709 34527 27767 34533
rect 27709 34524 27721 34527
rect 27488 34496 27721 34524
rect 27488 34484 27494 34496
rect 27709 34493 27721 34496
rect 27755 34493 27767 34527
rect 27709 34487 27767 34493
rect 28169 34527 28227 34533
rect 28169 34493 28181 34527
rect 28215 34524 28227 34527
rect 28215 34496 29040 34524
rect 28215 34493 28227 34496
rect 28169 34487 28227 34493
rect 29012 34468 29040 34496
rect 17512 34428 17632 34456
rect 11940 34360 14136 34388
rect 11940 34348 11946 34360
rect 14182 34348 14188 34400
rect 14240 34388 14246 34400
rect 17034 34388 17040 34400
rect 14240 34360 17040 34388
rect 14240 34348 14246 34360
rect 17034 34348 17040 34360
rect 17092 34348 17098 34400
rect 17402 34348 17408 34400
rect 17460 34388 17466 34400
rect 17497 34391 17555 34397
rect 17497 34388 17509 34391
rect 17460 34360 17509 34388
rect 17460 34348 17466 34360
rect 17497 34357 17509 34360
rect 17543 34357 17555 34391
rect 17604 34388 17632 34428
rect 17880 34428 18184 34456
rect 17880 34388 17908 34428
rect 18230 34416 18236 34468
rect 18288 34456 18294 34468
rect 20990 34456 20996 34468
rect 18288 34428 19555 34456
rect 20903 34428 20996 34456
rect 18288 34416 18294 34428
rect 17604 34360 17908 34388
rect 17957 34391 18015 34397
rect 17497 34351 17555 34357
rect 17957 34357 17969 34391
rect 18003 34388 18015 34391
rect 19426 34388 19432 34400
rect 18003 34360 19432 34388
rect 18003 34357 18015 34360
rect 17957 34351 18015 34357
rect 19426 34348 19432 34360
rect 19484 34348 19490 34400
rect 19527 34388 19555 34428
rect 20990 34416 20996 34428
rect 21048 34416 21054 34468
rect 22094 34456 22100 34468
rect 21100 34428 22100 34456
rect 21100 34388 21128 34428
rect 22094 34416 22100 34428
rect 22152 34416 22158 34468
rect 23566 34456 23572 34468
rect 23032 34428 23572 34456
rect 19527 34360 21128 34388
rect 21358 34348 21364 34400
rect 21416 34388 21422 34400
rect 23032 34388 23060 34428
rect 23566 34416 23572 34428
rect 23624 34416 23630 34468
rect 25148 34428 25452 34456
rect 21416 34360 23060 34388
rect 21416 34348 21422 34360
rect 23106 34348 23112 34400
rect 23164 34388 23170 34400
rect 25148 34388 25176 34428
rect 25314 34388 25320 34400
rect 23164 34360 25176 34388
rect 25275 34360 25320 34388
rect 23164 34348 23170 34360
rect 25314 34348 25320 34360
rect 25372 34348 25378 34400
rect 25424 34388 25452 34428
rect 25590 34416 25596 34468
rect 25648 34456 25654 34468
rect 27249 34459 27307 34465
rect 27249 34456 27261 34459
rect 25648 34428 27261 34456
rect 25648 34416 25654 34428
rect 27249 34425 27261 34428
rect 27295 34425 27307 34459
rect 27249 34419 27307 34425
rect 27522 34416 27528 34468
rect 27580 34456 27586 34468
rect 27985 34459 28043 34465
rect 27985 34456 27997 34459
rect 27580 34428 27997 34456
rect 27580 34416 27586 34428
rect 27985 34425 27997 34428
rect 28031 34425 28043 34459
rect 27985 34419 28043 34425
rect 28994 34416 29000 34468
rect 29052 34416 29058 34468
rect 28534 34388 28540 34400
rect 25424 34360 28540 34388
rect 28534 34348 28540 34360
rect 28592 34348 28598 34400
rect 28629 34391 28687 34397
rect 28629 34357 28641 34391
rect 28675 34388 28687 34391
rect 30282 34388 30288 34400
rect 28675 34360 30288 34388
rect 28675 34357 28687 34360
rect 28629 34351 28687 34357
rect 30282 34348 30288 34360
rect 30340 34348 30346 34400
rect 31018 34388 31024 34400
rect 30979 34360 31024 34388
rect 31018 34348 31024 34360
rect 31076 34348 31082 34400
rect 1104 34298 34868 34320
rect 1104 34246 6582 34298
rect 6634 34246 6646 34298
rect 6698 34246 6710 34298
rect 6762 34246 6774 34298
rect 6826 34246 6838 34298
rect 6890 34246 17846 34298
rect 17898 34246 17910 34298
rect 17962 34246 17974 34298
rect 18026 34246 18038 34298
rect 18090 34246 18102 34298
rect 18154 34246 29110 34298
rect 29162 34246 29174 34298
rect 29226 34246 29238 34298
rect 29290 34246 29302 34298
rect 29354 34246 29366 34298
rect 29418 34246 34868 34298
rect 1104 34224 34868 34246
rect 12894 34184 12900 34196
rect 12855 34156 12900 34184
rect 12894 34144 12900 34156
rect 12952 34144 12958 34196
rect 13078 34144 13084 34196
rect 13136 34184 13142 34196
rect 15746 34184 15752 34196
rect 13136 34156 15752 34184
rect 13136 34144 13142 34156
rect 15746 34144 15752 34156
rect 15804 34144 15810 34196
rect 15930 34144 15936 34196
rect 15988 34184 15994 34196
rect 16206 34184 16212 34196
rect 15988 34156 16212 34184
rect 15988 34144 15994 34156
rect 16206 34144 16212 34156
rect 16264 34144 16270 34196
rect 16298 34144 16304 34196
rect 16356 34184 16362 34196
rect 16574 34184 16580 34196
rect 16356 34156 16580 34184
rect 16356 34144 16362 34156
rect 16574 34144 16580 34156
rect 16632 34144 16638 34196
rect 16691 34156 20199 34184
rect 2498 34076 2504 34128
rect 2556 34116 2562 34128
rect 13357 34119 13415 34125
rect 2556 34088 6914 34116
rect 2556 34076 2562 34088
rect 2774 34048 2780 34060
rect 2735 34020 2780 34048
rect 2774 34008 2780 34020
rect 2832 34008 2838 34060
rect 6886 34048 6914 34088
rect 13357 34085 13369 34119
rect 13403 34085 13415 34119
rect 13357 34079 13415 34085
rect 13262 34048 13268 34060
rect 6886 34020 13268 34048
rect 13262 34008 13268 34020
rect 13320 34008 13326 34060
rect 13372 34048 13400 34079
rect 13446 34076 13452 34128
rect 13504 34116 13510 34128
rect 13504 34088 15025 34116
rect 13504 34076 13510 34088
rect 14550 34048 14556 34060
rect 13372 34020 14556 34048
rect 14550 34008 14556 34020
rect 14608 34008 14614 34060
rect 14997 34048 15025 34088
rect 15470 34076 15476 34128
rect 15528 34116 15534 34128
rect 16691 34116 16719 34156
rect 15528 34088 16719 34116
rect 18049 34119 18107 34125
rect 15528 34076 15534 34088
rect 18049 34085 18061 34119
rect 18095 34116 18107 34119
rect 18506 34116 18512 34128
rect 18095 34088 18512 34116
rect 18095 34085 18107 34088
rect 18049 34079 18107 34085
rect 18506 34076 18512 34088
rect 18564 34076 18570 34128
rect 18601 34119 18659 34125
rect 18601 34085 18613 34119
rect 18647 34116 18659 34119
rect 18966 34116 18972 34128
rect 18647 34088 18972 34116
rect 18647 34085 18659 34088
rect 18601 34079 18659 34085
rect 18966 34076 18972 34088
rect 19024 34076 19030 34128
rect 20171 34116 20199 34156
rect 20438 34144 20444 34196
rect 20496 34184 20502 34196
rect 20625 34187 20683 34193
rect 20625 34184 20637 34187
rect 20496 34156 20637 34184
rect 20496 34144 20502 34156
rect 20625 34153 20637 34156
rect 20671 34153 20683 34187
rect 20625 34147 20683 34153
rect 20714 34144 20720 34196
rect 20772 34184 20778 34196
rect 23382 34184 23388 34196
rect 20772 34156 23388 34184
rect 20772 34144 20778 34156
rect 23382 34144 23388 34156
rect 23440 34144 23446 34196
rect 23569 34187 23627 34193
rect 23569 34153 23581 34187
rect 23615 34184 23627 34187
rect 24670 34184 24676 34196
rect 23615 34156 24676 34184
rect 23615 34153 23627 34156
rect 23569 34147 23627 34153
rect 24670 34144 24676 34156
rect 24728 34144 24734 34196
rect 24762 34144 24768 34196
rect 24820 34184 24826 34196
rect 28626 34184 28632 34196
rect 24820 34156 28632 34184
rect 24820 34144 24826 34156
rect 28626 34144 28632 34156
rect 28684 34144 28690 34196
rect 30742 34184 30748 34196
rect 30703 34156 30748 34184
rect 30742 34144 30748 34156
rect 30800 34144 30806 34196
rect 31386 34144 31392 34196
rect 31444 34184 31450 34196
rect 32766 34184 32772 34196
rect 31444 34156 32772 34184
rect 31444 34144 31450 34156
rect 32766 34144 32772 34156
rect 32824 34144 32830 34196
rect 24857 34119 24915 34125
rect 24857 34116 24869 34119
rect 20171 34088 24869 34116
rect 24857 34085 24869 34088
rect 24903 34085 24915 34119
rect 31202 34116 31208 34128
rect 24857 34079 24915 34085
rect 30760 34088 31208 34116
rect 30760 34060 30788 34088
rect 31202 34076 31208 34088
rect 31260 34076 31266 34128
rect 14997 34020 16068 34048
rect 1394 33980 1400 33992
rect 1355 33952 1400 33980
rect 1394 33940 1400 33952
rect 1452 33940 1458 33992
rect 12253 33983 12311 33989
rect 12253 33949 12265 33983
rect 12299 33949 12311 33983
rect 12253 33943 12311 33949
rect 13541 33983 13599 33989
rect 13541 33949 13553 33983
rect 13587 33980 13599 33983
rect 13998 33980 14004 33992
rect 13587 33952 14004 33980
rect 13587 33949 13599 33952
rect 13541 33943 13599 33949
rect 1581 33915 1639 33921
rect 1581 33881 1593 33915
rect 1627 33912 1639 33915
rect 2590 33912 2596 33924
rect 1627 33884 2596 33912
rect 1627 33881 1639 33884
rect 1581 33875 1639 33881
rect 2590 33872 2596 33884
rect 2648 33872 2654 33924
rect 12268 33912 12296 33943
rect 13998 33940 14004 33952
rect 14056 33940 14062 33992
rect 14093 33983 14151 33989
rect 14093 33949 14105 33983
rect 14139 33980 14151 33983
rect 14182 33980 14188 33992
rect 14139 33952 14188 33980
rect 14139 33949 14151 33952
rect 14093 33943 14151 33949
rect 14182 33940 14188 33952
rect 14240 33940 14246 33992
rect 14277 33983 14335 33989
rect 14277 33949 14289 33983
rect 14323 33980 14335 33983
rect 14642 33980 14648 33992
rect 14323 33952 14648 33980
rect 14323 33949 14335 33952
rect 14277 33943 14335 33949
rect 14642 33940 14648 33952
rect 14700 33940 14706 33992
rect 14921 33983 14979 33989
rect 14921 33949 14933 33983
rect 14967 33980 14979 33983
rect 15470 33980 15476 33992
rect 14967 33952 15476 33980
rect 14967 33949 14979 33952
rect 14921 33943 14979 33949
rect 15470 33940 15476 33952
rect 15528 33940 15534 33992
rect 15565 33983 15623 33989
rect 15565 33949 15577 33983
rect 15611 33980 15623 33983
rect 15930 33980 15936 33992
rect 15611 33952 15936 33980
rect 15611 33949 15623 33952
rect 15565 33943 15623 33949
rect 15930 33940 15936 33952
rect 15988 33940 15994 33992
rect 16040 33989 16068 34020
rect 16206 34008 16212 34060
rect 16264 34048 16270 34060
rect 16264 34020 16574 34048
rect 16264 34008 16270 34020
rect 16025 33983 16083 33989
rect 16025 33949 16037 33983
rect 16071 33949 16083 33983
rect 16298 33980 16304 33992
rect 16025 33943 16083 33949
rect 16132 33952 16304 33980
rect 13262 33912 13268 33924
rect 12268 33884 13268 33912
rect 13262 33872 13268 33884
rect 13320 33872 13326 33924
rect 16132 33921 16160 33952
rect 16298 33940 16304 33952
rect 16356 33940 16362 33992
rect 16546 33980 16574 34020
rect 16666 34008 16672 34060
rect 16724 34048 16730 34060
rect 18690 34048 18696 34060
rect 16724 34020 16769 34048
rect 17696 34020 18696 34048
rect 16724 34008 16730 34020
rect 17696 33980 17724 34020
rect 18690 34008 18696 34020
rect 18748 34008 18754 34060
rect 18782 34008 18788 34060
rect 18840 34048 18846 34060
rect 18840 34020 19380 34048
rect 18840 34008 18846 34020
rect 16546 33952 17724 33980
rect 18509 33983 18567 33989
rect 18509 33949 18521 33983
rect 18555 33980 18567 33983
rect 18874 33980 18880 33992
rect 18555 33952 18880 33980
rect 18555 33949 18567 33952
rect 18509 33943 18567 33949
rect 18874 33940 18880 33952
rect 18932 33940 18938 33992
rect 19242 33980 19248 33992
rect 19203 33952 19248 33980
rect 19242 33940 19248 33952
rect 19300 33940 19306 33992
rect 19352 33980 19380 34020
rect 20254 34008 20260 34060
rect 20312 34048 20318 34060
rect 23106 34048 23112 34060
rect 20312 34020 23112 34048
rect 20312 34008 20318 34020
rect 23106 34008 23112 34020
rect 23164 34008 23170 34060
rect 23566 34008 23572 34060
rect 23624 34048 23630 34060
rect 23624 34020 24808 34048
rect 23624 34008 23630 34020
rect 21634 33980 21640 33992
rect 19352 33952 21640 33980
rect 21634 33940 21640 33952
rect 21692 33940 21698 33992
rect 21821 33983 21879 33989
rect 21821 33949 21833 33983
rect 21867 33980 21879 33983
rect 21910 33980 21916 33992
rect 21867 33952 21916 33980
rect 21867 33949 21879 33952
rect 21821 33943 21879 33949
rect 21910 33940 21916 33952
rect 21968 33940 21974 33992
rect 22097 33983 22155 33989
rect 22097 33949 22109 33983
rect 22143 33980 22155 33983
rect 22278 33980 22284 33992
rect 22143 33952 22284 33980
rect 22143 33949 22155 33952
rect 22097 33943 22155 33949
rect 22278 33940 22284 33952
rect 22336 33940 22342 33992
rect 22922 33940 22928 33992
rect 22980 33980 22986 33992
rect 23017 33983 23075 33989
rect 23017 33980 23029 33983
rect 22980 33952 23029 33980
rect 22980 33940 22986 33952
rect 23017 33949 23029 33952
rect 23063 33949 23075 33983
rect 23017 33943 23075 33949
rect 23293 33983 23351 33989
rect 23293 33949 23305 33983
rect 23339 33980 23351 33983
rect 23474 33980 23480 33992
rect 23339 33952 23480 33980
rect 23339 33949 23351 33952
rect 23293 33943 23351 33949
rect 23474 33940 23480 33952
rect 23532 33940 23538 33992
rect 23750 33940 23756 33992
rect 23808 33980 23814 33992
rect 24118 33980 24124 33992
rect 23808 33952 24124 33980
rect 23808 33940 23814 33952
rect 24118 33940 24124 33952
rect 24176 33940 24182 33992
rect 24578 33980 24584 33992
rect 24539 33952 24584 33980
rect 24578 33940 24584 33952
rect 24636 33940 24642 33992
rect 24673 33983 24731 33989
rect 24673 33949 24685 33983
rect 24719 33949 24731 33983
rect 24673 33943 24731 33949
rect 16117 33915 16175 33921
rect 14936 33884 15884 33912
rect 14277 33847 14335 33853
rect 14277 33813 14289 33847
rect 14323 33844 14335 33847
rect 14458 33844 14464 33856
rect 14323 33816 14464 33844
rect 14323 33813 14335 33816
rect 14277 33807 14335 33813
rect 14458 33804 14464 33816
rect 14516 33804 14522 33856
rect 14737 33847 14795 33853
rect 14737 33813 14749 33847
rect 14783 33844 14795 33847
rect 14936 33844 14964 33884
rect 14783 33816 14964 33844
rect 15381 33847 15439 33853
rect 14783 33813 14795 33816
rect 14737 33807 14795 33813
rect 15381 33813 15393 33847
rect 15427 33844 15439 33847
rect 15746 33844 15752 33856
rect 15427 33816 15752 33844
rect 15427 33813 15439 33816
rect 15381 33807 15439 33813
rect 15746 33804 15752 33816
rect 15804 33804 15810 33856
rect 15856 33844 15884 33884
rect 16117 33881 16129 33915
rect 16163 33881 16175 33915
rect 16117 33875 16175 33881
rect 16206 33872 16212 33924
rect 16264 33912 16270 33924
rect 16914 33915 16972 33921
rect 16914 33912 16926 33915
rect 16264 33884 16926 33912
rect 16264 33872 16270 33884
rect 16914 33881 16926 33884
rect 16960 33881 16972 33915
rect 16914 33875 16972 33881
rect 17236 33884 19295 33912
rect 17236 33844 17264 33884
rect 15856 33816 17264 33844
rect 17310 33804 17316 33856
rect 17368 33844 17374 33856
rect 17954 33844 17960 33856
rect 17368 33816 17960 33844
rect 17368 33804 17374 33816
rect 17954 33804 17960 33816
rect 18012 33804 18018 33856
rect 18046 33804 18052 33856
rect 18104 33844 18110 33856
rect 19150 33844 19156 33856
rect 18104 33816 19156 33844
rect 18104 33804 18110 33816
rect 19150 33804 19156 33816
rect 19208 33804 19214 33856
rect 19267 33844 19295 33884
rect 19334 33872 19340 33924
rect 19392 33912 19398 33924
rect 19490 33915 19548 33921
rect 19490 33912 19502 33915
rect 19392 33884 19502 33912
rect 19392 33872 19398 33884
rect 19490 33881 19502 33884
rect 19536 33881 19548 33915
rect 19490 33875 19548 33881
rect 20622 33872 20628 33924
rect 20680 33912 20686 33924
rect 24688 33912 24716 33943
rect 20680 33884 24716 33912
rect 24780 33912 24808 34020
rect 25130 34008 25136 34060
rect 25188 34048 25194 34060
rect 25317 34051 25375 34057
rect 25317 34048 25329 34051
rect 25188 34020 25329 34048
rect 25188 34008 25194 34020
rect 25317 34017 25329 34020
rect 25363 34017 25375 34051
rect 30742 34048 30748 34060
rect 25317 34011 25375 34017
rect 28184 34020 30748 34048
rect 24854 33940 24860 33992
rect 24912 33980 24918 33992
rect 25573 33983 25631 33989
rect 25573 33980 25585 33983
rect 24912 33952 25585 33980
rect 24912 33940 24918 33952
rect 25573 33949 25585 33952
rect 25619 33949 25631 33983
rect 25573 33943 25631 33949
rect 26510 33940 26516 33992
rect 26568 33980 26574 33992
rect 27157 33983 27215 33989
rect 27157 33980 27169 33983
rect 26568 33952 27169 33980
rect 26568 33940 26574 33952
rect 27157 33949 27169 33952
rect 27203 33949 27215 33983
rect 28184 33980 28212 34020
rect 30742 34008 30748 34020
rect 30800 34008 30806 34060
rect 32490 34048 32496 34060
rect 31128 34020 32496 34048
rect 27157 33943 27215 33949
rect 27244 33952 28212 33980
rect 27244 33912 27272 33952
rect 28534 33940 28540 33992
rect 28592 33940 28598 33992
rect 29638 33980 29644 33992
rect 29599 33952 29644 33980
rect 29638 33940 29644 33952
rect 29696 33940 29702 33992
rect 30098 33980 30104 33992
rect 30059 33952 30104 33980
rect 30098 33940 30104 33952
rect 30156 33940 30162 33992
rect 31018 33980 31024 33992
rect 30979 33952 31024 33980
rect 31018 33940 31024 33952
rect 31076 33940 31082 33992
rect 31128 33989 31156 34020
rect 32490 34008 32496 34020
rect 32548 34008 32554 34060
rect 34146 34048 34152 34060
rect 34107 34020 34152 34048
rect 34146 34008 34152 34020
rect 34204 34008 34210 34060
rect 31113 33983 31171 33989
rect 31113 33949 31125 33983
rect 31159 33949 31171 33983
rect 31113 33943 31171 33949
rect 24780 33884 27272 33912
rect 20680 33872 20686 33884
rect 27338 33872 27344 33924
rect 27396 33921 27402 33924
rect 27396 33915 27460 33921
rect 27396 33881 27414 33915
rect 27448 33881 27460 33915
rect 28442 33912 28448 33924
rect 27396 33875 27460 33881
rect 27724 33884 28448 33912
rect 27396 33872 27402 33875
rect 20530 33844 20536 33856
rect 19267 33816 20536 33844
rect 20530 33804 20536 33816
rect 20588 33804 20594 33856
rect 21450 33804 21456 33856
rect 21508 33844 21514 33856
rect 21637 33847 21695 33853
rect 21637 33844 21649 33847
rect 21508 33816 21649 33844
rect 21508 33804 21514 33816
rect 21637 33813 21649 33816
rect 21683 33813 21695 33847
rect 22002 33844 22008 33856
rect 21963 33816 22008 33844
rect 21637 33807 21695 33813
rect 22002 33804 22008 33816
rect 22060 33804 22066 33856
rect 22738 33804 22744 33856
rect 22796 33844 22802 33856
rect 23201 33847 23259 33853
rect 23201 33844 23213 33847
rect 22796 33816 23213 33844
rect 22796 33804 22802 33816
rect 23201 33813 23213 33816
rect 23247 33813 23259 33847
rect 23201 33807 23259 33813
rect 23290 33804 23296 33856
rect 23348 33844 23354 33856
rect 23385 33847 23443 33853
rect 23385 33844 23397 33847
rect 23348 33816 23397 33844
rect 23348 33804 23354 33816
rect 23385 33813 23397 33816
rect 23431 33813 23443 33847
rect 23385 33807 23443 33813
rect 23842 33804 23848 33856
rect 23900 33844 23906 33856
rect 26050 33844 26056 33856
rect 23900 33816 26056 33844
rect 23900 33804 23906 33816
rect 26050 33804 26056 33816
rect 26108 33844 26114 33856
rect 26697 33847 26755 33853
rect 26697 33844 26709 33847
rect 26108 33816 26709 33844
rect 26108 33804 26114 33816
rect 26697 33813 26709 33816
rect 26743 33813 26755 33847
rect 26697 33807 26755 33813
rect 27246 33804 27252 33856
rect 27304 33844 27310 33856
rect 27724 33844 27752 33884
rect 28442 33872 28448 33884
rect 28500 33872 28506 33924
rect 28552 33912 28580 33940
rect 28552 33884 28994 33912
rect 27304 33816 27752 33844
rect 27304 33804 27310 33816
rect 27798 33804 27804 33856
rect 27856 33844 27862 33856
rect 28537 33847 28595 33853
rect 28537 33844 28549 33847
rect 27856 33816 28549 33844
rect 27856 33804 27862 33816
rect 28537 33813 28549 33816
rect 28583 33813 28595 33847
rect 28966 33844 28994 33884
rect 30466 33872 30472 33924
rect 30524 33912 30530 33924
rect 31128 33912 31156 33943
rect 31202 33940 31208 33992
rect 31260 33980 31266 33992
rect 31260 33952 31305 33980
rect 31260 33940 31266 33952
rect 31386 33940 31392 33992
rect 31444 33980 31450 33992
rect 32309 33983 32367 33989
rect 31444 33952 31489 33980
rect 31444 33940 31450 33952
rect 32309 33949 32321 33983
rect 32355 33949 32367 33983
rect 32309 33943 32367 33949
rect 30524 33884 31156 33912
rect 30524 33872 30530 33884
rect 29638 33844 29644 33856
rect 28966 33816 29644 33844
rect 28537 33807 28595 33813
rect 29638 33804 29644 33816
rect 29696 33804 29702 33856
rect 32324 33844 32352 33943
rect 32490 33912 32496 33924
rect 32451 33884 32496 33912
rect 32490 33872 32496 33884
rect 32548 33872 32554 33924
rect 33226 33844 33232 33856
rect 32324 33816 33232 33844
rect 33226 33804 33232 33816
rect 33284 33804 33290 33856
rect 1104 33754 34868 33776
rect 1104 33702 12214 33754
rect 12266 33702 12278 33754
rect 12330 33702 12342 33754
rect 12394 33702 12406 33754
rect 12458 33702 12470 33754
rect 12522 33702 23478 33754
rect 23530 33702 23542 33754
rect 23594 33702 23606 33754
rect 23658 33702 23670 33754
rect 23722 33702 23734 33754
rect 23786 33702 34868 33754
rect 1104 33680 34868 33702
rect 2590 33640 2596 33652
rect 2551 33612 2596 33640
rect 2590 33600 2596 33612
rect 2648 33600 2654 33652
rect 12069 33643 12127 33649
rect 12069 33609 12081 33643
rect 12115 33640 12127 33643
rect 13170 33640 13176 33652
rect 12115 33612 13176 33640
rect 12115 33609 12127 33612
rect 12069 33603 12127 33609
rect 13170 33600 13176 33612
rect 13228 33600 13234 33652
rect 13541 33643 13599 33649
rect 13541 33609 13553 33643
rect 13587 33640 13599 33643
rect 13630 33640 13636 33652
rect 13587 33612 13636 33640
rect 13587 33609 13599 33612
rect 13541 33603 13599 33609
rect 13630 33600 13636 33612
rect 13688 33600 13694 33652
rect 18046 33640 18052 33652
rect 14108 33612 18052 33640
rect 1394 33464 1400 33516
rect 1452 33504 1458 33516
rect 2041 33507 2099 33513
rect 2041 33504 2053 33507
rect 1452 33476 2053 33504
rect 1452 33464 1458 33476
rect 2041 33473 2053 33476
rect 2087 33473 2099 33507
rect 2498 33504 2504 33516
rect 2459 33476 2504 33504
rect 2041 33467 2099 33473
rect 2498 33464 2504 33476
rect 2556 33464 2562 33516
rect 12253 33507 12311 33513
rect 12253 33504 12265 33507
rect 12084 33476 12265 33504
rect 12084 33368 12112 33476
rect 12253 33473 12265 33476
rect 12299 33473 12311 33507
rect 12710 33504 12716 33516
rect 12671 33476 12716 33504
rect 12253 33467 12311 33473
rect 12710 33464 12716 33476
rect 12768 33464 12774 33516
rect 12897 33507 12955 33513
rect 12897 33473 12909 33507
rect 12943 33504 12955 33507
rect 13078 33504 13084 33516
rect 12943 33476 13084 33504
rect 12943 33473 12955 33476
rect 12897 33467 12955 33473
rect 13078 33464 13084 33476
rect 13136 33464 13142 33516
rect 13354 33504 13360 33516
rect 13315 33476 13360 33504
rect 13354 33464 13360 33476
rect 13412 33464 13418 33516
rect 13446 33464 13452 33516
rect 13504 33504 13510 33516
rect 14108 33513 14136 33612
rect 18046 33600 18052 33612
rect 18104 33600 18110 33652
rect 18340 33612 19222 33640
rect 14458 33532 14464 33584
rect 14516 33572 14522 33584
rect 14982 33575 15040 33581
rect 14982 33572 14994 33575
rect 14516 33544 14994 33572
rect 14516 33532 14522 33544
rect 14982 33541 14994 33544
rect 15028 33541 15040 33575
rect 14982 33535 15040 33541
rect 15654 33532 15660 33584
rect 15712 33572 15718 33584
rect 16574 33572 16580 33584
rect 15712 33544 16580 33572
rect 15712 33532 15718 33544
rect 16574 33532 16580 33544
rect 16632 33532 16638 33584
rect 18340 33572 18368 33612
rect 16691 33544 18368 33572
rect 13541 33507 13599 33513
rect 13541 33504 13553 33507
rect 13504 33476 13553 33504
rect 13504 33464 13510 33476
rect 13541 33473 13553 33476
rect 13587 33473 13599 33507
rect 13541 33467 13599 33473
rect 14093 33507 14151 33513
rect 14093 33473 14105 33507
rect 14139 33473 14151 33507
rect 14093 33467 14151 33473
rect 14277 33507 14335 33513
rect 14277 33473 14289 33507
rect 14323 33504 14335 33507
rect 14550 33504 14556 33516
rect 14323 33476 14556 33504
rect 14323 33473 14335 33476
rect 14277 33467 14335 33473
rect 14550 33464 14556 33476
rect 14608 33464 14614 33516
rect 16691 33504 16719 33544
rect 18414 33532 18420 33584
rect 18472 33572 18478 33584
rect 18601 33575 18659 33581
rect 18601 33572 18613 33575
rect 18472 33544 18613 33572
rect 18472 33532 18478 33544
rect 18601 33541 18613 33544
rect 18647 33541 18659 33575
rect 18601 33535 18659 33541
rect 18690 33532 18696 33584
rect 18748 33532 18754 33584
rect 18817 33575 18875 33581
rect 18817 33541 18829 33575
rect 18863 33572 18875 33575
rect 18966 33572 18972 33584
rect 18863 33544 18972 33572
rect 18863 33541 18875 33544
rect 18817 33535 18875 33541
rect 18966 33532 18972 33544
rect 19024 33532 19030 33584
rect 16850 33504 16856 33516
rect 14660 33476 16719 33504
rect 16811 33476 16856 33504
rect 12158 33396 12164 33448
rect 12216 33436 12222 33448
rect 13906 33436 13912 33448
rect 12216 33408 13912 33436
rect 12216 33396 12222 33408
rect 13906 33396 13912 33408
rect 13964 33396 13970 33448
rect 14185 33439 14243 33445
rect 14185 33405 14197 33439
rect 14231 33436 14243 33439
rect 14660 33436 14688 33476
rect 16850 33464 16856 33476
rect 16908 33504 16914 33516
rect 17788 33513 17980 33514
rect 17788 33507 18015 33513
rect 17788 33504 17969 33507
rect 16908 33486 17969 33504
rect 16908 33476 17816 33486
rect 17952 33476 17969 33486
rect 16908 33464 16914 33476
rect 17957 33473 17969 33476
rect 18003 33473 18015 33507
rect 18138 33504 18144 33516
rect 18099 33476 18144 33504
rect 17957 33467 18015 33473
rect 18138 33464 18144 33476
rect 18196 33464 18202 33516
rect 18230 33464 18236 33516
rect 18288 33504 18294 33516
rect 18708 33504 18736 33532
rect 18288 33476 18736 33504
rect 19194 33504 19222 33612
rect 19334 33600 19340 33652
rect 19392 33640 19398 33652
rect 19392 33612 20668 33640
rect 19392 33600 19398 33612
rect 20438 33532 20444 33584
rect 20496 33572 20502 33584
rect 20533 33575 20591 33581
rect 20533 33572 20545 33575
rect 20496 33544 20545 33572
rect 20496 33532 20502 33544
rect 20533 33541 20545 33544
rect 20579 33541 20591 33575
rect 20640 33572 20668 33612
rect 21818 33600 21824 33652
rect 21876 33640 21882 33652
rect 21876 33612 21921 33640
rect 21876 33600 21882 33612
rect 22094 33600 22100 33652
rect 22152 33640 22158 33652
rect 23201 33643 23259 33649
rect 23201 33640 23213 33643
rect 22152 33612 23213 33640
rect 22152 33600 22158 33612
rect 23201 33609 23213 33612
rect 23247 33609 23259 33643
rect 23201 33603 23259 33609
rect 24578 33600 24584 33652
rect 24636 33640 24642 33652
rect 25314 33640 25320 33652
rect 24636 33612 25320 33640
rect 24636 33600 24642 33612
rect 25314 33600 25320 33612
rect 25372 33600 25378 33652
rect 25406 33600 25412 33652
rect 25464 33640 25470 33652
rect 25501 33643 25559 33649
rect 25501 33640 25513 33643
rect 25464 33612 25513 33640
rect 25464 33600 25470 33612
rect 25501 33609 25513 33612
rect 25547 33609 25559 33643
rect 27798 33640 27804 33652
rect 25501 33603 25559 33609
rect 26252 33612 27804 33640
rect 26252 33572 26280 33612
rect 27798 33600 27804 33612
rect 27856 33600 27862 33652
rect 28077 33643 28135 33649
rect 28077 33609 28089 33643
rect 28123 33640 28135 33643
rect 28810 33640 28816 33652
rect 28123 33612 28816 33640
rect 28123 33609 28135 33612
rect 28077 33603 28135 33609
rect 28810 33600 28816 33612
rect 28868 33600 28874 33652
rect 30285 33643 30343 33649
rect 30285 33609 30297 33643
rect 30331 33640 30343 33643
rect 31202 33640 31208 33652
rect 30331 33612 31208 33640
rect 30331 33609 30343 33612
rect 30285 33603 30343 33609
rect 31202 33600 31208 33612
rect 31260 33600 31266 33652
rect 31573 33643 31631 33649
rect 31573 33609 31585 33643
rect 31619 33640 31631 33643
rect 32674 33640 32680 33652
rect 31619 33612 32680 33640
rect 31619 33609 31631 33612
rect 31573 33603 31631 33609
rect 32674 33600 32680 33612
rect 32732 33600 32738 33652
rect 20640 33544 26280 33572
rect 20533 33535 20591 33541
rect 19610 33504 19616 33516
rect 19194 33476 19616 33504
rect 18288 33464 18294 33476
rect 19610 33464 19616 33476
rect 19668 33464 19674 33516
rect 19794 33504 19800 33516
rect 19755 33476 19800 33504
rect 19794 33464 19800 33476
rect 19852 33464 19858 33516
rect 19889 33507 19947 33513
rect 19889 33473 19901 33507
rect 19935 33473 19947 33507
rect 20070 33504 20076 33516
rect 20031 33476 20076 33504
rect 19889 33467 19947 33473
rect 14231 33408 14688 33436
rect 14737 33439 14795 33445
rect 14231 33405 14243 33408
rect 14185 33399 14243 33405
rect 14737 33405 14749 33439
rect 14783 33405 14795 33439
rect 14737 33399 14795 33405
rect 16669 33439 16727 33445
rect 16669 33405 16681 33439
rect 16715 33436 16727 33439
rect 17402 33436 17408 33448
rect 16715 33408 17408 33436
rect 16715 33405 16727 33408
rect 16669 33399 16727 33405
rect 14366 33368 14372 33380
rect 12084 33340 14372 33368
rect 14366 33328 14372 33340
rect 14424 33328 14430 33380
rect 14550 33328 14556 33380
rect 14608 33368 14614 33380
rect 14752 33368 14780 33399
rect 17402 33396 17408 33408
rect 17460 33396 17466 33448
rect 17773 33439 17831 33445
rect 17773 33405 17785 33439
rect 17819 33405 17831 33439
rect 17773 33399 17831 33405
rect 14608 33340 14780 33368
rect 14608 33328 14614 33340
rect 16390 33328 16396 33380
rect 16448 33368 16454 33380
rect 17037 33371 17095 33377
rect 17037 33368 17049 33371
rect 16448 33340 17049 33368
rect 16448 33328 16454 33340
rect 17037 33337 17049 33340
rect 17083 33337 17095 33371
rect 17037 33331 17095 33337
rect 17218 33328 17224 33380
rect 17276 33368 17282 33380
rect 17781 33368 17809 33399
rect 18046 33396 18052 33448
rect 18104 33436 18110 33448
rect 19518 33436 19524 33448
rect 18104 33408 19524 33436
rect 18104 33396 18110 33408
rect 19518 33396 19524 33408
rect 19576 33396 19582 33448
rect 19904 33436 19932 33467
rect 20070 33464 20076 33476
rect 20128 33464 20134 33516
rect 21634 33464 21640 33516
rect 21692 33504 21698 33516
rect 22005 33507 22063 33513
rect 22005 33504 22017 33507
rect 21692 33476 22017 33504
rect 21692 33464 21698 33476
rect 22005 33473 22017 33476
rect 22051 33473 22063 33507
rect 22005 33467 22063 33473
rect 22094 33464 22100 33516
rect 22152 33504 22158 33516
rect 22266 33507 22324 33513
rect 22152 33476 22197 33504
rect 22152 33464 22158 33476
rect 22266 33473 22278 33507
rect 22312 33473 22324 33507
rect 22266 33467 22324 33473
rect 22296 33436 22324 33467
rect 22370 33464 22376 33516
rect 22428 33504 22434 33516
rect 22428 33476 22473 33504
rect 22428 33464 22434 33476
rect 22646 33464 22652 33516
rect 22704 33504 22710 33516
rect 22704 33476 22968 33504
rect 22704 33464 22710 33476
rect 22738 33436 22744 33448
rect 19720 33408 22229 33436
rect 22296 33408 22744 33436
rect 17276 33340 17809 33368
rect 17276 33328 17282 33340
rect 18506 33328 18512 33380
rect 18564 33368 18570 33380
rect 19150 33368 19156 33380
rect 18564 33340 19156 33368
rect 18564 33328 18570 33340
rect 19150 33328 19156 33340
rect 19208 33328 19214 33380
rect 19720 33368 19748 33408
rect 19444 33340 19748 33368
rect 12802 33300 12808 33312
rect 12763 33272 12808 33300
rect 12802 33260 12808 33272
rect 12860 33260 12866 33312
rect 13170 33260 13176 33312
rect 13228 33300 13234 33312
rect 15930 33300 15936 33312
rect 13228 33272 15936 33300
rect 13228 33260 13234 33272
rect 15930 33260 15936 33272
rect 15988 33260 15994 33312
rect 16022 33260 16028 33312
rect 16080 33300 16086 33312
rect 16117 33303 16175 33309
rect 16117 33300 16129 33303
rect 16080 33272 16129 33300
rect 16080 33260 16086 33272
rect 16117 33269 16129 33272
rect 16163 33269 16175 33303
rect 16117 33263 16175 33269
rect 16206 33260 16212 33312
rect 16264 33300 16270 33312
rect 17310 33300 17316 33312
rect 16264 33272 17316 33300
rect 16264 33260 16270 33272
rect 17310 33260 17316 33272
rect 17368 33260 17374 33312
rect 17402 33260 17408 33312
rect 17460 33300 17466 33312
rect 18782 33300 18788 33312
rect 17460 33272 18788 33300
rect 17460 33260 17466 33272
rect 18782 33260 18788 33272
rect 18840 33260 18846 33312
rect 18874 33260 18880 33312
rect 18932 33300 18938 33312
rect 18969 33303 19027 33309
rect 18969 33300 18981 33303
rect 18932 33272 18981 33300
rect 18932 33260 18938 33272
rect 18969 33269 18981 33272
rect 19015 33269 19027 33303
rect 18969 33263 19027 33269
rect 19058 33260 19064 33312
rect 19116 33300 19122 33312
rect 19444 33300 19472 33340
rect 19794 33328 19800 33380
rect 19852 33368 19858 33380
rect 20809 33371 20867 33377
rect 20809 33368 20821 33371
rect 19852 33340 20821 33368
rect 19852 33328 19858 33340
rect 20809 33337 20821 33340
rect 20855 33337 20867 33371
rect 20809 33331 20867 33337
rect 20993 33371 21051 33377
rect 20993 33337 21005 33371
rect 21039 33368 21051 33371
rect 22094 33368 22100 33380
rect 21039 33340 22100 33368
rect 21039 33337 21051 33340
rect 20993 33331 21051 33337
rect 22094 33328 22100 33340
rect 22152 33328 22158 33380
rect 22201 33368 22229 33408
rect 22738 33396 22744 33408
rect 22796 33396 22802 33448
rect 22833 33439 22891 33445
rect 22833 33405 22845 33439
rect 22879 33405 22891 33439
rect 22940 33436 22968 33476
rect 23014 33464 23020 33516
rect 23072 33504 23078 33516
rect 23072 33476 23117 33504
rect 23072 33464 23078 33476
rect 23842 33464 23848 33516
rect 23900 33504 23906 33516
rect 24118 33504 24124 33516
rect 23900 33476 24124 33504
rect 23900 33464 23906 33476
rect 24118 33464 24124 33476
rect 24176 33464 24182 33516
rect 24377 33507 24435 33513
rect 24377 33504 24389 33507
rect 24219 33476 24389 33504
rect 23658 33436 23664 33448
rect 22940 33408 23664 33436
rect 22833 33399 22891 33405
rect 22646 33368 22652 33380
rect 22201 33340 22652 33368
rect 22646 33328 22652 33340
rect 22704 33328 22710 33380
rect 22848 33368 22876 33399
rect 23658 33396 23664 33408
rect 23716 33396 23722 33448
rect 24219 33436 24247 33476
rect 24377 33473 24389 33476
rect 24423 33473 24435 33507
rect 26050 33504 26056 33516
rect 26011 33476 26056 33504
rect 24377 33467 24435 33473
rect 26050 33464 26056 33476
rect 26108 33464 26114 33516
rect 26252 33513 26280 33544
rect 27246 33532 27252 33584
rect 27304 33572 27310 33584
rect 27522 33572 27528 33584
rect 27304 33544 27528 33572
rect 27304 33532 27310 33544
rect 27522 33532 27528 33544
rect 27580 33572 27586 33584
rect 27918 33575 27976 33581
rect 27918 33572 27930 33575
rect 27580 33544 27930 33572
rect 27580 33532 27586 33544
rect 27918 33541 27930 33544
rect 27964 33541 27976 33575
rect 27918 33535 27976 33541
rect 28442 33532 28448 33584
rect 28500 33572 28506 33584
rect 29362 33572 29368 33584
rect 28500 33544 29368 33572
rect 28500 33532 28506 33544
rect 29362 33532 29368 33544
rect 29420 33532 29426 33584
rect 29822 33532 29828 33584
rect 29880 33572 29886 33584
rect 30929 33575 30987 33581
rect 30929 33572 30941 33575
rect 29880 33544 30941 33572
rect 29880 33532 29886 33544
rect 30929 33541 30941 33544
rect 30975 33541 30987 33575
rect 30929 33535 30987 33541
rect 31846 33532 31852 33584
rect 31904 33572 31910 33584
rect 32493 33575 32551 33581
rect 32493 33572 32505 33575
rect 31904 33544 32505 33572
rect 31904 33532 31910 33544
rect 32493 33541 32505 33544
rect 32539 33541 32551 33575
rect 32493 33535 32551 33541
rect 26237 33507 26295 33513
rect 26237 33473 26249 33507
rect 26283 33473 26295 33507
rect 26237 33467 26295 33473
rect 26421 33507 26479 33513
rect 26421 33473 26433 33507
rect 26467 33504 26479 33507
rect 28721 33507 28779 33513
rect 28721 33504 28733 33507
rect 26467 33476 28733 33504
rect 26467 33473 26479 33476
rect 26421 33467 26479 33473
rect 28000 33448 28028 33476
rect 28721 33473 28733 33476
rect 28767 33473 28779 33507
rect 28721 33467 28779 33473
rect 28813 33507 28871 33513
rect 28813 33473 28825 33507
rect 28859 33504 28871 33507
rect 28902 33504 28908 33516
rect 28859 33476 28908 33504
rect 28859 33473 28871 33476
rect 28813 33467 28871 33473
rect 23768 33408 24247 33436
rect 22922 33368 22928 33380
rect 22848 33340 22928 33368
rect 22922 33328 22928 33340
rect 22980 33328 22986 33380
rect 23768 33377 23796 33408
rect 25314 33396 25320 33448
rect 25372 33436 25378 33448
rect 27430 33436 27436 33448
rect 25372 33408 27436 33436
rect 25372 33396 25378 33408
rect 27430 33396 27436 33408
rect 27488 33396 27494 33448
rect 27709 33439 27767 33445
rect 27709 33405 27721 33439
rect 27755 33405 27767 33439
rect 27709 33399 27767 33405
rect 23753 33371 23811 33377
rect 23753 33368 23765 33371
rect 23032 33340 23765 33368
rect 19116 33272 19472 33300
rect 19116 33260 19122 33272
rect 19518 33260 19524 33312
rect 19576 33300 19582 33312
rect 23032 33300 23060 33340
rect 23753 33337 23765 33340
rect 23799 33337 23811 33371
rect 23753 33331 23811 33337
rect 26050 33328 26056 33380
rect 26108 33368 26114 33380
rect 27724 33368 27752 33399
rect 27982 33396 27988 33448
rect 28040 33396 28046 33448
rect 28350 33396 28356 33448
rect 28408 33436 28414 33448
rect 28828 33436 28856 33467
rect 28902 33464 28908 33476
rect 28960 33464 28966 33516
rect 29089 33507 29147 33513
rect 29089 33473 29101 33507
rect 29135 33504 29147 33507
rect 29454 33504 29460 33516
rect 29135 33476 29460 33504
rect 29135 33473 29147 33476
rect 29089 33467 29147 33473
rect 29454 33464 29460 33476
rect 29512 33464 29518 33516
rect 30101 33507 30159 33513
rect 30101 33504 30113 33507
rect 29564 33476 30113 33504
rect 28994 33436 29000 33448
rect 28408 33408 28856 33436
rect 28955 33408 29000 33436
rect 28408 33396 28414 33408
rect 28994 33396 29000 33408
rect 29052 33396 29058 33448
rect 29270 33396 29276 33448
rect 29328 33436 29334 33448
rect 29564 33436 29592 33476
rect 30101 33473 30113 33476
rect 30147 33473 30159 33507
rect 31294 33504 31300 33516
rect 31255 33476 31300 33504
rect 30101 33467 30159 33473
rect 29328 33408 29592 33436
rect 29641 33439 29699 33445
rect 29328 33396 29334 33408
rect 29641 33405 29653 33439
rect 29687 33405 29699 33439
rect 30006 33436 30012 33448
rect 29967 33408 30012 33436
rect 29641 33399 29699 33405
rect 26108 33340 27752 33368
rect 26108 33328 26114 33340
rect 29454 33328 29460 33380
rect 29512 33368 29518 33380
rect 29656 33368 29684 33399
rect 30006 33396 30012 33408
rect 30064 33396 30070 33448
rect 29512 33340 29684 33368
rect 30116 33368 30144 33467
rect 31294 33464 31300 33476
rect 31352 33464 31358 33516
rect 32306 33504 32312 33516
rect 32267 33476 32312 33504
rect 32306 33464 32312 33476
rect 32364 33464 32370 33516
rect 30742 33396 30748 33448
rect 30800 33436 30806 33448
rect 31389 33439 31447 33445
rect 31389 33436 31401 33439
rect 30800 33408 31401 33436
rect 30800 33396 30806 33408
rect 31389 33405 31401 33408
rect 31435 33436 31447 33439
rect 33686 33436 33692 33448
rect 31435 33408 33692 33436
rect 31435 33405 31447 33408
rect 31389 33399 31447 33405
rect 33686 33396 33692 33408
rect 33744 33396 33750 33448
rect 34146 33436 34152 33448
rect 34107 33408 34152 33436
rect 34146 33396 34152 33408
rect 34204 33396 34210 33448
rect 31294 33368 31300 33380
rect 30116 33340 31300 33368
rect 29512 33328 29518 33340
rect 31294 33328 31300 33340
rect 31352 33328 31358 33380
rect 19576 33272 23060 33300
rect 19576 33260 19582 33272
rect 23106 33260 23112 33312
rect 23164 33300 23170 33312
rect 28350 33300 28356 33312
rect 23164 33272 28356 33300
rect 23164 33260 23170 33272
rect 28350 33260 28356 33272
rect 28408 33260 28414 33312
rect 28537 33303 28595 33309
rect 28537 33269 28549 33303
rect 28583 33300 28595 33303
rect 29822 33300 29828 33312
rect 28583 33272 29828 33300
rect 28583 33269 28595 33272
rect 28537 33263 28595 33269
rect 29822 33260 29828 33272
rect 29880 33260 29886 33312
rect 30282 33260 30288 33312
rect 30340 33300 30346 33312
rect 30742 33300 30748 33312
rect 30340 33272 30748 33300
rect 30340 33260 30346 33272
rect 30742 33260 30748 33272
rect 30800 33300 30806 33312
rect 32030 33300 32036 33312
rect 30800 33272 32036 33300
rect 30800 33260 30806 33272
rect 32030 33260 32036 33272
rect 32088 33260 32094 33312
rect 1104 33210 34868 33232
rect 1104 33158 6582 33210
rect 6634 33158 6646 33210
rect 6698 33158 6710 33210
rect 6762 33158 6774 33210
rect 6826 33158 6838 33210
rect 6890 33158 17846 33210
rect 17898 33158 17910 33210
rect 17962 33158 17974 33210
rect 18026 33158 18038 33210
rect 18090 33158 18102 33210
rect 18154 33158 29110 33210
rect 29162 33158 29174 33210
rect 29226 33158 29238 33210
rect 29290 33158 29302 33210
rect 29354 33158 29366 33210
rect 29418 33158 34868 33210
rect 1104 33136 34868 33158
rect 12069 33099 12127 33105
rect 12069 33065 12081 33099
rect 12115 33096 12127 33099
rect 12158 33096 12164 33108
rect 12115 33068 12164 33096
rect 12115 33065 12127 33068
rect 12069 33059 12127 33065
rect 12158 33056 12164 33068
rect 12216 33056 12222 33108
rect 16390 33096 16396 33108
rect 12268 33068 16396 33096
rect 12268 32901 12296 33068
rect 16390 33056 16396 33068
rect 16448 33056 16454 33108
rect 16482 33056 16488 33108
rect 16540 33096 16546 33108
rect 18506 33096 18512 33108
rect 16540 33068 18512 33096
rect 16540 33056 16546 33068
rect 18506 33056 18512 33068
rect 18564 33056 18570 33108
rect 18598 33056 18604 33108
rect 18656 33056 18662 33108
rect 18693 33099 18751 33105
rect 18693 33065 18705 33099
rect 18739 33096 18751 33099
rect 18782 33096 18788 33108
rect 18739 33068 18788 33096
rect 18739 33065 18751 33068
rect 18693 33059 18751 33065
rect 18782 33056 18788 33068
rect 18840 33096 18846 33108
rect 19058 33096 19064 33108
rect 18840 33068 19064 33096
rect 18840 33056 18846 33068
rect 19058 33056 19064 33068
rect 19116 33056 19122 33108
rect 19426 33056 19432 33108
rect 19484 33096 19490 33108
rect 22186 33096 22192 33108
rect 19484 33068 22192 33096
rect 19484 33056 19490 33068
rect 22186 33056 22192 33068
rect 22244 33056 22250 33108
rect 22370 33056 22376 33108
rect 22428 33096 22434 33108
rect 29641 33099 29699 33105
rect 22428 33068 29224 33096
rect 22428 33056 22434 33068
rect 12713 33031 12771 33037
rect 12713 32997 12725 33031
rect 12759 32997 12771 33031
rect 12713 32991 12771 32997
rect 13449 33031 13507 33037
rect 13449 32997 13461 33031
rect 13495 33028 13507 33031
rect 13538 33028 13544 33040
rect 13495 33000 13544 33028
rect 13495 32997 13507 33000
rect 13449 32991 13507 32997
rect 12728 32960 12756 32991
rect 13538 32988 13544 33000
rect 13596 32988 13602 33040
rect 14108 33000 15148 33028
rect 14108 32960 14136 33000
rect 14645 32963 14703 32969
rect 12728 32932 14136 32960
rect 14200 32932 14504 32960
rect 12253 32895 12311 32901
rect 12253 32861 12265 32895
rect 12299 32861 12311 32895
rect 12894 32892 12900 32904
rect 12855 32864 12900 32892
rect 12253 32855 12311 32861
rect 12894 32852 12900 32864
rect 12952 32852 12958 32904
rect 13170 32852 13176 32904
rect 13228 32892 13234 32904
rect 13357 32895 13415 32901
rect 13357 32892 13369 32895
rect 13228 32864 13369 32892
rect 13228 32852 13234 32864
rect 13357 32861 13369 32864
rect 13403 32861 13415 32895
rect 13357 32855 13415 32861
rect 13541 32895 13599 32901
rect 13541 32861 13553 32895
rect 13587 32892 13599 32895
rect 13630 32892 13636 32904
rect 13587 32864 13636 32892
rect 13587 32861 13599 32864
rect 13541 32855 13599 32861
rect 13630 32852 13636 32864
rect 13688 32852 13694 32904
rect 12802 32784 12808 32836
rect 12860 32824 12866 32836
rect 14200 32824 14228 32932
rect 14476 32904 14504 32932
rect 14645 32929 14657 32963
rect 14691 32960 14703 32963
rect 14734 32960 14740 32972
rect 14691 32932 14740 32960
rect 14691 32929 14703 32932
rect 14645 32923 14703 32929
rect 14734 32920 14740 32932
rect 14792 32920 14798 32972
rect 15120 32960 15148 33000
rect 16574 32988 16580 33040
rect 16632 33028 16638 33040
rect 18616 33028 18644 33056
rect 16632 33000 17356 33028
rect 16632 32988 16638 33000
rect 15120 32932 15240 32960
rect 14277 32895 14335 32901
rect 14277 32861 14289 32895
rect 14323 32861 14335 32895
rect 14458 32892 14464 32904
rect 14371 32864 14464 32892
rect 14277 32855 14335 32861
rect 12860 32796 14228 32824
rect 12860 32784 12866 32796
rect 14292 32756 14320 32855
rect 14458 32852 14464 32864
rect 14516 32852 14522 32904
rect 14550 32852 14556 32904
rect 14608 32892 14614 32904
rect 14918 32892 14924 32904
rect 14608 32864 14924 32892
rect 14608 32852 14614 32864
rect 14918 32852 14924 32864
rect 14976 32892 14982 32904
rect 15105 32895 15163 32901
rect 15105 32892 15117 32895
rect 14976 32864 15117 32892
rect 14976 32852 14982 32864
rect 15105 32861 15117 32864
rect 15151 32861 15163 32895
rect 15212 32892 15240 32932
rect 16114 32920 16120 32972
rect 16172 32960 16178 32972
rect 17126 32960 17132 32972
rect 16172 32932 17132 32960
rect 16172 32920 16178 32932
rect 17126 32920 17132 32932
rect 17184 32920 17190 32972
rect 17328 32960 17356 33000
rect 18331 33000 18644 33028
rect 17328 32932 17448 32960
rect 15212 32864 15516 32892
rect 15105 32855 15163 32861
rect 15194 32784 15200 32836
rect 15252 32824 15258 32836
rect 15350 32827 15408 32833
rect 15350 32824 15362 32827
rect 15252 32796 15362 32824
rect 15252 32784 15258 32796
rect 15350 32793 15362 32796
rect 15396 32793 15408 32827
rect 15488 32824 15516 32864
rect 15654 32852 15660 32904
rect 15712 32892 15718 32904
rect 16298 32892 16304 32904
rect 15712 32864 16304 32892
rect 15712 32852 15718 32864
rect 16298 32852 16304 32864
rect 16356 32892 16362 32904
rect 16850 32892 16856 32904
rect 16356 32864 16856 32892
rect 16356 32852 16362 32864
rect 16850 32852 16856 32864
rect 16908 32852 16914 32904
rect 16942 32852 16948 32904
rect 17000 32892 17006 32904
rect 17313 32895 17371 32901
rect 17313 32892 17325 32895
rect 17000 32864 17325 32892
rect 17000 32852 17006 32864
rect 17313 32861 17325 32864
rect 17359 32861 17371 32895
rect 17420 32892 17448 32932
rect 17420 32890 18092 32892
rect 18156 32890 18276 32892
rect 18331 32890 18359 33000
rect 18966 32988 18972 33040
rect 19024 33028 19030 33040
rect 19150 33028 19156 33040
rect 19024 33000 19156 33028
rect 19024 32988 19030 33000
rect 19150 32988 19156 33000
rect 19208 32988 19214 33040
rect 20714 32988 20720 33040
rect 20772 33028 20778 33040
rect 21910 33028 21916 33040
rect 20772 33000 21916 33028
rect 20772 32988 20778 33000
rect 21910 32988 21916 33000
rect 21968 33028 21974 33040
rect 22097 33031 22155 33037
rect 22097 33028 22109 33031
rect 21968 33000 22109 33028
rect 21968 32988 21974 33000
rect 22097 32997 22109 33000
rect 22143 32997 22155 33031
rect 22554 33028 22560 33040
rect 22515 33000 22560 33028
rect 22097 32991 22155 32997
rect 22554 32988 22560 33000
rect 22612 32988 22618 33040
rect 22646 32988 22652 33040
rect 22704 33028 22710 33040
rect 23845 33031 23903 33037
rect 23845 33028 23857 33031
rect 22704 33000 23857 33028
rect 22704 32988 22710 33000
rect 23845 32997 23857 33000
rect 23891 32997 23903 33031
rect 23845 32991 23903 32997
rect 24486 32988 24492 33040
rect 24544 33028 24550 33040
rect 24673 33031 24731 33037
rect 24673 33028 24685 33031
rect 24544 33000 24685 33028
rect 24544 32988 24550 33000
rect 24673 32997 24685 33000
rect 24719 32997 24731 33031
rect 24673 32991 24731 32997
rect 25593 33031 25651 33037
rect 25593 32997 25605 33031
rect 25639 33028 25651 33031
rect 25774 33028 25780 33040
rect 25639 33000 25780 33028
rect 25639 32997 25651 33000
rect 25593 32991 25651 32997
rect 25774 32988 25780 33000
rect 25832 32988 25838 33040
rect 27430 32988 27436 33040
rect 27488 33028 27494 33040
rect 27525 33031 27583 33037
rect 27525 33028 27537 33031
rect 27488 33000 27537 33028
rect 27488 32988 27494 33000
rect 27525 32997 27537 33000
rect 27571 32997 27583 33031
rect 27525 32991 27583 32997
rect 27709 33031 27767 33037
rect 27709 32997 27721 33031
rect 27755 33028 27767 33031
rect 27798 33028 27804 33040
rect 27755 33000 27804 33028
rect 27755 32997 27767 33000
rect 27709 32991 27767 32997
rect 27798 32988 27804 33000
rect 27856 32988 27862 33040
rect 28460 33000 28672 33028
rect 19242 32960 19248 32972
rect 17420 32864 18359 32890
rect 18064 32862 18184 32864
rect 18248 32862 18359 32864
rect 18432 32932 18670 32960
rect 19203 32932 19248 32960
rect 17313 32855 17371 32861
rect 17558 32827 17616 32833
rect 17558 32824 17570 32827
rect 15488 32796 17570 32824
rect 15350 32787 15408 32793
rect 17558 32793 17570 32796
rect 17604 32793 17616 32827
rect 17558 32787 17616 32793
rect 17678 32784 17684 32836
rect 17736 32824 17742 32836
rect 18432 32824 18460 32932
rect 18642 32892 18670 32932
rect 19242 32920 19248 32932
rect 19300 32920 19306 32972
rect 23106 32960 23112 32972
rect 20272 32932 23112 32960
rect 20272 32892 20300 32932
rect 23106 32920 23112 32932
rect 23164 32920 23170 32972
rect 23198 32920 23204 32972
rect 23256 32960 23262 32972
rect 23256 32932 23704 32960
rect 23256 32920 23262 32932
rect 21358 32892 21364 32904
rect 18642 32870 18722 32892
rect 18892 32870 20300 32892
rect 18642 32864 20300 32870
rect 21319 32864 21364 32892
rect 18694 32842 18920 32864
rect 21358 32852 21364 32864
rect 21416 32852 21422 32904
rect 21542 32892 21548 32904
rect 21503 32864 21548 32892
rect 21542 32852 21548 32864
rect 21600 32852 21606 32904
rect 21634 32852 21640 32904
rect 21692 32892 21698 32904
rect 21775 32895 21833 32901
rect 21692 32864 21737 32892
rect 21692 32852 21698 32864
rect 21775 32861 21787 32895
rect 21821 32861 21833 32895
rect 21775 32855 21833 32861
rect 21913 32895 21971 32901
rect 21913 32861 21925 32895
rect 21959 32892 21971 32895
rect 22094 32892 22100 32904
rect 21959 32864 22100 32892
rect 21959 32861 21971 32864
rect 21913 32855 21971 32861
rect 21805 32836 21833 32855
rect 22094 32852 22100 32864
rect 22152 32852 22158 32904
rect 22646 32892 22652 32904
rect 22201 32864 22652 32892
rect 17736 32796 18460 32824
rect 17736 32784 17742 32796
rect 18966 32784 18972 32836
rect 19024 32824 19030 32836
rect 19518 32833 19524 32836
rect 19024 32796 19472 32824
rect 19024 32784 19030 32796
rect 15470 32756 15476 32768
rect 14292 32728 15476 32756
rect 15470 32716 15476 32728
rect 15528 32716 15534 32768
rect 15562 32716 15568 32768
rect 15620 32756 15626 32768
rect 16390 32756 16396 32768
rect 15620 32728 16396 32756
rect 15620 32716 15626 32728
rect 16390 32716 16396 32728
rect 16448 32716 16454 32768
rect 16482 32716 16488 32768
rect 16540 32756 16546 32768
rect 16540 32728 16585 32756
rect 16540 32716 16546 32728
rect 17218 32716 17224 32768
rect 17276 32756 17282 32768
rect 18598 32756 18604 32768
rect 17276 32728 18604 32756
rect 17276 32716 17282 32728
rect 18598 32716 18604 32728
rect 18656 32716 18662 32768
rect 18782 32716 18788 32768
rect 18840 32756 18846 32768
rect 19150 32756 19156 32768
rect 18840 32728 19156 32756
rect 18840 32716 18846 32728
rect 19150 32716 19156 32728
rect 19208 32716 19214 32768
rect 19444 32756 19472 32796
rect 19512 32787 19524 32833
rect 19576 32824 19582 32836
rect 19576 32796 19612 32824
rect 19518 32784 19524 32787
rect 19576 32784 19582 32796
rect 19886 32784 19892 32836
rect 19944 32824 19950 32836
rect 21082 32824 21088 32836
rect 19944 32796 21088 32824
rect 19944 32784 19950 32796
rect 21082 32784 21088 32796
rect 21140 32784 21146 32836
rect 21805 32824 21824 32836
rect 21731 32796 21824 32824
rect 21818 32784 21824 32796
rect 21876 32824 21882 32836
rect 22201 32824 22229 32864
rect 22646 32852 22652 32864
rect 22704 32852 22710 32904
rect 22830 32901 22836 32904
rect 22787 32895 22836 32901
rect 22787 32861 22799 32895
rect 22833 32861 22836 32895
rect 22787 32855 22836 32861
rect 22830 32852 22836 32855
rect 22888 32852 22894 32904
rect 23014 32892 23020 32904
rect 22975 32864 23020 32892
rect 23014 32852 23020 32864
rect 23072 32852 23078 32904
rect 23676 32901 23704 32932
rect 23750 32920 23756 32972
rect 23808 32960 23814 32972
rect 24762 32960 24768 32972
rect 23808 32932 24768 32960
rect 23808 32920 23814 32932
rect 24504 32901 24532 32932
rect 24762 32920 24768 32932
rect 24820 32960 24826 32972
rect 26053 32963 26111 32969
rect 24820 32932 25820 32960
rect 24820 32920 24826 32932
rect 23477 32895 23535 32901
rect 23477 32861 23489 32895
rect 23523 32861 23535 32895
rect 23477 32855 23535 32861
rect 23661 32895 23719 32901
rect 23661 32861 23673 32895
rect 23707 32861 23719 32895
rect 23661 32855 23719 32861
rect 24489 32895 24547 32901
rect 24489 32861 24501 32895
rect 24535 32861 24547 32895
rect 25409 32895 25467 32901
rect 24489 32855 24547 32861
rect 24826 32864 25360 32892
rect 23492 32824 23520 32855
rect 21876 32796 22229 32824
rect 22399 32796 23520 32824
rect 21876 32784 21882 32796
rect 20625 32759 20683 32765
rect 20625 32756 20637 32759
rect 19444 32728 20637 32756
rect 20625 32725 20637 32728
rect 20671 32756 20683 32759
rect 20898 32756 20904 32768
rect 20671 32728 20904 32756
rect 20671 32725 20683 32728
rect 20625 32719 20683 32725
rect 20898 32716 20904 32728
rect 20956 32756 20962 32768
rect 22399 32756 22427 32796
rect 23566 32784 23572 32836
rect 23624 32824 23630 32836
rect 24026 32824 24032 32836
rect 23624 32796 24032 32824
rect 23624 32784 23630 32796
rect 24026 32784 24032 32796
rect 24084 32784 24090 32836
rect 20956 32728 22427 32756
rect 20956 32716 20962 32728
rect 22462 32716 22468 32768
rect 22520 32756 22526 32768
rect 22925 32759 22983 32765
rect 22925 32756 22937 32759
rect 22520 32728 22937 32756
rect 22520 32716 22526 32728
rect 22925 32725 22937 32728
rect 22971 32725 22983 32759
rect 22925 32719 22983 32725
rect 23106 32716 23112 32768
rect 23164 32756 23170 32768
rect 24826 32756 24854 32864
rect 25225 32827 25283 32833
rect 25225 32793 25237 32827
rect 25271 32793 25283 32827
rect 25332 32824 25360 32864
rect 25409 32861 25421 32895
rect 25455 32892 25467 32895
rect 25682 32892 25688 32904
rect 25455 32864 25688 32892
rect 25455 32861 25467 32864
rect 25409 32855 25467 32861
rect 25682 32852 25688 32864
rect 25740 32852 25746 32904
rect 25792 32892 25820 32932
rect 26053 32929 26065 32963
rect 26099 32960 26111 32963
rect 27246 32960 27252 32972
rect 26099 32932 27252 32960
rect 26099 32929 26111 32932
rect 26053 32923 26111 32929
rect 27246 32920 27252 32932
rect 27304 32920 27310 32972
rect 28460 32969 28488 33000
rect 28445 32963 28503 32969
rect 28445 32929 28457 32963
rect 28491 32929 28503 32963
rect 28644 32960 28672 33000
rect 28718 32988 28724 33040
rect 28776 33028 28782 33040
rect 29086 33028 29092 33040
rect 28776 33000 29092 33028
rect 28776 32988 28782 33000
rect 29086 32988 29092 33000
rect 29144 32988 29150 33040
rect 28994 32960 29000 32972
rect 28644 32932 29000 32960
rect 28445 32923 28503 32929
rect 28994 32920 29000 32932
rect 29052 32920 29058 32972
rect 26237 32895 26295 32901
rect 26237 32892 26249 32895
rect 25792 32864 26249 32892
rect 26237 32861 26249 32864
rect 26283 32861 26295 32895
rect 26237 32855 26295 32861
rect 28074 32852 28080 32904
rect 28132 32892 28138 32904
rect 28169 32895 28227 32901
rect 28169 32892 28181 32895
rect 28132 32864 28181 32892
rect 28132 32852 28138 32864
rect 28169 32861 28181 32864
rect 28215 32861 28227 32895
rect 28350 32892 28356 32904
rect 28311 32864 28356 32892
rect 28169 32855 28227 32861
rect 28350 32852 28356 32864
rect 28408 32852 28414 32904
rect 28537 32895 28595 32901
rect 28537 32890 28549 32895
rect 28460 32862 28549 32890
rect 26421 32827 26479 32833
rect 26421 32824 26433 32827
rect 25332 32796 26433 32824
rect 25225 32787 25283 32793
rect 26421 32793 26433 32796
rect 26467 32793 26479 32827
rect 26421 32787 26479 32793
rect 23164 32728 24854 32756
rect 25240 32756 25268 32787
rect 27982 32784 27988 32836
rect 28040 32824 28046 32836
rect 28460 32824 28488 32862
rect 28537 32861 28549 32862
rect 28583 32861 28595 32895
rect 28537 32855 28595 32861
rect 28704 32895 28762 32901
rect 28704 32861 28716 32895
rect 28750 32861 28762 32895
rect 28704 32855 28762 32861
rect 28040 32796 28488 32824
rect 28040 32784 28046 32796
rect 26142 32756 26148 32768
rect 25240 32728 26148 32756
rect 23164 32716 23170 32728
rect 26142 32716 26148 32728
rect 26200 32716 26206 32768
rect 27798 32716 27804 32768
rect 27856 32756 27862 32768
rect 28350 32756 28356 32768
rect 27856 32728 28356 32756
rect 27856 32716 27862 32728
rect 28350 32716 28356 32728
rect 28408 32756 28414 32768
rect 28722 32756 28750 32855
rect 29196 32824 29224 33068
rect 29641 33065 29653 33099
rect 29687 33096 29699 33099
rect 29730 33096 29736 33108
rect 29687 33068 29736 33096
rect 29687 33065 29699 33068
rect 29641 33059 29699 33065
rect 29730 33056 29736 33068
rect 29788 33056 29794 33108
rect 30098 33096 30104 33108
rect 29840 33068 30104 33096
rect 29270 32988 29276 33040
rect 29328 33028 29334 33040
rect 29546 33028 29552 33040
rect 29328 33000 29552 33028
rect 29328 32988 29334 33000
rect 29546 32988 29552 33000
rect 29604 32988 29610 33040
rect 29840 33028 29868 33068
rect 30098 33056 30104 33068
rect 30156 33056 30162 33108
rect 30561 33099 30619 33105
rect 30561 33065 30573 33099
rect 30607 33096 30619 33099
rect 31202 33096 31208 33108
rect 30607 33068 31208 33096
rect 30607 33065 30619 33068
rect 30561 33059 30619 33065
rect 31202 33056 31208 33068
rect 31260 33056 31266 33108
rect 29656 33000 29868 33028
rect 29546 32892 29552 32904
rect 29459 32864 29552 32892
rect 29546 32852 29552 32864
rect 29604 32892 29610 32904
rect 29656 32892 29684 33000
rect 29914 32988 29920 33040
rect 29972 33028 29978 33040
rect 29972 33000 30604 33028
rect 29972 32988 29978 33000
rect 29730 32920 29736 32972
rect 29788 32960 29794 32972
rect 30469 32963 30527 32969
rect 30469 32960 30481 32963
rect 29788 32932 30481 32960
rect 29788 32920 29794 32932
rect 30469 32929 30481 32932
rect 30515 32929 30527 32963
rect 30469 32923 30527 32929
rect 29604 32864 29684 32892
rect 29604 32852 29610 32864
rect 29822 32852 29828 32904
rect 29880 32892 29886 32904
rect 30193 32895 30251 32901
rect 30193 32892 30205 32895
rect 29880 32864 30205 32892
rect 29880 32852 29886 32864
rect 30193 32861 30205 32864
rect 30239 32861 30251 32895
rect 30576 32892 30604 33000
rect 31478 32988 31484 33040
rect 31536 33028 31542 33040
rect 31536 33000 31754 33028
rect 31536 32988 31542 33000
rect 31726 32960 31754 33000
rect 31938 32988 31944 33040
rect 31996 33028 32002 33040
rect 31996 33000 32720 33028
rect 31996 32988 32002 33000
rect 32692 32969 32720 33000
rect 31849 32963 31907 32969
rect 31849 32960 31861 32963
rect 31726 32932 31861 32960
rect 31849 32929 31861 32932
rect 31895 32960 31907 32963
rect 32677 32963 32735 32969
rect 31895 32932 32352 32960
rect 31895 32929 31907 32932
rect 31849 32923 31907 32929
rect 31481 32895 31539 32901
rect 31481 32892 31493 32895
rect 30576 32864 31493 32892
rect 30193 32855 30251 32861
rect 31481 32861 31493 32864
rect 31527 32861 31539 32895
rect 31662 32892 31668 32904
rect 31623 32864 31668 32892
rect 31481 32855 31539 32861
rect 31662 32852 31668 32864
rect 31720 32852 31726 32904
rect 31757 32895 31815 32901
rect 31757 32861 31769 32895
rect 31803 32861 31815 32895
rect 32030 32892 32036 32904
rect 31943 32864 32036 32892
rect 31757 32855 31815 32861
rect 31772 32824 31800 32855
rect 32030 32852 32036 32864
rect 32088 32852 32094 32904
rect 32324 32892 32352 32932
rect 32677 32929 32689 32963
rect 32723 32929 32735 32963
rect 32677 32923 32735 32929
rect 33318 32892 33324 32904
rect 32324 32864 33324 32892
rect 33318 32852 33324 32864
rect 33376 32852 33382 32904
rect 29196 32796 31800 32824
rect 28408 32728 28750 32756
rect 28408 32716 28414 32728
rect 28810 32716 28816 32768
rect 28868 32756 28874 32768
rect 28905 32759 28963 32765
rect 28905 32756 28917 32759
rect 28868 32728 28917 32756
rect 28868 32716 28874 32728
rect 28905 32725 28917 32728
rect 28951 32725 28963 32759
rect 28905 32719 28963 32725
rect 29454 32716 29460 32768
rect 29512 32756 29518 32768
rect 29822 32756 29828 32768
rect 29512 32728 29828 32756
rect 29512 32716 29518 32728
rect 29822 32716 29828 32728
rect 29880 32716 29886 32768
rect 30006 32716 30012 32768
rect 30064 32756 30070 32768
rect 30374 32756 30380 32768
rect 30064 32728 30380 32756
rect 30064 32716 30070 32728
rect 30374 32716 30380 32728
rect 30432 32716 30438 32768
rect 30745 32759 30803 32765
rect 30745 32725 30757 32759
rect 30791 32756 30803 32759
rect 31846 32756 31852 32768
rect 30791 32728 31852 32756
rect 30791 32725 30803 32728
rect 30745 32719 30803 32725
rect 31846 32716 31852 32728
rect 31904 32716 31910 32768
rect 32048 32756 32076 32852
rect 32217 32827 32275 32833
rect 32217 32793 32229 32827
rect 32263 32824 32275 32827
rect 32922 32827 32980 32833
rect 32922 32824 32934 32827
rect 32263 32796 32934 32824
rect 32263 32793 32275 32796
rect 32217 32787 32275 32793
rect 32922 32793 32934 32796
rect 32968 32793 32980 32827
rect 32922 32787 32980 32793
rect 33042 32756 33048 32768
rect 32048 32728 33048 32756
rect 33042 32716 33048 32728
rect 33100 32756 33106 32768
rect 34057 32759 34115 32765
rect 34057 32756 34069 32759
rect 33100 32728 34069 32756
rect 33100 32716 33106 32728
rect 34057 32725 34069 32728
rect 34103 32725 34115 32759
rect 34057 32719 34115 32725
rect 1104 32666 34868 32688
rect 1104 32614 12214 32666
rect 12266 32614 12278 32666
rect 12330 32614 12342 32666
rect 12394 32614 12406 32666
rect 12458 32614 12470 32666
rect 12522 32614 23478 32666
rect 23530 32614 23542 32666
rect 23594 32614 23606 32666
rect 23658 32614 23670 32666
rect 23722 32614 23734 32666
rect 23786 32614 34868 32666
rect 1104 32592 34868 32614
rect 12253 32555 12311 32561
rect 12253 32521 12265 32555
rect 12299 32552 12311 32555
rect 12802 32552 12808 32564
rect 12299 32524 12808 32552
rect 12299 32521 12311 32524
rect 12253 32515 12311 32521
rect 12802 32512 12808 32524
rect 12860 32512 12866 32564
rect 12894 32512 12900 32564
rect 12952 32552 12958 32564
rect 16206 32552 16212 32564
rect 12952 32524 16212 32552
rect 12952 32512 12958 32524
rect 16206 32512 16212 32524
rect 16264 32512 16270 32564
rect 16390 32512 16396 32564
rect 16448 32552 16454 32564
rect 16853 32555 16911 32561
rect 16853 32552 16865 32555
rect 16448 32524 16865 32552
rect 16448 32512 16454 32524
rect 16853 32521 16865 32524
rect 16899 32521 16911 32555
rect 16853 32515 16911 32521
rect 17310 32512 17316 32564
rect 17368 32552 17374 32564
rect 17862 32552 17868 32564
rect 17368 32524 17868 32552
rect 17368 32512 17374 32524
rect 17862 32512 17868 32524
rect 17920 32512 17926 32564
rect 17957 32555 18015 32561
rect 17957 32521 17969 32555
rect 18003 32552 18015 32555
rect 18322 32552 18328 32564
rect 18003 32524 18328 32552
rect 18003 32521 18015 32524
rect 17957 32515 18015 32521
rect 18322 32512 18328 32524
rect 18380 32512 18386 32564
rect 18432 32524 19555 32552
rect 12986 32484 12992 32496
rect 12947 32456 12992 32484
rect 12986 32444 12992 32456
rect 13044 32444 13050 32496
rect 14550 32484 14556 32496
rect 13556 32456 14556 32484
rect 12437 32419 12495 32425
rect 12437 32385 12449 32419
rect 12483 32416 12495 32419
rect 12618 32416 12624 32428
rect 12483 32388 12624 32416
rect 12483 32385 12495 32388
rect 12437 32379 12495 32385
rect 12618 32376 12624 32388
rect 12676 32376 12682 32428
rect 12894 32416 12900 32428
rect 12855 32388 12900 32416
rect 12894 32376 12900 32388
rect 12952 32376 12958 32428
rect 13078 32416 13084 32428
rect 13039 32388 13084 32416
rect 13078 32376 13084 32388
rect 13136 32376 13142 32428
rect 13556 32425 13584 32456
rect 14550 32444 14556 32456
rect 14608 32444 14614 32496
rect 14642 32444 14648 32496
rect 14700 32484 14706 32496
rect 14918 32484 14924 32496
rect 14700 32456 14924 32484
rect 14700 32444 14706 32456
rect 14918 32444 14924 32456
rect 14976 32444 14982 32496
rect 15657 32487 15715 32493
rect 15657 32453 15669 32487
rect 15703 32484 15715 32487
rect 16114 32484 16120 32496
rect 15703 32456 16120 32484
rect 15703 32453 15715 32456
rect 15657 32447 15715 32453
rect 16114 32444 16120 32456
rect 16172 32484 16178 32496
rect 16574 32484 16580 32496
rect 16172 32456 16580 32484
rect 16172 32444 16178 32456
rect 16574 32444 16580 32456
rect 16632 32444 16638 32496
rect 16761 32487 16819 32493
rect 16761 32453 16773 32487
rect 16807 32484 16819 32487
rect 17034 32484 17040 32496
rect 16807 32456 17040 32484
rect 16807 32453 16819 32456
rect 16761 32447 16819 32453
rect 17034 32444 17040 32456
rect 17092 32444 17098 32496
rect 17405 32487 17463 32493
rect 17405 32453 17417 32487
rect 17451 32484 17463 32487
rect 18432 32484 18460 32524
rect 19242 32484 19248 32496
rect 17451 32456 17908 32484
rect 17451 32453 17463 32456
rect 17405 32447 17463 32453
rect 13541 32419 13599 32425
rect 13541 32385 13553 32419
rect 13587 32385 13599 32419
rect 13541 32379 13599 32385
rect 14185 32419 14243 32425
rect 14185 32385 14197 32419
rect 14231 32385 14243 32419
rect 14185 32379 14243 32385
rect 11790 32348 11796 32360
rect 11751 32320 11796 32348
rect 11790 32308 11796 32320
rect 11848 32308 11854 32360
rect 14200 32348 14228 32379
rect 14458 32376 14464 32428
rect 14516 32416 14522 32428
rect 15013 32419 15071 32425
rect 15013 32416 15025 32419
rect 14516 32388 15025 32416
rect 14516 32376 14522 32388
rect 15013 32385 15025 32388
rect 15059 32416 15071 32419
rect 15562 32416 15568 32428
rect 15059 32388 15568 32416
rect 15059 32385 15071 32388
rect 15013 32379 15071 32385
rect 15562 32376 15568 32388
rect 15620 32376 15626 32428
rect 15933 32419 15991 32425
rect 15933 32416 15945 32419
rect 15764 32388 15945 32416
rect 14829 32351 14887 32357
rect 14200 32320 14780 32348
rect 12342 32240 12348 32292
rect 12400 32280 12406 32292
rect 14752 32280 14780 32320
rect 14829 32317 14841 32351
rect 14875 32348 14887 32351
rect 15764 32348 15792 32388
rect 15933 32385 15945 32388
rect 15979 32416 15991 32419
rect 16482 32416 16488 32428
rect 15979 32388 16488 32416
rect 15979 32385 15991 32388
rect 15933 32379 15991 32385
rect 16482 32376 16488 32388
rect 16540 32376 16546 32428
rect 17494 32416 17500 32428
rect 16592 32388 17500 32416
rect 14875 32320 15792 32348
rect 14875 32317 14887 32320
rect 14829 32311 14887 32317
rect 15838 32308 15844 32360
rect 15896 32348 15902 32360
rect 15896 32320 15941 32348
rect 15896 32308 15902 32320
rect 16206 32308 16212 32360
rect 16264 32348 16270 32360
rect 16592 32348 16620 32388
rect 17494 32376 17500 32388
rect 17552 32376 17558 32428
rect 17593 32419 17651 32425
rect 17593 32385 17605 32419
rect 17639 32416 17651 32419
rect 17770 32416 17776 32428
rect 17639 32388 17776 32416
rect 17639 32385 17651 32388
rect 17593 32379 17651 32385
rect 17770 32376 17776 32388
rect 17828 32376 17834 32428
rect 16264 32320 16620 32348
rect 16264 32308 16270 32320
rect 17034 32308 17040 32360
rect 17092 32348 17098 32360
rect 17681 32351 17739 32357
rect 17681 32348 17693 32351
rect 17092 32320 17693 32348
rect 17092 32308 17098 32320
rect 17681 32317 17693 32320
rect 17727 32317 17739 32351
rect 17880 32348 17908 32456
rect 17972 32456 18460 32484
rect 18524 32456 19248 32484
rect 17972 32428 18000 32456
rect 17954 32376 17960 32428
rect 18012 32376 18018 32428
rect 18049 32419 18107 32425
rect 18049 32385 18061 32419
rect 18095 32416 18107 32419
rect 18230 32416 18236 32428
rect 18095 32388 18236 32416
rect 18095 32385 18107 32388
rect 18049 32379 18107 32385
rect 18230 32376 18236 32388
rect 18288 32376 18294 32428
rect 18524 32425 18552 32456
rect 19242 32444 19248 32456
rect 19300 32444 19306 32496
rect 18509 32419 18567 32425
rect 18509 32385 18521 32419
rect 18555 32385 18567 32419
rect 18765 32419 18823 32425
rect 18765 32416 18777 32419
rect 18509 32379 18567 32385
rect 18616 32388 18777 32416
rect 18616 32348 18644 32388
rect 18765 32385 18777 32388
rect 18811 32385 18823 32419
rect 18765 32379 18823 32385
rect 19058 32376 19064 32428
rect 19116 32416 19122 32428
rect 19334 32416 19340 32428
rect 19116 32388 19340 32416
rect 19116 32376 19122 32388
rect 19334 32376 19340 32388
rect 19392 32376 19398 32428
rect 17880 32320 18644 32348
rect 19527 32348 19555 32524
rect 19794 32512 19800 32564
rect 19852 32552 19858 32564
rect 19889 32555 19947 32561
rect 19889 32552 19901 32555
rect 19852 32524 19901 32552
rect 19852 32512 19858 32524
rect 19889 32521 19901 32524
rect 19935 32552 19947 32555
rect 20898 32552 20904 32564
rect 19935 32524 20392 32552
rect 20859 32524 20904 32552
rect 19935 32521 19947 32524
rect 19889 32515 19947 32521
rect 20364 32416 20392 32524
rect 20898 32512 20904 32524
rect 20956 32512 20962 32564
rect 20990 32512 20996 32564
rect 21048 32552 21054 32564
rect 21269 32555 21327 32561
rect 21048 32524 21093 32552
rect 21048 32512 21054 32524
rect 21269 32521 21281 32555
rect 21315 32552 21327 32555
rect 22738 32552 22744 32564
rect 21315 32524 22744 32552
rect 21315 32521 21327 32524
rect 21269 32515 21327 32521
rect 22738 32512 22744 32524
rect 22796 32512 22802 32564
rect 22830 32512 22836 32564
rect 22888 32552 22894 32564
rect 29825 32555 29883 32561
rect 29825 32552 29837 32555
rect 22888 32524 29837 32552
rect 22888 32512 22894 32524
rect 29825 32521 29837 32524
rect 29871 32552 29883 32555
rect 30282 32552 30288 32564
rect 29871 32524 30288 32552
rect 29871 32521 29883 32524
rect 29825 32515 29883 32521
rect 30282 32512 30288 32524
rect 30340 32512 30346 32564
rect 30650 32512 30656 32564
rect 30708 32512 30714 32564
rect 20438 32444 20444 32496
rect 20496 32484 20502 32496
rect 21110 32487 21168 32493
rect 21110 32484 21122 32487
rect 20496 32456 21122 32484
rect 20496 32444 20502 32456
rect 21110 32453 21122 32456
rect 21156 32453 21168 32487
rect 21110 32447 21168 32453
rect 21542 32444 21548 32496
rect 21600 32484 21606 32496
rect 23014 32484 23020 32496
rect 21600 32456 23020 32484
rect 21600 32444 21606 32456
rect 20530 32416 20536 32428
rect 20364 32388 20536 32416
rect 20530 32376 20536 32388
rect 20588 32416 20594 32428
rect 20625 32419 20683 32425
rect 20625 32416 20637 32419
rect 20588 32388 20637 32416
rect 20588 32376 20594 32388
rect 20625 32385 20637 32388
rect 20671 32385 20683 32419
rect 20625 32379 20683 32385
rect 21818 32376 21824 32428
rect 21876 32416 21882 32428
rect 22112 32425 22140 32456
rect 23014 32444 23020 32456
rect 23072 32444 23078 32496
rect 23198 32444 23204 32496
rect 23256 32484 23262 32496
rect 23722 32487 23780 32493
rect 23722 32484 23734 32487
rect 23256 32456 23734 32484
rect 23256 32444 23262 32456
rect 23722 32453 23734 32456
rect 23768 32453 23780 32487
rect 23722 32447 23780 32453
rect 25501 32487 25559 32493
rect 25501 32453 25513 32487
rect 25547 32484 25559 32487
rect 25547 32456 30604 32484
rect 25547 32453 25559 32456
rect 25501 32447 25559 32453
rect 22005 32419 22063 32425
rect 22005 32416 22017 32419
rect 21876 32388 22017 32416
rect 21876 32376 21882 32388
rect 22005 32385 22017 32388
rect 22051 32385 22063 32419
rect 22005 32379 22063 32385
rect 22097 32419 22155 32425
rect 22097 32385 22109 32419
rect 22143 32385 22155 32419
rect 22097 32379 22155 32385
rect 22186 32376 22192 32428
rect 22244 32416 22250 32428
rect 22373 32419 22431 32425
rect 22373 32416 22385 32419
rect 22244 32388 22385 32416
rect 22244 32376 22250 32388
rect 22373 32385 22385 32388
rect 22419 32416 22431 32419
rect 22462 32416 22468 32428
rect 22419 32388 22468 32416
rect 22419 32385 22431 32388
rect 22373 32379 22431 32385
rect 22462 32376 22468 32388
rect 22520 32376 22526 32428
rect 22833 32419 22891 32425
rect 22833 32385 22845 32419
rect 22879 32416 22891 32419
rect 22922 32416 22928 32428
rect 22879 32388 22928 32416
rect 22879 32385 22891 32388
rect 22833 32379 22891 32385
rect 22922 32376 22928 32388
rect 22980 32376 22986 32428
rect 23474 32416 23480 32428
rect 23435 32388 23480 32416
rect 23474 32376 23480 32388
rect 23532 32376 23538 32428
rect 25317 32419 25375 32425
rect 25317 32385 25329 32419
rect 25363 32416 25375 32419
rect 25406 32416 25412 32428
rect 25363 32388 25412 32416
rect 25363 32385 25375 32388
rect 25317 32379 25375 32385
rect 25406 32376 25412 32388
rect 25464 32376 25470 32428
rect 25593 32419 25651 32425
rect 25593 32385 25605 32419
rect 25639 32416 25651 32419
rect 25774 32416 25780 32428
rect 25639 32388 25780 32416
rect 25639 32385 25651 32388
rect 25593 32379 25651 32385
rect 25774 32376 25780 32388
rect 25832 32376 25838 32428
rect 26237 32419 26295 32425
rect 26237 32416 26249 32419
rect 25884 32388 26249 32416
rect 23382 32348 23388 32360
rect 19527 32320 23388 32348
rect 17681 32311 17739 32317
rect 23382 32308 23388 32320
rect 23440 32308 23446 32360
rect 17954 32280 17960 32292
rect 12400 32252 14688 32280
rect 14752 32252 17960 32280
rect 12400 32240 12406 32252
rect 13630 32212 13636 32224
rect 13591 32184 13636 32212
rect 13630 32172 13636 32184
rect 13688 32172 13694 32224
rect 14277 32215 14335 32221
rect 14277 32181 14289 32215
rect 14323 32212 14335 32215
rect 14550 32212 14556 32224
rect 14323 32184 14556 32212
rect 14323 32181 14335 32184
rect 14277 32175 14335 32181
rect 14550 32172 14556 32184
rect 14608 32172 14614 32224
rect 14660 32212 14688 32252
rect 17954 32240 17960 32252
rect 18012 32240 18018 32292
rect 20714 32280 20720 32292
rect 20088 32252 20720 32280
rect 15197 32215 15255 32221
rect 15197 32212 15209 32215
rect 14660 32184 15209 32212
rect 15197 32181 15209 32184
rect 15243 32181 15255 32215
rect 15197 32175 15255 32181
rect 15470 32172 15476 32224
rect 15528 32212 15534 32224
rect 15933 32215 15991 32221
rect 15933 32212 15945 32215
rect 15528 32184 15945 32212
rect 15528 32172 15534 32184
rect 15933 32181 15945 32184
rect 15979 32212 15991 32215
rect 16022 32212 16028 32224
rect 15979 32184 16028 32212
rect 15979 32181 15991 32184
rect 15933 32175 15991 32181
rect 16022 32172 16028 32184
rect 16080 32172 16086 32224
rect 16117 32215 16175 32221
rect 16117 32181 16129 32215
rect 16163 32212 16175 32215
rect 17310 32212 17316 32224
rect 16163 32184 17316 32212
rect 16163 32181 16175 32184
rect 16117 32175 16175 32181
rect 17310 32172 17316 32184
rect 17368 32172 17374 32224
rect 17678 32172 17684 32224
rect 17736 32212 17742 32224
rect 20088 32212 20116 32252
rect 20714 32240 20720 32252
rect 20772 32240 20778 32292
rect 20990 32240 20996 32292
rect 21048 32280 21054 32292
rect 22646 32280 22652 32292
rect 21048 32252 22652 32280
rect 21048 32240 21054 32252
rect 22646 32240 22652 32252
rect 22704 32240 22710 32292
rect 23014 32280 23020 32292
rect 22747 32252 23020 32280
rect 17736 32184 20116 32212
rect 17736 32172 17742 32184
rect 20162 32172 20168 32224
rect 20220 32212 20226 32224
rect 21726 32212 21732 32224
rect 20220 32184 21732 32212
rect 20220 32172 20226 32184
rect 21726 32172 21732 32184
rect 21784 32172 21790 32224
rect 21821 32215 21879 32221
rect 21821 32181 21833 32215
rect 21867 32212 21879 32215
rect 22094 32212 22100 32224
rect 21867 32184 22100 32212
rect 21867 32181 21879 32184
rect 21821 32175 21879 32181
rect 22094 32172 22100 32184
rect 22152 32172 22158 32224
rect 22186 32172 22192 32224
rect 22244 32212 22250 32224
rect 22281 32215 22339 32221
rect 22281 32212 22293 32215
rect 22244 32184 22293 32212
rect 22244 32172 22250 32184
rect 22281 32181 22293 32184
rect 22327 32181 22339 32215
rect 22281 32175 22339 32181
rect 22370 32172 22376 32224
rect 22428 32212 22434 32224
rect 22747 32212 22775 32252
rect 23014 32240 23020 32252
rect 23072 32240 23078 32292
rect 24486 32240 24492 32292
rect 24544 32280 24550 32292
rect 25314 32280 25320 32292
rect 24544 32252 25176 32280
rect 25275 32252 25320 32280
rect 24544 32240 24550 32252
rect 22428 32184 22775 32212
rect 22925 32215 22983 32221
rect 22428 32172 22434 32184
rect 22925 32181 22937 32215
rect 22971 32212 22983 32215
rect 23290 32212 23296 32224
rect 22971 32184 23296 32212
rect 22971 32181 22983 32184
rect 22925 32175 22983 32181
rect 23290 32172 23296 32184
rect 23348 32172 23354 32224
rect 23382 32172 23388 32224
rect 23440 32212 23446 32224
rect 24854 32212 24860 32224
rect 23440 32184 24860 32212
rect 23440 32172 23446 32184
rect 24854 32172 24860 32184
rect 24912 32172 24918 32224
rect 25148 32212 25176 32252
rect 25314 32240 25320 32252
rect 25372 32240 25378 32292
rect 25884 32280 25912 32388
rect 26237 32385 26249 32388
rect 26283 32416 26295 32419
rect 27525 32419 27583 32425
rect 26283 32388 27476 32416
rect 26283 32385 26295 32388
rect 26237 32379 26295 32385
rect 26053 32351 26111 32357
rect 26053 32317 26065 32351
rect 26099 32348 26111 32351
rect 27246 32348 27252 32360
rect 26099 32320 27252 32348
rect 26099 32317 26111 32320
rect 26053 32311 26111 32317
rect 27246 32308 27252 32320
rect 27304 32308 27310 32360
rect 27448 32348 27476 32388
rect 27525 32385 27537 32419
rect 27571 32416 27583 32419
rect 27890 32416 27896 32428
rect 27571 32388 27896 32416
rect 27571 32385 27583 32388
rect 27525 32379 27583 32385
rect 27890 32376 27896 32388
rect 27948 32376 27954 32428
rect 28350 32376 28356 32428
rect 28408 32376 28414 32428
rect 28442 32376 28448 32428
rect 28500 32416 28506 32428
rect 28610 32419 28668 32425
rect 28500 32388 28545 32416
rect 28500 32376 28506 32388
rect 28610 32385 28622 32419
rect 28656 32385 28668 32419
rect 28610 32379 28668 32385
rect 28721 32419 28779 32425
rect 28721 32385 28733 32419
rect 28767 32385 28779 32419
rect 28721 32379 28779 32385
rect 27614 32348 27620 32360
rect 27448 32320 27620 32348
rect 27614 32308 27620 32320
rect 27672 32308 27678 32360
rect 27798 32348 27804 32360
rect 27759 32320 27804 32348
rect 27798 32308 27804 32320
rect 27856 32308 27862 32360
rect 28368 32348 28396 32376
rect 28625 32348 28653 32379
rect 28368 32320 28653 32348
rect 28736 32348 28764 32379
rect 28810 32376 28816 32428
rect 28868 32416 28874 32428
rect 29457 32419 29515 32425
rect 28868 32388 28913 32416
rect 28868 32376 28874 32388
rect 29457 32385 29469 32419
rect 29503 32416 29515 32419
rect 30006 32416 30012 32428
rect 29503 32388 30012 32416
rect 29503 32385 29515 32388
rect 29457 32379 29515 32385
rect 30006 32376 30012 32388
rect 30064 32376 30070 32428
rect 29549 32351 29607 32357
rect 28736 32320 28856 32348
rect 26418 32280 26424 32292
rect 25424 32252 25912 32280
rect 26379 32252 26424 32280
rect 25424 32212 25452 32252
rect 26418 32240 26424 32252
rect 26476 32240 26482 32292
rect 27341 32283 27399 32289
rect 27341 32249 27353 32283
rect 27387 32280 27399 32283
rect 27982 32280 27988 32292
rect 27387 32252 27988 32280
rect 27387 32249 27399 32252
rect 27341 32243 27399 32249
rect 27982 32240 27988 32252
rect 28040 32240 28046 32292
rect 28626 32280 28632 32292
rect 28184 32252 28632 32280
rect 25148 32184 25452 32212
rect 25498 32172 25504 32224
rect 25556 32212 25562 32224
rect 27709 32215 27767 32221
rect 27709 32212 27721 32215
rect 25556 32184 27721 32212
rect 25556 32172 25562 32184
rect 27709 32181 27721 32184
rect 27755 32212 27767 32215
rect 28184 32212 28212 32252
rect 28626 32240 28632 32252
rect 28684 32240 28690 32292
rect 28828 32280 28856 32320
rect 29549 32317 29561 32351
rect 29595 32317 29607 32351
rect 29549 32311 29607 32317
rect 28902 32280 28908 32292
rect 28828 32252 28908 32280
rect 28902 32240 28908 32252
rect 28960 32240 28966 32292
rect 27755 32184 28212 32212
rect 28261 32215 28319 32221
rect 27755 32181 27767 32184
rect 27709 32175 27767 32181
rect 28261 32181 28273 32215
rect 28307 32212 28319 32215
rect 28994 32212 29000 32224
rect 28307 32184 29000 32212
rect 28307 32181 28319 32184
rect 28261 32175 28319 32181
rect 28994 32172 29000 32184
rect 29052 32172 29058 32224
rect 29564 32212 29592 32311
rect 30576 32280 30604 32456
rect 30668 32416 30696 32512
rect 34146 32484 34152 32496
rect 34107 32456 34152 32484
rect 34146 32444 34152 32456
rect 34204 32444 34210 32496
rect 31021 32419 31079 32425
rect 31021 32416 31033 32419
rect 30668 32388 31033 32416
rect 31021 32385 31033 32388
rect 31067 32416 31079 32419
rect 31478 32416 31484 32428
rect 31067 32388 31484 32416
rect 31067 32385 31079 32388
rect 31021 32379 31079 32385
rect 31478 32376 31484 32388
rect 31536 32376 31542 32428
rect 32306 32416 32312 32428
rect 32267 32388 32312 32416
rect 32306 32376 32312 32388
rect 32364 32376 32370 32428
rect 30742 32348 30748 32360
rect 30703 32320 30748 32348
rect 30742 32308 30748 32320
rect 30800 32308 30806 32360
rect 31662 32308 31668 32360
rect 31720 32348 31726 32360
rect 32493 32351 32551 32357
rect 32493 32348 32505 32351
rect 31720 32320 32505 32348
rect 31720 32308 31726 32320
rect 32493 32317 32505 32320
rect 32539 32317 32551 32351
rect 32493 32311 32551 32317
rect 33778 32280 33784 32292
rect 30576 32252 33784 32280
rect 33778 32240 33784 32252
rect 33836 32240 33842 32292
rect 30098 32212 30104 32224
rect 29564 32184 30104 32212
rect 30098 32172 30104 32184
rect 30156 32212 30162 32224
rect 30742 32212 30748 32224
rect 30156 32184 30748 32212
rect 30156 32172 30162 32184
rect 30742 32172 30748 32184
rect 30800 32172 30806 32224
rect 1104 32122 34868 32144
rect 1104 32070 6582 32122
rect 6634 32070 6646 32122
rect 6698 32070 6710 32122
rect 6762 32070 6774 32122
rect 6826 32070 6838 32122
rect 6890 32070 17846 32122
rect 17898 32070 17910 32122
rect 17962 32070 17974 32122
rect 18026 32070 18038 32122
rect 18090 32070 18102 32122
rect 18154 32070 29110 32122
rect 29162 32070 29174 32122
rect 29226 32070 29238 32122
rect 29290 32070 29302 32122
rect 29354 32070 29366 32122
rect 29418 32070 34868 32122
rect 1104 32048 34868 32070
rect 12805 32011 12863 32017
rect 12805 31977 12817 32011
rect 12851 32008 12863 32011
rect 14734 32008 14740 32020
rect 12851 31980 14740 32008
rect 12851 31977 12863 31980
rect 12805 31971 12863 31977
rect 14734 31968 14740 31980
rect 14792 31968 14798 32020
rect 14918 31968 14924 32020
rect 14976 32008 14982 32020
rect 15654 32008 15660 32020
rect 14976 31980 15660 32008
rect 14976 31968 14982 31980
rect 15654 31968 15660 31980
rect 15712 32008 15718 32020
rect 16206 32008 16212 32020
rect 15712 31980 16212 32008
rect 15712 31968 15718 31980
rect 16206 31968 16212 31980
rect 16264 31968 16270 32020
rect 16390 31968 16396 32020
rect 16448 32008 16454 32020
rect 16574 32008 16580 32020
rect 16448 31980 16580 32008
rect 16448 31968 16454 31980
rect 16574 31968 16580 31980
rect 16632 32008 16638 32020
rect 16669 32011 16727 32017
rect 16669 32008 16681 32011
rect 16632 31980 16681 32008
rect 16632 31968 16638 31980
rect 16669 31977 16681 31980
rect 16715 31977 16727 32011
rect 16669 31971 16727 31977
rect 16758 31968 16764 32020
rect 16816 32008 16822 32020
rect 18230 32008 18236 32020
rect 16816 31980 18236 32008
rect 16816 31968 16822 31980
rect 18230 31968 18236 31980
rect 18288 31968 18294 32020
rect 18506 31968 18512 32020
rect 18564 32008 18570 32020
rect 18598 32008 18604 32020
rect 18564 31980 18604 32008
rect 18564 31968 18570 31980
rect 18598 31968 18604 31980
rect 18656 32008 18662 32020
rect 18966 32008 18972 32020
rect 18656 31980 18972 32008
rect 18656 31968 18662 31980
rect 18966 31968 18972 31980
rect 19024 31968 19030 32020
rect 19058 31968 19064 32020
rect 19116 32008 19122 32020
rect 20714 32008 20720 32020
rect 19116 31980 20720 32008
rect 19116 31968 19122 31980
rect 20714 31968 20720 31980
rect 20772 31968 20778 32020
rect 20993 32011 21051 32017
rect 20993 31977 21005 32011
rect 21039 32008 21051 32011
rect 21634 32008 21640 32020
rect 21039 31980 21640 32008
rect 21039 31977 21051 31980
rect 20993 31971 21051 31977
rect 21634 31968 21640 31980
rect 21692 32008 21698 32020
rect 22186 32008 22192 32020
rect 21692 31980 22192 32008
rect 21692 31968 21698 31980
rect 22186 31968 22192 31980
rect 22244 31968 22250 32020
rect 22278 31968 22284 32020
rect 22336 32008 22342 32020
rect 23198 32008 23204 32020
rect 22336 31980 22508 32008
rect 23159 31980 23204 32008
rect 22336 31968 22342 31980
rect 12161 31943 12219 31949
rect 12161 31909 12173 31943
rect 12207 31909 12219 31943
rect 12161 31903 12219 31909
rect 12176 31872 12204 31903
rect 14550 31900 14556 31952
rect 14608 31940 14614 31952
rect 14829 31943 14887 31949
rect 14829 31940 14841 31943
rect 14608 31912 14841 31940
rect 14608 31900 14614 31912
rect 14829 31909 14841 31912
rect 14875 31940 14887 31943
rect 14875 31912 15332 31940
rect 14875 31909 14887 31912
rect 14829 31903 14887 31909
rect 15304 31881 15332 31912
rect 16482 31900 16488 31952
rect 16540 31940 16546 31952
rect 17129 31943 17187 31949
rect 17129 31940 17141 31943
rect 16540 31912 17141 31940
rect 16540 31900 16546 31912
rect 17129 31909 17141 31912
rect 17175 31909 17187 31943
rect 17129 31903 17187 31909
rect 18693 31943 18751 31949
rect 18693 31909 18705 31943
rect 18739 31940 18751 31943
rect 19334 31940 19340 31952
rect 18739 31912 18819 31940
rect 18739 31909 18751 31912
rect 18693 31903 18751 31909
rect 15289 31875 15347 31881
rect 12176 31844 15240 31872
rect 1486 31764 1492 31816
rect 1544 31804 1550 31816
rect 1673 31807 1731 31813
rect 1673 31804 1685 31807
rect 1544 31776 1685 31804
rect 1544 31764 1550 31776
rect 1673 31773 1685 31776
rect 1719 31773 1731 31807
rect 1673 31767 1731 31773
rect 11701 31807 11759 31813
rect 11701 31773 11713 31807
rect 11747 31773 11759 31807
rect 12342 31804 12348 31816
rect 12303 31776 12348 31804
rect 11701 31767 11759 31773
rect 11716 31736 11744 31767
rect 12342 31764 12348 31776
rect 12400 31764 12406 31816
rect 12802 31804 12808 31816
rect 12763 31776 12808 31804
rect 12802 31764 12808 31776
rect 12860 31764 12866 31816
rect 12986 31764 12992 31816
rect 13044 31804 13050 31816
rect 13044 31776 13089 31804
rect 13044 31764 13050 31776
rect 14366 31764 14372 31816
rect 14424 31804 14430 31816
rect 14645 31807 14703 31813
rect 14424 31776 14596 31804
rect 14424 31764 14430 31776
rect 14458 31736 14464 31748
rect 11716 31708 14464 31736
rect 14458 31696 14464 31708
rect 14516 31696 14522 31748
rect 14568 31736 14596 31776
rect 14645 31773 14657 31807
rect 14691 31804 14703 31807
rect 14918 31804 14924 31816
rect 14691 31776 14924 31804
rect 14691 31773 14703 31776
rect 14645 31767 14703 31773
rect 14918 31764 14924 31776
rect 14976 31764 14982 31816
rect 15102 31736 15108 31748
rect 14568 31708 15108 31736
rect 15102 31696 15108 31708
rect 15160 31696 15166 31748
rect 15212 31736 15240 31844
rect 15289 31841 15301 31875
rect 15335 31841 15347 31875
rect 15289 31835 15347 31841
rect 15304 31804 15332 31835
rect 16574 31832 16580 31884
rect 16632 31872 16638 31884
rect 17681 31875 17739 31881
rect 16632 31844 17448 31872
rect 16632 31832 16638 31844
rect 15304 31776 15884 31804
rect 15534 31739 15592 31745
rect 15534 31736 15546 31739
rect 15212 31708 15546 31736
rect 15534 31705 15546 31708
rect 15580 31705 15592 31739
rect 15534 31699 15592 31705
rect 11517 31671 11575 31677
rect 11517 31637 11529 31671
rect 11563 31668 11575 31671
rect 12710 31668 12716 31680
rect 11563 31640 12716 31668
rect 11563 31637 11575 31640
rect 11517 31631 11575 31637
rect 12710 31628 12716 31640
rect 12768 31628 12774 31680
rect 13722 31628 13728 31680
rect 13780 31668 13786 31680
rect 15286 31668 15292 31680
rect 13780 31640 15292 31668
rect 13780 31628 13786 31640
rect 15286 31628 15292 31640
rect 15344 31628 15350 31680
rect 15856 31668 15884 31776
rect 16022 31764 16028 31816
rect 16080 31804 16086 31816
rect 17420 31813 17448 31844
rect 17681 31841 17693 31875
rect 17727 31872 17739 31875
rect 18138 31872 18144 31884
rect 17727 31844 18144 31872
rect 17727 31841 17739 31844
rect 17681 31835 17739 31841
rect 18138 31832 18144 31844
rect 18196 31832 18202 31884
rect 18417 31875 18475 31881
rect 18417 31841 18429 31875
rect 18463 31872 18475 31875
rect 18791 31872 18819 31912
rect 18984 31912 19340 31940
rect 18874 31872 18880 31884
rect 18463 31844 18736 31872
rect 18791 31844 18880 31872
rect 18463 31841 18475 31844
rect 18417 31835 18475 31841
rect 17313 31807 17371 31813
rect 17313 31804 17325 31807
rect 16080 31776 17325 31804
rect 16080 31764 16086 31776
rect 17313 31773 17325 31776
rect 17359 31773 17371 31807
rect 17313 31767 17371 31773
rect 17405 31807 17463 31813
rect 17405 31773 17417 31807
rect 17451 31773 17463 31807
rect 17405 31767 17463 31773
rect 17770 31764 17776 31816
rect 17828 31804 17834 31816
rect 18509 31807 18567 31813
rect 17828 31776 18276 31804
rect 17828 31764 17834 31776
rect 15930 31696 15936 31748
rect 15988 31736 15994 31748
rect 16574 31736 16580 31748
rect 15988 31708 16580 31736
rect 15988 31696 15994 31708
rect 16574 31696 16580 31708
rect 16632 31696 16638 31748
rect 16850 31696 16856 31748
rect 16908 31736 16914 31748
rect 18248 31745 18276 31776
rect 18509 31773 18521 31807
rect 18555 31804 18567 31807
rect 18598 31804 18604 31816
rect 18555 31776 18604 31804
rect 18555 31773 18567 31776
rect 18509 31767 18567 31773
rect 18598 31764 18604 31776
rect 18656 31764 18662 31816
rect 18708 31804 18736 31844
rect 18874 31832 18880 31844
rect 18932 31832 18938 31884
rect 18984 31804 19012 31912
rect 19334 31900 19340 31912
rect 19392 31900 19398 31952
rect 20438 31900 20444 31952
rect 20496 31940 20502 31952
rect 20809 31943 20867 31949
rect 20809 31940 20821 31943
rect 20496 31912 20821 31940
rect 20496 31900 20502 31912
rect 20809 31909 20821 31912
rect 20855 31909 20867 31943
rect 22480 31940 22508 31980
rect 23198 31968 23204 31980
rect 23256 31968 23262 32020
rect 23290 31968 23296 32020
rect 23348 32008 23354 32020
rect 23348 31980 24532 32008
rect 23348 31968 23354 31980
rect 24504 31940 24532 31980
rect 24854 31968 24860 32020
rect 24912 32008 24918 32020
rect 25869 32011 25927 32017
rect 25869 32008 25881 32011
rect 24912 31980 25881 32008
rect 24912 31968 24918 31980
rect 25869 31977 25881 31980
rect 25915 31977 25927 32011
rect 30558 32008 30564 32020
rect 25869 31971 25927 31977
rect 28276 31980 30564 32008
rect 25222 31940 25228 31952
rect 20809 31903 20867 31909
rect 20916 31912 22213 31940
rect 22480 31912 24440 31940
rect 24504 31912 25228 31940
rect 20916 31884 20944 31912
rect 19150 31832 19156 31884
rect 19208 31872 19214 31884
rect 19702 31872 19708 31884
rect 19208 31844 19708 31872
rect 19208 31832 19214 31844
rect 19702 31832 19708 31844
rect 19760 31832 19766 31884
rect 20530 31872 20536 31884
rect 20491 31844 20536 31872
rect 20530 31832 20536 31844
rect 20588 31832 20594 31884
rect 20898 31832 20904 31884
rect 20956 31832 20962 31884
rect 21450 31832 21456 31884
rect 21508 31872 21514 31884
rect 21818 31872 21824 31884
rect 21508 31844 21824 31872
rect 21508 31832 21514 31844
rect 21818 31832 21824 31844
rect 21876 31832 21882 31884
rect 21910 31832 21916 31884
rect 21968 31872 21974 31884
rect 22097 31875 22155 31881
rect 22097 31872 22109 31875
rect 21968 31844 22109 31872
rect 21968 31832 21974 31844
rect 22097 31841 22109 31844
rect 22143 31841 22155 31875
rect 22185 31872 22213 31912
rect 23290 31872 23296 31884
rect 22185 31844 23296 31872
rect 22097 31835 22155 31841
rect 23290 31832 23296 31844
rect 23348 31832 23354 31884
rect 24412 31881 24440 31912
rect 25222 31900 25228 31912
rect 25280 31900 25286 31952
rect 26326 31900 26332 31952
rect 26384 31940 26390 31952
rect 26384 31912 27614 31940
rect 26384 31900 26390 31912
rect 24397 31875 24455 31881
rect 23676 31844 24348 31872
rect 18708 31776 19012 31804
rect 19306 31776 21772 31804
rect 18233 31739 18291 31745
rect 16908 31708 17632 31736
rect 16908 31696 16914 31708
rect 16206 31668 16212 31680
rect 15856 31640 16212 31668
rect 16206 31628 16212 31640
rect 16264 31628 16270 31680
rect 16390 31628 16396 31680
rect 16448 31668 16454 31680
rect 17497 31671 17555 31677
rect 17497 31668 17509 31671
rect 16448 31640 17509 31668
rect 16448 31628 16454 31640
rect 17497 31637 17509 31640
rect 17543 31637 17555 31671
rect 17604 31668 17632 31708
rect 18233 31705 18245 31739
rect 18279 31736 18291 31739
rect 18279 31708 18644 31736
rect 18279 31705 18291 31708
rect 18233 31699 18291 31705
rect 18616 31680 18644 31708
rect 19058 31696 19064 31748
rect 19116 31736 19122 31748
rect 19306 31736 19334 31776
rect 19610 31736 19616 31748
rect 19116 31708 19334 31736
rect 19571 31708 19616 31736
rect 19116 31696 19122 31708
rect 19610 31696 19616 31708
rect 19668 31696 19674 31748
rect 19702 31696 19708 31748
rect 19760 31736 19766 31748
rect 19797 31739 19855 31745
rect 19797 31736 19809 31739
rect 19760 31708 19809 31736
rect 19760 31696 19766 31708
rect 19797 31705 19809 31708
rect 19843 31736 19855 31739
rect 21634 31736 21640 31748
rect 19843 31708 21640 31736
rect 19843 31705 19855 31708
rect 19797 31699 19855 31705
rect 21634 31696 21640 31708
rect 21692 31696 21698 31748
rect 21744 31736 21772 31776
rect 22002 31764 22008 31816
rect 22060 31804 22066 31816
rect 22189 31807 22247 31813
rect 22189 31804 22201 31807
rect 22060 31776 22201 31804
rect 22060 31764 22066 31776
rect 22189 31773 22201 31776
rect 22235 31773 22247 31807
rect 22830 31804 22836 31816
rect 22189 31767 22247 31773
rect 22281 31776 22836 31804
rect 22281 31736 22309 31776
rect 22830 31764 22836 31776
rect 22888 31764 22894 31816
rect 23382 31764 23388 31816
rect 23440 31804 23446 31816
rect 23676 31813 23704 31844
rect 23477 31807 23535 31813
rect 23477 31804 23489 31807
rect 23440 31776 23489 31804
rect 23440 31764 23446 31776
rect 23477 31773 23489 31776
rect 23523 31773 23535 31807
rect 23477 31767 23535 31773
rect 23569 31807 23627 31813
rect 23569 31773 23581 31807
rect 23615 31773 23627 31807
rect 23569 31767 23627 31773
rect 23661 31807 23719 31813
rect 23661 31773 23673 31807
rect 23707 31773 23719 31807
rect 23661 31767 23719 31773
rect 23845 31807 23903 31813
rect 23845 31773 23857 31807
rect 23891 31773 23903 31807
rect 23845 31767 23903 31773
rect 21744 31708 22309 31736
rect 22646 31696 22652 31748
rect 22704 31736 22710 31748
rect 23584 31736 23612 31767
rect 22704 31708 23612 31736
rect 22704 31696 22710 31708
rect 18506 31668 18512 31680
rect 17604 31640 18512 31668
rect 17497 31631 17555 31637
rect 18506 31628 18512 31640
rect 18564 31628 18570 31680
rect 18598 31628 18604 31680
rect 18656 31628 18662 31680
rect 18874 31628 18880 31680
rect 18932 31668 18938 31680
rect 19518 31668 19524 31680
rect 18932 31640 19524 31668
rect 18932 31628 18938 31640
rect 19518 31628 19524 31640
rect 19576 31628 19582 31680
rect 20070 31628 20076 31680
rect 20128 31668 20134 31680
rect 20622 31668 20628 31680
rect 20128 31640 20628 31668
rect 20128 31628 20134 31640
rect 20622 31628 20628 31640
rect 20680 31628 20686 31680
rect 20714 31628 20720 31680
rect 20772 31668 20778 31680
rect 22557 31671 22615 31677
rect 22557 31668 22569 31671
rect 20772 31640 22569 31668
rect 20772 31628 20778 31640
rect 22557 31637 22569 31640
rect 22603 31637 22615 31671
rect 22557 31631 22615 31637
rect 22738 31628 22744 31680
rect 22796 31668 22802 31680
rect 23860 31668 23888 31767
rect 24320 31736 24348 31844
rect 24397 31841 24409 31875
rect 24443 31841 24455 31875
rect 25041 31875 25099 31881
rect 25041 31872 25053 31875
rect 24397 31835 24455 31841
rect 24504 31844 25053 31872
rect 24504 31736 24532 31844
rect 25041 31841 25053 31844
rect 25087 31841 25099 31875
rect 25041 31835 25099 31841
rect 26142 31832 26148 31884
rect 26200 31872 26206 31884
rect 26200 31844 26832 31872
rect 26200 31832 26206 31844
rect 24578 31764 24584 31816
rect 24636 31804 24642 31816
rect 24765 31807 24823 31813
rect 24765 31804 24777 31807
rect 24636 31776 24777 31804
rect 24636 31764 24642 31776
rect 24765 31773 24777 31776
rect 24811 31773 24823 31807
rect 24765 31767 24823 31773
rect 24857 31807 24915 31813
rect 24857 31773 24869 31807
rect 24903 31773 24915 31807
rect 25498 31804 25504 31816
rect 25459 31776 25504 31804
rect 24857 31767 24915 31773
rect 24320 31708 24532 31736
rect 24670 31696 24676 31748
rect 24728 31736 24734 31748
rect 24872 31736 24900 31767
rect 25498 31764 25504 31776
rect 25556 31764 25562 31816
rect 25590 31764 25596 31816
rect 25648 31804 25654 31816
rect 26804 31813 26832 31844
rect 25685 31807 25743 31813
rect 25685 31804 25697 31807
rect 25648 31776 25697 31804
rect 25648 31764 25654 31776
rect 25685 31773 25697 31776
rect 25731 31773 25743 31807
rect 25685 31767 25743 31773
rect 25961 31807 26019 31813
rect 25961 31773 25973 31807
rect 26007 31773 26019 31807
rect 25961 31767 26019 31773
rect 26651 31807 26709 31813
rect 26651 31773 26663 31807
rect 26697 31773 26709 31807
rect 26651 31767 26709 31773
rect 26789 31807 26847 31813
rect 26789 31773 26801 31807
rect 26835 31773 26847 31807
rect 26789 31767 26847 31773
rect 25976 31736 26004 31767
rect 24728 31708 24900 31736
rect 25700 31708 26004 31736
rect 24728 31696 24734 31708
rect 25700 31680 25728 31708
rect 26050 31696 26056 31748
rect 26108 31736 26114 31748
rect 26666 31736 26694 31767
rect 26878 31764 26884 31816
rect 26936 31804 26942 31816
rect 27062 31804 27068 31816
rect 26936 31776 26981 31804
rect 27023 31776 27068 31804
rect 26936 31764 26942 31776
rect 27062 31764 27068 31776
rect 27120 31764 27126 31816
rect 27586 31804 27614 31912
rect 27798 31872 27804 31884
rect 27759 31844 27804 31872
rect 27798 31832 27804 31844
rect 27856 31832 27862 31884
rect 27890 31832 27896 31884
rect 27948 31832 27954 31884
rect 27709 31807 27767 31813
rect 27709 31804 27721 31807
rect 27586 31776 27721 31804
rect 27709 31773 27721 31776
rect 27755 31773 27767 31807
rect 27908 31804 27936 31832
rect 27908 31776 28028 31804
rect 27709 31767 27767 31773
rect 27890 31736 27896 31748
rect 26108 31708 27896 31736
rect 26108 31696 26114 31708
rect 27890 31696 27896 31708
rect 27948 31696 27954 31748
rect 28000 31736 28028 31776
rect 28074 31764 28080 31816
rect 28132 31804 28138 31816
rect 28276 31804 28304 31980
rect 30558 31968 30564 31980
rect 30616 31968 30622 32020
rect 30653 32011 30711 32017
rect 30653 31977 30665 32011
rect 30699 32008 30711 32011
rect 30926 32008 30932 32020
rect 30699 31980 30932 32008
rect 30699 31977 30711 31980
rect 30653 31971 30711 31977
rect 28626 31900 28632 31952
rect 28684 31940 28690 31952
rect 29270 31940 29276 31952
rect 28684 31912 29276 31940
rect 28684 31900 28690 31912
rect 29270 31900 29276 31912
rect 29328 31900 29334 31952
rect 30098 31832 30104 31884
rect 30156 31872 30162 31884
rect 30193 31875 30251 31881
rect 30193 31872 30205 31875
rect 30156 31844 30205 31872
rect 30156 31832 30162 31844
rect 30193 31841 30205 31844
rect 30239 31841 30251 31875
rect 30193 31835 30251 31841
rect 30374 31832 30380 31884
rect 30432 31872 30438 31884
rect 30668 31872 30696 31971
rect 30926 31968 30932 31980
rect 30984 31968 30990 32020
rect 31662 32008 31668 32020
rect 31036 31980 31668 32008
rect 30432 31844 30696 31872
rect 30432 31832 30438 31844
rect 28537 31807 28595 31813
rect 28537 31804 28549 31807
rect 28132 31776 28549 31804
rect 28132 31764 28138 31776
rect 28537 31773 28549 31776
rect 28583 31773 28595 31807
rect 28718 31804 28724 31816
rect 28679 31776 28724 31804
rect 28537 31767 28595 31773
rect 28718 31764 28724 31776
rect 28776 31764 28782 31816
rect 28994 31804 29000 31816
rect 28955 31776 29000 31804
rect 28994 31764 29000 31776
rect 29052 31764 29058 31816
rect 30285 31807 30343 31813
rect 30285 31804 30297 31807
rect 29748 31776 30297 31804
rect 29748 31736 29776 31776
rect 30285 31773 30297 31776
rect 30331 31804 30343 31807
rect 30650 31804 30656 31816
rect 30331 31776 30656 31804
rect 30331 31773 30343 31776
rect 30285 31767 30343 31773
rect 30650 31764 30656 31776
rect 30708 31764 30714 31816
rect 28000 31708 29776 31736
rect 29822 31696 29828 31748
rect 29880 31736 29886 31748
rect 30190 31736 30196 31748
rect 29880 31708 30196 31736
rect 29880 31696 29886 31708
rect 30190 31696 30196 31708
rect 30248 31696 30254 31748
rect 24210 31668 24216 31680
rect 22796 31640 24216 31668
rect 22796 31628 22802 31640
rect 24210 31628 24216 31640
rect 24268 31628 24274 31680
rect 25682 31628 25688 31680
rect 25740 31628 25746 31680
rect 26421 31671 26479 31677
rect 26421 31637 26433 31671
rect 26467 31668 26479 31671
rect 26602 31668 26608 31680
rect 26467 31640 26608 31668
rect 26467 31637 26479 31640
rect 26421 31631 26479 31637
rect 26602 31628 26608 31640
rect 26660 31628 26666 31680
rect 28074 31668 28080 31680
rect 28035 31640 28080 31668
rect 28074 31628 28080 31640
rect 28132 31628 28138 31680
rect 28626 31628 28632 31680
rect 28684 31668 28690 31680
rect 28905 31671 28963 31677
rect 28905 31668 28917 31671
rect 28684 31640 28917 31668
rect 28684 31628 28690 31640
rect 28905 31637 28917 31640
rect 28951 31637 28963 31671
rect 28905 31631 28963 31637
rect 28994 31628 29000 31680
rect 29052 31668 29058 31680
rect 31036 31668 31064 31980
rect 31662 31968 31668 31980
rect 31720 31968 31726 32020
rect 31478 31900 31484 31952
rect 31536 31900 31542 31952
rect 31849 31943 31907 31949
rect 31849 31909 31861 31943
rect 31895 31940 31907 31943
rect 32030 31940 32036 31952
rect 31895 31912 32036 31940
rect 31895 31909 31907 31912
rect 31849 31903 31907 31909
rect 32030 31900 32036 31912
rect 32088 31940 32094 31952
rect 33410 31940 33416 31952
rect 32088 31912 33416 31940
rect 32088 31900 32094 31912
rect 33410 31900 33416 31912
rect 33468 31900 33474 31952
rect 31389 31875 31447 31881
rect 31389 31841 31401 31875
rect 31435 31872 31447 31875
rect 31496 31872 31524 31900
rect 31938 31872 31944 31884
rect 31435 31844 31944 31872
rect 31435 31841 31447 31844
rect 31389 31835 31447 31841
rect 31938 31832 31944 31844
rect 31996 31832 32002 31884
rect 32306 31872 32312 31884
rect 32267 31844 32312 31872
rect 32306 31832 32312 31844
rect 32364 31832 32370 31884
rect 32493 31875 32551 31881
rect 32493 31841 32505 31875
rect 32539 31872 32551 31875
rect 32582 31872 32588 31884
rect 32539 31844 32588 31872
rect 32539 31841 32551 31844
rect 32493 31835 32551 31841
rect 32582 31832 32588 31844
rect 32640 31832 32646 31884
rect 34146 31872 34152 31884
rect 34107 31844 34152 31872
rect 34146 31832 34152 31844
rect 34204 31832 34210 31884
rect 31478 31804 31484 31816
rect 31439 31776 31484 31804
rect 31478 31764 31484 31776
rect 31536 31764 31542 31816
rect 29052 31640 31064 31668
rect 29052 31628 29058 31640
rect 1104 31578 34868 31600
rect 1104 31526 12214 31578
rect 12266 31526 12278 31578
rect 12330 31526 12342 31578
rect 12394 31526 12406 31578
rect 12458 31526 12470 31578
rect 12522 31526 23478 31578
rect 23530 31526 23542 31578
rect 23594 31526 23606 31578
rect 23658 31526 23670 31578
rect 23722 31526 23734 31578
rect 23786 31526 34868 31578
rect 1104 31504 34868 31526
rect 12897 31467 12955 31473
rect 12897 31433 12909 31467
rect 12943 31464 12955 31467
rect 12986 31464 12992 31476
rect 12943 31436 12992 31464
rect 12943 31433 12955 31436
rect 12897 31427 12955 31433
rect 12986 31424 12992 31436
rect 13044 31424 13050 31476
rect 13464 31436 18460 31464
rect 1486 31328 1492 31340
rect 1447 31300 1492 31328
rect 1486 31288 1492 31300
rect 1544 31288 1550 31340
rect 12250 31328 12256 31340
rect 12211 31300 12256 31328
rect 12250 31288 12256 31300
rect 12308 31288 12314 31340
rect 12805 31331 12863 31337
rect 12805 31297 12817 31331
rect 12851 31328 12863 31331
rect 12894 31328 12900 31340
rect 12851 31300 12900 31328
rect 12851 31297 12863 31300
rect 12805 31291 12863 31297
rect 12894 31288 12900 31300
rect 12952 31288 12958 31340
rect 13464 31337 13492 31436
rect 14642 31356 14648 31408
rect 14700 31396 14706 31408
rect 14982 31399 15040 31405
rect 14982 31396 14994 31399
rect 14700 31368 14994 31396
rect 14700 31356 14706 31368
rect 14982 31365 14994 31368
rect 15028 31365 15040 31399
rect 14982 31359 15040 31365
rect 15102 31356 15108 31408
rect 15160 31396 15166 31408
rect 16758 31396 16764 31408
rect 15160 31368 16620 31396
rect 16719 31368 16764 31396
rect 15160 31356 15166 31368
rect 12989 31331 13047 31337
rect 12989 31297 13001 31331
rect 13035 31297 13047 31331
rect 12989 31291 13047 31297
rect 13449 31331 13507 31337
rect 13449 31297 13461 31331
rect 13495 31297 13507 31331
rect 13449 31291 13507 31297
rect 13633 31331 13691 31337
rect 13633 31297 13645 31331
rect 13679 31328 13691 31331
rect 13722 31328 13728 31340
rect 13679 31300 13728 31328
rect 13679 31297 13691 31300
rect 13633 31291 13691 31297
rect 1673 31263 1731 31269
rect 1673 31229 1685 31263
rect 1719 31260 1731 31263
rect 1854 31260 1860 31272
rect 1719 31232 1860 31260
rect 1719 31229 1731 31232
rect 1673 31223 1731 31229
rect 1854 31220 1860 31232
rect 1912 31220 1918 31272
rect 1946 31220 1952 31272
rect 2004 31260 2010 31272
rect 13004 31260 13032 31291
rect 13722 31288 13728 31300
rect 13780 31288 13786 31340
rect 13814 31288 13820 31340
rect 13872 31328 13878 31340
rect 14093 31331 14151 31337
rect 14093 31328 14105 31331
rect 13872 31300 14105 31328
rect 13872 31288 13878 31300
rect 14093 31297 14105 31300
rect 14139 31297 14151 31331
rect 14093 31291 14151 31297
rect 14550 31288 14556 31340
rect 14608 31328 14614 31340
rect 14737 31331 14795 31337
rect 14737 31328 14749 31331
rect 14608 31300 14749 31328
rect 14608 31288 14614 31300
rect 14737 31297 14749 31300
rect 14783 31297 14795 31331
rect 16482 31328 16488 31340
rect 14737 31291 14795 31297
rect 14852 31300 16488 31328
rect 13998 31260 14004 31272
rect 2004 31232 2049 31260
rect 13004 31232 14004 31260
rect 2004 31220 2010 31232
rect 13998 31220 14004 31232
rect 14056 31220 14062 31272
rect 14185 31263 14243 31269
rect 14185 31229 14197 31263
rect 14231 31260 14243 31263
rect 14852 31260 14880 31300
rect 16482 31288 16488 31300
rect 16540 31288 16546 31340
rect 16592 31328 16620 31368
rect 16758 31356 16764 31368
rect 16816 31356 16822 31408
rect 16945 31399 17003 31405
rect 16945 31365 16957 31399
rect 16991 31396 17003 31399
rect 18230 31396 18236 31408
rect 16991 31368 17908 31396
rect 18191 31368 18236 31396
rect 16991 31365 17003 31368
rect 16945 31359 17003 31365
rect 17034 31328 17040 31340
rect 16592 31300 17040 31328
rect 17034 31288 17040 31300
rect 17092 31288 17098 31340
rect 17218 31288 17224 31340
rect 17276 31328 17282 31340
rect 17589 31331 17647 31337
rect 17589 31328 17601 31331
rect 17276 31300 17601 31328
rect 17276 31288 17282 31300
rect 17589 31297 17601 31300
rect 17635 31297 17647 31331
rect 17880 31328 17908 31368
rect 18230 31356 18236 31368
rect 18288 31356 18294 31408
rect 18432 31396 18460 31436
rect 18506 31424 18512 31476
rect 18564 31464 18570 31476
rect 18564 31436 19295 31464
rect 18564 31424 18570 31436
rect 18432 31368 19196 31396
rect 18046 31328 18052 31340
rect 17880 31300 18052 31328
rect 17589 31291 17647 31297
rect 18046 31288 18052 31300
rect 18104 31288 18110 31340
rect 18322 31288 18328 31340
rect 18380 31328 18386 31340
rect 18782 31338 18788 31340
rect 18694 31337 18788 31338
rect 18417 31331 18475 31337
rect 18417 31328 18429 31331
rect 18380 31300 18429 31328
rect 18380 31288 18386 31300
rect 18417 31297 18429 31300
rect 18463 31297 18475 31331
rect 18417 31291 18475 31297
rect 18673 31331 18788 31337
rect 18673 31297 18685 31331
rect 18719 31310 18788 31331
rect 18719 31297 18731 31310
rect 18673 31291 18731 31297
rect 14231 31232 14880 31260
rect 14231 31229 14243 31232
rect 14185 31223 14243 31229
rect 15838 31220 15844 31272
rect 15896 31260 15902 31272
rect 15896 31232 16979 31260
rect 15896 31220 15902 31232
rect 12069 31195 12127 31201
rect 12069 31161 12081 31195
rect 12115 31192 12127 31195
rect 12115 31164 14780 31192
rect 12115 31161 12127 31164
rect 12069 31155 12127 31161
rect 13538 31124 13544 31136
rect 13499 31096 13544 31124
rect 13538 31084 13544 31096
rect 13596 31084 13602 31136
rect 13998 31084 14004 31136
rect 14056 31124 14062 31136
rect 14550 31124 14556 31136
rect 14056 31096 14556 31124
rect 14056 31084 14062 31096
rect 14550 31084 14556 31096
rect 14608 31084 14614 31136
rect 14752 31124 14780 31164
rect 15930 31152 15936 31204
rect 15988 31192 15994 31204
rect 16117 31195 16175 31201
rect 16117 31192 16129 31195
rect 15988 31164 16129 31192
rect 15988 31152 15994 31164
rect 16117 31161 16129 31164
rect 16163 31161 16175 31195
rect 16117 31155 16175 31161
rect 16482 31152 16488 31204
rect 16540 31192 16546 31204
rect 16850 31192 16856 31204
rect 16540 31164 16856 31192
rect 16540 31152 16546 31164
rect 16850 31152 16856 31164
rect 16908 31152 16914 31204
rect 16951 31192 16979 31232
rect 17126 31220 17132 31272
rect 17184 31260 17190 31272
rect 17405 31263 17463 31269
rect 17405 31260 17417 31263
rect 17184 31232 17417 31260
rect 17184 31220 17190 31232
rect 17405 31229 17417 31232
rect 17451 31260 17463 31263
rect 17494 31260 17500 31272
rect 17451 31232 17500 31260
rect 17451 31229 17463 31232
rect 17405 31223 17463 31229
rect 17494 31220 17500 31232
rect 17552 31220 17558 31272
rect 17678 31220 17684 31272
rect 17736 31260 17742 31272
rect 18432 31260 18460 31291
rect 18782 31288 18788 31310
rect 18840 31288 18846 31340
rect 18874 31260 18880 31272
rect 17736 31232 18092 31260
rect 18432 31232 18880 31260
rect 17736 31220 17742 31232
rect 18064 31192 18092 31232
rect 18874 31220 18880 31232
rect 18932 31220 18938 31272
rect 18601 31195 18659 31201
rect 18601 31192 18613 31195
rect 16951 31164 17908 31192
rect 18064 31164 18613 31192
rect 16666 31124 16672 31136
rect 14752 31096 16672 31124
rect 16666 31084 16672 31096
rect 16724 31084 16730 31136
rect 16942 31084 16948 31136
rect 17000 31124 17006 31136
rect 17773 31127 17831 31133
rect 17773 31124 17785 31127
rect 17000 31096 17785 31124
rect 17000 31084 17006 31096
rect 17773 31093 17785 31096
rect 17819 31093 17831 31127
rect 17880 31124 17908 31164
rect 18601 31161 18613 31164
rect 18647 31161 18659 31195
rect 19168 31192 19196 31368
rect 19267 31260 19295 31436
rect 20824 31436 21312 31464
rect 19613 31399 19671 31405
rect 19613 31365 19625 31399
rect 19659 31396 19671 31399
rect 20349 31399 20407 31405
rect 20349 31396 20361 31399
rect 19659 31368 20361 31396
rect 19659 31365 19671 31368
rect 19613 31359 19671 31365
rect 20349 31365 20361 31368
rect 20395 31396 20407 31399
rect 20824 31396 20852 31436
rect 21284 31425 21312 31436
rect 21284 31397 21404 31425
rect 21450 31424 21456 31476
rect 21508 31464 21514 31476
rect 24118 31464 24124 31476
rect 21508 31436 24124 31464
rect 21508 31424 21514 31436
rect 24118 31424 24124 31436
rect 24176 31424 24182 31476
rect 24210 31424 24216 31476
rect 24268 31464 24274 31476
rect 27062 31464 27068 31476
rect 24268 31436 27068 31464
rect 24268 31424 24274 31436
rect 27062 31424 27068 31436
rect 27120 31464 27126 31476
rect 27430 31464 27436 31476
rect 27120 31436 27436 31464
rect 27120 31424 27126 31436
rect 27430 31424 27436 31436
rect 27488 31424 27494 31476
rect 27982 31424 27988 31476
rect 28040 31464 28046 31476
rect 28258 31464 28264 31476
rect 28040 31436 28264 31464
rect 28040 31424 28046 31436
rect 28258 31424 28264 31436
rect 28316 31424 28322 31476
rect 28534 31424 28540 31476
rect 28592 31464 28598 31476
rect 28592 31436 28994 31464
rect 28592 31424 28598 31436
rect 20395 31368 20852 31396
rect 21376 31396 21404 31397
rect 22094 31396 22100 31408
rect 21376 31368 22100 31396
rect 20395 31365 20407 31368
rect 20349 31359 20407 31365
rect 19334 31288 19340 31340
rect 19392 31328 19398 31340
rect 20162 31328 20168 31340
rect 19392 31300 20168 31328
rect 19392 31288 19398 31300
rect 20162 31288 20168 31300
rect 20220 31328 20226 31340
rect 20533 31331 20591 31337
rect 20533 31328 20545 31331
rect 20220 31300 20545 31328
rect 20220 31288 20226 31300
rect 20533 31297 20545 31300
rect 20579 31297 20591 31331
rect 20533 31291 20591 31297
rect 20993 31331 21051 31337
rect 20993 31297 21005 31331
rect 21039 31328 21051 31331
rect 21542 31328 21548 31340
rect 21039 31300 21548 31328
rect 21039 31297 21051 31300
rect 20993 31291 21051 31297
rect 21542 31288 21548 31300
rect 21600 31288 21606 31340
rect 21836 31337 21864 31368
rect 22094 31356 22100 31368
rect 22152 31356 22158 31408
rect 22738 31356 22744 31408
rect 22796 31396 22802 31408
rect 24489 31399 24547 31405
rect 24489 31396 24501 31399
rect 22796 31368 24501 31396
rect 22796 31356 22802 31368
rect 24489 31365 24501 31368
rect 24535 31396 24547 31399
rect 24670 31396 24676 31408
rect 24535 31368 24676 31396
rect 24535 31365 24547 31368
rect 24489 31359 24547 31365
rect 24670 31356 24676 31368
rect 24728 31356 24734 31408
rect 28966 31396 28994 31436
rect 29638 31424 29644 31476
rect 29696 31464 29702 31476
rect 30190 31464 30196 31476
rect 29696 31436 30196 31464
rect 29696 31424 29702 31436
rect 30190 31424 30196 31436
rect 30248 31424 30254 31476
rect 32122 31464 32128 31476
rect 30484 31436 32128 31464
rect 30484 31396 30512 31436
rect 32122 31424 32128 31436
rect 32180 31424 32186 31476
rect 31389 31399 31447 31405
rect 31389 31396 31401 31399
rect 28966 31368 30512 31396
rect 30576 31368 31401 31396
rect 30576 31340 30604 31368
rect 31389 31365 31401 31368
rect 31435 31365 31447 31399
rect 31389 31359 31447 31365
rect 21821 31331 21879 31337
rect 21821 31297 21833 31331
rect 21867 31297 21879 31331
rect 21821 31291 21879 31297
rect 22833 31331 22891 31337
rect 22833 31297 22845 31331
rect 22879 31328 22891 31331
rect 22922 31328 22928 31340
rect 22879 31300 22928 31328
rect 22879 31297 22891 31300
rect 22833 31291 22891 31297
rect 22922 31288 22928 31300
rect 22980 31288 22986 31340
rect 23106 31288 23112 31340
rect 23164 31328 23170 31340
rect 23474 31328 23480 31340
rect 23164 31300 23480 31328
rect 23164 31288 23170 31300
rect 23474 31288 23480 31300
rect 23532 31328 23538 31340
rect 23750 31337 23756 31340
rect 23739 31331 23756 31337
rect 23532 31300 23704 31328
rect 23532 31288 23538 31300
rect 21082 31260 21088 31272
rect 19267 31232 21088 31260
rect 21082 31220 21088 31232
rect 21140 31220 21146 31272
rect 21269 31263 21327 31269
rect 21269 31229 21281 31263
rect 21315 31229 21327 31263
rect 21269 31223 21327 31229
rect 20622 31192 20628 31204
rect 19168 31164 20628 31192
rect 18601 31155 18659 31161
rect 20622 31152 20628 31164
rect 20680 31152 20686 31204
rect 20714 31152 20720 31204
rect 20772 31192 20778 31204
rect 21177 31195 21235 31201
rect 21177 31192 21189 31195
rect 20772 31164 21189 31192
rect 20772 31152 20778 31164
rect 21177 31161 21189 31164
rect 21223 31161 21235 31195
rect 21284 31192 21312 31223
rect 21450 31220 21456 31272
rect 21508 31260 21514 31272
rect 22097 31263 22155 31269
rect 22097 31260 22109 31263
rect 21508 31232 22109 31260
rect 21508 31220 21514 31232
rect 22097 31229 22109 31232
rect 22143 31229 22155 31263
rect 23566 31260 23572 31272
rect 22097 31223 22155 31229
rect 22184 31232 23572 31260
rect 21358 31192 21364 31204
rect 21284 31164 21364 31192
rect 21177 31155 21235 31161
rect 21358 31152 21364 31164
rect 21416 31152 21422 31204
rect 21634 31152 21640 31204
rect 21692 31192 21698 31204
rect 22184 31192 22212 31232
rect 23566 31220 23572 31232
rect 23624 31220 23630 31272
rect 23676 31269 23704 31300
rect 23739 31297 23751 31331
rect 23808 31328 23814 31340
rect 24394 31328 24400 31340
rect 23808 31300 24400 31328
rect 23739 31291 23756 31297
rect 23750 31288 23756 31291
rect 23808 31288 23814 31300
rect 24394 31288 24400 31300
rect 24452 31288 24458 31340
rect 24854 31328 24860 31340
rect 24815 31300 24860 31328
rect 24854 31288 24860 31300
rect 24912 31288 24918 31340
rect 25406 31288 25412 31340
rect 25464 31328 25470 31340
rect 25777 31331 25835 31337
rect 25777 31328 25789 31331
rect 25464 31300 25789 31328
rect 25464 31288 25470 31300
rect 25777 31297 25789 31300
rect 25823 31297 25835 31331
rect 30374 31328 30380 31340
rect 30335 31300 30380 31328
rect 25777 31291 25835 31297
rect 30374 31288 30380 31300
rect 30432 31288 30438 31340
rect 30558 31328 30564 31340
rect 30519 31300 30564 31328
rect 30558 31288 30564 31300
rect 30616 31288 30622 31340
rect 30653 31331 30711 31337
rect 30653 31297 30665 31331
rect 30699 31328 30711 31331
rect 30834 31328 30840 31340
rect 30699 31300 30840 31328
rect 30699 31297 30711 31300
rect 30653 31291 30711 31297
rect 30834 31288 30840 31300
rect 30892 31288 30898 31340
rect 31205 31331 31263 31337
rect 31205 31328 31217 31331
rect 30944 31300 31217 31328
rect 23661 31263 23719 31269
rect 23661 31229 23673 31263
rect 23707 31229 23719 31263
rect 23661 31223 23719 31229
rect 23842 31220 23848 31272
rect 23900 31260 23906 31272
rect 24949 31263 25007 31269
rect 24949 31260 24961 31263
rect 23900 31232 24961 31260
rect 23900 31220 23906 31232
rect 24949 31229 24961 31232
rect 24995 31260 25007 31263
rect 25038 31260 25044 31272
rect 24995 31232 25044 31260
rect 24995 31229 25007 31232
rect 24949 31223 25007 31229
rect 25038 31220 25044 31232
rect 25096 31220 25102 31272
rect 25133 31263 25191 31269
rect 25133 31229 25145 31263
rect 25179 31260 25191 31263
rect 25685 31263 25743 31269
rect 25685 31260 25697 31263
rect 25179 31232 25697 31260
rect 25179 31229 25191 31232
rect 25133 31223 25191 31229
rect 25685 31229 25697 31232
rect 25731 31229 25743 31263
rect 27522 31260 27528 31272
rect 27483 31232 27528 31260
rect 25685 31223 25743 31229
rect 27522 31220 27528 31232
rect 27580 31220 27586 31272
rect 27709 31263 27767 31269
rect 27709 31229 27721 31263
rect 27755 31229 27767 31263
rect 27982 31260 27988 31272
rect 27943 31232 27988 31260
rect 27709 31223 27767 31229
rect 22370 31192 22376 31204
rect 21692 31164 22212 31192
rect 22331 31164 22376 31192
rect 21692 31152 21698 31164
rect 22370 31152 22376 31164
rect 22428 31152 22434 31204
rect 22925 31195 22983 31201
rect 22925 31161 22937 31195
rect 22971 31192 22983 31195
rect 27724 31192 27752 31223
rect 27982 31220 27988 31232
rect 28040 31220 28046 31272
rect 29730 31260 29736 31272
rect 28092 31232 29736 31260
rect 22971 31164 27752 31192
rect 22971 31161 22983 31164
rect 22925 31155 22983 31161
rect 18782 31124 18788 31136
rect 17880 31096 18788 31124
rect 17773 31087 17831 31093
rect 18782 31084 18788 31096
rect 18840 31084 18846 31136
rect 18874 31084 18880 31136
rect 18932 31124 18938 31136
rect 19426 31124 19432 31136
rect 18932 31096 19432 31124
rect 18932 31084 18938 31096
rect 19426 31084 19432 31096
rect 19484 31084 19490 31136
rect 19610 31084 19616 31136
rect 19668 31124 19674 31136
rect 19705 31127 19763 31133
rect 19705 31124 19717 31127
rect 19668 31096 19717 31124
rect 19668 31084 19674 31096
rect 19705 31093 19717 31096
rect 19751 31093 19763 31127
rect 19705 31087 19763 31093
rect 21082 31084 21088 31136
rect 21140 31124 21146 31136
rect 21140 31096 21185 31124
rect 21140 31084 21146 31096
rect 21266 31084 21272 31136
rect 21324 31124 21330 31136
rect 22002 31124 22008 31136
rect 21324 31096 22008 31124
rect 21324 31084 21330 31096
rect 22002 31084 22008 31096
rect 22060 31084 22066 31136
rect 22189 31127 22247 31133
rect 22189 31093 22201 31127
rect 22235 31124 22247 31127
rect 23842 31124 23848 31136
rect 22235 31096 23848 31124
rect 22235 31093 22247 31096
rect 22189 31087 22247 31093
rect 23842 31084 23848 31096
rect 23900 31084 23906 31136
rect 23937 31127 23995 31133
rect 23937 31093 23949 31127
rect 23983 31124 23995 31127
rect 24118 31124 24124 31136
rect 23983 31096 24124 31124
rect 23983 31093 23995 31096
rect 23937 31087 23995 31093
rect 24118 31084 24124 31096
rect 24176 31084 24182 31136
rect 24210 31084 24216 31136
rect 24268 31124 24274 31136
rect 26053 31127 26111 31133
rect 26053 31124 26065 31127
rect 24268 31096 26065 31124
rect 24268 31084 24274 31096
rect 26053 31093 26065 31096
rect 26099 31093 26111 31127
rect 26053 31087 26111 31093
rect 26234 31084 26240 31136
rect 26292 31124 26298 31136
rect 27246 31124 27252 31136
rect 26292 31096 27252 31124
rect 26292 31084 26298 31096
rect 27246 31084 27252 31096
rect 27304 31124 27310 31136
rect 28092 31124 28120 31232
rect 29730 31220 29736 31232
rect 29788 31220 29794 31272
rect 30282 31220 30288 31272
rect 30340 31260 30346 31272
rect 30469 31263 30527 31269
rect 30469 31260 30481 31263
rect 30340 31232 30481 31260
rect 30340 31220 30346 31232
rect 30469 31229 30481 31232
rect 30515 31260 30527 31263
rect 30944 31260 30972 31300
rect 31205 31297 31217 31300
rect 31251 31297 31263 31331
rect 34146 31328 34152 31340
rect 34107 31300 34152 31328
rect 31205 31291 31263 31297
rect 34146 31288 34152 31300
rect 34204 31288 34210 31340
rect 31573 31263 31631 31269
rect 31573 31260 31585 31263
rect 30515 31232 30972 31260
rect 31312 31232 31585 31260
rect 30515 31229 30527 31232
rect 30469 31223 30527 31229
rect 30558 31152 30564 31204
rect 30616 31192 30622 31204
rect 31312 31192 31340 31232
rect 31573 31229 31585 31232
rect 31619 31229 31631 31263
rect 32306 31260 32312 31272
rect 32267 31232 32312 31260
rect 31573 31223 31631 31229
rect 32306 31220 32312 31232
rect 32364 31220 32370 31272
rect 32493 31263 32551 31269
rect 32493 31229 32505 31263
rect 32539 31260 32551 31263
rect 34054 31260 34060 31272
rect 32539 31232 34060 31260
rect 32539 31229 32551 31232
rect 32493 31223 32551 31229
rect 34054 31220 34060 31232
rect 34112 31220 34118 31272
rect 30616 31164 31340 31192
rect 30616 31152 30622 31164
rect 27304 31096 28120 31124
rect 27304 31084 27310 31096
rect 28994 31084 29000 31136
rect 29052 31124 29058 31136
rect 31570 31124 31576 31136
rect 29052 31096 31576 31124
rect 29052 31084 29058 31096
rect 31570 31084 31576 31096
rect 31628 31084 31634 31136
rect 1104 31034 34868 31056
rect 1104 30982 6582 31034
rect 6634 30982 6646 31034
rect 6698 30982 6710 31034
rect 6762 30982 6774 31034
rect 6826 30982 6838 31034
rect 6890 30982 17846 31034
rect 17898 30982 17910 31034
rect 17962 30982 17974 31034
rect 18026 30982 18038 31034
rect 18090 30982 18102 31034
rect 18154 30982 29110 31034
rect 29162 30982 29174 31034
rect 29226 30982 29238 31034
rect 29290 30982 29302 31034
rect 29354 30982 29366 31034
rect 29418 30982 34868 31034
rect 1104 30960 34868 30982
rect 1854 30920 1860 30932
rect 1815 30892 1860 30920
rect 1854 30880 1860 30892
rect 1912 30880 1918 30932
rect 12066 30920 12072 30932
rect 12027 30892 12072 30920
rect 12066 30880 12072 30892
rect 12124 30880 12130 30932
rect 13078 30880 13084 30932
rect 13136 30920 13142 30932
rect 13357 30923 13415 30929
rect 13357 30920 13369 30923
rect 13136 30892 13369 30920
rect 13136 30880 13142 30892
rect 13357 30889 13369 30892
rect 13403 30889 13415 30923
rect 13357 30883 13415 30889
rect 13538 30880 13544 30932
rect 13596 30920 13602 30932
rect 15194 30920 15200 30932
rect 13596 30892 15200 30920
rect 13596 30880 13602 30892
rect 15194 30880 15200 30892
rect 15252 30880 15258 30932
rect 15286 30880 15292 30932
rect 15344 30920 15350 30932
rect 15344 30892 15853 30920
rect 15344 30880 15350 30892
rect 12250 30812 12256 30864
rect 12308 30852 12314 30864
rect 12308 30824 15608 30852
rect 12308 30812 12314 30824
rect 12802 30784 12808 30796
rect 12763 30756 12808 30784
rect 12802 30744 12808 30756
rect 12860 30744 12866 30796
rect 15580 30784 15608 30824
rect 15654 30812 15660 30864
rect 15712 30852 15718 30864
rect 15825 30852 15853 30892
rect 15930 30880 15936 30932
rect 15988 30920 15994 30932
rect 15988 30892 18644 30920
rect 15988 30880 15994 30892
rect 17126 30852 17132 30864
rect 15712 30824 15757 30852
rect 15825 30824 17132 30852
rect 15712 30812 15718 30824
rect 17126 30812 17132 30824
rect 17184 30812 17190 30864
rect 18616 30852 18644 30892
rect 18690 30880 18696 30932
rect 18748 30920 18754 30932
rect 23017 30923 23075 30929
rect 23017 30920 23029 30923
rect 18748 30892 18793 30920
rect 19536 30892 23029 30920
rect 18748 30880 18754 30892
rect 19536 30852 19564 30892
rect 23017 30889 23029 30892
rect 23063 30920 23075 30923
rect 24670 30920 24676 30932
rect 23063 30892 24676 30920
rect 23063 30889 23075 30892
rect 23017 30883 23075 30889
rect 24670 30880 24676 30892
rect 24728 30880 24734 30932
rect 25222 30880 25228 30932
rect 25280 30920 25286 30932
rect 27890 30920 27896 30932
rect 25280 30892 27614 30920
rect 27851 30892 27896 30920
rect 25280 30880 25286 30892
rect 18616 30824 19564 30852
rect 20254 30812 20260 30864
rect 20312 30852 20318 30864
rect 21450 30852 21456 30864
rect 20312 30824 21456 30852
rect 20312 30812 20318 30824
rect 21450 30812 21456 30824
rect 21508 30812 21514 30864
rect 23382 30852 23388 30864
rect 21928 30824 23388 30852
rect 15838 30784 15844 30796
rect 12912 30756 15516 30784
rect 15580 30756 15844 30784
rect 1762 30716 1768 30728
rect 1723 30688 1768 30716
rect 1762 30676 1768 30688
rect 1820 30676 1826 30728
rect 11609 30719 11667 30725
rect 11609 30685 11621 30719
rect 11655 30716 11667 30719
rect 11974 30716 11980 30728
rect 11655 30688 11980 30716
rect 11655 30685 11667 30688
rect 11609 30679 11667 30685
rect 11974 30676 11980 30688
rect 12032 30676 12038 30728
rect 12253 30719 12311 30725
rect 12253 30685 12265 30719
rect 12299 30716 12311 30719
rect 12618 30716 12624 30728
rect 12299 30688 12624 30716
rect 12299 30685 12311 30688
rect 12253 30679 12311 30685
rect 12618 30676 12624 30688
rect 12676 30676 12682 30728
rect 12912 30725 12940 30756
rect 12713 30719 12771 30725
rect 12713 30685 12725 30719
rect 12759 30685 12771 30719
rect 12713 30679 12771 30685
rect 12897 30719 12955 30725
rect 12897 30685 12909 30719
rect 12943 30685 12955 30719
rect 12897 30679 12955 30685
rect 12728 30648 12756 30679
rect 12986 30676 12992 30728
rect 13044 30716 13050 30728
rect 13357 30719 13415 30725
rect 13357 30716 13369 30719
rect 13044 30688 13369 30716
rect 13044 30676 13050 30688
rect 13357 30685 13369 30688
rect 13403 30685 13415 30719
rect 13538 30716 13544 30728
rect 13499 30688 13544 30716
rect 13357 30679 13415 30685
rect 13170 30648 13176 30660
rect 12728 30620 13176 30648
rect 13170 30608 13176 30620
rect 13228 30608 13234 30660
rect 13372 30648 13400 30679
rect 13538 30676 13544 30688
rect 13596 30676 13602 30728
rect 14737 30719 14795 30725
rect 14737 30685 14749 30719
rect 14783 30716 14795 30719
rect 15102 30716 15108 30728
rect 14783 30688 15108 30716
rect 14783 30685 14795 30688
rect 14737 30679 14795 30685
rect 15102 30676 15108 30688
rect 15160 30676 15166 30728
rect 15488 30716 15516 30756
rect 15838 30744 15844 30756
rect 15896 30744 15902 30796
rect 16022 30744 16028 30796
rect 16080 30784 16086 30796
rect 16117 30787 16175 30793
rect 16117 30784 16129 30787
rect 16080 30756 16129 30784
rect 16080 30744 16086 30756
rect 16117 30753 16129 30756
rect 16163 30753 16175 30787
rect 16117 30747 16175 30753
rect 16390 30744 16396 30796
rect 16448 30784 16454 30796
rect 17310 30784 17316 30796
rect 16448 30756 16804 30784
rect 17271 30756 17316 30784
rect 16448 30744 16454 30756
rect 15930 30716 15936 30728
rect 15488 30688 15936 30716
rect 15930 30676 15936 30688
rect 15988 30676 15994 30728
rect 16298 30716 16304 30728
rect 16259 30688 16304 30716
rect 16298 30676 16304 30688
rect 16356 30676 16362 30728
rect 16666 30676 16672 30728
rect 16724 30676 16730 30728
rect 16776 30716 16804 30756
rect 17310 30744 17316 30756
rect 17368 30744 17374 30796
rect 19610 30784 19616 30796
rect 18331 30756 19616 30784
rect 16776 30712 17356 30716
rect 17512 30712 17724 30716
rect 16776 30688 17724 30712
rect 17328 30684 17540 30688
rect 14642 30648 14648 30660
rect 13372 30620 14648 30648
rect 14642 30608 14648 30620
rect 14700 30648 14706 30660
rect 14826 30648 14832 30660
rect 14700 30620 14832 30648
rect 14700 30608 14706 30620
rect 14826 30608 14832 30620
rect 14884 30608 14890 30660
rect 14921 30651 14979 30657
rect 14921 30617 14933 30651
rect 14967 30648 14979 30651
rect 15286 30648 15292 30660
rect 14967 30620 15292 30648
rect 14967 30617 14979 30620
rect 14921 30611 14979 30617
rect 15286 30608 15292 30620
rect 15344 30608 15350 30660
rect 15470 30648 15476 30660
rect 15431 30620 15476 30648
rect 15470 30608 15476 30620
rect 15528 30608 15534 30660
rect 15838 30608 15844 30660
rect 15896 30648 15902 30660
rect 16684 30648 16712 30676
rect 17558 30651 17616 30657
rect 17558 30648 17570 30651
rect 15896 30620 16620 30648
rect 16684 30620 17570 30648
rect 15896 30608 15902 30620
rect 14458 30540 14464 30592
rect 14516 30580 14522 30592
rect 16485 30583 16543 30589
rect 16485 30580 16497 30583
rect 14516 30552 16497 30580
rect 14516 30540 14522 30552
rect 16485 30549 16497 30552
rect 16531 30549 16543 30583
rect 16592 30580 16620 30620
rect 17558 30617 17570 30620
rect 17604 30617 17616 30651
rect 17696 30648 17724 30688
rect 18138 30676 18144 30728
rect 18196 30716 18202 30728
rect 18331 30716 18359 30756
rect 19610 30744 19616 30756
rect 19668 30784 19674 30796
rect 19668 30756 20944 30784
rect 19668 30744 19674 30756
rect 18196 30688 18359 30716
rect 18196 30676 18202 30688
rect 18414 30676 18420 30728
rect 18472 30716 18478 30728
rect 18690 30716 18696 30728
rect 18472 30688 18696 30716
rect 18472 30676 18478 30688
rect 18690 30676 18696 30688
rect 18748 30676 18754 30728
rect 18966 30676 18972 30728
rect 19024 30716 19030 30728
rect 19245 30719 19303 30725
rect 19245 30716 19257 30719
rect 19024 30688 19257 30716
rect 19024 30676 19030 30688
rect 19245 30685 19257 30688
rect 19291 30685 19303 30719
rect 19245 30679 19303 30685
rect 19334 30676 19340 30728
rect 19392 30716 19398 30728
rect 19429 30719 19487 30725
rect 19429 30716 19441 30719
rect 19392 30688 19441 30716
rect 19392 30676 19398 30688
rect 19429 30685 19441 30688
rect 19475 30685 19487 30719
rect 19429 30679 19487 30685
rect 19794 30676 19800 30728
rect 19852 30716 19858 30728
rect 20806 30716 20812 30728
rect 19852 30688 20812 30716
rect 19852 30676 19858 30688
rect 20806 30676 20812 30688
rect 20864 30676 20870 30728
rect 20916 30716 20944 30756
rect 20990 30744 20996 30796
rect 21048 30784 21054 30796
rect 21361 30787 21419 30793
rect 21361 30784 21373 30787
rect 21048 30756 21373 30784
rect 21048 30744 21054 30756
rect 21361 30753 21373 30756
rect 21407 30753 21419 30787
rect 21361 30747 21419 30753
rect 21545 30787 21603 30793
rect 21545 30753 21557 30787
rect 21591 30784 21603 30787
rect 21726 30784 21732 30796
rect 21591 30756 21732 30784
rect 21591 30753 21603 30756
rect 21545 30747 21603 30753
rect 21174 30716 21180 30728
rect 20916 30688 21180 30716
rect 21174 30676 21180 30688
rect 21232 30676 21238 30728
rect 21269 30719 21327 30725
rect 21269 30685 21281 30719
rect 21315 30685 21327 30719
rect 21376 30716 21404 30747
rect 21726 30744 21732 30756
rect 21784 30744 21790 30796
rect 21928 30716 21956 30824
rect 23382 30812 23388 30824
rect 23440 30812 23446 30864
rect 25130 30852 25136 30864
rect 25043 30824 25136 30852
rect 25130 30812 25136 30824
rect 25188 30852 25194 30864
rect 25406 30852 25412 30864
rect 25188 30824 25412 30852
rect 25188 30812 25194 30824
rect 25406 30812 25412 30824
rect 25464 30812 25470 30864
rect 25774 30812 25780 30864
rect 25832 30852 25838 30864
rect 25958 30852 25964 30864
rect 25832 30824 25964 30852
rect 25832 30812 25838 30824
rect 25958 30812 25964 30824
rect 26016 30812 26022 30864
rect 27586 30852 27614 30892
rect 27890 30880 27896 30892
rect 27948 30880 27954 30932
rect 28258 30880 28264 30932
rect 28316 30920 28322 30932
rect 30834 30920 30840 30932
rect 28316 30892 30840 30920
rect 28316 30880 28322 30892
rect 30834 30880 30840 30892
rect 30892 30880 30898 30932
rect 33873 30923 33931 30929
rect 33873 30920 33885 30923
rect 31404 30892 33885 30920
rect 28997 30855 29055 30861
rect 28997 30852 29009 30855
rect 27586 30824 29009 30852
rect 28997 30821 29009 30824
rect 29043 30821 29055 30855
rect 28997 30815 29055 30821
rect 22094 30784 22100 30796
rect 22055 30756 22100 30784
rect 22094 30744 22100 30756
rect 22152 30744 22158 30796
rect 22830 30744 22836 30796
rect 22888 30784 22894 30796
rect 23477 30787 23535 30793
rect 23477 30784 23489 30787
rect 22888 30756 23489 30784
rect 22888 30744 22894 30756
rect 23477 30753 23489 30756
rect 23523 30753 23535 30787
rect 23477 30747 23535 30753
rect 23566 30744 23572 30796
rect 23624 30784 23630 30796
rect 24673 30787 24731 30793
rect 24673 30784 24685 30787
rect 23624 30756 24685 30784
rect 23624 30744 23630 30756
rect 24673 30753 24685 30756
rect 24719 30784 24731 30787
rect 25590 30784 25596 30796
rect 24719 30756 25596 30784
rect 24719 30753 24731 30756
rect 24673 30747 24731 30753
rect 25590 30744 25596 30756
rect 25648 30744 25654 30796
rect 26326 30784 26332 30796
rect 25976 30756 26332 30784
rect 21376 30688 21956 30716
rect 21269 30679 21327 30685
rect 19702 30648 19708 30660
rect 17696 30620 19708 30648
rect 17558 30611 17616 30617
rect 19702 30608 19708 30620
rect 19760 30608 19766 30660
rect 20162 30608 20168 30660
rect 20220 30648 20226 30660
rect 20257 30651 20315 30657
rect 20257 30648 20269 30651
rect 20220 30620 20269 30648
rect 20220 30608 20226 30620
rect 20257 30617 20269 30620
rect 20303 30617 20315 30651
rect 20257 30611 20315 30617
rect 20441 30651 20499 30657
rect 20441 30617 20453 30651
rect 20487 30648 20499 30651
rect 21284 30648 21312 30679
rect 22002 30648 22008 30660
rect 20487 30620 21220 30648
rect 21284 30620 22008 30648
rect 20487 30617 20499 30620
rect 20441 30611 20499 30617
rect 19613 30583 19671 30589
rect 19613 30580 19625 30583
rect 16592 30552 19625 30580
rect 16485 30543 16543 30549
rect 19613 30549 19625 30552
rect 19659 30549 19671 30583
rect 20272 30580 20300 30611
rect 20901 30583 20959 30589
rect 20901 30580 20913 30583
rect 20272 30552 20913 30580
rect 19613 30543 19671 30549
rect 20901 30549 20913 30552
rect 20947 30549 20959 30583
rect 21192 30580 21220 30620
rect 22002 30608 22008 30620
rect 22060 30608 22066 30660
rect 22112 30648 22140 30744
rect 22189 30719 22247 30725
rect 22189 30685 22201 30719
rect 22235 30716 22247 30719
rect 22922 30716 22928 30728
rect 22235 30688 22928 30716
rect 22235 30685 22247 30688
rect 22189 30679 22247 30685
rect 22922 30676 22928 30688
rect 22980 30676 22986 30728
rect 23198 30716 23204 30728
rect 23159 30688 23204 30716
rect 23198 30676 23204 30688
rect 23256 30676 23262 30728
rect 23293 30719 23351 30725
rect 23293 30685 23305 30719
rect 23339 30685 23351 30719
rect 23293 30679 23351 30685
rect 23385 30719 23443 30725
rect 23385 30685 23397 30719
rect 23431 30716 23443 30719
rect 24302 30716 24308 30728
rect 23431 30688 24308 30716
rect 23431 30685 23443 30688
rect 23385 30679 23443 30685
rect 22370 30648 22376 30660
rect 22112 30620 22376 30648
rect 22370 30608 22376 30620
rect 22428 30608 22434 30660
rect 23308 30648 23336 30679
rect 24302 30676 24308 30688
rect 24360 30676 24366 30728
rect 24765 30719 24823 30725
rect 24765 30685 24777 30719
rect 24811 30685 24823 30719
rect 24765 30679 24823 30685
rect 22572 30620 23336 30648
rect 24781 30648 24809 30679
rect 24946 30676 24952 30728
rect 25004 30716 25010 30728
rect 25774 30716 25780 30728
rect 25004 30688 25780 30716
rect 25004 30676 25010 30688
rect 25774 30676 25780 30688
rect 25832 30676 25838 30728
rect 25976 30725 26004 30756
rect 26326 30744 26332 30756
rect 26384 30744 26390 30796
rect 28534 30784 28540 30796
rect 28495 30756 28540 30784
rect 28534 30744 28540 30756
rect 28592 30744 28598 30796
rect 29730 30784 29736 30796
rect 28644 30756 29736 30784
rect 25961 30719 26019 30725
rect 25961 30685 25973 30719
rect 26007 30685 26019 30719
rect 25961 30679 26019 30685
rect 26053 30719 26111 30725
rect 26053 30685 26065 30719
rect 26099 30685 26111 30719
rect 26510 30716 26516 30728
rect 26471 30688 26516 30716
rect 26053 30679 26111 30685
rect 25314 30648 25320 30660
rect 24781 30620 25320 30648
rect 22186 30580 22192 30592
rect 21192 30552 22192 30580
rect 20901 30543 20959 30549
rect 22186 30540 22192 30552
rect 22244 30540 22250 30592
rect 22462 30540 22468 30592
rect 22520 30580 22526 30592
rect 22572 30589 22600 30620
rect 25314 30608 25320 30620
rect 25372 30608 25378 30660
rect 25406 30608 25412 30660
rect 25464 30648 25470 30660
rect 26068 30648 26096 30679
rect 26510 30676 26516 30688
rect 26568 30676 26574 30728
rect 26602 30676 26608 30728
rect 26660 30716 26666 30728
rect 26769 30719 26827 30725
rect 26769 30716 26781 30719
rect 26660 30688 26781 30716
rect 26660 30676 26666 30688
rect 26769 30685 26781 30688
rect 26815 30685 26827 30719
rect 26769 30679 26827 30685
rect 27154 30676 27160 30728
rect 27212 30716 27218 30728
rect 28644 30716 28672 30756
rect 29730 30744 29736 30756
rect 29788 30784 29794 30796
rect 30006 30784 30012 30796
rect 29788 30756 30012 30784
rect 29788 30744 29794 30756
rect 30006 30744 30012 30756
rect 30064 30744 30070 30796
rect 31404 30784 31432 30892
rect 33873 30889 33885 30892
rect 33919 30889 33931 30923
rect 33873 30883 33931 30889
rect 31938 30812 31944 30864
rect 31996 30852 32002 30864
rect 31996 30824 33088 30852
rect 31996 30812 32002 30824
rect 31404 30756 31524 30784
rect 31496 30728 31524 30756
rect 32030 30744 32036 30796
rect 32088 30784 32094 30796
rect 32125 30787 32183 30793
rect 32125 30784 32137 30787
rect 32088 30756 32137 30784
rect 32088 30744 32094 30756
rect 32125 30753 32137 30756
rect 32171 30753 32183 30787
rect 32125 30747 32183 30753
rect 32214 30744 32220 30796
rect 32272 30784 32278 30796
rect 32272 30756 32317 30784
rect 32272 30744 32278 30756
rect 28718 30725 28724 30728
rect 27212 30688 28672 30716
rect 28707 30719 28724 30725
rect 27212 30676 27218 30688
rect 28707 30685 28719 30719
rect 28707 30679 28724 30685
rect 28718 30676 28724 30679
rect 28776 30676 28782 30728
rect 30098 30716 30104 30728
rect 30059 30688 30104 30716
rect 30098 30676 30104 30688
rect 30156 30676 30162 30728
rect 31478 30676 31484 30728
rect 31536 30676 31542 30728
rect 31570 30676 31576 30728
rect 31628 30716 31634 30728
rect 31938 30716 31944 30728
rect 31628 30688 31944 30716
rect 31628 30676 31634 30688
rect 31938 30676 31944 30688
rect 31996 30676 32002 30728
rect 32306 30716 32312 30728
rect 32267 30688 32312 30716
rect 32306 30676 32312 30688
rect 32364 30676 32370 30728
rect 32401 30719 32459 30725
rect 32401 30685 32413 30719
rect 32447 30716 32459 30719
rect 32953 30719 33011 30725
rect 32953 30716 32965 30719
rect 32447 30688 32965 30716
rect 32447 30685 32459 30688
rect 32401 30679 32459 30685
rect 32953 30685 32965 30688
rect 32999 30685 33011 30719
rect 33060 30716 33088 30824
rect 33321 30787 33379 30793
rect 33321 30753 33333 30787
rect 33367 30784 33379 30787
rect 33502 30784 33508 30796
rect 33367 30756 33508 30784
rect 33367 30753 33379 30756
rect 33321 30747 33379 30753
rect 33502 30744 33508 30756
rect 33560 30784 33566 30796
rect 34238 30784 34244 30796
rect 33560 30756 34244 30784
rect 33560 30744 33566 30756
rect 34238 30744 34244 30756
rect 34296 30744 34302 30796
rect 33137 30719 33195 30725
rect 33137 30716 33149 30719
rect 33060 30688 33149 30716
rect 32953 30679 33011 30685
rect 33137 30685 33149 30688
rect 33183 30685 33195 30719
rect 33137 30679 33195 30685
rect 33413 30719 33471 30725
rect 33413 30685 33425 30719
rect 33459 30685 33471 30719
rect 33870 30716 33876 30728
rect 33831 30688 33876 30716
rect 33413 30679 33471 30685
rect 27798 30648 27804 30660
rect 25464 30620 27804 30648
rect 25464 30608 25470 30620
rect 27798 30608 27804 30620
rect 27856 30608 27862 30660
rect 27890 30608 27896 30660
rect 27948 30648 27954 30660
rect 28902 30648 28908 30660
rect 27948 30620 28908 30648
rect 27948 30608 27954 30620
rect 28902 30608 28908 30620
rect 28960 30608 28966 30660
rect 29638 30608 29644 30660
rect 29696 30648 29702 30660
rect 30346 30651 30404 30657
rect 30346 30648 30358 30651
rect 29696 30620 30358 30648
rect 29696 30608 29702 30620
rect 30346 30617 30358 30620
rect 30392 30617 30404 30651
rect 30346 30611 30404 30617
rect 30484 30620 32076 30648
rect 22557 30583 22615 30589
rect 22557 30580 22569 30583
rect 22520 30552 22569 30580
rect 22520 30540 22526 30552
rect 22557 30549 22569 30552
rect 22603 30549 22615 30583
rect 22557 30543 22615 30549
rect 22830 30540 22836 30592
rect 22888 30580 22894 30592
rect 24394 30580 24400 30592
rect 22888 30552 24400 30580
rect 22888 30540 22894 30552
rect 24394 30540 24400 30552
rect 24452 30540 24458 30592
rect 25593 30583 25651 30589
rect 25593 30549 25605 30583
rect 25639 30580 25651 30583
rect 27338 30580 27344 30592
rect 25639 30552 27344 30580
rect 25639 30549 25651 30552
rect 25593 30543 25651 30549
rect 27338 30540 27344 30552
rect 27396 30540 27402 30592
rect 27982 30540 27988 30592
rect 28040 30580 28046 30592
rect 30484 30580 30512 30620
rect 28040 30552 30512 30580
rect 28040 30540 28046 30552
rect 30650 30540 30656 30592
rect 30708 30580 30714 30592
rect 31018 30580 31024 30592
rect 30708 30552 31024 30580
rect 30708 30540 30714 30552
rect 31018 30540 31024 30552
rect 31076 30580 31082 30592
rect 31481 30583 31539 30589
rect 31481 30580 31493 30583
rect 31076 30552 31493 30580
rect 31076 30540 31082 30552
rect 31481 30549 31493 30552
rect 31527 30549 31539 30583
rect 31938 30580 31944 30592
rect 31899 30552 31944 30580
rect 31481 30543 31539 30549
rect 31938 30540 31944 30552
rect 31996 30540 32002 30592
rect 32048 30580 32076 30620
rect 33042 30608 33048 30660
rect 33100 30648 33106 30660
rect 33428 30648 33456 30679
rect 33870 30676 33876 30688
rect 33928 30676 33934 30728
rect 33962 30676 33968 30728
rect 34020 30716 34026 30728
rect 34149 30719 34207 30725
rect 34149 30716 34161 30719
rect 34020 30688 34161 30716
rect 34020 30676 34026 30688
rect 34149 30685 34161 30688
rect 34195 30685 34207 30719
rect 34149 30679 34207 30685
rect 33100 30620 33456 30648
rect 33100 30608 33106 30620
rect 34057 30583 34115 30589
rect 34057 30580 34069 30583
rect 32048 30552 34069 30580
rect 34057 30549 34069 30552
rect 34103 30549 34115 30583
rect 34057 30543 34115 30549
rect 1104 30490 34868 30512
rect 1104 30438 12214 30490
rect 12266 30438 12278 30490
rect 12330 30438 12342 30490
rect 12394 30438 12406 30490
rect 12458 30438 12470 30490
rect 12522 30438 23478 30490
rect 23530 30438 23542 30490
rect 23594 30438 23606 30490
rect 23658 30438 23670 30490
rect 23722 30438 23734 30490
rect 23786 30438 34868 30490
rect 1104 30416 34868 30438
rect 13814 30336 13820 30388
rect 13872 30376 13878 30388
rect 16942 30376 16948 30388
rect 13872 30348 16948 30376
rect 13872 30336 13878 30348
rect 16942 30336 16948 30348
rect 17000 30336 17006 30388
rect 17043 30379 17101 30385
rect 17043 30345 17055 30379
rect 17089 30376 17101 30379
rect 17678 30376 17684 30388
rect 17089 30348 17684 30376
rect 17089 30345 17101 30348
rect 17043 30339 17101 30345
rect 17678 30336 17684 30348
rect 17736 30336 17742 30388
rect 20990 30376 20996 30388
rect 17781 30348 20996 30376
rect 14826 30308 14832 30320
rect 12544 30280 14832 30308
rect 11790 30200 11796 30252
rect 11848 30240 11854 30252
rect 11885 30243 11943 30249
rect 11885 30240 11897 30243
rect 11848 30212 11897 30240
rect 11848 30200 11854 30212
rect 11885 30209 11897 30212
rect 11931 30209 11943 30243
rect 11885 30203 11943 30209
rect 12069 30243 12127 30249
rect 12069 30209 12081 30243
rect 12115 30240 12127 30243
rect 12434 30240 12440 30252
rect 12115 30212 12440 30240
rect 12115 30209 12127 30212
rect 12069 30203 12127 30209
rect 12434 30200 12440 30212
rect 12492 30200 12498 30252
rect 12544 30249 12572 30280
rect 14826 30268 14832 30280
rect 14884 30268 14890 30320
rect 15197 30311 15255 30317
rect 15197 30277 15209 30311
rect 15243 30308 15255 30311
rect 15470 30308 15476 30320
rect 15243 30280 15476 30308
rect 15243 30277 15255 30280
rect 15197 30271 15255 30277
rect 15470 30268 15476 30280
rect 15528 30308 15534 30320
rect 16117 30311 16175 30317
rect 16117 30308 16129 30311
rect 15528 30280 16129 30308
rect 15528 30268 15534 30280
rect 16117 30277 16129 30280
rect 16163 30277 16175 30311
rect 16117 30271 16175 30277
rect 16574 30268 16580 30320
rect 16632 30308 16638 30320
rect 17781 30308 17809 30348
rect 20990 30336 20996 30348
rect 21048 30336 21054 30388
rect 21100 30348 21576 30376
rect 18414 30308 18420 30320
rect 16632 30280 17809 30308
rect 17880 30280 18420 30308
rect 16632 30268 16638 30280
rect 12529 30243 12587 30249
rect 12529 30209 12541 30243
rect 12575 30209 12587 30243
rect 12529 30203 12587 30209
rect 12618 30200 12624 30252
rect 12676 30240 12682 30252
rect 12713 30243 12771 30249
rect 12713 30240 12725 30243
rect 12676 30212 12725 30240
rect 12676 30200 12682 30212
rect 12713 30209 12725 30212
rect 12759 30240 12771 30243
rect 12802 30240 12808 30252
rect 12759 30212 12808 30240
rect 12759 30209 12771 30212
rect 12713 30203 12771 30209
rect 12802 30200 12808 30212
rect 12860 30200 12866 30252
rect 13173 30243 13231 30249
rect 13173 30209 13185 30243
rect 13219 30240 13231 30243
rect 13262 30240 13268 30252
rect 13219 30212 13268 30240
rect 13219 30209 13231 30212
rect 13173 30203 13231 30209
rect 13262 30200 13268 30212
rect 13320 30200 13326 30252
rect 13357 30243 13415 30249
rect 13357 30209 13369 30243
rect 13403 30240 13415 30243
rect 13722 30240 13728 30252
rect 13403 30212 13728 30240
rect 13403 30209 13415 30212
rect 13357 30203 13415 30209
rect 13722 30200 13728 30212
rect 13780 30200 13786 30252
rect 13817 30243 13875 30249
rect 13817 30209 13829 30243
rect 13863 30240 13875 30243
rect 14274 30240 14280 30252
rect 13863 30212 14280 30240
rect 13863 30209 13875 30212
rect 13817 30203 13875 30209
rect 14274 30200 14280 30212
rect 14332 30200 14338 30252
rect 14461 30243 14519 30249
rect 14461 30209 14473 30243
rect 14507 30240 14519 30243
rect 14550 30240 14556 30252
rect 14507 30212 14556 30240
rect 14507 30209 14519 30212
rect 14461 30203 14519 30209
rect 14550 30200 14556 30212
rect 14608 30200 14614 30252
rect 15102 30200 15108 30252
rect 15160 30240 15166 30252
rect 15381 30243 15439 30249
rect 15381 30240 15393 30243
rect 15160 30212 15393 30240
rect 15160 30200 15166 30212
rect 15381 30209 15393 30212
rect 15427 30209 15439 30243
rect 15381 30203 15439 30209
rect 15838 30200 15844 30252
rect 15896 30240 15902 30252
rect 15933 30243 15991 30249
rect 15933 30240 15945 30243
rect 15896 30212 15945 30240
rect 15896 30200 15902 30212
rect 15933 30209 15945 30212
rect 15979 30209 15991 30243
rect 15933 30203 15991 30209
rect 16022 30200 16028 30252
rect 16080 30240 16086 30252
rect 16298 30240 16304 30252
rect 16080 30212 16304 30240
rect 16080 30200 16086 30212
rect 16298 30200 16304 30212
rect 16356 30200 16362 30252
rect 16850 30200 16856 30252
rect 16908 30240 16914 30252
rect 16945 30243 17003 30249
rect 16945 30240 16957 30243
rect 16908 30212 16957 30240
rect 16908 30200 16914 30212
rect 16945 30209 16957 30212
rect 16991 30209 17003 30243
rect 17126 30240 17132 30252
rect 17087 30212 17132 30240
rect 16945 30203 17003 30209
rect 17126 30200 17132 30212
rect 17184 30200 17190 30252
rect 17236 30249 17264 30280
rect 17221 30243 17279 30249
rect 17221 30209 17233 30243
rect 17267 30209 17279 30243
rect 17221 30203 17279 30209
rect 17310 30200 17316 30252
rect 17368 30240 17374 30252
rect 17586 30240 17592 30252
rect 17368 30212 17592 30240
rect 17368 30200 17374 30212
rect 17586 30200 17592 30212
rect 17644 30200 17650 30252
rect 17681 30243 17739 30249
rect 17681 30209 17693 30243
rect 17727 30240 17739 30243
rect 17880 30240 17908 30280
rect 18414 30268 18420 30280
rect 18472 30308 18478 30320
rect 19788 30311 19846 30317
rect 18472 30280 19288 30308
rect 18472 30268 18478 30280
rect 19260 30252 19288 30280
rect 19788 30277 19800 30311
rect 19834 30308 19846 30311
rect 21100 30308 21128 30348
rect 19834 30280 21128 30308
rect 21548 30308 21576 30348
rect 21726 30336 21732 30388
rect 21784 30376 21790 30388
rect 21784 30348 22324 30376
rect 21784 30336 21790 30348
rect 21821 30311 21879 30317
rect 21821 30308 21833 30311
rect 21548 30280 21833 30308
rect 19834 30277 19846 30280
rect 19788 30271 19846 30277
rect 21821 30277 21833 30280
rect 21867 30277 21879 30311
rect 21821 30271 21879 30277
rect 17954 30249 17960 30252
rect 17727 30212 17908 30240
rect 17937 30243 17960 30249
rect 17727 30209 17739 30212
rect 17681 30203 17739 30209
rect 17937 30209 17949 30243
rect 17937 30203 17960 30209
rect 17954 30200 17960 30203
rect 18012 30200 18018 30252
rect 18322 30200 18328 30252
rect 18380 30240 18386 30252
rect 18380 30212 18722 30240
rect 18380 30200 18386 30212
rect 11977 30175 12035 30181
rect 11977 30141 11989 30175
rect 12023 30172 12035 30175
rect 18694 30172 18722 30212
rect 19242 30200 19248 30252
rect 19300 30240 19306 30252
rect 19518 30240 19524 30252
rect 19300 30212 19524 30240
rect 19300 30200 19306 30212
rect 19518 30200 19524 30212
rect 19576 30200 19582 30252
rect 20254 30240 20260 30252
rect 19628 30212 20260 30240
rect 19628 30172 19656 30212
rect 20254 30200 20260 30212
rect 20312 30200 20318 30252
rect 20530 30200 20536 30252
rect 20588 30240 20594 30252
rect 22051 30243 22109 30249
rect 22051 30240 22063 30243
rect 20588 30212 22063 30240
rect 20588 30200 20594 30212
rect 22051 30209 22063 30212
rect 22097 30209 22109 30243
rect 22051 30203 22109 30209
rect 12023 30144 17632 30172
rect 18694 30144 19656 30172
rect 12023 30141 12035 30144
rect 11977 30135 12035 30141
rect 12621 30107 12679 30113
rect 12621 30073 12633 30107
rect 12667 30104 12679 30107
rect 17034 30104 17040 30116
rect 12667 30076 17040 30104
rect 12667 30073 12679 30076
rect 12621 30067 12679 30073
rect 17034 30064 17040 30076
rect 17092 30064 17098 30116
rect 17494 30064 17500 30116
rect 17552 30064 17558 30116
rect 13170 29996 13176 30048
rect 13228 30036 13234 30048
rect 13265 30039 13323 30045
rect 13265 30036 13277 30039
rect 13228 30008 13277 30036
rect 13228 29996 13234 30008
rect 13265 30005 13277 30008
rect 13311 30005 13323 30039
rect 13265 29999 13323 30005
rect 13909 30039 13967 30045
rect 13909 30005 13921 30039
rect 13955 30036 13967 30039
rect 14182 30036 14188 30048
rect 13955 30008 14188 30036
rect 13955 30005 13967 30008
rect 13909 29999 13967 30005
rect 14182 29996 14188 30008
rect 14240 29996 14246 30048
rect 14553 30039 14611 30045
rect 14553 30005 14565 30039
rect 14599 30036 14611 30039
rect 14918 30036 14924 30048
rect 14599 30008 14924 30036
rect 14599 30005 14611 30008
rect 14553 29999 14611 30005
rect 14918 29996 14924 30008
rect 14976 29996 14982 30048
rect 15470 29996 15476 30048
rect 15528 30036 15534 30048
rect 16206 30036 16212 30048
rect 15528 30008 16212 30036
rect 15528 29996 15534 30008
rect 16206 29996 16212 30008
rect 16264 29996 16270 30048
rect 16298 29996 16304 30048
rect 16356 30036 16362 30048
rect 17512 30036 17540 30064
rect 16356 30008 17540 30036
rect 17604 30036 17632 30144
rect 20990 30132 20996 30184
rect 21048 30172 21054 30184
rect 22066 30172 22094 30203
rect 22167 30200 22173 30252
rect 22225 30246 22244 30252
rect 22296 30249 22324 30348
rect 22370 30336 22376 30388
rect 22428 30376 22434 30388
rect 30006 30376 30012 30388
rect 22428 30348 22968 30376
rect 22428 30336 22434 30348
rect 22554 30268 22560 30320
rect 22612 30308 22618 30320
rect 22738 30308 22744 30320
rect 22612 30280 22744 30308
rect 22612 30268 22618 30280
rect 22738 30268 22744 30280
rect 22796 30268 22802 30320
rect 22232 30212 22244 30246
rect 22225 30206 22244 30212
rect 22281 30243 22339 30249
rect 22281 30209 22293 30243
rect 22327 30209 22339 30243
rect 22225 30200 22231 30206
rect 22281 30203 22339 30209
rect 22465 30243 22523 30249
rect 22465 30209 22477 30243
rect 22511 30240 22523 30243
rect 22646 30240 22652 30252
rect 22511 30212 22652 30240
rect 22511 30209 22523 30212
rect 22465 30203 22523 30209
rect 22646 30200 22652 30212
rect 22704 30200 22710 30252
rect 22830 30172 22836 30184
rect 21048 30144 21833 30172
rect 22066 30144 22836 30172
rect 21048 30132 21054 30144
rect 21805 30104 21833 30144
rect 22830 30132 22836 30144
rect 22888 30132 22894 30184
rect 22940 30172 22968 30348
rect 23584 30348 30012 30376
rect 23109 30243 23167 30249
rect 23109 30209 23121 30243
rect 23155 30240 23167 30243
rect 23474 30240 23480 30252
rect 23155 30212 23480 30240
rect 23155 30209 23167 30212
rect 23109 30203 23167 30209
rect 23474 30200 23480 30212
rect 23532 30200 23538 30252
rect 23017 30175 23075 30181
rect 23017 30172 23029 30175
rect 22940 30144 23029 30172
rect 23017 30141 23029 30144
rect 23063 30141 23075 30175
rect 23584 30172 23612 30348
rect 25130 30308 25136 30320
rect 24781 30280 25136 30308
rect 23934 30240 23940 30252
rect 23895 30212 23940 30240
rect 23934 30200 23940 30212
rect 23992 30200 23998 30252
rect 24118 30200 24124 30252
rect 24176 30240 24182 30252
rect 24781 30249 24809 30280
rect 25130 30268 25136 30280
rect 25188 30268 25194 30320
rect 25774 30268 25780 30320
rect 25832 30308 25838 30320
rect 27448 30317 27476 30348
rect 30006 30336 30012 30348
rect 30064 30336 30070 30388
rect 30558 30376 30564 30388
rect 30208 30348 30564 30376
rect 26421 30311 26479 30317
rect 26421 30308 26433 30311
rect 25832 30280 26433 30308
rect 25832 30268 25838 30280
rect 26421 30277 26433 30280
rect 26467 30277 26479 30311
rect 26421 30271 26479 30277
rect 27433 30311 27491 30317
rect 27433 30277 27445 30311
rect 27479 30277 27491 30311
rect 28994 30308 29000 30320
rect 27433 30271 27491 30277
rect 27540 30280 29000 30308
rect 24765 30243 24823 30249
rect 24176 30212 24716 30240
rect 24176 30200 24182 30212
rect 23017 30135 23075 30141
rect 23121 30144 23612 30172
rect 24688 30172 24716 30212
rect 24765 30209 24777 30243
rect 24811 30209 24823 30243
rect 24765 30203 24823 30209
rect 25041 30243 25099 30249
rect 25041 30209 25053 30243
rect 25087 30240 25099 30243
rect 25498 30240 25504 30252
rect 25087 30212 25504 30240
rect 25087 30209 25099 30212
rect 25041 30203 25099 30209
rect 25498 30200 25504 30212
rect 25556 30200 25562 30252
rect 25590 30200 25596 30252
rect 25648 30240 25654 30252
rect 27540 30249 27568 30280
rect 28994 30268 29000 30280
rect 29052 30268 29058 30320
rect 29638 30268 29644 30320
rect 29696 30308 29702 30320
rect 29917 30311 29975 30317
rect 29917 30308 29929 30311
rect 29696 30280 29929 30308
rect 29696 30268 29702 30280
rect 29917 30277 29929 30280
rect 29963 30277 29975 30311
rect 29917 30271 29975 30277
rect 28258 30249 28264 30252
rect 26237 30243 26295 30249
rect 26237 30240 26249 30243
rect 25648 30212 26249 30240
rect 25648 30200 25654 30212
rect 26237 30209 26249 30212
rect 26283 30209 26295 30243
rect 27249 30243 27307 30249
rect 27249 30240 27261 30243
rect 26237 30203 26295 30209
rect 26344 30212 27261 30240
rect 24857 30175 24915 30181
rect 24857 30172 24869 30175
rect 24688 30144 24869 30172
rect 23121 30104 23149 30144
rect 24857 30141 24869 30144
rect 24903 30141 24915 30175
rect 24857 30135 24915 30141
rect 24946 30132 24952 30184
rect 25004 30172 25010 30184
rect 26050 30172 26056 30184
rect 25004 30144 25049 30172
rect 26011 30144 26056 30172
rect 25004 30132 25010 30144
rect 26050 30132 26056 30144
rect 26108 30132 26114 30184
rect 18616 30076 19196 30104
rect 18616 30036 18644 30076
rect 17604 30008 18644 30036
rect 16356 29996 16362 30008
rect 18690 29996 18696 30048
rect 18748 30036 18754 30048
rect 19061 30039 19119 30045
rect 19061 30036 19073 30039
rect 18748 30008 19073 30036
rect 18748 29996 18754 30008
rect 19061 30005 19073 30008
rect 19107 30005 19119 30039
rect 19168 30036 19196 30076
rect 20456 30076 21036 30104
rect 21805 30076 23149 30104
rect 20456 30036 20484 30076
rect 19168 30008 20484 30036
rect 19061 29999 19119 30005
rect 20530 29996 20536 30048
rect 20588 30036 20594 30048
rect 20901 30039 20959 30045
rect 20901 30036 20913 30039
rect 20588 30008 20913 30036
rect 20588 29996 20594 30008
rect 20901 30005 20913 30008
rect 20947 30005 20959 30039
rect 21008 30036 21036 30076
rect 23290 30064 23296 30116
rect 23348 30104 23354 30116
rect 23477 30107 23535 30113
rect 23477 30104 23489 30107
rect 23348 30076 23489 30104
rect 23348 30064 23354 30076
rect 23477 30073 23489 30076
rect 23523 30073 23535 30107
rect 23477 30067 23535 30073
rect 24581 30107 24639 30113
rect 24581 30073 24593 30107
rect 24627 30104 24639 30107
rect 25406 30104 25412 30116
rect 24627 30076 25412 30104
rect 24627 30073 24639 30076
rect 24581 30067 24639 30073
rect 25406 30064 25412 30076
rect 25464 30064 25470 30116
rect 25866 30064 25872 30116
rect 25924 30104 25930 30116
rect 26344 30104 26372 30212
rect 27249 30209 27261 30212
rect 27295 30209 27307 30243
rect 27249 30203 27307 30209
rect 27525 30243 27583 30249
rect 27525 30209 27537 30243
rect 27571 30209 27583 30243
rect 27525 30203 27583 30209
rect 28252 30203 28264 30249
rect 28316 30240 28322 30252
rect 28316 30212 28352 30240
rect 28258 30200 28264 30203
rect 28316 30200 28322 30212
rect 28534 30200 28540 30252
rect 28592 30240 28598 30252
rect 30208 30249 30236 30348
rect 30558 30336 30564 30348
rect 30616 30336 30622 30388
rect 30650 30336 30656 30388
rect 30708 30376 30714 30388
rect 31363 30379 31421 30385
rect 31363 30376 31375 30379
rect 30708 30348 31375 30376
rect 30708 30336 30714 30348
rect 31363 30345 31375 30348
rect 31409 30345 31421 30379
rect 31363 30339 31421 30345
rect 30742 30308 30748 30320
rect 30570 30280 30748 30308
rect 30193 30243 30251 30249
rect 28592 30212 29500 30240
rect 28592 30200 28598 30212
rect 26510 30132 26516 30184
rect 26568 30172 26574 30184
rect 27154 30172 27160 30184
rect 26568 30144 27160 30172
rect 26568 30132 26574 30144
rect 27154 30132 27160 30144
rect 27212 30172 27218 30184
rect 27985 30175 28043 30181
rect 27985 30172 27997 30175
rect 27212 30144 27997 30172
rect 27212 30132 27218 30144
rect 27985 30141 27997 30144
rect 28031 30141 28043 30175
rect 27985 30135 28043 30141
rect 27890 30104 27896 30116
rect 25924 30076 26372 30104
rect 26528 30076 27896 30104
rect 25924 30064 25930 30076
rect 23934 30036 23940 30048
rect 21008 30008 23940 30036
rect 20901 29999 20959 30005
rect 23934 29996 23940 30008
rect 23992 29996 23998 30048
rect 24029 30039 24087 30045
rect 24029 30005 24041 30039
rect 24075 30036 24087 30039
rect 26528 30036 26556 30076
rect 27890 30064 27896 30076
rect 27948 30064 27954 30116
rect 28994 30064 29000 30116
rect 29052 30104 29058 30116
rect 29365 30107 29423 30113
rect 29365 30104 29377 30107
rect 29052 30076 29377 30104
rect 29052 30064 29058 30076
rect 29365 30073 29377 30076
rect 29411 30073 29423 30107
rect 29472 30104 29500 30212
rect 30193 30209 30205 30243
rect 30239 30209 30251 30243
rect 30193 30203 30251 30209
rect 30282 30243 30340 30249
rect 30282 30209 30294 30243
rect 30328 30209 30340 30243
rect 30282 30203 30340 30209
rect 30398 30246 30456 30252
rect 30570 30249 30598 30280
rect 30742 30268 30748 30280
rect 30800 30268 30806 30320
rect 30834 30268 30840 30320
rect 30892 30308 30898 30320
rect 31573 30311 31631 30317
rect 31573 30308 31585 30311
rect 30892 30280 31585 30308
rect 30892 30268 30898 30280
rect 31573 30277 31585 30280
rect 31619 30277 31631 30311
rect 31573 30271 31631 30277
rect 31662 30268 31668 30320
rect 31720 30308 31726 30320
rect 33870 30308 33876 30320
rect 31720 30280 33876 30308
rect 31720 30268 31726 30280
rect 33870 30268 33876 30280
rect 33928 30268 33934 30320
rect 30398 30212 30410 30246
rect 30444 30243 30456 30246
rect 30561 30243 30619 30249
rect 30444 30215 30512 30243
rect 30444 30212 30456 30215
rect 30398 30206 30456 30212
rect 30297 30116 30325 30203
rect 30484 30172 30512 30215
rect 30561 30209 30573 30243
rect 30607 30209 30619 30243
rect 30561 30203 30619 30209
rect 30650 30200 30656 30252
rect 30708 30240 30714 30252
rect 32493 30243 32551 30249
rect 32493 30240 32505 30243
rect 30708 30212 32505 30240
rect 30708 30200 30714 30212
rect 32493 30209 32505 30212
rect 32539 30209 32551 30243
rect 32493 30203 32551 30209
rect 33134 30200 33140 30252
rect 33192 30240 33198 30252
rect 33505 30243 33563 30249
rect 33505 30240 33517 30243
rect 33192 30212 33517 30240
rect 33192 30200 33198 30212
rect 33505 30209 33517 30212
rect 33551 30209 33563 30243
rect 33778 30240 33784 30252
rect 33739 30212 33784 30240
rect 33505 30203 33563 30209
rect 33778 30200 33784 30212
rect 33836 30200 33842 30252
rect 31846 30172 31852 30184
rect 30484 30144 31852 30172
rect 31846 30132 31852 30144
rect 31904 30132 31910 30184
rect 31938 30132 31944 30184
rect 31996 30172 32002 30184
rect 32401 30175 32459 30181
rect 32401 30172 32413 30175
rect 31996 30144 32413 30172
rect 31996 30132 32002 30144
rect 32401 30141 32413 30144
rect 32447 30141 32459 30175
rect 32401 30135 32459 30141
rect 29638 30104 29644 30116
rect 29472 30076 29644 30104
rect 29365 30067 29423 30073
rect 29638 30064 29644 30076
rect 29696 30064 29702 30116
rect 30282 30064 30288 30116
rect 30340 30064 30346 30116
rect 31202 30104 31208 30116
rect 31163 30076 31208 30104
rect 31202 30064 31208 30076
rect 31260 30064 31266 30116
rect 24075 30008 26556 30036
rect 27065 30039 27123 30045
rect 24075 30005 24087 30008
rect 24029 29999 24087 30005
rect 27065 30005 27077 30039
rect 27111 30036 27123 30039
rect 30374 30036 30380 30048
rect 27111 30008 30380 30036
rect 27111 30005 27123 30008
rect 27065 29999 27123 30005
rect 30374 29996 30380 30008
rect 30432 29996 30438 30048
rect 30834 30036 30840 30048
rect 30795 30008 30840 30036
rect 30834 29996 30840 30008
rect 30892 29996 30898 30048
rect 31294 29996 31300 30048
rect 31352 30036 31358 30048
rect 31389 30039 31447 30045
rect 31389 30036 31401 30039
rect 31352 30008 31401 30036
rect 31352 29996 31358 30008
rect 31389 30005 31401 30008
rect 31435 30005 31447 30039
rect 31389 29999 31447 30005
rect 31478 29996 31484 30048
rect 31536 30036 31542 30048
rect 32769 30039 32827 30045
rect 32769 30036 32781 30039
rect 31536 30008 32781 30036
rect 31536 29996 31542 30008
rect 32769 30005 32781 30008
rect 32815 30005 32827 30039
rect 32769 29999 32827 30005
rect 33134 29996 33140 30048
rect 33192 30036 33198 30048
rect 33321 30039 33379 30045
rect 33321 30036 33333 30039
rect 33192 30008 33333 30036
rect 33192 29996 33198 30008
rect 33321 30005 33333 30008
rect 33367 30005 33379 30039
rect 33321 29999 33379 30005
rect 33410 29996 33416 30048
rect 33468 30036 33474 30048
rect 33689 30039 33747 30045
rect 33689 30036 33701 30039
rect 33468 30008 33701 30036
rect 33468 29996 33474 30008
rect 33689 30005 33701 30008
rect 33735 30005 33747 30039
rect 33689 29999 33747 30005
rect 1104 29946 34868 29968
rect 1104 29894 6582 29946
rect 6634 29894 6646 29946
rect 6698 29894 6710 29946
rect 6762 29894 6774 29946
rect 6826 29894 6838 29946
rect 6890 29894 17846 29946
rect 17898 29894 17910 29946
rect 17962 29894 17974 29946
rect 18026 29894 18038 29946
rect 18090 29894 18102 29946
rect 18154 29894 29110 29946
rect 29162 29894 29174 29946
rect 29226 29894 29238 29946
rect 29290 29894 29302 29946
rect 29354 29894 29366 29946
rect 29418 29894 34868 29946
rect 1104 29872 34868 29894
rect 15286 29792 15292 29844
rect 15344 29832 15350 29844
rect 20438 29832 20444 29844
rect 15344 29804 20444 29832
rect 15344 29792 15350 29804
rect 20438 29792 20444 29804
rect 20496 29792 20502 29844
rect 22830 29832 22836 29844
rect 20548 29804 22600 29832
rect 22791 29804 22836 29832
rect 11790 29724 11796 29776
rect 11848 29764 11854 29776
rect 15930 29764 15936 29776
rect 11848 29736 15936 29764
rect 11848 29724 11854 29736
rect 15930 29724 15936 29736
rect 15988 29724 15994 29776
rect 16022 29724 16028 29776
rect 16080 29724 16086 29776
rect 17034 29724 17040 29776
rect 17092 29764 17098 29776
rect 19426 29764 19432 29776
rect 17092 29736 19432 29764
rect 17092 29724 17098 29736
rect 19426 29724 19432 29736
rect 19484 29724 19490 29776
rect 12805 29699 12863 29705
rect 12805 29665 12817 29699
rect 12851 29696 12863 29699
rect 16040 29696 16068 29724
rect 12851 29668 16068 29696
rect 12851 29665 12863 29668
rect 12805 29659 12863 29665
rect 17126 29656 17132 29708
rect 17184 29696 17190 29708
rect 19518 29696 19524 29708
rect 17184 29668 19222 29696
rect 19479 29668 19524 29696
rect 17184 29656 17190 29668
rect 11882 29588 11888 29640
rect 11940 29628 11946 29640
rect 12253 29631 12311 29637
rect 12253 29628 12265 29631
rect 11940 29600 12265 29628
rect 11940 29588 11946 29600
rect 12253 29597 12265 29600
rect 12299 29597 12311 29631
rect 12710 29628 12716 29640
rect 12671 29600 12716 29628
rect 12253 29591 12311 29597
rect 12710 29588 12716 29600
rect 12768 29588 12774 29640
rect 12894 29628 12900 29640
rect 12855 29600 12900 29628
rect 12894 29588 12900 29600
rect 12952 29588 12958 29640
rect 13354 29628 13360 29640
rect 13315 29600 13360 29628
rect 13354 29588 13360 29600
rect 13412 29588 13418 29640
rect 13541 29631 13599 29637
rect 13541 29597 13553 29631
rect 13587 29628 13599 29631
rect 13998 29628 14004 29640
rect 13587 29600 14004 29628
rect 13587 29597 13599 29600
rect 13541 29591 13599 29597
rect 13998 29588 14004 29600
rect 14056 29588 14062 29640
rect 14093 29631 14151 29637
rect 14093 29597 14105 29631
rect 14139 29628 14151 29631
rect 14182 29628 14188 29640
rect 14139 29600 14188 29628
rect 14139 29597 14151 29600
rect 14093 29591 14151 29597
rect 14182 29588 14188 29600
rect 14240 29588 14246 29640
rect 14277 29631 14335 29637
rect 14277 29597 14289 29631
rect 14323 29628 14335 29631
rect 14366 29628 14372 29640
rect 14323 29600 14372 29628
rect 14323 29597 14335 29600
rect 14277 29591 14335 29597
rect 14366 29588 14372 29600
rect 14424 29588 14430 29640
rect 14737 29631 14795 29637
rect 14737 29597 14749 29631
rect 14783 29628 14795 29631
rect 14826 29628 14832 29640
rect 14783 29600 14832 29628
rect 14783 29597 14795 29600
rect 14737 29591 14795 29597
rect 14826 29588 14832 29600
rect 14884 29588 14890 29640
rect 15378 29628 15384 29640
rect 15339 29600 15384 29628
rect 15378 29588 15384 29600
rect 15436 29588 15442 29640
rect 15470 29588 15476 29640
rect 15528 29628 15534 29640
rect 15528 29600 15573 29628
rect 15528 29588 15534 29600
rect 15746 29588 15752 29640
rect 15804 29628 15810 29640
rect 15930 29628 15936 29640
rect 15804 29600 15936 29628
rect 15804 29588 15810 29600
rect 15930 29588 15936 29600
rect 15988 29588 15994 29640
rect 16025 29631 16083 29637
rect 16025 29597 16037 29631
rect 16071 29628 16083 29631
rect 17310 29628 17316 29640
rect 16071 29600 17316 29628
rect 16071 29597 16083 29600
rect 16025 29591 16083 29597
rect 16408 29572 16436 29600
rect 17310 29588 17316 29600
rect 17368 29588 17374 29640
rect 17770 29588 17776 29640
rect 17828 29628 17834 29640
rect 17865 29631 17923 29637
rect 17865 29628 17877 29631
rect 17828 29600 17877 29628
rect 17828 29588 17834 29600
rect 17865 29597 17877 29600
rect 17911 29597 17923 29631
rect 18046 29628 18052 29640
rect 18007 29600 18052 29628
rect 17865 29591 17923 29597
rect 18046 29588 18052 29600
rect 18104 29588 18110 29640
rect 18138 29588 18144 29640
rect 18196 29628 18202 29640
rect 18196 29600 18552 29628
rect 18196 29588 18202 29600
rect 16270 29563 16328 29569
rect 16270 29560 16282 29563
rect 12084 29532 16282 29560
rect 12084 29501 12112 29532
rect 16270 29529 16282 29532
rect 16316 29529 16328 29563
rect 16270 29523 16328 29529
rect 16390 29520 16396 29572
rect 16448 29520 16454 29572
rect 16666 29520 16672 29572
rect 16724 29560 16730 29572
rect 17034 29560 17040 29572
rect 16724 29532 17040 29560
rect 16724 29520 16730 29532
rect 17034 29520 17040 29532
rect 17092 29520 17098 29572
rect 17954 29560 17960 29572
rect 17144 29532 17960 29560
rect 12069 29495 12127 29501
rect 12069 29461 12081 29495
rect 12115 29461 12127 29495
rect 12069 29455 12127 29461
rect 13262 29452 13268 29504
rect 13320 29492 13326 29504
rect 13449 29495 13507 29501
rect 13449 29492 13461 29495
rect 13320 29464 13461 29492
rect 13320 29452 13326 29464
rect 13449 29461 13461 29464
rect 13495 29461 13507 29495
rect 13449 29455 13507 29461
rect 14277 29495 14335 29501
rect 14277 29461 14289 29495
rect 14323 29492 14335 29495
rect 14642 29492 14648 29504
rect 14323 29464 14648 29492
rect 14323 29461 14335 29464
rect 14277 29455 14335 29461
rect 14642 29452 14648 29464
rect 14700 29452 14706 29504
rect 14829 29495 14887 29501
rect 14829 29461 14841 29495
rect 14875 29492 14887 29495
rect 15746 29492 15752 29504
rect 14875 29464 15752 29492
rect 14875 29461 14887 29464
rect 14829 29455 14887 29461
rect 15746 29452 15752 29464
rect 15804 29452 15810 29504
rect 16022 29452 16028 29504
rect 16080 29492 16086 29504
rect 17144 29492 17172 29532
rect 17954 29520 17960 29532
rect 18012 29520 18018 29572
rect 18524 29560 18552 29600
rect 18598 29588 18604 29640
rect 18656 29628 18662 29640
rect 18966 29628 18972 29640
rect 18656 29600 18972 29628
rect 18656 29588 18662 29600
rect 18966 29588 18972 29600
rect 19024 29588 19030 29640
rect 19194 29628 19222 29668
rect 19518 29656 19524 29668
rect 19576 29656 19582 29708
rect 20548 29628 20576 29804
rect 20622 29724 20628 29776
rect 20680 29764 20686 29776
rect 20901 29767 20959 29773
rect 20901 29764 20913 29767
rect 20680 29736 20913 29764
rect 20680 29724 20686 29736
rect 20901 29733 20913 29736
rect 20947 29733 20959 29767
rect 20901 29727 20959 29733
rect 21818 29724 21824 29776
rect 21876 29764 21882 29776
rect 22278 29764 22284 29776
rect 21876 29736 22284 29764
rect 21876 29724 21882 29736
rect 22278 29724 22284 29736
rect 22336 29724 22342 29776
rect 22462 29764 22468 29776
rect 22423 29736 22468 29764
rect 22462 29724 22468 29736
rect 22520 29724 22526 29776
rect 22572 29764 22600 29804
rect 22830 29792 22836 29804
rect 22888 29792 22894 29844
rect 23382 29792 23388 29844
rect 23440 29832 23446 29844
rect 23569 29835 23627 29841
rect 23569 29832 23581 29835
rect 23440 29804 23581 29832
rect 23440 29792 23446 29804
rect 23569 29801 23581 29804
rect 23615 29801 23627 29835
rect 23569 29795 23627 29801
rect 23753 29835 23811 29841
rect 23753 29801 23765 29835
rect 23799 29832 23811 29835
rect 23842 29832 23848 29844
rect 23799 29804 23848 29832
rect 23799 29801 23811 29804
rect 23753 29795 23811 29801
rect 23842 29792 23848 29804
rect 23900 29792 23906 29844
rect 24578 29792 24584 29844
rect 24636 29832 24642 29844
rect 24765 29835 24823 29841
rect 24765 29832 24777 29835
rect 24636 29804 24777 29832
rect 24636 29792 24642 29804
rect 24765 29801 24777 29804
rect 24811 29801 24823 29835
rect 24765 29795 24823 29801
rect 26206 29804 27384 29832
rect 26206 29764 26234 29804
rect 22572 29736 26234 29764
rect 26697 29767 26755 29773
rect 26697 29733 26709 29767
rect 26743 29764 26755 29767
rect 26743 29736 27292 29764
rect 26743 29733 26755 29736
rect 26697 29727 26755 29733
rect 21910 29656 21916 29708
rect 21968 29696 21974 29708
rect 21968 29668 22048 29696
rect 21968 29656 21974 29668
rect 19194 29600 20576 29628
rect 20622 29588 20628 29640
rect 20680 29628 20686 29640
rect 21637 29631 21695 29637
rect 21637 29630 21649 29631
rect 21468 29628 21649 29630
rect 20680 29602 21649 29628
rect 20680 29600 21496 29602
rect 21632 29600 21649 29602
rect 20680 29588 20686 29600
rect 21637 29597 21649 29600
rect 21683 29597 21695 29631
rect 21637 29591 21695 29597
rect 21729 29631 21787 29637
rect 21729 29597 21741 29631
rect 21775 29597 21787 29631
rect 21729 29591 21787 29597
rect 19788 29563 19846 29569
rect 18062 29532 18359 29560
rect 18524 29532 19739 29560
rect 16080 29464 17172 29492
rect 16080 29452 16086 29464
rect 17218 29452 17224 29504
rect 17276 29492 17282 29504
rect 17405 29495 17463 29501
rect 17405 29492 17417 29495
rect 17276 29464 17417 29492
rect 17276 29452 17282 29464
rect 17405 29461 17417 29464
rect 17451 29461 17463 29495
rect 17405 29455 17463 29461
rect 17494 29452 17500 29504
rect 17552 29492 17558 29504
rect 18062 29492 18090 29532
rect 18230 29492 18236 29504
rect 17552 29464 18090 29492
rect 18191 29464 18236 29492
rect 17552 29452 17558 29464
rect 18230 29452 18236 29464
rect 18288 29452 18294 29504
rect 18331 29492 18359 29532
rect 19610 29492 19616 29504
rect 18331 29464 19616 29492
rect 19610 29452 19616 29464
rect 19668 29452 19674 29504
rect 19711 29492 19739 29532
rect 19788 29529 19800 29563
rect 19834 29560 19846 29563
rect 21361 29563 21419 29569
rect 21361 29560 21373 29563
rect 19834 29532 21373 29560
rect 19834 29529 19846 29532
rect 19788 29523 19846 29529
rect 21361 29529 21373 29532
rect 21407 29529 21419 29563
rect 21361 29523 21419 29529
rect 20990 29492 20996 29504
rect 19711 29464 20996 29492
rect 20990 29452 20996 29464
rect 21048 29452 21054 29504
rect 21082 29452 21088 29504
rect 21140 29492 21146 29504
rect 21450 29492 21456 29504
rect 21140 29464 21456 29492
rect 21140 29452 21146 29464
rect 21450 29452 21456 29464
rect 21508 29452 21514 29504
rect 21652 29492 21680 29591
rect 21744 29560 21772 29591
rect 21818 29588 21824 29640
rect 21876 29628 21882 29640
rect 22020 29637 22048 29668
rect 25038 29656 25044 29708
rect 25096 29696 25102 29708
rect 27264 29705 27292 29736
rect 26237 29699 26295 29705
rect 26237 29696 26249 29699
rect 25096 29668 26249 29696
rect 25096 29656 25102 29668
rect 26237 29665 26249 29668
rect 26283 29665 26295 29699
rect 26237 29659 26295 29665
rect 27249 29699 27307 29705
rect 27249 29665 27261 29699
rect 27295 29665 27307 29699
rect 27356 29696 27384 29804
rect 27614 29792 27620 29844
rect 27672 29832 27678 29844
rect 27890 29832 27896 29844
rect 27672 29804 27896 29832
rect 27672 29792 27678 29804
rect 27890 29792 27896 29804
rect 27948 29792 27954 29844
rect 28258 29792 28264 29844
rect 28316 29832 28322 29844
rect 28353 29835 28411 29841
rect 28353 29832 28365 29835
rect 28316 29804 28365 29832
rect 28316 29792 28322 29804
rect 28353 29801 28365 29804
rect 28399 29801 28411 29835
rect 28353 29795 28411 29801
rect 28718 29792 28724 29844
rect 28776 29832 28782 29844
rect 30282 29832 30288 29844
rect 28776 29804 30288 29832
rect 28776 29792 28782 29804
rect 30282 29792 30288 29804
rect 30340 29832 30346 29844
rect 32030 29832 32036 29844
rect 30340 29804 32036 29832
rect 30340 29792 30346 29804
rect 32030 29792 32036 29804
rect 32088 29792 32094 29844
rect 32217 29835 32275 29841
rect 32217 29801 32229 29835
rect 32263 29832 32275 29835
rect 32490 29832 32496 29844
rect 32263 29804 32496 29832
rect 32263 29801 32275 29804
rect 32217 29795 32275 29801
rect 32490 29792 32496 29804
rect 32548 29792 32554 29844
rect 33042 29792 33048 29844
rect 33100 29832 33106 29844
rect 34149 29835 34207 29841
rect 34149 29832 34161 29835
rect 33100 29804 34161 29832
rect 33100 29792 33106 29804
rect 34149 29801 34161 29804
rect 34195 29801 34207 29835
rect 34149 29795 34207 29801
rect 27430 29724 27436 29776
rect 27488 29764 27494 29776
rect 27488 29736 28994 29764
rect 27488 29724 27494 29736
rect 28966 29696 28994 29736
rect 29638 29724 29644 29776
rect 29696 29724 29702 29776
rect 30190 29724 30196 29776
rect 30248 29764 30254 29776
rect 30248 29736 32812 29764
rect 30248 29724 30254 29736
rect 29656 29696 29684 29724
rect 30009 29699 30067 29705
rect 27356 29668 28856 29696
rect 28966 29668 29040 29696
rect 29656 29668 29869 29696
rect 27249 29659 27307 29665
rect 22005 29631 22063 29637
rect 21876 29600 21921 29628
rect 21876 29588 21882 29600
rect 22005 29597 22017 29631
rect 22051 29597 22063 29631
rect 22005 29591 22063 29597
rect 22370 29588 22376 29640
rect 22428 29628 22434 29640
rect 22649 29631 22707 29637
rect 22649 29628 22661 29631
rect 22428 29600 22661 29628
rect 22428 29588 22434 29600
rect 22649 29597 22661 29600
rect 22695 29597 22707 29631
rect 22649 29591 22707 29597
rect 22738 29588 22744 29640
rect 22796 29628 22802 29640
rect 22925 29631 22983 29637
rect 22925 29628 22937 29631
rect 22796 29600 22937 29628
rect 22796 29588 22802 29600
rect 22925 29597 22937 29600
rect 22971 29597 22983 29631
rect 25406 29628 25412 29640
rect 22925 29591 22983 29597
rect 23012 29600 25066 29628
rect 25367 29600 25412 29628
rect 22186 29560 22192 29572
rect 21744 29532 22192 29560
rect 22186 29520 22192 29532
rect 22244 29520 22250 29572
rect 22554 29520 22560 29572
rect 22612 29560 22618 29572
rect 23012 29560 23040 29600
rect 22612 29532 23040 29560
rect 23385 29563 23443 29569
rect 22612 29520 22618 29532
rect 23385 29529 23397 29563
rect 23431 29560 23443 29563
rect 23474 29560 23480 29572
rect 23431 29532 23480 29560
rect 23431 29529 23443 29532
rect 23385 29523 23443 29529
rect 23474 29520 23480 29532
rect 23532 29520 23538 29572
rect 24118 29520 24124 29572
rect 24176 29560 24182 29572
rect 24397 29563 24455 29569
rect 24397 29560 24409 29563
rect 24176 29532 24409 29560
rect 24176 29520 24182 29532
rect 24397 29529 24409 29532
rect 24443 29529 24455 29563
rect 24397 29523 24455 29529
rect 24581 29563 24639 29569
rect 24581 29529 24593 29563
rect 24627 29560 24639 29563
rect 24670 29560 24676 29572
rect 24627 29532 24676 29560
rect 24627 29529 24639 29532
rect 24581 29523 24639 29529
rect 24670 29520 24676 29532
rect 24728 29560 24734 29572
rect 24946 29560 24952 29572
rect 24728 29532 24952 29560
rect 24728 29520 24734 29532
rect 24946 29520 24952 29532
rect 25004 29520 25010 29572
rect 25038 29560 25066 29600
rect 25406 29588 25412 29600
rect 25464 29588 25470 29640
rect 25498 29588 25504 29640
rect 25556 29628 25562 29640
rect 25556 29600 26234 29628
rect 25556 29588 25562 29600
rect 25685 29563 25743 29569
rect 25685 29560 25697 29563
rect 25038 29532 25697 29560
rect 25685 29529 25697 29532
rect 25731 29560 25743 29563
rect 25866 29560 25872 29572
rect 25731 29532 25872 29560
rect 25731 29529 25743 29532
rect 25685 29523 25743 29529
rect 25866 29520 25872 29532
rect 25924 29520 25930 29572
rect 26206 29560 26234 29600
rect 26326 29588 26332 29640
rect 26384 29628 26390 29640
rect 27062 29628 27068 29640
rect 26384 29600 26429 29628
rect 26804 29600 27068 29628
rect 26384 29588 26390 29600
rect 26804 29560 26832 29600
rect 27062 29588 27068 29600
rect 27120 29588 27126 29640
rect 27338 29628 27344 29640
rect 27299 29600 27344 29628
rect 27338 29588 27344 29600
rect 27396 29588 27402 29640
rect 28442 29588 28448 29640
rect 28500 29628 28506 29640
rect 28583 29631 28641 29637
rect 28583 29628 28595 29631
rect 28500 29600 28595 29628
rect 28500 29588 28506 29600
rect 28583 29597 28595 29600
rect 28629 29597 28641 29631
rect 28718 29628 28724 29640
rect 28679 29600 28724 29628
rect 28583 29591 28641 29597
rect 28718 29588 28724 29600
rect 28776 29588 28782 29640
rect 28828 29634 28856 29668
rect 29012 29637 29040 29668
rect 28813 29628 28871 29634
rect 28813 29594 28825 29628
rect 28859 29594 28871 29628
rect 28813 29588 28871 29594
rect 28997 29631 29055 29637
rect 28997 29597 29009 29631
rect 29043 29597 29055 29631
rect 28997 29591 29055 29597
rect 29362 29588 29368 29640
rect 29420 29628 29426 29640
rect 29841 29637 29869 29668
rect 30009 29665 30021 29699
rect 30055 29696 30067 29699
rect 30466 29696 30472 29708
rect 30055 29668 30472 29696
rect 30055 29665 30067 29668
rect 30009 29659 30067 29665
rect 30466 29656 30472 29668
rect 30524 29656 30530 29708
rect 30834 29656 30840 29708
rect 30892 29696 30898 29708
rect 32784 29705 32812 29736
rect 31205 29699 31263 29705
rect 31205 29696 31217 29699
rect 30892 29668 31217 29696
rect 30892 29656 30898 29668
rect 31205 29665 31217 29668
rect 31251 29665 31263 29699
rect 31205 29659 31263 29665
rect 32769 29699 32827 29705
rect 32769 29665 32781 29699
rect 32815 29665 32827 29699
rect 32769 29659 32827 29665
rect 29733 29631 29791 29637
rect 29733 29630 29745 29631
rect 29656 29628 29745 29630
rect 29420 29602 29745 29628
rect 29420 29600 29684 29602
rect 29420 29588 29426 29600
rect 29733 29597 29745 29602
rect 29779 29597 29791 29631
rect 29733 29591 29791 29597
rect 29826 29631 29884 29637
rect 29826 29597 29838 29631
rect 29872 29597 29884 29631
rect 29826 29591 29884 29597
rect 30101 29631 30159 29637
rect 30101 29597 30113 29631
rect 30147 29628 30159 29631
rect 30650 29628 30656 29640
rect 30147 29600 30656 29628
rect 30147 29597 30159 29600
rect 30101 29591 30159 29597
rect 30650 29588 30656 29600
rect 30708 29588 30714 29640
rect 31375 29631 31433 29637
rect 31375 29597 31387 29631
rect 31421 29628 31433 29631
rect 31421 29600 32076 29628
rect 31421 29597 31433 29600
rect 31375 29591 31433 29597
rect 26206 29532 26832 29560
rect 26878 29520 26884 29572
rect 26936 29560 26942 29572
rect 29270 29560 29276 29572
rect 26936 29532 29276 29560
rect 26936 29520 26942 29532
rect 29270 29520 29276 29532
rect 29328 29520 29334 29572
rect 22738 29492 22744 29504
rect 21652 29464 22744 29492
rect 22738 29452 22744 29464
rect 22796 29452 22802 29504
rect 23290 29452 23296 29504
rect 23348 29492 23354 29504
rect 23585 29495 23643 29501
rect 23585 29492 23597 29495
rect 23348 29464 23597 29492
rect 23348 29452 23354 29464
rect 23585 29461 23597 29464
rect 23631 29461 23643 29495
rect 23585 29455 23643 29461
rect 25958 29452 25964 29504
rect 26016 29492 26022 29504
rect 27709 29495 27767 29501
rect 27709 29492 27721 29495
rect 26016 29464 27721 29492
rect 26016 29452 26022 29464
rect 27709 29461 27721 29464
rect 27755 29461 27767 29495
rect 27709 29455 27767 29461
rect 27798 29452 27804 29504
rect 27856 29492 27862 29504
rect 29362 29492 29368 29504
rect 27856 29464 29368 29492
rect 27856 29452 27862 29464
rect 29362 29452 29368 29464
rect 29420 29452 29426 29504
rect 29549 29495 29607 29501
rect 29549 29461 29561 29495
rect 29595 29492 29607 29495
rect 30006 29492 30012 29504
rect 29595 29464 30012 29492
rect 29595 29461 29607 29464
rect 29549 29455 29607 29461
rect 30006 29452 30012 29464
rect 30064 29452 30070 29504
rect 31294 29452 31300 29504
rect 31352 29492 31358 29504
rect 31665 29495 31723 29501
rect 31665 29492 31677 29495
rect 31352 29464 31677 29492
rect 31352 29452 31358 29464
rect 31665 29461 31677 29464
rect 31711 29461 31723 29495
rect 32048 29492 32076 29600
rect 32122 29588 32128 29640
rect 32180 29628 32186 29640
rect 34146 29628 34152 29640
rect 32180 29600 34152 29628
rect 32180 29588 32186 29600
rect 34146 29588 34152 29600
rect 34204 29588 34210 29640
rect 32858 29520 32864 29572
rect 32916 29560 32922 29572
rect 33014 29563 33072 29569
rect 33014 29560 33026 29563
rect 32916 29532 33026 29560
rect 32916 29520 32922 29532
rect 33014 29529 33026 29532
rect 33060 29529 33072 29563
rect 33014 29523 33072 29529
rect 33686 29492 33692 29504
rect 32048 29464 33692 29492
rect 31665 29455 31723 29461
rect 33686 29452 33692 29464
rect 33744 29452 33750 29504
rect 1104 29402 34868 29424
rect 1104 29350 12214 29402
rect 12266 29350 12278 29402
rect 12330 29350 12342 29402
rect 12394 29350 12406 29402
rect 12458 29350 12470 29402
rect 12522 29350 23478 29402
rect 23530 29350 23542 29402
rect 23594 29350 23606 29402
rect 23658 29350 23670 29402
rect 23722 29350 23734 29402
rect 23786 29350 34868 29402
rect 1104 29328 34868 29350
rect 12986 29288 12992 29300
rect 12947 29260 12992 29288
rect 12986 29248 12992 29260
rect 13044 29248 13050 29300
rect 14182 29248 14188 29300
rect 14240 29288 14246 29300
rect 14240 29260 15608 29288
rect 14240 29248 14246 29260
rect 13814 29220 13820 29232
rect 11992 29192 12434 29220
rect 11992 29161 12020 29192
rect 11977 29155 12035 29161
rect 11977 29121 11989 29155
rect 12023 29121 12035 29155
rect 11977 29115 12035 29121
rect 12406 29084 12434 29192
rect 13188 29192 13820 29220
rect 13188 29161 13216 29192
rect 13814 29180 13820 29192
rect 13872 29180 13878 29232
rect 14642 29220 14648 29232
rect 14603 29192 14648 29220
rect 14642 29180 14648 29192
rect 14700 29180 14706 29232
rect 15580 29220 15608 29260
rect 15654 29248 15660 29300
rect 15712 29288 15718 29300
rect 22554 29288 22560 29300
rect 15712 29260 22560 29288
rect 15712 29248 15718 29260
rect 22554 29248 22560 29260
rect 22612 29248 22618 29300
rect 24302 29288 24308 29300
rect 22664 29260 24308 29288
rect 16574 29220 16580 29232
rect 15580 29192 16580 29220
rect 16574 29180 16580 29192
rect 16632 29180 16638 29232
rect 16675 29192 17356 29220
rect 13173 29155 13231 29161
rect 13173 29121 13185 29155
rect 13219 29121 13231 29155
rect 13173 29115 13231 29121
rect 13262 29112 13268 29164
rect 13320 29152 13326 29164
rect 13449 29155 13507 29161
rect 13320 29124 13365 29152
rect 13320 29112 13326 29124
rect 13449 29121 13461 29155
rect 13495 29152 13507 29155
rect 13630 29152 13636 29164
rect 13495 29124 13636 29152
rect 13495 29121 13507 29124
rect 13449 29115 13507 29121
rect 13630 29112 13636 29124
rect 13688 29112 13694 29164
rect 13909 29155 13967 29161
rect 13909 29152 13921 29155
rect 13832 29124 13921 29152
rect 13832 29096 13860 29124
rect 13909 29121 13921 29124
rect 13955 29121 13967 29155
rect 13909 29115 13967 29121
rect 14093 29155 14151 29161
rect 14093 29121 14105 29155
rect 14139 29121 14151 29155
rect 14550 29152 14556 29164
rect 14511 29124 14556 29152
rect 14093 29115 14151 29121
rect 12529 29087 12587 29093
rect 12529 29084 12541 29087
rect 12406 29056 12541 29084
rect 12529 29053 12541 29056
rect 12575 29084 12587 29087
rect 12897 29087 12955 29093
rect 12897 29084 12909 29087
rect 12575 29056 12909 29084
rect 12575 29053 12587 29056
rect 12529 29047 12587 29053
rect 12897 29053 12909 29056
rect 12943 29084 12955 29087
rect 13722 29084 13728 29096
rect 12943 29056 13728 29084
rect 12943 29053 12955 29056
rect 12897 29047 12955 29053
rect 13722 29044 13728 29056
rect 13780 29044 13786 29096
rect 13814 29044 13820 29096
rect 13872 29044 13878 29096
rect 13998 29084 14004 29096
rect 13959 29056 14004 29084
rect 13998 29044 14004 29056
rect 14056 29044 14062 29096
rect 14108 29084 14136 29115
rect 14550 29112 14556 29124
rect 14608 29112 14614 29164
rect 14737 29155 14795 29161
rect 14737 29121 14749 29155
rect 14783 29152 14795 29155
rect 15102 29152 15108 29164
rect 14783 29124 15108 29152
rect 14783 29121 14795 29124
rect 14737 29115 14795 29121
rect 15102 29112 15108 29124
rect 15160 29112 15166 29164
rect 15197 29155 15255 29161
rect 15197 29121 15209 29155
rect 15243 29152 15255 29155
rect 15470 29152 15476 29164
rect 15243 29124 15476 29152
rect 15243 29121 15255 29124
rect 15197 29115 15255 29121
rect 15470 29112 15476 29124
rect 15528 29112 15534 29164
rect 15654 29112 15660 29164
rect 15712 29152 15718 29164
rect 15841 29155 15899 29161
rect 15841 29152 15853 29155
rect 15712 29124 15853 29152
rect 15712 29112 15718 29124
rect 15841 29121 15853 29124
rect 15887 29121 15899 29155
rect 15841 29115 15899 29121
rect 16025 29155 16083 29161
rect 16025 29121 16037 29155
rect 16071 29121 16083 29155
rect 16025 29115 16083 29121
rect 14826 29084 14832 29096
rect 14108 29056 14832 29084
rect 14826 29044 14832 29056
rect 14884 29044 14890 29096
rect 15562 29044 15568 29096
rect 15620 29084 15626 29096
rect 16040 29084 16068 29115
rect 16114 29112 16120 29164
rect 16172 29152 16178 29164
rect 16172 29124 16217 29152
rect 16172 29112 16178 29124
rect 16675 29084 16703 29192
rect 17201 29155 17259 29161
rect 17201 29152 17213 29155
rect 15620 29056 16703 29084
rect 16776 29124 17213 29152
rect 15620 29044 15626 29056
rect 15286 28976 15292 29028
rect 15344 29016 15350 29028
rect 16114 29016 16120 29028
rect 15344 28988 15389 29016
rect 15672 28988 16120 29016
rect 15344 28976 15350 28988
rect 12158 28948 12164 28960
rect 12119 28920 12164 28948
rect 12158 28908 12164 28920
rect 12216 28908 12222 28960
rect 13446 28948 13452 28960
rect 13407 28920 13452 28948
rect 13446 28908 13452 28920
rect 13504 28908 13510 28960
rect 13630 28908 13636 28960
rect 13688 28948 13694 28960
rect 13725 28951 13783 28957
rect 13725 28948 13737 28951
rect 13688 28920 13737 28948
rect 13688 28908 13694 28920
rect 13725 28917 13737 28920
rect 13771 28917 13783 28951
rect 13725 28911 13783 28917
rect 13998 28908 14004 28960
rect 14056 28948 14062 28960
rect 15010 28948 15016 28960
rect 14056 28920 15016 28948
rect 14056 28908 14062 28920
rect 15010 28908 15016 28920
rect 15068 28948 15074 28960
rect 15672 28948 15700 28988
rect 16114 28976 16120 28988
rect 16172 28976 16178 29028
rect 16206 28976 16212 29028
rect 16264 29016 16270 29028
rect 16776 29016 16804 29124
rect 17201 29121 17213 29124
rect 17247 29121 17259 29155
rect 17328 29152 17356 29192
rect 17402 29180 17408 29232
rect 17460 29220 17466 29232
rect 18322 29220 18328 29232
rect 17460 29192 18328 29220
rect 17460 29180 17466 29192
rect 18322 29180 18328 29192
rect 18380 29180 18386 29232
rect 18506 29180 18512 29232
rect 18564 29220 18570 29232
rect 19981 29223 20039 29229
rect 19981 29220 19993 29223
rect 18564 29192 19993 29220
rect 18564 29180 18570 29192
rect 19981 29189 19993 29192
rect 20027 29189 20039 29223
rect 19981 29183 20039 29189
rect 20438 29180 20444 29232
rect 20496 29220 20502 29232
rect 21818 29220 21824 29232
rect 20496 29192 21683 29220
rect 21779 29192 21824 29220
rect 20496 29180 20502 29192
rect 17328 29124 17991 29152
rect 17201 29115 17259 29121
rect 16942 29084 16948 29096
rect 16903 29056 16948 29084
rect 16942 29044 16948 29056
rect 17000 29044 17006 29096
rect 17963 29084 17991 29124
rect 18046 29112 18052 29164
rect 18104 29152 18110 29164
rect 18598 29152 18604 29164
rect 18104 29124 18604 29152
rect 18104 29112 18110 29124
rect 18598 29112 18604 29124
rect 18656 29112 18662 29164
rect 18708 29124 18920 29152
rect 18708 29084 18736 29124
rect 17963 29056 18736 29084
rect 18785 29087 18843 29093
rect 18785 29053 18797 29087
rect 18831 29053 18843 29087
rect 18892 29084 18920 29124
rect 18966 29112 18972 29164
rect 19024 29152 19030 29164
rect 19797 29155 19855 29161
rect 19797 29152 19809 29155
rect 19024 29124 19809 29152
rect 19024 29112 19030 29124
rect 19797 29121 19809 29124
rect 19843 29121 19855 29155
rect 20990 29152 20996 29164
rect 20951 29124 20996 29152
rect 19797 29115 19855 29121
rect 20990 29112 20996 29124
rect 21048 29112 21054 29164
rect 21269 29155 21327 29161
rect 21269 29121 21281 29155
rect 21315 29152 21327 29155
rect 21358 29152 21364 29164
rect 21315 29124 21364 29152
rect 21315 29121 21327 29124
rect 21269 29115 21327 29121
rect 21358 29112 21364 29124
rect 21416 29112 21422 29164
rect 21655 29152 21683 29192
rect 21818 29180 21824 29192
rect 21876 29180 21882 29232
rect 22002 29220 22008 29232
rect 21963 29192 22008 29220
rect 22002 29180 22008 29192
rect 22060 29220 22066 29232
rect 22664 29220 22692 29260
rect 24302 29248 24308 29260
rect 24360 29248 24366 29300
rect 25406 29248 25412 29300
rect 25464 29288 25470 29300
rect 31662 29288 31668 29300
rect 25464 29260 31668 29288
rect 25464 29248 25470 29260
rect 31662 29248 31668 29260
rect 31720 29248 31726 29300
rect 32858 29288 32864 29300
rect 32819 29260 32864 29288
rect 32858 29248 32864 29260
rect 32916 29248 32922 29300
rect 33318 29248 33324 29300
rect 33376 29248 33382 29300
rect 34054 29288 34060 29300
rect 34015 29260 34060 29288
rect 34054 29248 34060 29260
rect 34112 29248 34118 29300
rect 22060 29192 22692 29220
rect 22060 29180 22066 29192
rect 22738 29180 22744 29232
rect 22796 29220 22802 29232
rect 27062 29220 27068 29232
rect 22796 29192 22841 29220
rect 22940 29192 23149 29220
rect 22796 29180 22802 29192
rect 22462 29152 22468 29164
rect 21655 29124 22468 29152
rect 22462 29112 22468 29124
rect 22520 29112 22526 29164
rect 22830 29112 22836 29164
rect 22888 29152 22894 29164
rect 22940 29152 22968 29192
rect 23014 29161 23020 29164
rect 22888 29124 22968 29152
rect 22997 29155 23020 29161
rect 22888 29112 22894 29124
rect 22997 29121 23009 29155
rect 22997 29115 23020 29121
rect 23014 29112 23020 29115
rect 23072 29112 23078 29164
rect 23121 29161 23149 29192
rect 24136 29192 27068 29220
rect 23244 29161 23250 29164
rect 23121 29155 23180 29161
rect 23121 29124 23134 29155
rect 23122 29121 23134 29124
rect 23168 29121 23180 29155
rect 23122 29115 23180 29121
rect 23222 29155 23250 29161
rect 23222 29121 23234 29155
rect 23222 29115 23250 29121
rect 23244 29112 23250 29115
rect 23302 29112 23308 29164
rect 23385 29155 23443 29161
rect 23385 29121 23397 29155
rect 23431 29152 23443 29155
rect 23474 29152 23480 29164
rect 23431 29124 23480 29152
rect 23431 29121 23443 29124
rect 23385 29115 23443 29121
rect 23474 29112 23480 29124
rect 23532 29112 23538 29164
rect 24136 29161 24164 29192
rect 24394 29161 24400 29164
rect 24121 29155 24179 29161
rect 24121 29121 24133 29155
rect 24167 29121 24179 29155
rect 24388 29152 24400 29161
rect 24355 29124 24400 29152
rect 24121 29115 24179 29121
rect 24388 29115 24400 29124
rect 19610 29084 19616 29096
rect 18892 29056 19380 29084
rect 19571 29056 19616 29084
rect 18785 29047 18843 29053
rect 16264 28988 16804 29016
rect 18325 29019 18383 29025
rect 16264 28976 16270 28988
rect 18325 28985 18337 29019
rect 18371 29016 18383 29019
rect 18800 29016 18828 29047
rect 18966 29016 18972 29028
rect 18371 28988 18972 29016
rect 18371 28985 18383 28988
rect 18325 28979 18383 28985
rect 18966 28976 18972 28988
rect 19024 28976 19030 29028
rect 19153 29019 19211 29025
rect 19153 28985 19165 29019
rect 19199 29016 19211 29019
rect 19242 29016 19248 29028
rect 19199 28988 19248 29016
rect 19199 28985 19211 28988
rect 19153 28979 19211 28985
rect 19242 28976 19248 28988
rect 19300 28976 19306 29028
rect 19352 29016 19380 29056
rect 19610 29044 19616 29056
rect 19668 29044 19674 29096
rect 19711 29056 21956 29084
rect 19711 29016 19739 29056
rect 19352 28988 19739 29016
rect 20162 28976 20168 29028
rect 20220 29016 20226 29028
rect 20993 29019 21051 29025
rect 20993 29016 21005 29019
rect 20220 28988 21005 29016
rect 20220 28976 20226 28988
rect 20993 28985 21005 28988
rect 21039 28985 21051 29019
rect 20993 28979 21051 28985
rect 21085 29019 21143 29025
rect 21085 28985 21097 29019
rect 21131 29016 21143 29019
rect 21818 29016 21824 29028
rect 21131 28988 21824 29016
rect 21131 28985 21143 28988
rect 21085 28979 21143 28985
rect 21818 28976 21824 28988
rect 21876 28976 21882 29028
rect 21928 29016 21956 29056
rect 22094 29044 22100 29096
rect 22152 29084 22158 29096
rect 22189 29087 22247 29093
rect 22189 29084 22201 29087
rect 22152 29056 22201 29084
rect 22152 29044 22158 29056
rect 22189 29053 22201 29056
rect 22235 29053 22247 29087
rect 22480 29084 22508 29112
rect 24136 29084 24164 29115
rect 24394 29112 24400 29115
rect 24452 29112 24458 29164
rect 24670 29112 24676 29164
rect 24728 29152 24734 29164
rect 25958 29152 25964 29164
rect 24728 29124 25176 29152
rect 25919 29124 25964 29152
rect 24728 29112 24734 29124
rect 22480 29056 24164 29084
rect 25148 29084 25176 29124
rect 25958 29112 25964 29124
rect 26016 29112 26022 29164
rect 26142 29152 26148 29164
rect 26103 29124 26148 29152
rect 26142 29112 26148 29124
rect 26200 29112 26206 29164
rect 26329 29155 26387 29161
rect 26329 29121 26341 29155
rect 26375 29152 26387 29155
rect 26602 29152 26608 29164
rect 26375 29124 26608 29152
rect 26375 29121 26387 29124
rect 26329 29115 26387 29121
rect 26602 29112 26608 29124
rect 26660 29112 26666 29164
rect 26988 29161 27016 29192
rect 27062 29180 27068 29192
rect 27120 29220 27126 29232
rect 30098 29220 30104 29232
rect 27120 29192 30104 29220
rect 27120 29180 27126 29192
rect 28828 29161 28856 29192
rect 30098 29180 30104 29192
rect 30156 29180 30162 29232
rect 32217 29223 32275 29229
rect 32217 29220 32229 29223
rect 30208 29192 31432 29220
rect 29086 29161 29092 29164
rect 26973 29155 27031 29161
rect 26973 29121 26985 29155
rect 27019 29121 27031 29155
rect 27229 29155 27287 29161
rect 27229 29152 27241 29155
rect 26973 29115 27031 29121
rect 27080 29124 27241 29152
rect 26237 29087 26295 29093
rect 26237 29084 26249 29087
rect 25148 29056 26249 29084
rect 22189 29047 22247 29053
rect 26237 29053 26249 29056
rect 26283 29053 26295 29087
rect 26237 29047 26295 29053
rect 26421 29087 26479 29093
rect 26421 29053 26433 29087
rect 26467 29084 26479 29087
rect 27080 29084 27108 29124
rect 27229 29121 27241 29124
rect 27275 29121 27287 29155
rect 27229 29115 27287 29121
rect 28813 29155 28871 29161
rect 28813 29121 28825 29155
rect 28859 29121 28871 29155
rect 28813 29115 28871 29121
rect 29080 29115 29092 29161
rect 29144 29152 29150 29164
rect 29144 29124 29180 29152
rect 29086 29112 29092 29115
rect 29144 29112 29150 29124
rect 29362 29112 29368 29164
rect 29420 29152 29426 29164
rect 30208 29152 30236 29192
rect 29420 29124 30236 29152
rect 29420 29112 29426 29124
rect 30374 29112 30380 29164
rect 30432 29152 30438 29164
rect 31205 29155 31263 29161
rect 31205 29152 31217 29155
rect 30432 29124 31217 29152
rect 30432 29112 30438 29124
rect 31205 29121 31217 29124
rect 31251 29121 31263 29155
rect 31205 29115 31263 29121
rect 31294 29084 31300 29096
rect 26467 29056 27108 29084
rect 31255 29056 31300 29084
rect 26467 29053 26479 29056
rect 26421 29047 26479 29053
rect 31294 29044 31300 29056
rect 31352 29044 31358 29096
rect 31404 29084 31432 29192
rect 31726 29192 32229 29220
rect 31726 29164 31754 29192
rect 32217 29189 32229 29192
rect 32263 29189 32275 29223
rect 33336 29220 33364 29248
rect 33594 29220 33600 29232
rect 32217 29183 32275 29189
rect 33244 29192 33600 29220
rect 31662 29112 31668 29164
rect 31720 29124 31754 29164
rect 31720 29112 31726 29124
rect 31846 29112 31852 29164
rect 31904 29152 31910 29164
rect 33042 29152 33048 29164
rect 31904 29124 33048 29152
rect 31904 29112 31910 29124
rect 33042 29112 33048 29124
rect 33100 29152 33106 29164
rect 33244 29161 33272 29192
rect 33594 29180 33600 29192
rect 33652 29180 33658 29232
rect 33137 29155 33195 29161
rect 33137 29152 33149 29155
rect 33100 29124 33149 29152
rect 33100 29112 33106 29124
rect 33137 29121 33149 29124
rect 33183 29121 33195 29155
rect 33137 29115 33195 29121
rect 33229 29155 33287 29161
rect 33229 29121 33241 29155
rect 33275 29121 33287 29155
rect 33229 29115 33287 29121
rect 33321 29155 33379 29161
rect 33321 29121 33333 29155
rect 33367 29121 33379 29155
rect 33502 29152 33508 29164
rect 33463 29124 33508 29152
rect 33321 29115 33379 29121
rect 33336 29084 33364 29115
rect 33502 29112 33508 29124
rect 33560 29112 33566 29164
rect 33870 29112 33876 29164
rect 33928 29152 33934 29164
rect 33965 29155 34023 29161
rect 33965 29152 33977 29155
rect 33928 29124 33977 29152
rect 33928 29112 33934 29124
rect 33965 29121 33977 29124
rect 34011 29121 34023 29155
rect 33965 29115 34023 29121
rect 31404 29056 33364 29084
rect 22554 29016 22560 29028
rect 21928 28988 22560 29016
rect 22554 28976 22560 28988
rect 22612 28976 22618 29028
rect 22646 28976 22652 29028
rect 22704 29016 22710 29028
rect 28353 29019 28411 29025
rect 28353 29016 28365 29019
rect 22704 28988 24063 29016
rect 22704 28976 22710 28988
rect 15068 28920 15700 28948
rect 15841 28951 15899 28957
rect 15068 28908 15074 28920
rect 15841 28917 15853 28951
rect 15887 28948 15899 28951
rect 22094 28948 22100 28960
rect 15887 28920 22100 28948
rect 15887 28917 15899 28920
rect 15841 28911 15899 28917
rect 22094 28908 22100 28920
rect 22152 28908 22158 28960
rect 22278 28908 22284 28960
rect 22336 28948 22342 28960
rect 23934 28948 23940 28960
rect 22336 28920 23940 28948
rect 22336 28908 22342 28920
rect 23934 28908 23940 28920
rect 23992 28908 23998 28960
rect 24035 28948 24063 28988
rect 25056 28988 26372 29016
rect 25056 28948 25084 28988
rect 24035 28920 25084 28948
rect 25501 28951 25559 28957
rect 25501 28917 25513 28951
rect 25547 28948 25559 28951
rect 25682 28948 25688 28960
rect 25547 28920 25688 28948
rect 25547 28917 25559 28920
rect 25501 28911 25559 28917
rect 25682 28908 25688 28920
rect 25740 28908 25746 28960
rect 26344 28948 26372 28988
rect 27908 28988 28365 29016
rect 27908 28948 27936 28988
rect 28353 28985 28365 28988
rect 28399 28985 28411 29019
rect 31573 29019 31631 29025
rect 31573 29016 31585 29019
rect 28353 28979 28411 28985
rect 29748 28988 31585 29016
rect 26344 28920 27936 28948
rect 28718 28908 28724 28960
rect 28776 28948 28782 28960
rect 29748 28948 29776 28988
rect 31573 28985 31585 28988
rect 31619 28985 31631 29019
rect 31573 28979 31631 28985
rect 32401 29019 32459 29025
rect 32401 28985 32413 29019
rect 32447 29016 32459 29019
rect 32490 29016 32496 29028
rect 32447 28988 32496 29016
rect 32447 28985 32459 28988
rect 32401 28979 32459 28985
rect 32490 28976 32496 28988
rect 32548 28976 32554 29028
rect 30190 28948 30196 28960
rect 28776 28920 29776 28948
rect 30151 28920 30196 28948
rect 28776 28908 28782 28920
rect 30190 28908 30196 28920
rect 30248 28908 30254 28960
rect 1104 28858 34868 28880
rect 1104 28806 6582 28858
rect 6634 28806 6646 28858
rect 6698 28806 6710 28858
rect 6762 28806 6774 28858
rect 6826 28806 6838 28858
rect 6890 28806 17846 28858
rect 17898 28806 17910 28858
rect 17962 28806 17974 28858
rect 18026 28806 18038 28858
rect 18090 28806 18102 28858
rect 18154 28806 29110 28858
rect 29162 28806 29174 28858
rect 29226 28806 29238 28858
rect 29290 28806 29302 28858
rect 29354 28806 29366 28858
rect 29418 28806 34868 28858
rect 1104 28784 34868 28806
rect 12713 28747 12771 28753
rect 12713 28713 12725 28747
rect 12759 28744 12771 28747
rect 16574 28744 16580 28756
rect 12759 28716 16580 28744
rect 12759 28713 12771 28716
rect 12713 28707 12771 28713
rect 16574 28704 16580 28716
rect 16632 28704 16638 28756
rect 16666 28704 16672 28756
rect 16724 28744 16730 28756
rect 19058 28744 19064 28756
rect 16724 28716 19064 28744
rect 16724 28704 16730 28716
rect 19058 28704 19064 28716
rect 19116 28704 19122 28756
rect 19518 28744 19524 28756
rect 19260 28716 19524 28744
rect 13357 28679 13415 28685
rect 13357 28645 13369 28679
rect 13403 28676 13415 28679
rect 16206 28676 16212 28688
rect 13403 28648 16212 28676
rect 13403 28645 13415 28648
rect 13357 28639 13415 28645
rect 16206 28636 16212 28648
rect 16264 28636 16270 28688
rect 17494 28636 17500 28688
rect 17552 28676 17558 28688
rect 18506 28676 18512 28688
rect 17552 28648 18512 28676
rect 17552 28636 17558 28648
rect 18506 28636 18512 28648
rect 18564 28636 18570 28688
rect 18598 28636 18604 28688
rect 18656 28676 18662 28688
rect 18874 28676 18880 28688
rect 18656 28648 18880 28676
rect 18656 28636 18662 28648
rect 18874 28636 18880 28648
rect 18932 28636 18938 28688
rect 12158 28568 12164 28620
rect 12216 28608 12222 28620
rect 16114 28608 16120 28620
rect 12216 28580 16120 28608
rect 12216 28568 12222 28580
rect 16114 28568 16120 28580
rect 16172 28568 16178 28620
rect 18141 28611 18199 28617
rect 18141 28577 18153 28611
rect 18187 28608 18199 28611
rect 18966 28608 18972 28620
rect 18187 28580 18972 28608
rect 18187 28577 18199 28580
rect 18141 28571 18199 28577
rect 18966 28568 18972 28580
rect 19024 28568 19030 28620
rect 19260 28617 19288 28716
rect 19518 28704 19524 28716
rect 19576 28704 19582 28756
rect 19610 28704 19616 28756
rect 19668 28744 19674 28756
rect 20625 28747 20683 28753
rect 20625 28744 20637 28747
rect 19668 28716 20637 28744
rect 19668 28704 19674 28716
rect 20625 28713 20637 28716
rect 20671 28713 20683 28747
rect 22002 28744 22008 28756
rect 20625 28707 20683 28713
rect 20916 28716 22008 28744
rect 20254 28636 20260 28688
rect 20312 28636 20318 28688
rect 20438 28636 20444 28688
rect 20496 28676 20502 28688
rect 20916 28676 20944 28716
rect 22002 28704 22008 28716
rect 22060 28704 22066 28756
rect 22094 28704 22100 28756
rect 22152 28744 22158 28756
rect 22152 28716 23520 28744
rect 22152 28704 22158 28716
rect 21082 28676 21088 28688
rect 20496 28648 20944 28676
rect 21043 28648 21088 28676
rect 20496 28636 20502 28648
rect 21082 28636 21088 28648
rect 21140 28636 21146 28688
rect 21453 28679 21511 28685
rect 21453 28645 21465 28679
rect 21499 28676 21511 28679
rect 22186 28676 22192 28688
rect 21499 28648 22192 28676
rect 21499 28645 21511 28648
rect 21453 28639 21511 28645
rect 22186 28636 22192 28648
rect 22244 28636 22250 28688
rect 19245 28611 19303 28617
rect 19245 28577 19257 28611
rect 19291 28577 19303 28611
rect 20272 28608 20300 28636
rect 20272 28580 22416 28608
rect 19245 28571 19303 28577
rect 12897 28543 12955 28549
rect 12897 28509 12909 28543
rect 12943 28540 12955 28543
rect 13446 28540 13452 28552
rect 12943 28512 13452 28540
rect 12943 28509 12955 28512
rect 12897 28503 12955 28509
rect 13446 28500 13452 28512
rect 13504 28500 13510 28552
rect 13541 28543 13599 28549
rect 13541 28509 13553 28543
rect 13587 28540 13599 28543
rect 13722 28540 13728 28552
rect 13587 28512 13728 28540
rect 13587 28509 13599 28512
rect 13541 28503 13599 28509
rect 13722 28500 13728 28512
rect 13780 28500 13786 28552
rect 14642 28540 14648 28552
rect 14603 28512 14648 28540
rect 14642 28500 14648 28512
rect 14700 28500 14706 28552
rect 14737 28543 14795 28549
rect 14737 28509 14749 28543
rect 14783 28540 14795 28543
rect 14826 28540 14832 28552
rect 14783 28512 14832 28540
rect 14783 28509 14795 28512
rect 14737 28503 14795 28509
rect 14826 28500 14832 28512
rect 14884 28500 14890 28552
rect 15102 28500 15108 28552
rect 15160 28540 15166 28552
rect 15286 28540 15292 28552
rect 15160 28512 15292 28540
rect 15160 28500 15166 28512
rect 15286 28500 15292 28512
rect 15344 28500 15350 28552
rect 15381 28543 15439 28549
rect 15381 28509 15393 28543
rect 15427 28540 15439 28543
rect 15470 28540 15476 28552
rect 15427 28512 15476 28540
rect 15427 28509 15439 28512
rect 15381 28503 15439 28509
rect 15470 28500 15476 28512
rect 15528 28500 15534 28552
rect 16301 28543 16359 28549
rect 16301 28509 16313 28543
rect 16347 28540 16359 28543
rect 16942 28540 16948 28552
rect 16347 28512 16948 28540
rect 16347 28509 16359 28512
rect 16301 28503 16359 28509
rect 16942 28500 16948 28512
rect 17000 28540 17006 28552
rect 17310 28540 17316 28552
rect 17000 28512 17316 28540
rect 17000 28500 17006 28512
rect 17310 28500 17316 28512
rect 17368 28500 17374 28552
rect 17512 28512 19831 28540
rect 13262 28432 13268 28484
rect 13320 28472 13326 28484
rect 16557 28475 16615 28481
rect 16557 28472 16569 28475
rect 13320 28444 16569 28472
rect 13320 28432 13326 28444
rect 16557 28441 16569 28444
rect 16603 28441 16615 28475
rect 16557 28435 16615 28441
rect 16850 28364 16856 28416
rect 16908 28404 16914 28416
rect 17512 28404 17540 28512
rect 17770 28432 17776 28484
rect 17828 28432 17834 28484
rect 18417 28475 18475 28481
rect 18417 28441 18429 28475
rect 18463 28472 18475 28475
rect 19334 28472 19340 28484
rect 18463 28444 19340 28472
rect 18463 28441 18475 28444
rect 18417 28435 18475 28441
rect 19334 28432 19340 28444
rect 19392 28432 19398 28484
rect 19512 28475 19570 28481
rect 19512 28441 19524 28475
rect 19558 28472 19570 28475
rect 19702 28472 19708 28484
rect 19558 28444 19708 28472
rect 19558 28441 19570 28444
rect 19512 28435 19570 28441
rect 19702 28432 19708 28444
rect 19760 28432 19766 28484
rect 19803 28472 19831 28512
rect 20254 28500 20260 28552
rect 20312 28540 20318 28552
rect 21269 28543 21327 28549
rect 21269 28540 21281 28543
rect 20312 28512 21281 28540
rect 20312 28500 20318 28512
rect 21269 28509 21281 28512
rect 21315 28509 21327 28543
rect 21269 28503 21327 28509
rect 21358 28500 21364 28552
rect 21416 28540 21422 28552
rect 21545 28543 21603 28549
rect 21545 28540 21557 28543
rect 21416 28512 21557 28540
rect 21416 28500 21422 28512
rect 21545 28509 21557 28512
rect 21591 28509 21603 28543
rect 22388 28540 22416 28580
rect 22462 28568 22468 28620
rect 22520 28608 22526 28620
rect 23492 28608 23520 28716
rect 23566 28704 23572 28756
rect 23624 28744 23630 28756
rect 28074 28744 28080 28756
rect 23624 28716 28080 28744
rect 23624 28704 23630 28716
rect 28074 28704 28080 28716
rect 28132 28704 28138 28756
rect 28537 28747 28595 28753
rect 28537 28713 28549 28747
rect 28583 28744 28595 28747
rect 28994 28744 29000 28756
rect 28583 28716 29000 28744
rect 28583 28713 28595 28716
rect 28537 28707 28595 28713
rect 28994 28704 29000 28716
rect 29052 28704 29058 28756
rect 29104 28716 31064 28744
rect 23842 28636 23848 28688
rect 23900 28676 23906 28688
rect 24210 28676 24216 28688
rect 23900 28648 24216 28676
rect 23900 28636 23906 28648
rect 24210 28636 24216 28648
rect 24268 28636 24274 28688
rect 27065 28679 27123 28685
rect 27065 28645 27077 28679
rect 27111 28676 27123 28679
rect 27522 28676 27528 28688
rect 27111 28648 27528 28676
rect 27111 28645 27123 28648
rect 27065 28639 27123 28645
rect 27522 28636 27528 28648
rect 27580 28636 27586 28688
rect 28626 28636 28632 28688
rect 28684 28676 28690 28688
rect 28905 28679 28963 28685
rect 28905 28676 28917 28679
rect 28684 28648 28917 28676
rect 28684 28636 28690 28648
rect 28905 28645 28917 28648
rect 28951 28645 28963 28679
rect 28905 28639 28963 28645
rect 22520 28580 22565 28608
rect 23492 28580 28120 28608
rect 22520 28568 22526 28580
rect 22554 28540 22560 28552
rect 22388 28512 22560 28540
rect 21545 28503 21603 28509
rect 22554 28500 22560 28512
rect 22612 28500 22618 28552
rect 22738 28549 22744 28552
rect 22732 28503 22744 28549
rect 22796 28540 22802 28552
rect 26329 28543 26387 28549
rect 26329 28540 26341 28543
rect 22796 28512 22832 28540
rect 22940 28512 26341 28540
rect 22738 28500 22744 28503
rect 22796 28500 22802 28512
rect 22940 28472 22968 28512
rect 26329 28509 26341 28512
rect 26375 28509 26387 28543
rect 26329 28503 26387 28509
rect 26973 28543 27031 28549
rect 26973 28509 26985 28543
rect 27019 28509 27031 28543
rect 27246 28540 27252 28552
rect 27207 28512 27252 28540
rect 26973 28503 27031 28509
rect 19803 28444 22968 28472
rect 23014 28432 23020 28484
rect 23072 28472 23078 28484
rect 23566 28472 23572 28484
rect 23072 28444 23572 28472
rect 23072 28432 23078 28444
rect 23566 28432 23572 28444
rect 23624 28432 23630 28484
rect 24762 28472 24768 28484
rect 24723 28444 24768 28472
rect 24762 28432 24768 28444
rect 24820 28432 24826 28484
rect 16908 28376 17540 28404
rect 17681 28407 17739 28413
rect 16908 28364 16914 28376
rect 17681 28373 17693 28407
rect 17727 28404 17739 28407
rect 17788 28404 17816 28432
rect 18322 28404 18328 28416
rect 17727 28376 18328 28404
rect 17727 28373 17739 28376
rect 17681 28367 17739 28373
rect 18322 28364 18328 28376
rect 18380 28364 18386 28416
rect 18506 28404 18512 28416
rect 18467 28376 18512 28404
rect 18506 28364 18512 28376
rect 18564 28364 18570 28416
rect 18690 28364 18696 28416
rect 18748 28404 18754 28416
rect 18748 28376 18793 28404
rect 18748 28364 18754 28376
rect 18874 28364 18880 28416
rect 18932 28404 18938 28416
rect 19150 28404 19156 28416
rect 18932 28376 19156 28404
rect 18932 28364 18938 28376
rect 19150 28364 19156 28376
rect 19208 28404 19214 28416
rect 19610 28404 19616 28416
rect 19208 28376 19616 28404
rect 19208 28364 19214 28376
rect 19610 28364 19616 28376
rect 19668 28364 19674 28416
rect 19794 28364 19800 28416
rect 19852 28404 19858 28416
rect 22278 28404 22284 28416
rect 19852 28376 22284 28404
rect 19852 28364 19858 28376
rect 22278 28364 22284 28376
rect 22336 28364 22342 28416
rect 22370 28364 22376 28416
rect 22428 28404 22434 28416
rect 23106 28404 23112 28416
rect 22428 28376 23112 28404
rect 22428 28364 22434 28376
rect 23106 28364 23112 28376
rect 23164 28364 23170 28416
rect 23198 28364 23204 28416
rect 23256 28404 23262 28416
rect 23845 28407 23903 28413
rect 23845 28404 23857 28407
rect 23256 28376 23857 28404
rect 23256 28364 23262 28376
rect 23845 28373 23857 28376
rect 23891 28373 23903 28407
rect 23845 28367 23903 28373
rect 24210 28364 24216 28416
rect 24268 28404 24274 28416
rect 24670 28404 24676 28416
rect 24268 28376 24676 28404
rect 24268 28364 24274 28376
rect 24670 28364 24676 28376
rect 24728 28364 24734 28416
rect 26988 28404 27016 28503
rect 27246 28500 27252 28512
rect 27304 28500 27310 28552
rect 27430 28540 27436 28552
rect 27391 28512 27436 28540
rect 27430 28500 27436 28512
rect 27488 28500 27494 28552
rect 27801 28543 27859 28549
rect 27801 28509 27813 28543
rect 27847 28509 27859 28543
rect 27982 28540 27988 28552
rect 27943 28512 27988 28540
rect 27801 28503 27859 28509
rect 27062 28432 27068 28484
rect 27120 28472 27126 28484
rect 27522 28472 27528 28484
rect 27120 28444 27528 28472
rect 27120 28432 27126 28444
rect 27522 28432 27528 28444
rect 27580 28472 27586 28484
rect 27816 28472 27844 28503
rect 27982 28500 27988 28512
rect 28040 28500 28046 28552
rect 28092 28540 28120 28580
rect 28258 28568 28264 28620
rect 28316 28608 28322 28620
rect 29104 28608 29132 28716
rect 31036 28676 31064 28716
rect 33137 28679 33195 28685
rect 31036 28648 33088 28676
rect 30098 28608 30104 28620
rect 28316 28580 29132 28608
rect 30059 28580 30104 28608
rect 28316 28568 28322 28580
rect 30098 28568 30104 28580
rect 30156 28568 30162 28620
rect 31570 28568 31576 28620
rect 31628 28608 31634 28620
rect 32950 28608 32956 28620
rect 31628 28580 32076 28608
rect 31628 28568 31634 28580
rect 28721 28543 28779 28549
rect 28721 28540 28733 28543
rect 28092 28512 28733 28540
rect 28721 28509 28733 28512
rect 28767 28509 28779 28543
rect 28994 28540 29000 28552
rect 28955 28512 29000 28540
rect 28721 28503 28779 28509
rect 28994 28500 29000 28512
rect 29052 28540 29058 28552
rect 30190 28540 30196 28552
rect 29052 28512 30196 28540
rect 29052 28500 29058 28512
rect 30190 28500 30196 28512
rect 30248 28500 30254 28552
rect 31938 28540 31944 28552
rect 31899 28512 31944 28540
rect 31938 28500 31944 28512
rect 31996 28500 32002 28552
rect 32048 28549 32076 28580
rect 32508 28580 32956 28608
rect 32034 28543 32092 28549
rect 32034 28509 32046 28543
rect 32080 28540 32092 28543
rect 32122 28540 32128 28552
rect 32080 28512 32128 28540
rect 32080 28509 32092 28512
rect 32034 28503 32092 28509
rect 32122 28500 32128 28512
rect 32180 28500 32186 28552
rect 32406 28543 32464 28549
rect 32406 28509 32418 28543
rect 32452 28540 32464 28543
rect 32508 28540 32536 28580
rect 32950 28568 32956 28580
rect 33008 28568 33014 28620
rect 32452 28512 32536 28540
rect 32452 28509 32464 28512
rect 32406 28503 32464 28509
rect 32582 28500 32588 28552
rect 32640 28500 32646 28552
rect 33060 28549 33088 28648
rect 33137 28645 33149 28679
rect 33183 28676 33195 28679
rect 33226 28676 33232 28688
rect 33183 28648 33232 28676
rect 33183 28645 33195 28648
rect 33137 28639 33195 28645
rect 33226 28636 33232 28648
rect 33284 28636 33290 28688
rect 33045 28543 33103 28549
rect 33045 28509 33057 28543
rect 33091 28509 33103 28543
rect 33318 28540 33324 28552
rect 33279 28512 33324 28540
rect 33045 28503 33103 28509
rect 27580 28444 27844 28472
rect 27580 28432 27586 28444
rect 29454 28432 29460 28484
rect 29512 28472 29518 28484
rect 30346 28475 30404 28481
rect 30346 28472 30358 28475
rect 29512 28444 30358 28472
rect 29512 28432 29518 28444
rect 30346 28441 30358 28444
rect 30392 28441 30404 28475
rect 30346 28435 30404 28441
rect 32217 28475 32275 28481
rect 32217 28441 32229 28475
rect 32263 28441 32275 28475
rect 32217 28435 32275 28441
rect 32309 28475 32367 28481
rect 32309 28441 32321 28475
rect 32355 28472 32367 28475
rect 32600 28472 32628 28500
rect 32355 28444 32628 28472
rect 32355 28441 32367 28444
rect 32309 28435 32367 28441
rect 27982 28404 27988 28416
rect 26988 28376 27988 28404
rect 27982 28364 27988 28376
rect 28040 28404 28046 28416
rect 28902 28404 28908 28416
rect 28040 28376 28908 28404
rect 28040 28364 28046 28376
rect 28902 28364 28908 28376
rect 28960 28364 28966 28416
rect 28994 28364 29000 28416
rect 29052 28404 29058 28416
rect 29914 28404 29920 28416
rect 29052 28376 29920 28404
rect 29052 28364 29058 28376
rect 29914 28364 29920 28376
rect 29972 28364 29978 28416
rect 31386 28364 31392 28416
rect 31444 28404 31450 28416
rect 31481 28407 31539 28413
rect 31481 28404 31493 28407
rect 31444 28376 31493 28404
rect 31444 28364 31450 28376
rect 31481 28373 31493 28376
rect 31527 28373 31539 28407
rect 31481 28367 31539 28373
rect 32030 28364 32036 28416
rect 32088 28404 32094 28416
rect 32232 28404 32260 28435
rect 32088 28376 32260 28404
rect 32585 28407 32643 28413
rect 32088 28364 32094 28376
rect 32585 28373 32597 28407
rect 32631 28404 32643 28407
rect 32766 28404 32772 28416
rect 32631 28376 32772 28404
rect 32631 28373 32643 28376
rect 32585 28367 32643 28373
rect 32766 28364 32772 28376
rect 32824 28364 32830 28416
rect 33060 28404 33088 28503
rect 33318 28500 33324 28512
rect 33376 28500 33382 28552
rect 33597 28543 33655 28549
rect 33597 28509 33609 28543
rect 33643 28509 33655 28543
rect 33778 28540 33784 28552
rect 33739 28512 33784 28540
rect 33597 28503 33655 28509
rect 33612 28472 33640 28503
rect 33778 28500 33784 28512
rect 33836 28500 33842 28552
rect 33686 28472 33692 28484
rect 33612 28444 33692 28472
rect 33686 28432 33692 28444
rect 33744 28432 33750 28484
rect 33502 28404 33508 28416
rect 33060 28376 33508 28404
rect 33502 28364 33508 28376
rect 33560 28364 33566 28416
rect 1104 28314 34868 28336
rect 1104 28262 12214 28314
rect 12266 28262 12278 28314
rect 12330 28262 12342 28314
rect 12394 28262 12406 28314
rect 12458 28262 12470 28314
rect 12522 28262 23478 28314
rect 23530 28262 23542 28314
rect 23594 28262 23606 28314
rect 23658 28262 23670 28314
rect 23722 28262 23734 28314
rect 23786 28262 34868 28314
rect 1104 28240 34868 28262
rect 13262 28200 13268 28212
rect 13223 28172 13268 28200
rect 13262 28160 13268 28172
rect 13320 28160 13326 28212
rect 17313 28203 17371 28209
rect 17313 28200 17325 28203
rect 13740 28172 17325 28200
rect 13449 28067 13507 28073
rect 13449 28033 13461 28067
rect 13495 28064 13507 28067
rect 13740 28064 13768 28172
rect 17313 28169 17325 28172
rect 17359 28169 17371 28203
rect 17313 28163 17371 28169
rect 17402 28160 17408 28212
rect 17460 28200 17466 28212
rect 20254 28200 20260 28212
rect 17460 28172 20260 28200
rect 17460 28160 17466 28172
rect 20254 28160 20260 28172
rect 20312 28160 20318 28212
rect 21266 28200 21272 28212
rect 21227 28172 21272 28200
rect 21266 28160 21272 28172
rect 21324 28160 21330 28212
rect 21910 28160 21916 28212
rect 21968 28200 21974 28212
rect 22370 28200 22376 28212
rect 21968 28172 22376 28200
rect 21968 28160 21974 28172
rect 22370 28160 22376 28172
rect 22428 28160 22434 28212
rect 23014 28200 23020 28212
rect 22480 28172 23020 28200
rect 22480 28144 22508 28172
rect 23014 28160 23020 28172
rect 23072 28160 23078 28212
rect 23934 28200 23940 28212
rect 23895 28172 23940 28200
rect 23934 28160 23940 28172
rect 23992 28200 23998 28212
rect 26142 28200 26148 28212
rect 23992 28172 26148 28200
rect 23992 28160 23998 28172
rect 26142 28160 26148 28172
rect 26200 28160 26206 28212
rect 26326 28200 26332 28212
rect 26287 28172 26332 28200
rect 26326 28160 26332 28172
rect 26384 28160 26390 28212
rect 26973 28203 27031 28209
rect 26973 28169 26985 28203
rect 27019 28200 27031 28203
rect 27246 28200 27252 28212
rect 27019 28172 27252 28200
rect 27019 28169 27031 28172
rect 26973 28163 27031 28169
rect 27246 28160 27252 28172
rect 27304 28160 27310 28212
rect 27338 28160 27344 28212
rect 27396 28200 27402 28212
rect 31386 28200 31392 28212
rect 27396 28172 31392 28200
rect 27396 28160 27402 28172
rect 31386 28160 31392 28172
rect 31444 28160 31450 28212
rect 13814 28092 13820 28144
rect 13872 28132 13878 28144
rect 13872 28104 14596 28132
rect 13872 28092 13878 28104
rect 14568 28076 14596 28104
rect 14642 28092 14648 28144
rect 14700 28132 14706 28144
rect 14700 28104 14745 28132
rect 14700 28092 14706 28104
rect 15102 28092 15108 28144
rect 15160 28132 15166 28144
rect 16025 28135 16083 28141
rect 15160 28104 15884 28132
rect 15160 28092 15166 28104
rect 13495 28036 13768 28064
rect 13909 28067 13967 28073
rect 13495 28033 13507 28036
rect 13449 28027 13507 28033
rect 13909 28033 13921 28067
rect 13955 28064 13967 28067
rect 13998 28064 14004 28076
rect 13955 28036 14004 28064
rect 13955 28033 13967 28036
rect 13909 28027 13967 28033
rect 13998 28024 14004 28036
rect 14056 28024 14062 28076
rect 14093 28067 14151 28073
rect 14093 28033 14105 28067
rect 14139 28064 14151 28067
rect 14458 28064 14464 28076
rect 14139 28036 14464 28064
rect 14139 28033 14151 28036
rect 14093 28027 14151 28033
rect 14458 28024 14464 28036
rect 14516 28024 14522 28076
rect 14550 28024 14556 28076
rect 14608 28064 14614 28076
rect 14737 28067 14795 28073
rect 14608 28036 14701 28064
rect 14608 28024 14614 28036
rect 14737 28033 14749 28067
rect 14783 28064 14795 28067
rect 14918 28064 14924 28076
rect 14783 28036 14924 28064
rect 14783 28033 14795 28036
rect 14737 28027 14795 28033
rect 14918 28024 14924 28036
rect 14976 28024 14982 28076
rect 15194 28064 15200 28076
rect 15155 28036 15200 28064
rect 15194 28024 15200 28036
rect 15252 28024 15258 28076
rect 15289 28067 15347 28073
rect 15289 28033 15301 28067
rect 15335 28064 15347 28067
rect 15746 28064 15752 28076
rect 15335 28036 15752 28064
rect 15335 28033 15347 28036
rect 15289 28027 15347 28033
rect 15746 28024 15752 28036
rect 15804 28024 15810 28076
rect 15856 28073 15884 28104
rect 16025 28101 16037 28135
rect 16071 28132 16083 28135
rect 16206 28132 16212 28144
rect 16071 28104 16212 28132
rect 16071 28101 16083 28104
rect 16025 28095 16083 28101
rect 16206 28092 16212 28104
rect 16264 28092 16270 28144
rect 16666 28092 16672 28144
rect 16724 28132 16730 28144
rect 18294 28135 18352 28141
rect 18294 28132 18306 28135
rect 16724 28104 18306 28132
rect 16724 28092 16730 28104
rect 18294 28101 18306 28104
rect 18340 28101 18352 28135
rect 18294 28095 18352 28101
rect 18506 28092 18512 28144
rect 18564 28132 18570 28144
rect 18874 28132 18880 28144
rect 18564 28104 18880 28132
rect 18564 28092 18570 28104
rect 18874 28092 18880 28104
rect 18932 28092 18938 28144
rect 19058 28092 19064 28144
rect 19116 28132 19122 28144
rect 20156 28135 20214 28141
rect 19116 28104 20024 28132
rect 19116 28092 19122 28104
rect 15841 28067 15899 28073
rect 15841 28033 15853 28067
rect 15887 28033 15899 28067
rect 16114 28064 16120 28076
rect 16027 28036 16120 28064
rect 15841 28027 15899 28033
rect 16108 28024 16120 28036
rect 16172 28024 16178 28076
rect 16298 28024 16304 28076
rect 16356 28064 16362 28076
rect 16356 28036 17080 28064
rect 16356 28024 16362 28036
rect 14182 27956 14188 28008
rect 14240 27996 14246 28008
rect 15212 27996 15240 28024
rect 14240 27968 15240 27996
rect 14240 27956 14246 27968
rect 14550 27888 14556 27940
rect 14608 27928 14614 27940
rect 16108 27928 16136 28024
rect 16758 27956 16764 28008
rect 16816 27996 16822 28008
rect 16945 27999 17003 28005
rect 16945 27996 16957 27999
rect 16816 27968 16957 27996
rect 16816 27956 16822 27968
rect 16945 27965 16957 27968
rect 16991 27965 17003 27999
rect 17052 27996 17080 28036
rect 17126 28024 17132 28076
rect 17184 28064 17190 28076
rect 17184 28036 17229 28064
rect 17184 28024 17190 28036
rect 17310 28024 17316 28076
rect 17368 28064 17374 28076
rect 18046 28064 18052 28076
rect 17368 28036 18052 28064
rect 17368 28024 17374 28036
rect 18046 28024 18052 28036
rect 18104 28024 18110 28076
rect 18156 28036 19104 28064
rect 17954 27996 17960 28008
rect 17052 27968 17960 27996
rect 16945 27959 17003 27965
rect 17954 27956 17960 27968
rect 18012 27956 18018 28008
rect 18156 27996 18184 28036
rect 18064 27968 18184 27996
rect 19076 27996 19104 28036
rect 19518 28024 19524 28076
rect 19576 28064 19582 28076
rect 19889 28067 19947 28073
rect 19889 28064 19901 28067
rect 19576 28036 19901 28064
rect 19576 28024 19582 28036
rect 19889 28033 19901 28036
rect 19935 28033 19947 28067
rect 19996 28064 20024 28104
rect 20156 28101 20168 28135
rect 20202 28132 20214 28135
rect 21082 28132 21088 28144
rect 20202 28104 21088 28132
rect 20202 28101 20214 28104
rect 20156 28095 20214 28101
rect 21082 28092 21088 28104
rect 21140 28092 21146 28144
rect 22005 28135 22063 28141
rect 22005 28101 22017 28135
rect 22051 28132 22063 28135
rect 22462 28132 22468 28144
rect 22051 28104 22468 28132
rect 22051 28101 22063 28104
rect 22005 28095 22063 28101
rect 22462 28092 22468 28104
rect 22520 28092 22526 28144
rect 22554 28092 22560 28144
rect 22612 28132 22618 28144
rect 24118 28132 24124 28144
rect 22612 28104 24124 28132
rect 22612 28092 22618 28104
rect 24118 28092 24124 28104
rect 24176 28092 24182 28144
rect 24305 28135 24363 28141
rect 24305 28101 24317 28135
rect 24351 28132 24363 28135
rect 24394 28132 24400 28144
rect 24351 28104 24400 28132
rect 24351 28101 24363 28104
rect 24305 28095 24363 28101
rect 24394 28092 24400 28104
rect 24452 28092 24458 28144
rect 24486 28092 24492 28144
rect 24544 28132 24550 28144
rect 24544 28104 25084 28132
rect 24544 28092 24550 28104
rect 19996 28036 22031 28064
rect 19889 28027 19947 28033
rect 19794 27996 19800 28008
rect 19076 27968 19800 27996
rect 14608 27900 16136 27928
rect 14608 27888 14614 27900
rect 16390 27888 16396 27940
rect 16448 27928 16454 27940
rect 16448 27900 17448 27928
rect 16448 27888 16454 27900
rect 13909 27863 13967 27869
rect 13909 27829 13921 27863
rect 13955 27860 13967 27863
rect 15746 27860 15752 27872
rect 13955 27832 15752 27860
rect 13955 27829 13967 27832
rect 13909 27823 13967 27829
rect 15746 27820 15752 27832
rect 15804 27820 15810 27872
rect 15841 27863 15899 27869
rect 15841 27829 15853 27863
rect 15887 27860 15899 27863
rect 17310 27860 17316 27872
rect 15887 27832 17316 27860
rect 15887 27829 15899 27832
rect 15841 27823 15899 27829
rect 17310 27820 17316 27832
rect 17368 27820 17374 27872
rect 17420 27860 17448 27900
rect 17586 27888 17592 27940
rect 17644 27928 17650 27940
rect 18064 27928 18092 27968
rect 19794 27956 19800 27968
rect 19852 27956 19858 28008
rect 21174 27956 21180 28008
rect 21232 27996 21238 28008
rect 21910 27996 21916 28008
rect 21232 27968 21916 27996
rect 21232 27956 21238 27968
rect 21910 27956 21916 27968
rect 21968 27956 21974 28008
rect 22003 27996 22031 28036
rect 22094 28024 22100 28076
rect 22152 28064 22158 28076
rect 22189 28067 22247 28073
rect 22189 28064 22201 28067
rect 22152 28036 22201 28064
rect 22152 28024 22158 28036
rect 22189 28033 22201 28036
rect 22235 28033 22247 28067
rect 22189 28027 22247 28033
rect 22278 28024 22284 28076
rect 22336 28064 22342 28076
rect 22738 28064 22744 28076
rect 22336 28036 22381 28064
rect 22699 28036 22744 28064
rect 22336 28024 22342 28036
rect 22738 28024 22744 28036
rect 22796 28024 22802 28076
rect 22830 28024 22836 28076
rect 22888 28064 22894 28076
rect 23014 28064 23020 28076
rect 22888 28036 22933 28064
rect 22975 28036 23020 28064
rect 22888 28024 22894 28036
rect 23014 28024 23020 28036
rect 23072 28024 23078 28076
rect 23106 28024 23112 28076
rect 23164 28064 23170 28076
rect 23247 28067 23305 28073
rect 23164 28036 23209 28064
rect 23164 28024 23170 28036
rect 23247 28033 23259 28067
rect 23293 28064 23305 28067
rect 23474 28064 23480 28076
rect 23293 28036 23480 28064
rect 23293 28033 23305 28036
rect 23247 28027 23305 28033
rect 23474 28024 23480 28036
rect 23532 28024 23538 28076
rect 23842 28064 23848 28076
rect 23803 28036 23848 28064
rect 23842 28024 23848 28036
rect 23900 28024 23906 28076
rect 24578 28064 24584 28076
rect 23952 28036 24584 28064
rect 23952 27996 23980 28036
rect 24578 28024 24584 28036
rect 24636 28024 24642 28076
rect 24670 28024 24676 28076
rect 24728 28064 24734 28076
rect 24765 28067 24823 28073
rect 24765 28064 24777 28067
rect 24728 28036 24777 28064
rect 24728 28024 24734 28036
rect 24765 28033 24777 28036
rect 24811 28033 24823 28067
rect 24946 28064 24952 28076
rect 24907 28036 24952 28064
rect 24765 28027 24823 28033
rect 24946 28024 24952 28036
rect 25004 28024 25010 28076
rect 25056 28073 25084 28104
rect 28074 28092 28080 28144
rect 28132 28132 28138 28144
rect 28132 28104 29316 28132
rect 28132 28092 28138 28104
rect 25041 28067 25099 28073
rect 25041 28033 25053 28067
rect 25087 28033 25099 28067
rect 25314 28064 25320 28076
rect 25275 28036 25320 28064
rect 25041 28027 25099 28033
rect 25314 28024 25320 28036
rect 25372 28024 25378 28076
rect 26145 28067 26203 28073
rect 26145 28033 26157 28067
rect 26191 28033 26203 28067
rect 26145 28027 26203 28033
rect 22003 27968 23980 27996
rect 24213 27999 24271 28005
rect 24213 27965 24225 27999
rect 24259 27996 24271 27999
rect 24302 27996 24308 28008
rect 24259 27968 24308 27996
rect 24259 27965 24271 27968
rect 24213 27959 24271 27965
rect 24302 27956 24308 27968
rect 24360 27956 24366 28008
rect 25130 27956 25136 28008
rect 25188 27996 25194 28008
rect 25188 27968 25233 27996
rect 25188 27956 25194 27968
rect 25406 27956 25412 28008
rect 25464 27996 25470 28008
rect 25961 27999 26019 28005
rect 25961 27996 25973 27999
rect 25464 27968 25973 27996
rect 25464 27956 25470 27968
rect 25961 27965 25973 27968
rect 26007 27965 26019 27999
rect 25961 27959 26019 27965
rect 17644 27900 18092 27928
rect 17644 27888 17650 27900
rect 19334 27888 19340 27940
rect 19392 27928 19398 27940
rect 19429 27931 19487 27937
rect 19429 27928 19441 27931
rect 19392 27900 19441 27928
rect 19392 27888 19398 27900
rect 19429 27897 19441 27900
rect 19475 27897 19487 27931
rect 19429 27891 19487 27897
rect 21818 27888 21824 27940
rect 21876 27928 21882 27940
rect 22005 27931 22063 27937
rect 22005 27928 22017 27931
rect 21876 27900 22017 27928
rect 21876 27888 21882 27900
rect 22005 27897 22017 27900
rect 22051 27897 22063 27931
rect 26160 27928 26188 28027
rect 26326 28024 26332 28076
rect 26384 28064 26390 28076
rect 27157 28067 27215 28073
rect 27157 28064 27169 28067
rect 26384 28036 27169 28064
rect 26384 28024 26390 28036
rect 27157 28033 27169 28036
rect 27203 28033 27215 28067
rect 27157 28027 27215 28033
rect 27249 28067 27307 28073
rect 27249 28033 27261 28067
rect 27295 28033 27307 28067
rect 27522 28064 27528 28076
rect 27483 28036 27528 28064
rect 27249 28027 27307 28033
rect 26234 27956 26240 28008
rect 26292 27996 26298 28008
rect 27264 27996 27292 28027
rect 27522 28024 27528 28036
rect 27580 28024 27586 28076
rect 28528 28067 28586 28073
rect 28528 28033 28540 28067
rect 28574 28064 28586 28067
rect 28810 28064 28816 28076
rect 28574 28036 28816 28064
rect 28574 28033 28586 28036
rect 28528 28027 28586 28033
rect 28810 28024 28816 28036
rect 28868 28024 28874 28076
rect 26292 27968 27292 27996
rect 26292 27956 26298 27968
rect 27706 27956 27712 28008
rect 27764 27996 27770 28008
rect 28261 27999 28319 28005
rect 28261 27996 28273 27999
rect 27764 27968 28273 27996
rect 27764 27956 27770 27968
rect 28261 27965 28273 27968
rect 28307 27965 28319 27999
rect 29288 27996 29316 28104
rect 29638 28092 29644 28144
rect 29696 28132 29702 28144
rect 32493 28135 32551 28141
rect 32493 28132 32505 28135
rect 29696 28104 30604 28132
rect 29696 28092 29702 28104
rect 29914 28024 29920 28076
rect 29972 28064 29978 28076
rect 30285 28067 30343 28073
rect 30285 28064 30297 28067
rect 29972 28036 30297 28064
rect 29972 28024 29978 28036
rect 30285 28033 30297 28036
rect 30331 28033 30343 28067
rect 30285 28027 30343 28033
rect 30374 28024 30380 28076
rect 30432 28064 30438 28076
rect 30576 28073 30604 28104
rect 31726 28104 32505 28132
rect 30561 28067 30619 28073
rect 30432 28036 30477 28064
rect 30432 28024 30438 28036
rect 30561 28033 30573 28067
rect 30607 28033 30619 28067
rect 30561 28027 30619 28033
rect 30653 28067 30711 28073
rect 30653 28033 30665 28067
rect 30699 28033 30711 28067
rect 30653 28027 30711 28033
rect 30668 27996 30696 28027
rect 30742 28024 30748 28076
rect 30800 28064 30806 28076
rect 31018 28064 31024 28076
rect 30800 28036 31024 28064
rect 30800 28024 30806 28036
rect 31018 28024 31024 28036
rect 31076 28064 31082 28076
rect 31113 28067 31171 28073
rect 31113 28064 31125 28067
rect 31076 28036 31125 28064
rect 31076 28024 31082 28036
rect 31113 28033 31125 28036
rect 31159 28033 31171 28067
rect 31113 28027 31171 28033
rect 29288 27968 30696 27996
rect 28261 27959 28319 27965
rect 22005 27891 22063 27897
rect 22103 27900 26188 27928
rect 27433 27931 27491 27937
rect 22103 27860 22131 27900
rect 27433 27897 27445 27931
rect 27479 27928 27491 27931
rect 27890 27928 27896 27940
rect 27479 27900 27896 27928
rect 27479 27897 27491 27900
rect 27433 27891 27491 27897
rect 27890 27888 27896 27900
rect 27948 27888 27954 27940
rect 29546 27888 29552 27940
rect 29604 27928 29610 27940
rect 29641 27931 29699 27937
rect 29641 27928 29653 27931
rect 29604 27900 29653 27928
rect 29604 27888 29610 27900
rect 29641 27897 29653 27900
rect 29687 27928 29699 27931
rect 29914 27928 29920 27940
rect 29687 27900 29920 27928
rect 29687 27897 29699 27900
rect 29641 27891 29699 27897
rect 29914 27888 29920 27900
rect 29972 27888 29978 27940
rect 30101 27931 30159 27937
rect 30101 27897 30113 27931
rect 30147 27928 30159 27931
rect 30190 27928 30196 27940
rect 30147 27900 30196 27928
rect 30147 27897 30159 27900
rect 30101 27891 30159 27897
rect 30190 27888 30196 27900
rect 30248 27888 30254 27940
rect 31726 27928 31754 28104
rect 32493 28101 32505 28104
rect 32539 28101 32551 28135
rect 32493 28095 32551 28101
rect 32306 28064 32312 28076
rect 32267 28036 32312 28064
rect 32306 28024 32312 28036
rect 32364 28024 32370 28076
rect 34146 27996 34152 28008
rect 34107 27968 34152 27996
rect 34146 27956 34152 27968
rect 34204 27956 34210 28008
rect 30760 27900 31754 27928
rect 23382 27860 23388 27872
rect 17420 27832 22131 27860
rect 23343 27832 23388 27860
rect 23382 27820 23388 27832
rect 23440 27820 23446 27872
rect 24118 27860 24124 27872
rect 24079 27832 24124 27860
rect 24118 27820 24124 27832
rect 24176 27820 24182 27872
rect 25501 27863 25559 27869
rect 25501 27829 25513 27863
rect 25547 27860 25559 27863
rect 25866 27860 25872 27872
rect 25547 27832 25872 27860
rect 25547 27829 25559 27832
rect 25501 27823 25559 27829
rect 25866 27820 25872 27832
rect 25924 27820 25930 27872
rect 27798 27820 27804 27872
rect 27856 27860 27862 27872
rect 30760 27860 30788 27900
rect 31294 27860 31300 27872
rect 27856 27832 30788 27860
rect 31255 27832 31300 27860
rect 27856 27820 27862 27832
rect 31294 27820 31300 27832
rect 31352 27820 31358 27872
rect 31478 27820 31484 27872
rect 31536 27860 31542 27872
rect 31573 27863 31631 27869
rect 31573 27860 31585 27863
rect 31536 27832 31585 27860
rect 31536 27820 31542 27832
rect 31573 27829 31585 27832
rect 31619 27829 31631 27863
rect 31573 27823 31631 27829
rect 31754 27820 31760 27872
rect 31812 27860 31818 27872
rect 32858 27860 32864 27872
rect 31812 27832 32864 27860
rect 31812 27820 31818 27832
rect 32858 27820 32864 27832
rect 32916 27820 32922 27872
rect 1104 27770 34868 27792
rect 1104 27718 6582 27770
rect 6634 27718 6646 27770
rect 6698 27718 6710 27770
rect 6762 27718 6774 27770
rect 6826 27718 6838 27770
rect 6890 27718 17846 27770
rect 17898 27718 17910 27770
rect 17962 27718 17974 27770
rect 18026 27718 18038 27770
rect 18090 27718 18102 27770
rect 18154 27718 29110 27770
rect 29162 27718 29174 27770
rect 29226 27718 29238 27770
rect 29290 27718 29302 27770
rect 29354 27718 29366 27770
rect 29418 27718 34868 27770
rect 1104 27696 34868 27718
rect 14458 27616 14464 27668
rect 14516 27656 14522 27668
rect 14516 27628 18368 27656
rect 14516 27616 14522 27628
rect 13357 27591 13415 27597
rect 13357 27557 13369 27591
rect 13403 27588 13415 27591
rect 15010 27588 15016 27600
rect 13403 27560 15016 27588
rect 13403 27557 13415 27560
rect 13357 27551 13415 27557
rect 15010 27548 15016 27560
rect 15068 27548 15074 27600
rect 15746 27548 15752 27600
rect 15804 27588 15810 27600
rect 18046 27588 18052 27600
rect 15804 27560 18052 27588
rect 15804 27548 15810 27560
rect 18046 27548 18052 27560
rect 18104 27548 18110 27600
rect 18340 27588 18368 27628
rect 18414 27616 18420 27668
rect 18472 27656 18478 27668
rect 19245 27659 19303 27665
rect 19245 27656 19257 27659
rect 18472 27628 19257 27656
rect 18472 27616 18478 27628
rect 19245 27625 19257 27628
rect 19291 27625 19303 27659
rect 19245 27619 19303 27625
rect 19886 27616 19892 27668
rect 19944 27656 19950 27668
rect 22186 27656 22192 27668
rect 19944 27628 22192 27656
rect 19944 27616 19950 27628
rect 22186 27616 22192 27628
rect 22244 27616 22250 27668
rect 22370 27616 22376 27668
rect 22428 27656 22434 27668
rect 26234 27656 26240 27668
rect 22428 27628 26240 27656
rect 22428 27616 22434 27628
rect 26234 27616 26240 27628
rect 26292 27616 26298 27668
rect 26513 27659 26571 27665
rect 26513 27625 26525 27659
rect 26559 27656 26571 27659
rect 27430 27656 27436 27668
rect 26559 27628 27436 27656
rect 26559 27625 26571 27628
rect 26513 27619 26571 27625
rect 27430 27616 27436 27628
rect 27488 27616 27494 27668
rect 28258 27656 28264 27668
rect 28092 27628 28264 27656
rect 18506 27588 18512 27600
rect 18340 27560 18512 27588
rect 18506 27548 18512 27560
rect 18564 27548 18570 27600
rect 19705 27591 19763 27597
rect 19705 27588 19717 27591
rect 18616 27560 19717 27588
rect 14737 27523 14795 27529
rect 14737 27489 14749 27523
rect 14783 27520 14795 27523
rect 15930 27520 15936 27532
rect 14783 27492 15936 27520
rect 14783 27489 14795 27492
rect 14737 27483 14795 27489
rect 15930 27480 15936 27492
rect 15988 27480 15994 27532
rect 16117 27523 16175 27529
rect 16117 27489 16129 27523
rect 16163 27520 16175 27523
rect 16669 27523 16727 27529
rect 16163 27492 16589 27520
rect 16163 27489 16175 27492
rect 16117 27483 16175 27489
rect 13541 27455 13599 27461
rect 13541 27421 13553 27455
rect 13587 27421 13599 27455
rect 13541 27415 13599 27421
rect 13556 27316 13584 27415
rect 14366 27412 14372 27464
rect 14424 27452 14430 27464
rect 14645 27455 14703 27461
rect 14645 27452 14657 27455
rect 14424 27424 14657 27452
rect 14424 27412 14430 27424
rect 14645 27421 14657 27424
rect 14691 27421 14703 27455
rect 14645 27415 14703 27421
rect 14829 27455 14887 27461
rect 14829 27421 14841 27455
rect 14875 27452 14887 27455
rect 14918 27452 14924 27464
rect 14875 27424 14924 27452
rect 14875 27421 14887 27424
rect 14829 27415 14887 27421
rect 14918 27412 14924 27424
rect 14976 27412 14982 27464
rect 15194 27412 15200 27464
rect 15252 27452 15258 27464
rect 15289 27455 15347 27461
rect 15289 27452 15301 27455
rect 15252 27424 15301 27452
rect 15252 27412 15258 27424
rect 15289 27421 15301 27424
rect 15335 27421 15347 27455
rect 15289 27415 15347 27421
rect 15473 27455 15531 27461
rect 15473 27421 15485 27455
rect 15519 27452 15531 27455
rect 15562 27452 15568 27464
rect 15519 27424 15568 27452
rect 15519 27421 15531 27424
rect 15473 27415 15531 27421
rect 15562 27412 15568 27424
rect 15620 27452 15626 27464
rect 15746 27452 15752 27464
rect 15620 27424 15752 27452
rect 15620 27412 15626 27424
rect 15746 27412 15752 27424
rect 15804 27412 15810 27464
rect 16025 27455 16083 27461
rect 16025 27421 16037 27455
rect 16071 27452 16083 27455
rect 16206 27452 16212 27464
rect 16071 27424 16212 27452
rect 16071 27421 16083 27424
rect 16025 27415 16083 27421
rect 16206 27412 16212 27424
rect 16264 27412 16270 27464
rect 13722 27344 13728 27396
rect 13780 27384 13786 27396
rect 16298 27384 16304 27396
rect 13780 27356 16304 27384
rect 13780 27344 13786 27356
rect 16298 27344 16304 27356
rect 16356 27344 16362 27396
rect 15286 27316 15292 27328
rect 13556 27288 15292 27316
rect 15286 27276 15292 27288
rect 15344 27276 15350 27328
rect 15381 27319 15439 27325
rect 15381 27285 15393 27319
rect 15427 27316 15439 27319
rect 15654 27316 15660 27328
rect 15427 27288 15660 27316
rect 15427 27285 15439 27288
rect 15381 27279 15439 27285
rect 15654 27276 15660 27288
rect 15712 27276 15718 27328
rect 16561 27316 16589 27492
rect 16669 27489 16681 27523
rect 16715 27520 16727 27523
rect 17402 27520 17408 27532
rect 16715 27492 17408 27520
rect 16715 27489 16727 27492
rect 16669 27483 16727 27489
rect 17402 27480 17408 27492
rect 17460 27480 17466 27532
rect 17497 27523 17555 27529
rect 17497 27489 17509 27523
rect 17543 27520 17555 27523
rect 17586 27520 17592 27532
rect 17543 27492 17592 27520
rect 17543 27489 17555 27492
rect 17497 27483 17555 27489
rect 17586 27480 17592 27492
rect 17644 27480 17650 27532
rect 18414 27520 18420 27532
rect 17696 27492 18420 27520
rect 16853 27455 16911 27461
rect 16853 27421 16865 27455
rect 16899 27452 16911 27455
rect 17126 27452 17132 27464
rect 16899 27424 17132 27452
rect 16899 27421 16911 27424
rect 16853 27415 16911 27421
rect 17126 27412 17132 27424
rect 17184 27452 17190 27464
rect 17696 27461 17724 27492
rect 18414 27480 18420 27492
rect 18472 27480 18478 27532
rect 17681 27455 17739 27461
rect 17681 27452 17693 27455
rect 17184 27424 17693 27452
rect 17184 27412 17190 27424
rect 17681 27421 17693 27424
rect 17727 27421 17739 27455
rect 17681 27415 17739 27421
rect 18325 27455 18383 27461
rect 18325 27421 18337 27455
rect 18371 27452 18383 27455
rect 18616 27452 18644 27560
rect 19705 27557 19717 27560
rect 19751 27557 19763 27591
rect 19705 27551 19763 27557
rect 20806 27548 20812 27600
rect 20864 27548 20870 27600
rect 22646 27588 22652 27600
rect 21560 27560 22652 27588
rect 19426 27520 19432 27532
rect 19387 27492 19432 27520
rect 19426 27480 19432 27492
rect 19484 27480 19490 27532
rect 19610 27480 19616 27532
rect 19668 27520 19674 27532
rect 20824 27520 20852 27548
rect 21560 27520 21588 27560
rect 22646 27548 22652 27560
rect 22704 27548 22710 27600
rect 23474 27588 23480 27600
rect 23387 27560 23480 27588
rect 21726 27520 21732 27532
rect 19668 27492 20852 27520
rect 21192 27492 21588 27520
rect 21687 27492 21732 27520
rect 19668 27480 19674 27492
rect 18371 27424 18644 27452
rect 18371 27421 18383 27424
rect 18325 27415 18383 27421
rect 18966 27412 18972 27464
rect 19024 27452 19030 27464
rect 19521 27455 19579 27461
rect 19521 27452 19533 27455
rect 19024 27424 19533 27452
rect 19024 27412 19030 27424
rect 19521 27421 19533 27424
rect 19567 27421 19579 27455
rect 19521 27415 19579 27421
rect 20806 27412 20812 27464
rect 20864 27448 20870 27464
rect 20901 27455 20959 27461
rect 20901 27448 20913 27455
rect 20864 27421 20913 27448
rect 20947 27421 20959 27455
rect 20864 27420 20959 27421
rect 20864 27412 20870 27420
rect 20901 27415 20959 27420
rect 20990 27412 20996 27464
rect 21048 27452 21054 27464
rect 21192 27461 21220 27492
rect 21726 27480 21732 27492
rect 21784 27480 21790 27532
rect 23014 27520 23020 27532
rect 21836 27492 23020 27520
rect 21177 27455 21235 27461
rect 21048 27424 21093 27452
rect 21048 27412 21054 27424
rect 21177 27421 21189 27455
rect 21223 27421 21235 27455
rect 21177 27415 21235 27421
rect 21266 27412 21272 27464
rect 21324 27452 21330 27464
rect 21324 27424 21369 27452
rect 21324 27412 21330 27424
rect 16666 27344 16672 27396
rect 16724 27384 16730 27396
rect 17037 27387 17095 27393
rect 17037 27384 17049 27387
rect 16724 27356 17049 27384
rect 16724 27344 16730 27356
rect 17037 27353 17049 27356
rect 17083 27353 17095 27387
rect 17037 27347 17095 27353
rect 17586 27344 17592 27396
rect 17644 27384 17650 27396
rect 17865 27387 17923 27393
rect 17865 27384 17877 27387
rect 17644 27356 17877 27384
rect 17644 27344 17650 27356
rect 17865 27353 17877 27356
rect 17911 27353 17923 27387
rect 18506 27384 18512 27396
rect 18467 27356 18512 27384
rect 17865 27347 17923 27353
rect 18506 27344 18512 27356
rect 18564 27344 18570 27396
rect 18616 27356 19104 27384
rect 17954 27316 17960 27328
rect 16561 27288 17960 27316
rect 17954 27276 17960 27288
rect 18012 27276 18018 27328
rect 18046 27276 18052 27328
rect 18104 27316 18110 27328
rect 18616 27316 18644 27356
rect 18104 27288 18644 27316
rect 18693 27319 18751 27325
rect 18104 27276 18110 27288
rect 18693 27285 18705 27319
rect 18739 27316 18751 27319
rect 18966 27316 18972 27328
rect 18739 27288 18972 27316
rect 18739 27285 18751 27288
rect 18693 27279 18751 27285
rect 18966 27276 18972 27288
rect 19024 27276 19030 27328
rect 19076 27316 19104 27356
rect 19150 27344 19156 27396
rect 19208 27384 19214 27396
rect 19245 27387 19303 27393
rect 19245 27384 19257 27387
rect 19208 27356 19257 27384
rect 19208 27344 19214 27356
rect 19245 27353 19257 27356
rect 19291 27353 19303 27387
rect 21836 27384 21864 27492
rect 23014 27480 23020 27492
rect 23072 27480 23078 27532
rect 21910 27412 21916 27464
rect 21968 27412 21974 27464
rect 22005 27455 22063 27461
rect 22005 27421 22017 27455
rect 22051 27452 22063 27455
rect 22094 27452 22100 27464
rect 22051 27424 22100 27452
rect 22051 27421 22063 27424
rect 22005 27415 22063 27421
rect 22094 27412 22100 27424
rect 22152 27412 22158 27464
rect 22554 27412 22560 27464
rect 22612 27452 22618 27464
rect 23198 27452 23204 27464
rect 22612 27424 23204 27452
rect 22612 27412 22618 27424
rect 23198 27412 23204 27424
rect 23256 27412 23262 27464
rect 23405 27452 23433 27560
rect 23474 27548 23480 27560
rect 23532 27588 23538 27600
rect 24118 27588 24124 27600
rect 23532 27560 24124 27588
rect 23532 27548 23538 27560
rect 24118 27548 24124 27560
rect 24176 27548 24182 27600
rect 24670 27548 24676 27600
rect 24728 27588 24734 27600
rect 24949 27591 25007 27597
rect 24949 27588 24961 27591
rect 24728 27560 24961 27588
rect 24728 27548 24734 27560
rect 24949 27557 24961 27560
rect 24995 27557 25007 27591
rect 24949 27551 25007 27557
rect 26142 27548 26148 27600
rect 26200 27588 26206 27600
rect 28092 27588 28120 27628
rect 28258 27616 28264 27628
rect 28316 27616 28322 27668
rect 28828 27628 29592 27656
rect 26200 27560 28120 27588
rect 26200 27548 26206 27560
rect 28166 27548 28172 27600
rect 28224 27588 28230 27600
rect 28828 27588 28856 27628
rect 28224 27560 28856 27588
rect 28905 27591 28963 27597
rect 28224 27548 28230 27560
rect 28905 27557 28917 27591
rect 28951 27588 28963 27591
rect 29454 27588 29460 27600
rect 28951 27560 29460 27588
rect 28951 27557 28963 27560
rect 28905 27551 28963 27557
rect 29454 27548 29460 27560
rect 29512 27548 29518 27600
rect 29564 27588 29592 27628
rect 31938 27616 31944 27668
rect 31996 27656 32002 27668
rect 32309 27659 32367 27665
rect 32309 27656 32321 27659
rect 31996 27628 32321 27656
rect 31996 27616 32002 27628
rect 32309 27625 32321 27628
rect 32355 27625 32367 27659
rect 32309 27619 32367 27625
rect 33778 27616 33784 27668
rect 33836 27656 33842 27668
rect 34149 27659 34207 27665
rect 34149 27656 34161 27659
rect 33836 27628 34161 27656
rect 33836 27616 33842 27628
rect 34149 27625 34161 27628
rect 34195 27625 34207 27659
rect 34149 27619 34207 27625
rect 31662 27588 31668 27600
rect 29564 27560 31668 27588
rect 31662 27548 31668 27560
rect 31720 27548 31726 27600
rect 23750 27480 23756 27532
rect 23808 27520 23814 27532
rect 28813 27523 28871 27529
rect 28813 27520 28825 27523
rect 23808 27492 28825 27520
rect 23808 27480 23814 27492
rect 28813 27489 28825 27492
rect 28859 27489 28871 27523
rect 29546 27520 29552 27532
rect 29507 27492 29552 27520
rect 28813 27483 28871 27489
rect 29546 27480 29552 27492
rect 29604 27480 29610 27532
rect 29914 27480 29920 27532
rect 29972 27520 29978 27532
rect 30929 27523 30987 27529
rect 30929 27520 30941 27523
rect 29972 27492 30941 27520
rect 29972 27480 29978 27492
rect 30929 27489 30941 27492
rect 30975 27489 30987 27523
rect 30929 27483 30987 27489
rect 31018 27480 31024 27532
rect 31076 27520 31082 27532
rect 31113 27523 31171 27529
rect 31113 27520 31125 27523
rect 31076 27492 31125 27520
rect 31076 27480 31082 27492
rect 31113 27489 31125 27492
rect 31159 27489 31171 27523
rect 31113 27483 31171 27489
rect 31202 27480 31208 27532
rect 31260 27520 31266 27532
rect 31849 27523 31907 27529
rect 31849 27520 31861 27523
rect 31260 27492 31861 27520
rect 31260 27480 31266 27492
rect 31849 27489 31861 27492
rect 31895 27489 31907 27523
rect 31849 27483 31907 27489
rect 31941 27523 31999 27529
rect 31941 27489 31953 27523
rect 31987 27520 31999 27523
rect 32030 27520 32036 27532
rect 31987 27492 32036 27520
rect 31987 27489 31999 27492
rect 31941 27483 31999 27489
rect 32030 27480 32036 27492
rect 32088 27480 32094 27532
rect 23477 27455 23535 27461
rect 23477 27452 23489 27455
rect 23405 27424 23489 27452
rect 23477 27421 23489 27424
rect 23523 27421 23535 27455
rect 23477 27415 23535 27421
rect 23566 27412 23572 27464
rect 23624 27452 23630 27464
rect 24397 27455 24455 27461
rect 24397 27452 24409 27455
rect 23624 27424 24409 27452
rect 23624 27412 23630 27424
rect 24397 27421 24409 27424
rect 24443 27421 24455 27455
rect 24397 27415 24455 27421
rect 24486 27412 24492 27464
rect 24544 27452 24550 27464
rect 24673 27455 24731 27461
rect 24673 27452 24685 27455
rect 24544 27424 24685 27452
rect 24544 27412 24550 27424
rect 24673 27421 24685 27424
rect 24719 27421 24731 27455
rect 24673 27415 24731 27421
rect 24765 27455 24823 27461
rect 24765 27421 24777 27455
rect 24811 27452 24823 27455
rect 24946 27452 24952 27464
rect 24811 27424 24952 27452
rect 24811 27421 24823 27424
rect 24765 27415 24823 27421
rect 24946 27412 24952 27424
rect 25004 27412 25010 27464
rect 25866 27452 25872 27464
rect 25827 27424 25872 27452
rect 25866 27412 25872 27424
rect 25924 27412 25930 27464
rect 25958 27412 25964 27464
rect 26016 27452 26022 27464
rect 26234 27452 26240 27464
rect 26016 27424 26061 27452
rect 26195 27424 26240 27452
rect 26016 27412 26022 27424
rect 26234 27412 26240 27424
rect 26292 27412 26298 27464
rect 26326 27412 26332 27464
rect 26384 27461 26390 27464
rect 26384 27452 26392 27461
rect 26384 27424 26429 27452
rect 26384 27415 26392 27424
rect 26384 27412 26390 27415
rect 27246 27412 27252 27464
rect 27304 27452 27310 27464
rect 27304 27424 27349 27452
rect 27304 27412 27310 27424
rect 27430 27412 27436 27464
rect 27488 27452 27494 27464
rect 27709 27455 27767 27461
rect 27709 27452 27721 27455
rect 27488 27424 27721 27452
rect 27488 27412 27494 27424
rect 27709 27421 27721 27424
rect 27755 27421 27767 27455
rect 27709 27415 27767 27421
rect 28537 27455 28595 27461
rect 28537 27421 28549 27455
rect 28583 27452 28595 27455
rect 28718 27452 28724 27464
rect 28583 27424 28724 27452
rect 28583 27421 28595 27424
rect 28537 27415 28595 27421
rect 28718 27412 28724 27424
rect 28776 27412 28782 27464
rect 28902 27452 28908 27464
rect 28863 27424 28908 27452
rect 28902 27412 28908 27424
rect 28960 27412 28966 27464
rect 29270 27412 29276 27464
rect 29328 27452 29334 27464
rect 29825 27455 29883 27461
rect 29825 27452 29837 27455
rect 29328 27424 29837 27452
rect 29328 27412 29334 27424
rect 29825 27421 29837 27424
rect 29871 27452 29883 27455
rect 30098 27452 30104 27464
rect 29871 27424 30104 27452
rect 29871 27421 29883 27424
rect 29825 27415 29883 27421
rect 30098 27412 30104 27424
rect 30156 27412 30162 27464
rect 30282 27412 30288 27464
rect 30340 27452 30346 27464
rect 30837 27455 30895 27461
rect 30837 27452 30849 27455
rect 30340 27424 30849 27452
rect 30340 27412 30346 27424
rect 30837 27421 30849 27424
rect 30883 27421 30895 27455
rect 31570 27452 31576 27464
rect 31531 27424 31576 27452
rect 30837 27415 30895 27421
rect 31570 27412 31576 27424
rect 31628 27412 31634 27464
rect 31754 27412 31760 27464
rect 31812 27452 31818 27464
rect 32122 27452 32128 27464
rect 31812 27424 31857 27452
rect 32083 27424 32128 27452
rect 31812 27412 31818 27424
rect 32122 27412 32128 27424
rect 32180 27412 32186 27464
rect 32306 27412 32312 27464
rect 32364 27452 32370 27464
rect 32769 27455 32827 27461
rect 32769 27452 32781 27455
rect 32364 27424 32781 27452
rect 32364 27412 32370 27424
rect 32769 27421 32781 27424
rect 32815 27421 32827 27455
rect 32769 27415 32827 27421
rect 19245 27347 19303 27353
rect 20640 27356 21864 27384
rect 21928 27384 21956 27412
rect 21928 27356 22048 27384
rect 20640 27316 20668 27356
rect 19076 27288 20668 27316
rect 20717 27319 20775 27325
rect 20717 27285 20729 27319
rect 20763 27316 20775 27319
rect 21910 27316 21916 27328
rect 20763 27288 21916 27316
rect 20763 27285 20775 27288
rect 20717 27279 20775 27285
rect 21910 27276 21916 27288
rect 21968 27276 21974 27328
rect 22020 27316 22048 27356
rect 23106 27344 23112 27396
rect 23164 27384 23170 27396
rect 23661 27387 23719 27393
rect 23661 27384 23673 27387
rect 23164 27356 23673 27384
rect 23164 27344 23170 27356
rect 23661 27353 23673 27356
rect 23707 27353 23719 27387
rect 23661 27347 23719 27353
rect 23845 27387 23903 27393
rect 23845 27353 23857 27387
rect 23891 27384 23903 27387
rect 24581 27387 24639 27393
rect 24581 27384 24593 27387
rect 23891 27356 24593 27384
rect 23891 27353 23903 27356
rect 23845 27347 23903 27353
rect 24581 27353 24593 27356
rect 24627 27353 24639 27387
rect 24581 27347 24639 27353
rect 25130 27344 25136 27396
rect 25188 27384 25194 27396
rect 25774 27384 25780 27396
rect 25188 27356 25780 27384
rect 25188 27344 25194 27356
rect 25774 27344 25780 27356
rect 25832 27384 25838 27396
rect 26145 27387 26203 27393
rect 26145 27384 26157 27387
rect 25832 27356 26157 27384
rect 25832 27344 25838 27356
rect 26145 27353 26157 27356
rect 26191 27353 26203 27387
rect 26145 27347 26203 27353
rect 26970 27344 26976 27396
rect 27028 27384 27034 27396
rect 27065 27387 27123 27393
rect 27065 27384 27077 27387
rect 27028 27356 27077 27384
rect 27028 27344 27034 27356
rect 27065 27353 27077 27356
rect 27111 27353 27123 27387
rect 31113 27387 31171 27393
rect 31113 27384 31125 27387
rect 27065 27347 27123 27353
rect 27172 27356 31125 27384
rect 27172 27316 27200 27356
rect 31113 27353 31125 27356
rect 31159 27353 31171 27387
rect 31113 27347 31171 27353
rect 33036 27387 33094 27393
rect 33036 27353 33048 27387
rect 33082 27384 33094 27387
rect 33134 27384 33140 27396
rect 33082 27356 33140 27384
rect 33082 27353 33094 27356
rect 33036 27347 33094 27353
rect 33134 27344 33140 27356
rect 33192 27344 33198 27396
rect 22020 27288 27200 27316
rect 27893 27319 27951 27325
rect 27893 27285 27905 27319
rect 27939 27316 27951 27319
rect 28442 27316 28448 27328
rect 27939 27288 28448 27316
rect 27939 27285 27951 27288
rect 27893 27279 27951 27285
rect 28442 27276 28448 27288
rect 28500 27276 28506 27328
rect 28626 27316 28632 27328
rect 28587 27288 28632 27316
rect 28626 27276 28632 27288
rect 28684 27316 28690 27328
rect 33594 27316 33600 27328
rect 28684 27288 33600 27316
rect 28684 27276 28690 27288
rect 33594 27276 33600 27288
rect 33652 27276 33658 27328
rect 1104 27226 34868 27248
rect 1104 27174 12214 27226
rect 12266 27174 12278 27226
rect 12330 27174 12342 27226
rect 12394 27174 12406 27226
rect 12458 27174 12470 27226
rect 12522 27174 23478 27226
rect 23530 27174 23542 27226
rect 23594 27174 23606 27226
rect 23658 27174 23670 27226
rect 23722 27174 23734 27226
rect 23786 27174 34868 27226
rect 1104 27152 34868 27174
rect 15381 27115 15439 27121
rect 15381 27081 15393 27115
rect 15427 27112 15439 27115
rect 16942 27112 16948 27124
rect 15427 27084 16948 27112
rect 15427 27081 15439 27084
rect 15381 27075 15439 27081
rect 16942 27072 16948 27084
rect 17000 27072 17006 27124
rect 17402 27072 17408 27124
rect 17460 27112 17466 27124
rect 17589 27115 17647 27121
rect 17589 27112 17601 27115
rect 17460 27084 17601 27112
rect 17460 27072 17466 27084
rect 17589 27081 17601 27084
rect 17635 27081 17647 27115
rect 17589 27075 17647 27081
rect 17678 27072 17684 27124
rect 17736 27112 17742 27124
rect 17773 27115 17831 27121
rect 17773 27112 17785 27115
rect 17736 27084 17785 27112
rect 17736 27072 17742 27084
rect 17773 27081 17785 27084
rect 17819 27081 17831 27115
rect 17773 27075 17831 27081
rect 17862 27072 17868 27124
rect 17920 27112 17926 27124
rect 18782 27112 18788 27124
rect 17920 27084 18788 27112
rect 17920 27072 17926 27084
rect 18782 27072 18788 27084
rect 18840 27072 18846 27124
rect 19978 27112 19984 27124
rect 19076 27084 19984 27112
rect 16574 27044 16580 27056
rect 14844 27016 16580 27044
rect 13538 26976 13544 26988
rect 13499 26948 13544 26976
rect 13538 26936 13544 26948
rect 13596 26936 13602 26988
rect 14182 26976 14188 26988
rect 14143 26948 14188 26976
rect 14182 26936 14188 26948
rect 14240 26936 14246 26988
rect 14844 26985 14872 27016
rect 16574 27004 16580 27016
rect 16632 27004 16638 27056
rect 17218 27044 17224 27056
rect 16684 27016 17224 27044
rect 14829 26979 14887 26985
rect 14829 26945 14841 26979
rect 14875 26945 14887 26979
rect 14829 26939 14887 26945
rect 15289 26979 15347 26985
rect 15289 26945 15301 26979
rect 15335 26945 15347 26979
rect 15470 26976 15476 26988
rect 15431 26948 15476 26976
rect 15289 26939 15347 26945
rect 15304 26908 15332 26939
rect 15470 26936 15476 26948
rect 15528 26936 15534 26988
rect 15562 26936 15568 26988
rect 15620 26976 15626 26988
rect 15930 26976 15936 26988
rect 15620 26948 15936 26976
rect 15620 26936 15626 26948
rect 15930 26936 15936 26948
rect 15988 26936 15994 26988
rect 16025 26979 16083 26985
rect 16025 26945 16037 26979
rect 16071 26976 16083 26979
rect 16684 26976 16712 27016
rect 17218 27004 17224 27016
rect 17276 27004 17282 27056
rect 18690 27004 18696 27056
rect 18748 27044 18754 27056
rect 19076 27053 19104 27084
rect 19978 27072 19984 27084
rect 20036 27072 20042 27124
rect 20806 27072 20812 27124
rect 20864 27112 20870 27124
rect 21269 27115 21327 27121
rect 21269 27112 21281 27115
rect 20864 27084 21281 27112
rect 20864 27072 20870 27084
rect 21269 27081 21281 27084
rect 21315 27112 21327 27115
rect 21726 27112 21732 27124
rect 21315 27084 21732 27112
rect 21315 27081 21327 27084
rect 21269 27075 21327 27081
rect 21726 27072 21732 27084
rect 21784 27072 21790 27124
rect 22649 27115 22707 27121
rect 22649 27081 22661 27115
rect 22695 27112 22707 27115
rect 22738 27112 22744 27124
rect 22695 27084 22744 27112
rect 22695 27081 22707 27084
rect 22649 27075 22707 27081
rect 22738 27072 22744 27084
rect 22796 27072 22802 27124
rect 23216 27084 23428 27112
rect 18969 27047 19027 27053
rect 18969 27044 18981 27047
rect 18748 27016 18981 27044
rect 18748 27004 18754 27016
rect 18969 27013 18981 27016
rect 19015 27013 19027 27047
rect 18969 27007 19027 27013
rect 19061 27047 19119 27053
rect 19061 27013 19073 27047
rect 19107 27013 19119 27047
rect 19702 27044 19708 27056
rect 19061 27007 19119 27013
rect 19352 27016 19708 27044
rect 16071 26948 16712 26976
rect 16071 26945 16083 26948
rect 16025 26939 16083 26945
rect 16758 26936 16764 26988
rect 16816 26976 16822 26988
rect 17681 26979 17739 26985
rect 17681 26976 17693 26979
rect 16816 26948 16861 26976
rect 17144 26948 17693 26976
rect 16816 26936 16822 26948
rect 15304 26880 16712 26908
rect 14001 26843 14059 26849
rect 14001 26809 14013 26843
rect 14047 26840 14059 26843
rect 16574 26840 16580 26852
rect 14047 26812 16580 26840
rect 14047 26809 14059 26812
rect 14001 26803 14059 26809
rect 16574 26800 16580 26812
rect 16632 26800 16638 26852
rect 16684 26840 16712 26880
rect 16850 26868 16856 26920
rect 16908 26908 16914 26920
rect 17144 26908 17172 26948
rect 17681 26945 17693 26948
rect 17727 26945 17739 26979
rect 17681 26939 17739 26945
rect 17957 26979 18015 26985
rect 17957 26945 17969 26979
rect 18003 26976 18015 26979
rect 18877 26979 18935 26985
rect 18877 26976 18889 26979
rect 18003 26948 18889 26976
rect 18003 26945 18015 26948
rect 17957 26939 18015 26945
rect 18877 26945 18889 26948
rect 18923 26945 18935 26979
rect 18877 26939 18935 26945
rect 16908 26880 17172 26908
rect 16908 26868 16914 26880
rect 17218 26868 17224 26920
rect 17276 26908 17282 26920
rect 17405 26911 17463 26917
rect 17405 26908 17417 26911
rect 17276 26880 17417 26908
rect 17276 26868 17282 26880
rect 17405 26877 17417 26880
rect 17451 26877 17463 26911
rect 17405 26871 17463 26877
rect 17696 26840 17724 26939
rect 19150 26936 19156 26988
rect 19208 26985 19214 26988
rect 19352 26985 19380 27016
rect 19702 27004 19708 27016
rect 19760 27004 19766 27056
rect 21174 27044 21180 27056
rect 19812 27016 21180 27044
rect 19208 26979 19237 26985
rect 19225 26945 19237 26979
rect 19208 26939 19237 26945
rect 19337 26979 19395 26985
rect 19337 26945 19349 26979
rect 19383 26945 19395 26979
rect 19812 26976 19840 27016
rect 21174 27004 21180 27016
rect 21232 27004 21238 27056
rect 21450 27004 21456 27056
rect 21508 27044 21514 27056
rect 23216 27044 23244 27084
rect 21508 27016 23244 27044
rect 23400 27044 23428 27084
rect 24394 27072 24400 27124
rect 24452 27112 24458 27124
rect 24946 27112 24952 27124
rect 24452 27084 24952 27112
rect 24452 27072 24458 27084
rect 24946 27072 24952 27084
rect 25004 27112 25010 27124
rect 25225 27115 25283 27121
rect 25225 27112 25237 27115
rect 25004 27084 25237 27112
rect 25004 27072 25010 27084
rect 25225 27081 25237 27084
rect 25271 27081 25283 27115
rect 25225 27075 25283 27081
rect 27890 27072 27896 27124
rect 27948 27112 27954 27124
rect 28353 27115 28411 27121
rect 28353 27112 28365 27115
rect 27948 27084 28365 27112
rect 27948 27072 27954 27084
rect 28353 27081 28365 27084
rect 28399 27081 28411 27115
rect 28810 27112 28816 27124
rect 28771 27084 28816 27112
rect 28353 27075 28411 27081
rect 28810 27072 28816 27084
rect 28868 27072 28874 27124
rect 29914 27072 29920 27124
rect 29972 27072 29978 27124
rect 30098 27072 30104 27124
rect 30156 27112 30162 27124
rect 30374 27112 30380 27124
rect 30156 27084 30380 27112
rect 30156 27072 30162 27084
rect 30374 27072 30380 27084
rect 30432 27112 30438 27124
rect 30558 27112 30564 27124
rect 30432 27084 30564 27112
rect 30432 27072 30438 27084
rect 30558 27072 30564 27084
rect 30616 27072 30622 27124
rect 30926 27072 30932 27124
rect 30984 27112 30990 27124
rect 31570 27112 31576 27124
rect 30984 27084 31156 27112
rect 31531 27084 31576 27112
rect 30984 27072 30990 27084
rect 24090 27047 24148 27053
rect 24090 27044 24102 27047
rect 23400 27016 24102 27044
rect 21508 27004 21514 27016
rect 24090 27013 24102 27016
rect 24136 27013 24148 27047
rect 24090 27007 24148 27013
rect 24302 27004 24308 27056
rect 24360 27044 24366 27056
rect 29932 27044 29960 27072
rect 30190 27044 30196 27056
rect 24360 27016 29960 27044
rect 30151 27016 30196 27044
rect 24360 27004 24366 27016
rect 30190 27004 30196 27016
rect 30248 27004 30254 27056
rect 30285 27047 30343 27053
rect 30285 27013 30297 27047
rect 30331 27044 30343 27047
rect 30650 27044 30656 27056
rect 30331 27016 30656 27044
rect 30331 27013 30343 27016
rect 30285 27007 30343 27013
rect 30650 27004 30656 27016
rect 30708 27004 30714 27056
rect 19337 26939 19395 26945
rect 19444 26948 19840 26976
rect 20156 26979 20214 26985
rect 19208 26936 19214 26939
rect 18046 26868 18052 26920
rect 18104 26908 18110 26920
rect 19444 26908 19472 26948
rect 20156 26945 20168 26979
rect 20202 26976 20214 26979
rect 21082 26976 21088 26988
rect 20202 26948 21088 26976
rect 20202 26945 20214 26948
rect 20156 26939 20214 26945
rect 21082 26936 21088 26948
rect 21140 26936 21146 26988
rect 21910 26976 21916 26988
rect 21871 26948 21916 26976
rect 21910 26936 21916 26948
rect 21968 26936 21974 26988
rect 22094 26976 22100 26988
rect 22055 26948 22100 26976
rect 22094 26936 22100 26948
rect 22152 26976 22158 26988
rect 22465 26979 22523 26985
rect 22152 26948 22427 26976
rect 22152 26936 22158 26948
rect 18104 26880 19472 26908
rect 18104 26868 18110 26880
rect 19518 26868 19524 26920
rect 19576 26908 19582 26920
rect 19886 26908 19892 26920
rect 19576 26880 19892 26908
rect 19576 26868 19582 26880
rect 19886 26868 19892 26880
rect 19944 26868 19950 26920
rect 20990 26868 20996 26920
rect 21048 26908 21054 26920
rect 22189 26911 22247 26917
rect 22189 26908 22201 26911
rect 21048 26880 22201 26908
rect 21048 26868 21054 26880
rect 22189 26877 22201 26880
rect 22235 26877 22247 26911
rect 22189 26871 22247 26877
rect 22281 26911 22339 26917
rect 22281 26877 22293 26911
rect 22327 26877 22339 26911
rect 22399 26908 22427 26948
rect 22465 26945 22477 26979
rect 22511 26976 22523 26979
rect 22830 26976 22836 26988
rect 22511 26948 22836 26976
rect 22511 26945 22523 26948
rect 22465 26939 22523 26945
rect 22830 26936 22836 26948
rect 22888 26936 22894 26988
rect 22922 26936 22928 26988
rect 22980 26976 22986 26988
rect 23109 26979 23167 26985
rect 23109 26976 23121 26979
rect 22980 26948 23121 26976
rect 22980 26936 22986 26948
rect 23109 26945 23121 26948
rect 23155 26945 23167 26979
rect 23293 26979 23351 26985
rect 23293 26976 23305 26979
rect 23109 26939 23167 26945
rect 23216 26948 23305 26976
rect 23216 26920 23244 26948
rect 23293 26945 23305 26948
rect 23339 26945 23351 26979
rect 23293 26939 23351 26945
rect 23382 26936 23388 26988
rect 23440 26976 23446 26988
rect 25774 26976 25780 26988
rect 23440 26948 23485 26976
rect 25735 26948 25780 26976
rect 23440 26936 23446 26948
rect 25774 26936 25780 26948
rect 25832 26936 25838 26988
rect 25869 26979 25927 26985
rect 25869 26945 25881 26979
rect 25915 26976 25927 26979
rect 25958 26976 25964 26988
rect 25915 26948 25964 26976
rect 25915 26945 25927 26948
rect 25869 26939 25927 26945
rect 25958 26936 25964 26948
rect 26016 26936 26022 26988
rect 27062 26936 27068 26988
rect 27120 26976 27126 26988
rect 27229 26979 27287 26985
rect 27229 26976 27241 26979
rect 27120 26948 27241 26976
rect 27120 26936 27126 26948
rect 27229 26945 27241 26948
rect 27275 26945 27287 26979
rect 27229 26939 27287 26945
rect 28997 26979 29055 26985
rect 28997 26945 29009 26979
rect 29043 26945 29055 26979
rect 29914 26976 29920 26988
rect 29875 26948 29920 26976
rect 28997 26939 29055 26945
rect 23198 26908 23204 26920
rect 22399 26880 23204 26908
rect 22281 26871 22339 26877
rect 18230 26840 18236 26852
rect 16684 26812 17540 26840
rect 17696 26812 18236 26840
rect 14642 26772 14648 26784
rect 14603 26744 14648 26772
rect 14642 26732 14648 26744
rect 14700 26732 14706 26784
rect 15654 26732 15660 26784
rect 15712 26772 15718 26784
rect 16666 26772 16672 26784
rect 15712 26744 16672 26772
rect 15712 26732 15718 26744
rect 16666 26732 16672 26744
rect 16724 26732 16730 26784
rect 16850 26772 16856 26784
rect 16811 26744 16856 26772
rect 16850 26732 16856 26744
rect 16908 26732 16914 26784
rect 17512 26772 17540 26812
rect 18230 26800 18236 26812
rect 18288 26800 18294 26852
rect 21818 26840 21824 26852
rect 18331 26812 19932 26840
rect 18331 26772 18359 26812
rect 17512 26744 18359 26772
rect 18693 26775 18751 26781
rect 18693 26741 18705 26775
rect 18739 26772 18751 26775
rect 19518 26772 19524 26784
rect 18739 26744 19524 26772
rect 18739 26741 18751 26744
rect 18693 26735 18751 26741
rect 19518 26732 19524 26744
rect 19576 26732 19582 26784
rect 19904 26772 19932 26812
rect 21468 26812 21824 26840
rect 21468 26772 21496 26812
rect 21818 26800 21824 26812
rect 21876 26800 21882 26852
rect 22296 26840 22324 26871
rect 23198 26868 23204 26880
rect 23256 26868 23262 26920
rect 23842 26908 23848 26920
rect 23803 26880 23848 26908
rect 23842 26868 23848 26880
rect 23900 26868 23906 26920
rect 26973 26911 27031 26917
rect 26973 26877 26985 26911
rect 27019 26877 27031 26911
rect 26973 26871 27031 26877
rect 22462 26840 22468 26852
rect 22296 26812 22468 26840
rect 22462 26800 22468 26812
rect 22520 26800 22526 26852
rect 19904 26744 21496 26772
rect 21542 26732 21548 26784
rect 21600 26772 21606 26784
rect 23109 26775 23167 26781
rect 23109 26772 23121 26775
rect 21600 26744 23121 26772
rect 21600 26732 21606 26744
rect 23109 26741 23121 26744
rect 23155 26741 23167 26775
rect 23109 26735 23167 26741
rect 23474 26732 23480 26784
rect 23532 26772 23538 26784
rect 26053 26775 26111 26781
rect 26053 26772 26065 26775
rect 23532 26744 26065 26772
rect 23532 26732 23538 26744
rect 26053 26741 26065 26744
rect 26099 26772 26111 26775
rect 26786 26772 26792 26784
rect 26099 26744 26792 26772
rect 26099 26741 26111 26744
rect 26053 26735 26111 26741
rect 26786 26732 26792 26744
rect 26844 26732 26850 26784
rect 26988 26772 27016 26871
rect 29012 26840 29040 26939
rect 29914 26936 29920 26948
rect 29972 26936 29978 26988
rect 30006 26936 30012 26988
rect 30064 26976 30070 26988
rect 30466 26985 30472 26988
rect 30423 26979 30472 26985
rect 30064 26948 30109 26976
rect 30064 26936 30070 26948
rect 30423 26945 30435 26979
rect 30469 26945 30472 26979
rect 30423 26939 30472 26945
rect 30466 26936 30472 26939
rect 30524 26936 30530 26988
rect 31021 26979 31079 26985
rect 31021 26976 31033 26979
rect 30576 26948 31033 26976
rect 29270 26908 29276 26920
rect 29231 26880 29276 26908
rect 29270 26868 29276 26880
rect 29328 26868 29334 26920
rect 30576 26849 30604 26948
rect 31021 26945 31033 26948
rect 31067 26945 31079 26979
rect 31021 26939 31079 26945
rect 30561 26843 30619 26849
rect 29012 26812 29859 26840
rect 27706 26772 27712 26784
rect 26988 26744 27712 26772
rect 27706 26732 27712 26744
rect 27764 26732 27770 26784
rect 28258 26732 28264 26784
rect 28316 26772 28322 26784
rect 28902 26772 28908 26784
rect 28316 26744 28908 26772
rect 28316 26732 28322 26744
rect 28902 26732 28908 26744
rect 28960 26732 28966 26784
rect 29181 26775 29239 26781
rect 29181 26741 29193 26775
rect 29227 26772 29239 26775
rect 29730 26772 29736 26784
rect 29227 26744 29736 26772
rect 29227 26741 29239 26744
rect 29181 26735 29239 26741
rect 29730 26732 29736 26744
rect 29788 26732 29794 26784
rect 29831 26772 29859 26812
rect 30561 26809 30573 26843
rect 30607 26809 30619 26843
rect 31128 26840 31156 27084
rect 31570 27072 31576 27084
rect 31628 27072 31634 27124
rect 32217 27115 32275 27121
rect 32217 27081 32229 27115
rect 32263 27112 32275 27115
rect 32398 27112 32404 27124
rect 32263 27084 32404 27112
rect 32263 27081 32275 27084
rect 32217 27075 32275 27081
rect 32398 27072 32404 27084
rect 32456 27072 32462 27124
rect 32950 27072 32956 27124
rect 33008 27112 33014 27124
rect 33008 27084 33180 27112
rect 33008 27072 33014 27084
rect 31205 27047 31263 27053
rect 31205 27013 31217 27047
rect 31251 27044 31263 27047
rect 31478 27044 31484 27056
rect 31251 27016 31484 27044
rect 31251 27013 31263 27016
rect 31205 27007 31263 27013
rect 31478 27004 31484 27016
rect 31536 27004 31542 27056
rect 31662 27004 31668 27056
rect 31720 27044 31726 27056
rect 32674 27044 32680 27056
rect 31720 27016 32680 27044
rect 31720 27004 31726 27016
rect 31297 26979 31355 26985
rect 31297 26945 31309 26979
rect 31343 26945 31355 26979
rect 31297 26939 31355 26945
rect 31389 26979 31447 26985
rect 31389 26945 31401 26979
rect 31435 26976 31447 26979
rect 31754 26976 31760 26988
rect 31435 26948 31760 26976
rect 31435 26945 31447 26948
rect 31389 26939 31447 26945
rect 31202 26868 31208 26920
rect 31260 26908 31266 26920
rect 31312 26908 31340 26939
rect 31754 26936 31760 26948
rect 31812 26936 31818 26988
rect 32140 26985 32168 27016
rect 32674 27004 32680 27016
rect 32732 27004 32738 27056
rect 32125 26979 32183 26985
rect 32125 26945 32137 26979
rect 32171 26945 32183 26979
rect 32766 26976 32772 26988
rect 32727 26948 32772 26976
rect 32125 26939 32183 26945
rect 32766 26936 32772 26948
rect 32824 26936 32830 26988
rect 32957 26977 33015 26983
rect 32957 26943 32969 26977
rect 33003 26974 33015 26977
rect 33152 26976 33180 27084
rect 33318 27072 33324 27124
rect 33376 27112 33382 27124
rect 33505 27115 33563 27121
rect 33505 27112 33517 27115
rect 33376 27084 33517 27112
rect 33376 27072 33382 27084
rect 33505 27081 33517 27084
rect 33551 27081 33563 27115
rect 33505 27075 33563 27081
rect 33060 26974 33180 26976
rect 33003 26948 33180 26974
rect 33321 26979 33379 26985
rect 33003 26946 33088 26948
rect 33003 26943 33015 26946
rect 32957 26937 33015 26943
rect 33321 26945 33333 26979
rect 33367 26976 33379 26979
rect 33594 26976 33600 26988
rect 33367 26948 33600 26976
rect 33367 26945 33379 26948
rect 33321 26939 33379 26945
rect 33594 26936 33600 26948
rect 33652 26936 33658 26988
rect 33965 26979 34023 26985
rect 33965 26945 33977 26979
rect 34011 26945 34023 26979
rect 33965 26939 34023 26945
rect 31260 26880 31340 26908
rect 31260 26868 31266 26880
rect 32582 26868 32588 26920
rect 32640 26908 32646 26920
rect 33045 26911 33103 26917
rect 33045 26908 33057 26911
rect 32640 26880 33057 26908
rect 32640 26868 32646 26880
rect 33045 26877 33057 26880
rect 33091 26877 33103 26911
rect 33045 26871 33103 26877
rect 33137 26911 33195 26917
rect 33137 26877 33149 26911
rect 33183 26908 33195 26911
rect 33778 26908 33784 26920
rect 33183 26880 33784 26908
rect 33183 26877 33195 26880
rect 33137 26871 33195 26877
rect 33778 26868 33784 26880
rect 33836 26868 33842 26920
rect 33980 26840 34008 26939
rect 31128 26812 34008 26840
rect 30561 26803 30619 26809
rect 31754 26772 31760 26784
rect 29831 26744 31760 26772
rect 31754 26732 31760 26744
rect 31812 26732 31818 26784
rect 33134 26732 33140 26784
rect 33192 26772 33198 26784
rect 34057 26775 34115 26781
rect 34057 26772 34069 26775
rect 33192 26744 34069 26772
rect 33192 26732 33198 26744
rect 34057 26741 34069 26744
rect 34103 26741 34115 26775
rect 34057 26735 34115 26741
rect 1104 26682 34868 26704
rect 1104 26630 6582 26682
rect 6634 26630 6646 26682
rect 6698 26630 6710 26682
rect 6762 26630 6774 26682
rect 6826 26630 6838 26682
rect 6890 26630 17846 26682
rect 17898 26630 17910 26682
rect 17962 26630 17974 26682
rect 18026 26630 18038 26682
rect 18090 26630 18102 26682
rect 18154 26630 29110 26682
rect 29162 26630 29174 26682
rect 29226 26630 29238 26682
rect 29290 26630 29302 26682
rect 29354 26630 29366 26682
rect 29418 26630 34868 26682
rect 1104 26608 34868 26630
rect 14277 26571 14335 26577
rect 14277 26537 14289 26571
rect 14323 26568 14335 26571
rect 14323 26540 16528 26568
rect 14323 26537 14335 26540
rect 14277 26531 14335 26537
rect 16500 26500 16528 26540
rect 16666 26528 16672 26580
rect 16724 26568 16730 26580
rect 16945 26571 17003 26577
rect 16945 26568 16957 26571
rect 16724 26540 16957 26568
rect 16724 26528 16730 26540
rect 16945 26537 16957 26540
rect 16991 26537 17003 26571
rect 16945 26531 17003 26537
rect 17216 26540 17428 26568
rect 17216 26500 17244 26540
rect 16500 26472 17244 26500
rect 17400 26500 17428 26540
rect 17494 26528 17500 26580
rect 17552 26568 17558 26580
rect 17865 26571 17923 26577
rect 17552 26540 17597 26568
rect 17552 26528 17558 26540
rect 17865 26537 17877 26571
rect 17911 26568 17923 26571
rect 18506 26568 18512 26580
rect 17911 26540 18512 26568
rect 17911 26537 17923 26540
rect 17865 26531 17923 26537
rect 18506 26528 18512 26540
rect 18564 26528 18570 26580
rect 18690 26528 18696 26580
rect 18748 26568 18754 26580
rect 21082 26568 21088 26580
rect 18748 26540 20208 26568
rect 21043 26540 21088 26568
rect 18748 26528 18754 26540
rect 17400 26472 18276 26500
rect 14642 26392 14648 26444
rect 14700 26432 14706 26444
rect 17126 26432 17132 26444
rect 14700 26404 15700 26432
rect 14700 26392 14706 26404
rect 14461 26367 14519 26373
rect 14461 26333 14473 26367
rect 14507 26364 14519 26367
rect 14826 26364 14832 26376
rect 14507 26336 14832 26364
rect 14507 26333 14519 26336
rect 14461 26327 14519 26333
rect 14826 26324 14832 26336
rect 14884 26324 14890 26376
rect 14921 26367 14979 26373
rect 14921 26333 14933 26367
rect 14967 26333 14979 26367
rect 14921 26327 14979 26333
rect 15105 26367 15163 26373
rect 15105 26333 15117 26367
rect 15151 26364 15163 26367
rect 15562 26364 15568 26376
rect 15151 26336 15424 26364
rect 15523 26336 15568 26364
rect 15151 26333 15163 26336
rect 15105 26327 15163 26333
rect 14936 26296 14964 26327
rect 15286 26296 15292 26308
rect 14936 26268 15292 26296
rect 15286 26256 15292 26268
rect 15344 26256 15350 26308
rect 15396 26296 15424 26336
rect 15562 26324 15568 26336
rect 15620 26324 15626 26376
rect 15672 26364 15700 26404
rect 16592 26404 17132 26432
rect 15821 26367 15879 26373
rect 15821 26364 15833 26367
rect 15672 26336 15833 26364
rect 15821 26333 15833 26336
rect 15867 26333 15879 26367
rect 16592 26364 16620 26404
rect 17126 26392 17132 26404
rect 17184 26392 17190 26444
rect 17589 26435 17647 26441
rect 17589 26401 17601 26435
rect 17635 26432 17647 26435
rect 18138 26432 18144 26444
rect 17635 26404 18144 26432
rect 17635 26401 17647 26404
rect 17589 26395 17647 26401
rect 18138 26392 18144 26404
rect 18196 26392 18202 26444
rect 18248 26432 18276 26472
rect 18322 26460 18328 26512
rect 18380 26500 18386 26512
rect 20180 26500 20208 26540
rect 21082 26528 21088 26540
rect 21140 26528 21146 26580
rect 21358 26528 21364 26580
rect 21416 26568 21422 26580
rect 21416 26540 23152 26568
rect 21416 26528 21422 26540
rect 23124 26512 23152 26540
rect 23198 26528 23204 26580
rect 23256 26568 23262 26580
rect 23477 26571 23535 26577
rect 23477 26568 23489 26571
rect 23256 26540 23489 26568
rect 23256 26528 23262 26540
rect 23477 26537 23489 26540
rect 23523 26537 23535 26571
rect 23477 26531 23535 26537
rect 23661 26571 23719 26577
rect 23661 26537 23673 26571
rect 23707 26568 23719 26571
rect 24302 26568 24308 26580
rect 23707 26540 24308 26568
rect 23707 26537 23719 26540
rect 23661 26531 23719 26537
rect 21450 26500 21456 26512
rect 18380 26472 19288 26500
rect 20180 26472 21456 26500
rect 18380 26460 18386 26472
rect 18248 26404 18920 26432
rect 15821 26327 15879 26333
rect 16500 26336 16620 26364
rect 16500 26308 16528 26336
rect 16666 26324 16672 26376
rect 16724 26364 16730 26376
rect 17218 26364 17224 26376
rect 16724 26336 17224 26364
rect 16724 26324 16730 26336
rect 17218 26324 17224 26336
rect 17276 26364 17282 26376
rect 17681 26367 17739 26373
rect 17276 26340 17540 26364
rect 17276 26336 17632 26340
rect 17276 26324 17282 26336
rect 17512 26312 17632 26336
rect 17681 26333 17693 26367
rect 17727 26333 17739 26367
rect 18325 26367 18383 26373
rect 18325 26364 18337 26367
rect 17681 26327 17739 26333
rect 17880 26336 18337 26364
rect 16298 26296 16304 26308
rect 15396 26268 16304 26296
rect 16298 26256 16304 26268
rect 16356 26256 16362 26308
rect 16482 26256 16488 26308
rect 16540 26256 16546 26308
rect 17310 26256 17316 26308
rect 17368 26296 17374 26308
rect 17405 26299 17463 26305
rect 17405 26296 17417 26299
rect 17368 26268 17417 26296
rect 17368 26256 17374 26268
rect 17405 26265 17417 26268
rect 17451 26265 17463 26299
rect 17604 26296 17632 26312
rect 17696 26296 17724 26327
rect 17880 26296 17908 26336
rect 18325 26333 18337 26336
rect 18371 26333 18383 26367
rect 18325 26327 18383 26333
rect 18414 26324 18420 26376
rect 18472 26364 18478 26376
rect 18509 26367 18567 26373
rect 18509 26364 18521 26367
rect 18472 26336 18521 26364
rect 18472 26324 18478 26336
rect 18509 26333 18521 26336
rect 18555 26333 18567 26367
rect 18509 26327 18567 26333
rect 18892 26296 18920 26404
rect 19260 26373 19288 26472
rect 21450 26460 21456 26472
rect 21508 26460 21514 26512
rect 23106 26500 23112 26512
rect 23019 26472 23112 26500
rect 23106 26460 23112 26472
rect 23164 26500 23170 26512
rect 23676 26500 23704 26531
rect 24302 26528 24308 26540
rect 24360 26528 24366 26580
rect 25774 26528 25780 26580
rect 25832 26568 25838 26580
rect 26050 26568 26056 26580
rect 25832 26540 26056 26568
rect 25832 26528 25838 26540
rect 26050 26528 26056 26540
rect 26108 26568 26114 26580
rect 26237 26571 26295 26577
rect 26237 26568 26249 26571
rect 26108 26540 26249 26568
rect 26108 26528 26114 26540
rect 26237 26537 26249 26540
rect 26283 26537 26295 26571
rect 26237 26531 26295 26537
rect 28718 26528 28724 26580
rect 28776 26568 28782 26580
rect 28813 26571 28871 26577
rect 28813 26568 28825 26571
rect 28776 26540 28825 26568
rect 28776 26528 28782 26540
rect 28813 26537 28825 26540
rect 28859 26537 28871 26571
rect 28813 26531 28871 26537
rect 28902 26528 28908 26580
rect 28960 26568 28966 26580
rect 28997 26571 29055 26577
rect 28997 26568 29009 26571
rect 28960 26540 29009 26568
rect 28960 26528 28966 26540
rect 28997 26537 29009 26540
rect 29043 26568 29055 26571
rect 29546 26568 29552 26580
rect 29043 26540 29552 26568
rect 29043 26537 29055 26540
rect 28997 26531 29055 26537
rect 29546 26528 29552 26540
rect 29604 26528 29610 26580
rect 29914 26528 29920 26580
rect 29972 26568 29978 26580
rect 31389 26571 31447 26577
rect 31389 26568 31401 26571
rect 29972 26540 31401 26568
rect 29972 26528 29978 26540
rect 31389 26537 31401 26540
rect 31435 26537 31447 26571
rect 33689 26571 33747 26577
rect 33689 26568 33701 26571
rect 31389 26531 31447 26537
rect 33612 26540 33701 26568
rect 23164 26472 23704 26500
rect 23164 26460 23170 26472
rect 28166 26460 28172 26512
rect 28224 26500 28230 26512
rect 30282 26500 30288 26512
rect 28224 26472 30288 26500
rect 28224 26460 28230 26472
rect 30282 26460 30288 26472
rect 30340 26460 30346 26512
rect 30374 26460 30380 26512
rect 30432 26500 30438 26512
rect 31294 26500 31300 26512
rect 30432 26472 31064 26500
rect 31207 26472 31300 26500
rect 30432 26460 30438 26472
rect 22005 26435 22063 26441
rect 22005 26401 22017 26435
rect 22051 26432 22063 26435
rect 22186 26432 22192 26444
rect 22051 26404 22192 26432
rect 22051 26401 22063 26404
rect 22005 26395 22063 26401
rect 22186 26392 22192 26404
rect 22244 26432 22250 26444
rect 22646 26432 22652 26444
rect 22244 26404 22652 26432
rect 22244 26392 22250 26404
rect 22646 26392 22652 26404
rect 22704 26392 22710 26444
rect 29638 26432 29644 26444
rect 29599 26404 29644 26432
rect 29638 26392 29644 26404
rect 29696 26392 29702 26444
rect 29730 26392 29736 26444
rect 29788 26432 29794 26444
rect 29917 26435 29975 26441
rect 29917 26432 29929 26435
rect 29788 26404 29929 26432
rect 29788 26392 29794 26404
rect 29917 26401 29929 26404
rect 29963 26432 29975 26435
rect 30650 26432 30656 26444
rect 29963 26404 30656 26432
rect 29963 26401 29975 26404
rect 29917 26395 29975 26401
rect 30650 26392 30656 26404
rect 30708 26392 30714 26444
rect 30742 26392 30748 26444
rect 30800 26432 30806 26444
rect 30929 26435 30987 26441
rect 30929 26432 30941 26435
rect 30800 26404 30941 26432
rect 30800 26392 30806 26404
rect 30929 26401 30941 26404
rect 30975 26401 30987 26435
rect 31036 26432 31064 26472
rect 31294 26460 31300 26472
rect 31352 26500 31358 26512
rect 31662 26500 31668 26512
rect 31352 26472 31668 26500
rect 31352 26460 31358 26472
rect 31662 26460 31668 26472
rect 31720 26460 31726 26512
rect 31036 26404 32444 26432
rect 30929 26395 30987 26401
rect 19245 26367 19303 26373
rect 19245 26333 19257 26367
rect 19291 26364 19303 26367
rect 19334 26364 19340 26376
rect 19291 26336 19340 26364
rect 19291 26333 19303 26336
rect 19245 26327 19303 26333
rect 19334 26324 19340 26336
rect 19392 26324 19398 26376
rect 19518 26373 19524 26376
rect 19512 26364 19524 26373
rect 19479 26336 19524 26364
rect 19512 26327 19524 26336
rect 19518 26324 19524 26327
rect 19576 26324 19582 26376
rect 19886 26324 19892 26376
rect 19944 26364 19950 26376
rect 20806 26364 20812 26376
rect 19944 26336 20812 26364
rect 19944 26324 19950 26336
rect 20806 26324 20812 26336
rect 20864 26324 20870 26376
rect 21269 26367 21327 26373
rect 21269 26333 21281 26367
rect 21315 26364 21327 26367
rect 21358 26364 21364 26376
rect 21315 26336 21364 26364
rect 21315 26333 21327 26336
rect 21269 26327 21327 26333
rect 21358 26324 21364 26336
rect 21416 26324 21422 26376
rect 21453 26367 21511 26373
rect 21453 26333 21465 26367
rect 21499 26333 21511 26367
rect 21453 26327 21511 26333
rect 21545 26367 21603 26373
rect 21545 26333 21557 26367
rect 21591 26364 21603 26367
rect 22094 26364 22100 26376
rect 21591 26336 22100 26364
rect 21591 26333 21603 26336
rect 21545 26327 21603 26333
rect 19702 26296 19708 26308
rect 17604 26268 17908 26296
rect 18524 26268 18828 26296
rect 18892 26268 19708 26296
rect 17405 26259 17463 26265
rect 15010 26228 15016 26240
rect 14971 26200 15016 26228
rect 15010 26188 15016 26200
rect 15068 26188 15074 26240
rect 15102 26188 15108 26240
rect 15160 26228 15166 26240
rect 18524 26228 18552 26268
rect 18690 26228 18696 26240
rect 15160 26200 18552 26228
rect 18651 26200 18696 26228
rect 15160 26188 15166 26200
rect 18690 26188 18696 26200
rect 18748 26188 18754 26240
rect 18800 26228 18828 26268
rect 19702 26256 19708 26268
rect 19760 26256 19766 26308
rect 21468 26296 21496 26327
rect 22094 26324 22100 26336
rect 22152 26324 22158 26376
rect 22278 26324 22284 26376
rect 22336 26364 22342 26376
rect 23382 26364 23388 26376
rect 22336 26336 23388 26364
rect 22336 26324 22342 26336
rect 23382 26324 23388 26336
rect 23440 26364 23446 26376
rect 24857 26367 24915 26373
rect 23440 26339 23536 26364
rect 23440 26336 23581 26339
rect 23440 26324 23446 26336
rect 23508 26333 23581 26336
rect 22296 26296 22324 26324
rect 20548 26268 22324 26296
rect 20548 26228 20576 26268
rect 22462 26256 22468 26308
rect 22520 26296 22526 26308
rect 23290 26296 23296 26308
rect 22520 26268 23296 26296
rect 22520 26256 22526 26268
rect 23290 26256 23296 26268
rect 23348 26256 23354 26308
rect 23508 26302 23535 26333
rect 23523 26299 23535 26302
rect 23569 26299 23581 26333
rect 24857 26333 24869 26367
rect 24903 26364 24915 26367
rect 26697 26367 26755 26373
rect 26697 26364 26709 26367
rect 24903 26336 26709 26364
rect 24903 26333 24915 26336
rect 24857 26327 24915 26333
rect 26697 26333 26709 26336
rect 26743 26364 26755 26367
rect 27706 26364 27712 26376
rect 26743 26336 27712 26364
rect 26743 26333 26755 26336
rect 26697 26327 26755 26333
rect 27706 26324 27712 26336
rect 27764 26364 27770 26376
rect 28350 26364 28356 26376
rect 27764 26336 28356 26364
rect 27764 26324 27770 26336
rect 28350 26324 28356 26336
rect 28408 26324 28414 26376
rect 30208 26336 31064 26364
rect 23523 26293 23581 26299
rect 25124 26299 25182 26305
rect 25124 26265 25136 26299
rect 25170 26296 25182 26299
rect 25590 26296 25596 26308
rect 25170 26268 25596 26296
rect 25170 26265 25182 26268
rect 25124 26259 25182 26265
rect 25590 26256 25596 26268
rect 25648 26256 25654 26308
rect 26942 26299 27000 26305
rect 26942 26265 26954 26299
rect 26988 26265 27000 26299
rect 26942 26259 27000 26265
rect 28629 26299 28687 26305
rect 28629 26265 28641 26299
rect 28675 26296 28687 26299
rect 30208 26296 30236 26336
rect 28675 26268 30236 26296
rect 31036 26296 31064 26336
rect 32122 26324 32128 26376
rect 32180 26364 32186 26376
rect 32306 26364 32312 26376
rect 32180 26336 32312 26364
rect 32180 26324 32186 26336
rect 32306 26324 32312 26336
rect 32364 26324 32370 26376
rect 32416 26364 32444 26404
rect 32565 26367 32623 26373
rect 32565 26364 32577 26367
rect 32416 26336 32577 26364
rect 32565 26333 32577 26336
rect 32611 26333 32623 26367
rect 32565 26327 32623 26333
rect 32766 26296 32772 26308
rect 31036 26268 31984 26296
rect 28675 26265 28687 26268
rect 28629 26259 28687 26265
rect 18800 26200 20576 26228
rect 20622 26188 20628 26240
rect 20680 26228 20686 26240
rect 20680 26200 20725 26228
rect 20680 26188 20686 26200
rect 23934 26188 23940 26240
rect 23992 26228 23998 26240
rect 26957 26228 26985 26259
rect 23992 26200 26985 26228
rect 23992 26188 23998 26200
rect 27430 26188 27436 26240
rect 27488 26228 27494 26240
rect 27706 26228 27712 26240
rect 27488 26200 27712 26228
rect 27488 26188 27494 26200
rect 27706 26188 27712 26200
rect 27764 26188 27770 26240
rect 28077 26231 28135 26237
rect 28077 26197 28089 26231
rect 28123 26228 28135 26231
rect 28258 26228 28264 26240
rect 28123 26200 28264 26228
rect 28123 26197 28135 26200
rect 28077 26191 28135 26197
rect 28258 26188 28264 26200
rect 28316 26188 28322 26240
rect 28810 26188 28816 26240
rect 28868 26237 28874 26240
rect 28868 26231 28887 26237
rect 28875 26197 28887 26231
rect 31956 26228 31984 26268
rect 32692 26268 32772 26296
rect 32692 26228 32720 26268
rect 32766 26256 32772 26268
rect 32824 26296 32830 26308
rect 32950 26296 32956 26308
rect 32824 26268 32956 26296
rect 32824 26256 32830 26268
rect 32950 26256 32956 26268
rect 33008 26296 33014 26308
rect 33612 26296 33640 26540
rect 33689 26537 33701 26540
rect 33735 26537 33747 26571
rect 33689 26531 33747 26537
rect 33008 26268 33640 26296
rect 33008 26256 33014 26268
rect 31956 26200 32720 26228
rect 28868 26191 28887 26197
rect 28868 26188 28874 26191
rect 1104 26138 34868 26160
rect 1104 26086 12214 26138
rect 12266 26086 12278 26138
rect 12330 26086 12342 26138
rect 12394 26086 12406 26138
rect 12458 26086 12470 26138
rect 12522 26086 23478 26138
rect 23530 26086 23542 26138
rect 23594 26086 23606 26138
rect 23658 26086 23670 26138
rect 23722 26086 23734 26138
rect 23786 26086 34868 26138
rect 1104 26064 34868 26086
rect 18690 26024 18696 26036
rect 14384 25996 18696 26024
rect 14001 25891 14059 25897
rect 14001 25857 14013 25891
rect 14047 25888 14059 25891
rect 14384 25888 14412 25996
rect 18690 25984 18696 25996
rect 18748 25984 18754 26036
rect 18782 25984 18788 26036
rect 18840 26024 18846 26036
rect 25590 26024 25596 26036
rect 18840 25996 24072 26024
rect 25551 25996 25596 26024
rect 18840 25984 18846 25996
rect 15102 25956 15108 25968
rect 14476 25928 15108 25956
rect 14476 25897 14504 25928
rect 15102 25916 15108 25928
rect 15160 25916 15166 25968
rect 15381 25959 15439 25965
rect 15381 25925 15393 25959
rect 15427 25956 15439 25959
rect 15654 25956 15660 25968
rect 15427 25928 15660 25956
rect 15427 25925 15439 25928
rect 15381 25919 15439 25925
rect 15654 25916 15660 25928
rect 15712 25956 15718 25968
rect 16758 25956 16764 25968
rect 15712 25928 16764 25956
rect 15712 25916 15718 25928
rect 16758 25916 16764 25928
rect 16816 25916 16822 25968
rect 16942 25916 16948 25968
rect 17000 25956 17006 25968
rect 17000 25928 18348 25956
rect 17000 25916 17006 25928
rect 14047 25860 14412 25888
rect 14461 25891 14519 25897
rect 14047 25857 14059 25860
rect 14001 25851 14059 25857
rect 14461 25857 14473 25891
rect 14507 25857 14519 25891
rect 14461 25851 14519 25857
rect 14645 25891 14703 25897
rect 14645 25857 14657 25891
rect 14691 25857 14703 25891
rect 14645 25851 14703 25857
rect 15197 25891 15255 25897
rect 15197 25857 15209 25891
rect 15243 25888 15255 25891
rect 15286 25888 15292 25900
rect 15243 25860 15292 25888
rect 15243 25857 15255 25860
rect 15197 25851 15255 25857
rect 14660 25820 14688 25851
rect 15286 25848 15292 25860
rect 15344 25848 15350 25900
rect 15933 25891 15991 25897
rect 15933 25857 15945 25891
rect 15979 25888 15991 25891
rect 16390 25888 16396 25900
rect 15979 25860 16396 25888
rect 15979 25857 15991 25860
rect 15933 25851 15991 25857
rect 16390 25848 16396 25860
rect 16448 25848 16454 25900
rect 16574 25848 16580 25900
rect 16632 25888 16638 25900
rect 17385 25891 17443 25897
rect 17385 25888 17397 25891
rect 16632 25860 17397 25888
rect 16632 25848 16638 25860
rect 17385 25857 17397 25860
rect 17431 25857 17443 25891
rect 18320 25888 18348 25928
rect 18414 25916 18420 25968
rect 18472 25956 18478 25968
rect 19702 25965 19708 25968
rect 19696 25956 19708 25965
rect 18472 25928 19564 25956
rect 19663 25928 19708 25956
rect 18472 25916 18478 25928
rect 18782 25888 18788 25900
rect 18320 25860 18788 25888
rect 17385 25851 17443 25857
rect 18782 25848 18788 25860
rect 18840 25848 18846 25900
rect 19426 25888 19432 25900
rect 19387 25860 19432 25888
rect 19426 25848 19432 25860
rect 19484 25848 19490 25900
rect 19536 25888 19564 25928
rect 19696 25919 19708 25928
rect 19702 25916 19708 25919
rect 19760 25916 19766 25968
rect 19794 25916 19800 25968
rect 19852 25956 19858 25968
rect 20622 25956 20628 25968
rect 19852 25928 20628 25956
rect 19852 25916 19858 25928
rect 20622 25916 20628 25928
rect 20680 25916 20686 25968
rect 23842 25956 23848 25968
rect 21928 25928 23848 25956
rect 19536 25860 20576 25888
rect 15470 25820 15476 25832
rect 14660 25792 15476 25820
rect 15470 25780 15476 25792
rect 15528 25780 15534 25832
rect 15562 25780 15568 25832
rect 15620 25820 15626 25832
rect 16850 25820 16856 25832
rect 15620 25792 16856 25820
rect 15620 25780 15626 25792
rect 16850 25780 16856 25792
rect 16908 25820 16914 25832
rect 17129 25823 17187 25829
rect 17129 25820 17141 25823
rect 16908 25792 17141 25820
rect 16908 25780 16914 25792
rect 17129 25789 17141 25792
rect 17175 25789 17187 25823
rect 17129 25783 17187 25789
rect 18230 25780 18236 25832
rect 18288 25780 18294 25832
rect 14461 25755 14519 25761
rect 14461 25721 14473 25755
rect 14507 25752 14519 25755
rect 18248 25752 18276 25780
rect 18509 25755 18567 25761
rect 18509 25752 18521 25755
rect 14507 25724 17172 25752
rect 18248 25724 18521 25752
rect 14507 25721 14519 25724
rect 14461 25715 14519 25721
rect 13814 25684 13820 25696
rect 13775 25656 13820 25684
rect 13814 25644 13820 25656
rect 13872 25644 13878 25696
rect 16025 25687 16083 25693
rect 16025 25653 16037 25687
rect 16071 25684 16083 25687
rect 16666 25684 16672 25696
rect 16071 25656 16672 25684
rect 16071 25653 16083 25656
rect 16025 25647 16083 25653
rect 16666 25644 16672 25656
rect 16724 25644 16730 25696
rect 17144 25684 17172 25724
rect 18509 25721 18521 25724
rect 18555 25721 18567 25755
rect 20548 25752 20576 25860
rect 20806 25848 20812 25900
rect 20864 25888 20870 25900
rect 21928 25897 21956 25928
rect 21913 25891 21971 25897
rect 21913 25888 21925 25891
rect 20864 25860 21925 25888
rect 20864 25848 20870 25860
rect 21913 25857 21925 25860
rect 21959 25857 21971 25891
rect 21913 25851 21971 25857
rect 22002 25848 22008 25900
rect 22060 25888 22066 25900
rect 23768 25897 23796 25928
rect 23842 25916 23848 25928
rect 23900 25916 23906 25968
rect 24044 25965 24072 25996
rect 25590 25984 25596 25996
rect 25648 25984 25654 26036
rect 26973 26027 27031 26033
rect 26973 25993 26985 26027
rect 27019 26024 27031 26027
rect 27062 26024 27068 26036
rect 27019 25996 27068 26024
rect 27019 25993 27031 25996
rect 26973 25987 27031 25993
rect 27062 25984 27068 25996
rect 27120 25984 27126 26036
rect 28534 26024 28540 26036
rect 27264 25996 28540 26024
rect 24020 25959 24078 25965
rect 24020 25925 24032 25959
rect 24066 25925 24078 25959
rect 24020 25919 24078 25925
rect 22169 25891 22227 25897
rect 22169 25888 22181 25891
rect 22060 25860 22181 25888
rect 22060 25848 22066 25860
rect 22169 25857 22181 25860
rect 22215 25857 22227 25891
rect 22169 25851 22227 25857
rect 23753 25891 23811 25897
rect 23753 25857 23765 25891
rect 23799 25857 23811 25891
rect 25777 25891 25835 25897
rect 25777 25888 25789 25891
rect 23753 25851 23811 25857
rect 23860 25860 25789 25888
rect 23860 25820 23888 25860
rect 25777 25857 25789 25860
rect 25823 25857 25835 25891
rect 26050 25888 26056 25900
rect 26011 25860 26056 25888
rect 25777 25851 25835 25857
rect 26050 25848 26056 25860
rect 26108 25848 26114 25900
rect 27157 25891 27215 25897
rect 27157 25857 27169 25891
rect 27203 25888 27215 25891
rect 27264 25888 27292 25996
rect 28534 25984 28540 25996
rect 28592 25984 28598 26036
rect 29638 25984 29644 26036
rect 29696 26024 29702 26036
rect 29733 26027 29791 26033
rect 29733 26024 29745 26027
rect 29696 25996 29745 26024
rect 29696 25984 29702 25996
rect 29733 25993 29745 25996
rect 29779 25993 29791 26027
rect 33962 26024 33968 26036
rect 29733 25987 29791 25993
rect 29840 25996 33968 26024
rect 29840 25956 29868 25996
rect 33962 25984 33968 25996
rect 34020 25984 34026 26036
rect 27356 25928 29868 25956
rect 30193 25959 30251 25965
rect 27356 25900 27384 25928
rect 30193 25925 30205 25959
rect 30239 25925 30251 25959
rect 30193 25919 30251 25925
rect 30409 25959 30467 25965
rect 30409 25925 30421 25959
rect 30455 25956 30467 25959
rect 30650 25956 30656 25968
rect 30455 25928 30656 25956
rect 30455 25925 30467 25928
rect 30409 25919 30467 25925
rect 27203 25860 27292 25888
rect 27203 25857 27215 25860
rect 27157 25851 27215 25857
rect 27338 25848 27344 25900
rect 27396 25888 27402 25900
rect 28620 25891 28678 25897
rect 27396 25860 27489 25888
rect 27396 25848 27402 25860
rect 28620 25857 28632 25891
rect 28666 25888 28678 25891
rect 28902 25888 28908 25900
rect 28666 25860 28908 25888
rect 28666 25857 28678 25860
rect 28620 25851 28678 25857
rect 28902 25848 28908 25860
rect 28960 25848 28966 25900
rect 30208 25888 30236 25919
rect 30650 25916 30656 25928
rect 30708 25916 30714 25968
rect 30558 25888 30564 25900
rect 30208 25860 30564 25888
rect 30558 25848 30564 25860
rect 30616 25888 30622 25900
rect 30926 25888 30932 25900
rect 30616 25860 30932 25888
rect 30616 25848 30622 25860
rect 30926 25848 30932 25860
rect 30984 25848 30990 25900
rect 31297 25891 31355 25897
rect 31297 25857 31309 25891
rect 31343 25888 31355 25891
rect 31938 25888 31944 25900
rect 31343 25860 31944 25888
rect 31343 25857 31355 25860
rect 31297 25851 31355 25857
rect 31938 25848 31944 25860
rect 31996 25848 32002 25900
rect 32030 25848 32036 25900
rect 32088 25848 32094 25900
rect 34146 25888 34152 25900
rect 34107 25860 34152 25888
rect 34146 25848 34152 25860
rect 34204 25848 34210 25900
rect 23216 25792 23888 25820
rect 27433 25823 27491 25829
rect 20548 25724 21956 25752
rect 18509 25715 18567 25721
rect 20714 25684 20720 25696
rect 17144 25656 20720 25684
rect 20714 25644 20720 25656
rect 20772 25644 20778 25696
rect 20809 25687 20867 25693
rect 20809 25653 20821 25687
rect 20855 25684 20867 25687
rect 21818 25684 21824 25696
rect 20855 25656 21824 25684
rect 20855 25653 20867 25656
rect 20809 25647 20867 25653
rect 21818 25644 21824 25656
rect 21876 25644 21882 25696
rect 21928 25684 21956 25724
rect 23216 25684 23244 25792
rect 27433 25789 27445 25823
rect 27479 25820 27491 25823
rect 27890 25820 27896 25832
rect 27479 25792 27896 25820
rect 27479 25789 27491 25792
rect 27433 25783 27491 25789
rect 27890 25780 27896 25792
rect 27948 25780 27954 25832
rect 28350 25820 28356 25832
rect 28311 25792 28356 25820
rect 28350 25780 28356 25792
rect 28408 25780 28414 25832
rect 29730 25780 29736 25832
rect 29788 25820 29794 25832
rect 31481 25823 31539 25829
rect 31481 25820 31493 25823
rect 29788 25792 31493 25820
rect 29788 25780 29794 25792
rect 31481 25789 31493 25792
rect 31527 25789 31539 25823
rect 31481 25783 31539 25789
rect 31573 25823 31631 25829
rect 31573 25789 31585 25823
rect 31619 25820 31631 25823
rect 32048 25820 32076 25848
rect 31619 25792 32168 25820
rect 31619 25789 31631 25792
rect 31573 25783 31631 25789
rect 23290 25712 23296 25764
rect 23348 25752 23354 25764
rect 25130 25752 25136 25764
rect 23348 25724 23393 25752
rect 25043 25724 25136 25752
rect 23348 25712 23354 25724
rect 25130 25712 25136 25724
rect 25188 25752 25194 25764
rect 28166 25752 28172 25764
rect 25188 25724 28172 25752
rect 25188 25712 25194 25724
rect 28166 25712 28172 25724
rect 28224 25712 28230 25764
rect 31113 25755 31171 25761
rect 31113 25721 31125 25755
rect 31159 25752 31171 25755
rect 32030 25752 32036 25764
rect 31159 25724 32036 25752
rect 31159 25721 31171 25724
rect 31113 25715 31171 25721
rect 32030 25712 32036 25724
rect 32088 25712 32094 25764
rect 32140 25752 32168 25792
rect 32214 25780 32220 25832
rect 32272 25820 32278 25832
rect 32309 25823 32367 25829
rect 32309 25820 32321 25823
rect 32272 25792 32321 25820
rect 32272 25780 32278 25792
rect 32309 25789 32321 25792
rect 32355 25789 32367 25823
rect 32309 25783 32367 25789
rect 32493 25823 32551 25829
rect 32493 25789 32505 25823
rect 32539 25820 32551 25823
rect 34054 25820 34060 25832
rect 32539 25792 34060 25820
rect 32539 25789 32551 25792
rect 32493 25783 32551 25789
rect 34054 25780 34060 25792
rect 34112 25780 34118 25832
rect 32140 25724 32352 25752
rect 32324 25696 32352 25724
rect 25958 25684 25964 25696
rect 21928 25656 23244 25684
rect 25919 25656 25964 25684
rect 25958 25644 25964 25656
rect 26016 25644 26022 25696
rect 30377 25687 30435 25693
rect 30377 25653 30389 25687
rect 30423 25684 30435 25687
rect 30466 25684 30472 25696
rect 30423 25656 30472 25684
rect 30423 25653 30435 25656
rect 30377 25647 30435 25653
rect 30466 25644 30472 25656
rect 30524 25644 30530 25696
rect 30561 25687 30619 25693
rect 30561 25653 30573 25687
rect 30607 25684 30619 25687
rect 31018 25684 31024 25696
rect 30607 25656 31024 25684
rect 30607 25653 30619 25656
rect 30561 25647 30619 25653
rect 31018 25644 31024 25656
rect 31076 25644 31082 25696
rect 32306 25644 32312 25696
rect 32364 25644 32370 25696
rect 1104 25594 34868 25616
rect 1104 25542 6582 25594
rect 6634 25542 6646 25594
rect 6698 25542 6710 25594
rect 6762 25542 6774 25594
rect 6826 25542 6838 25594
rect 6890 25542 17846 25594
rect 17898 25542 17910 25594
rect 17962 25542 17974 25594
rect 18026 25542 18038 25594
rect 18090 25542 18102 25594
rect 18154 25542 29110 25594
rect 29162 25542 29174 25594
rect 29226 25542 29238 25594
rect 29290 25542 29302 25594
rect 29354 25542 29366 25594
rect 29418 25542 34868 25594
rect 1104 25520 34868 25542
rect 14369 25483 14427 25489
rect 14369 25449 14381 25483
rect 14415 25480 14427 25483
rect 16942 25480 16948 25492
rect 14415 25452 16948 25480
rect 14415 25449 14427 25452
rect 14369 25443 14427 25449
rect 16942 25440 16948 25452
rect 17000 25440 17006 25492
rect 17129 25483 17187 25489
rect 17129 25449 17141 25483
rect 17175 25480 17187 25483
rect 17310 25480 17316 25492
rect 17175 25452 17316 25480
rect 17175 25449 17187 25452
rect 17129 25443 17187 25449
rect 17310 25440 17316 25452
rect 17368 25480 17374 25492
rect 17494 25480 17500 25492
rect 17368 25452 17500 25480
rect 17368 25440 17374 25452
rect 17494 25440 17500 25452
rect 17552 25440 17558 25492
rect 21726 25480 21732 25492
rect 17604 25452 21732 25480
rect 17604 25412 17632 25452
rect 21726 25440 21732 25452
rect 21784 25440 21790 25492
rect 22002 25440 22008 25492
rect 22060 25480 22066 25492
rect 23845 25483 23903 25489
rect 23845 25480 23857 25483
rect 22060 25452 23857 25480
rect 22060 25440 22066 25452
rect 23845 25449 23857 25452
rect 23891 25449 23903 25483
rect 23845 25443 23903 25449
rect 24581 25483 24639 25489
rect 24581 25449 24593 25483
rect 24627 25480 24639 25483
rect 25130 25480 25136 25492
rect 24627 25452 25136 25480
rect 24627 25449 24639 25452
rect 24581 25443 24639 25449
rect 17144 25384 17632 25412
rect 1854 25344 1860 25356
rect 1815 25316 1860 25344
rect 1854 25304 1860 25316
rect 1912 25304 1918 25356
rect 13814 25304 13820 25356
rect 13872 25344 13878 25356
rect 13872 25316 14964 25344
rect 13872 25304 13878 25316
rect 1394 25276 1400 25288
rect 1355 25248 1400 25276
rect 1394 25236 1400 25248
rect 1452 25236 1458 25288
rect 14550 25276 14556 25288
rect 14511 25248 14556 25276
rect 14550 25236 14556 25248
rect 14608 25236 14614 25288
rect 14936 25276 14964 25316
rect 15562 25304 15568 25356
rect 15620 25344 15626 25356
rect 15749 25347 15807 25353
rect 15749 25344 15761 25347
rect 15620 25316 15761 25344
rect 15620 25304 15626 25316
rect 15749 25313 15761 25316
rect 15795 25313 15807 25347
rect 15749 25307 15807 25313
rect 16005 25279 16063 25285
rect 16005 25276 16017 25279
rect 14936 25248 16017 25276
rect 16005 25245 16017 25248
rect 16051 25245 16063 25279
rect 16005 25239 16063 25245
rect 16390 25236 16396 25288
rect 16448 25276 16454 25288
rect 17144 25276 17172 25384
rect 17678 25372 17684 25424
rect 17736 25412 17742 25424
rect 20073 25415 20131 25421
rect 20073 25412 20085 25415
rect 17736 25384 20085 25412
rect 17736 25372 17742 25384
rect 20073 25381 20085 25384
rect 20119 25381 20131 25415
rect 22186 25412 22192 25424
rect 22147 25384 22192 25412
rect 20073 25375 20131 25381
rect 22186 25372 22192 25384
rect 22244 25372 22250 25424
rect 17402 25304 17408 25356
rect 17460 25344 17466 25356
rect 18322 25344 18328 25356
rect 17460 25316 18328 25344
rect 17460 25304 17466 25316
rect 18322 25304 18328 25316
rect 18380 25304 18386 25356
rect 20806 25344 20812 25356
rect 18432 25316 19334 25344
rect 20767 25316 20812 25344
rect 18432 25285 18460 25316
rect 16448 25248 17172 25276
rect 18417 25279 18475 25285
rect 16448 25236 16454 25248
rect 18417 25245 18429 25279
rect 18463 25245 18475 25279
rect 18417 25239 18475 25245
rect 18509 25279 18567 25285
rect 18509 25245 18521 25279
rect 18555 25276 18567 25279
rect 18782 25276 18788 25288
rect 18555 25248 18788 25276
rect 18555 25245 18567 25248
rect 18509 25239 18567 25245
rect 18782 25236 18788 25248
rect 18840 25236 18846 25288
rect 19306 25276 19334 25316
rect 20806 25304 20812 25316
rect 20864 25304 20870 25356
rect 23106 25304 23112 25356
rect 23164 25344 23170 25356
rect 23477 25347 23535 25353
rect 23164 25316 23433 25344
rect 23164 25304 23170 25316
rect 19426 25276 19432 25288
rect 19306 25248 19432 25276
rect 19426 25236 19432 25248
rect 19484 25236 19490 25288
rect 19794 25276 19800 25288
rect 19755 25248 19800 25276
rect 19794 25236 19800 25248
rect 19852 25236 19858 25288
rect 19889 25279 19947 25285
rect 19889 25245 19901 25279
rect 19935 25276 19947 25279
rect 20070 25276 20076 25288
rect 19935 25248 20076 25276
rect 19935 25245 19947 25248
rect 19889 25239 19947 25245
rect 20070 25236 20076 25248
rect 20128 25236 20134 25288
rect 20714 25236 20720 25288
rect 20772 25276 20778 25288
rect 21065 25279 21123 25285
rect 21065 25276 21077 25279
rect 20772 25248 21077 25276
rect 20772 25236 20778 25248
rect 21065 25245 21077 25248
rect 21111 25245 21123 25279
rect 23198 25276 23204 25288
rect 21065 25239 21123 25245
rect 22480 25248 23204 25276
rect 1578 25208 1584 25220
rect 1539 25180 1584 25208
rect 1578 25168 1584 25180
rect 1636 25168 1642 25220
rect 15102 25208 15108 25220
rect 15063 25180 15108 25208
rect 15102 25168 15108 25180
rect 15160 25168 15166 25220
rect 15289 25211 15347 25217
rect 15289 25177 15301 25211
rect 15335 25208 15347 25211
rect 16206 25208 16212 25220
rect 15335 25180 16212 25208
rect 15335 25177 15347 25180
rect 15289 25171 15347 25177
rect 16206 25168 16212 25180
rect 16264 25168 16270 25220
rect 17034 25168 17040 25220
rect 17092 25208 17098 25220
rect 17678 25208 17684 25220
rect 17092 25180 17684 25208
rect 17092 25168 17098 25180
rect 17678 25168 17684 25180
rect 17736 25168 17742 25220
rect 17865 25211 17923 25217
rect 17865 25177 17877 25211
rect 17911 25208 17923 25211
rect 22480 25208 22508 25248
rect 23198 25236 23204 25248
rect 23256 25236 23262 25288
rect 23405 25276 23433 25316
rect 23477 25313 23489 25347
rect 23523 25344 23535 25347
rect 24118 25344 24124 25356
rect 23523 25316 24124 25344
rect 23523 25313 23535 25316
rect 23477 25307 23535 25313
rect 24118 25304 24124 25316
rect 24176 25344 24182 25356
rect 24596 25344 24624 25443
rect 25130 25440 25136 25452
rect 25188 25440 25194 25492
rect 25498 25480 25504 25492
rect 25459 25452 25504 25480
rect 25498 25440 25504 25452
rect 25556 25440 25562 25492
rect 26050 25440 26056 25492
rect 26108 25480 26114 25492
rect 26237 25483 26295 25489
rect 26237 25480 26249 25483
rect 26108 25452 26249 25480
rect 26108 25440 26114 25452
rect 26237 25449 26249 25452
rect 26283 25449 26295 25483
rect 26237 25443 26295 25449
rect 26418 25440 26424 25492
rect 26476 25480 26482 25492
rect 27338 25480 27344 25492
rect 26476 25452 27344 25480
rect 26476 25440 26482 25452
rect 27338 25440 27344 25452
rect 27396 25440 27402 25492
rect 27982 25480 27988 25492
rect 27943 25452 27988 25480
rect 27982 25440 27988 25452
rect 28040 25480 28046 25492
rect 28442 25480 28448 25492
rect 28040 25452 28448 25480
rect 28040 25440 28046 25452
rect 28442 25440 28448 25452
rect 28500 25440 28506 25492
rect 28997 25483 29055 25489
rect 28997 25449 29009 25483
rect 29043 25480 29055 25483
rect 31478 25480 31484 25492
rect 29043 25452 31484 25480
rect 29043 25449 29055 25452
rect 28997 25443 29055 25449
rect 31478 25440 31484 25452
rect 31536 25440 31542 25492
rect 24670 25372 24676 25424
rect 24728 25412 24734 25424
rect 24765 25415 24823 25421
rect 24765 25412 24777 25415
rect 24728 25384 24777 25412
rect 24728 25372 24734 25384
rect 24765 25381 24777 25384
rect 24811 25412 24823 25415
rect 25958 25412 25964 25424
rect 24811 25384 25964 25412
rect 24811 25381 24823 25384
rect 24765 25375 24823 25381
rect 25958 25372 25964 25384
rect 26016 25372 26022 25424
rect 26602 25372 26608 25424
rect 26660 25412 26666 25424
rect 27249 25415 27307 25421
rect 27249 25412 27261 25415
rect 26660 25384 27261 25412
rect 26660 25372 26666 25384
rect 27249 25381 27261 25384
rect 27295 25381 27307 25415
rect 27249 25375 27307 25381
rect 24176 25316 24624 25344
rect 24176 25304 24182 25316
rect 23661 25279 23719 25285
rect 23661 25276 23673 25279
rect 23405 25248 23673 25276
rect 23661 25245 23673 25248
rect 23707 25276 23719 25279
rect 23707 25251 24640 25276
rect 23707 25248 24685 25251
rect 23707 25245 23719 25248
rect 23661 25239 23719 25245
rect 24612 25245 24685 25248
rect 22646 25208 22652 25220
rect 17911 25180 22508 25208
rect 22607 25180 22652 25208
rect 17911 25177 17923 25180
rect 17865 25171 17923 25177
rect 22646 25168 22652 25180
rect 22704 25168 22710 25220
rect 22833 25211 22891 25217
rect 22833 25177 22845 25211
rect 22879 25208 22891 25211
rect 22879 25180 23536 25208
rect 22879 25177 22891 25180
rect 22833 25171 22891 25177
rect 15470 25100 15476 25152
rect 15528 25140 15534 25152
rect 18138 25140 18144 25152
rect 15528 25112 18144 25140
rect 15528 25100 15534 25112
rect 18138 25100 18144 25112
rect 18196 25100 18202 25152
rect 18230 25100 18236 25152
rect 18288 25140 18294 25152
rect 18693 25143 18751 25149
rect 18693 25140 18705 25143
rect 18288 25112 18705 25140
rect 18288 25100 18294 25112
rect 18693 25109 18705 25112
rect 18739 25109 18751 25143
rect 18693 25103 18751 25109
rect 18782 25100 18788 25152
rect 18840 25140 18846 25152
rect 20070 25140 20076 25152
rect 18840 25112 20076 25140
rect 18840 25100 18846 25112
rect 20070 25100 20076 25112
rect 20128 25100 20134 25152
rect 23017 25143 23075 25149
rect 23017 25109 23029 25143
rect 23063 25140 23075 25143
rect 23382 25140 23388 25152
rect 23063 25112 23388 25140
rect 23063 25109 23075 25112
rect 23017 25103 23075 25109
rect 23382 25100 23388 25112
rect 23440 25100 23446 25152
rect 23508 25140 23536 25180
rect 24394 25168 24400 25220
rect 24452 25208 24458 25220
rect 24612 25214 24639 25245
rect 24627 25211 24639 25214
rect 24673 25211 24685 25245
rect 25314 25236 25320 25288
rect 25372 25276 25378 25288
rect 25409 25279 25467 25285
rect 25409 25276 25421 25279
rect 25372 25248 25421 25276
rect 25372 25236 25378 25248
rect 25409 25245 25421 25248
rect 25455 25245 25467 25279
rect 25976 25276 26004 25372
rect 26050 25304 26056 25356
rect 26108 25344 26114 25356
rect 26326 25344 26332 25356
rect 26108 25316 26332 25344
rect 26108 25304 26114 25316
rect 26326 25304 26332 25316
rect 26384 25344 26390 25356
rect 28166 25344 28172 25356
rect 26384 25316 28172 25344
rect 26384 25304 26390 25316
rect 28166 25304 28172 25316
rect 28224 25304 28230 25356
rect 28350 25304 28356 25356
rect 28408 25344 28414 25356
rect 28408 25316 29592 25344
rect 28408 25304 28414 25316
rect 25976 25251 26296 25276
rect 25976 25248 26341 25251
rect 25409 25239 25467 25245
rect 26268 25245 26341 25248
rect 24452 25180 24497 25208
rect 24627 25205 24685 25211
rect 24452 25168 24458 25180
rect 24118 25140 24124 25152
rect 23508 25112 24124 25140
rect 24118 25100 24124 25112
rect 24176 25100 24182 25152
rect 25424 25140 25452 25239
rect 26050 25208 26056 25220
rect 26011 25180 26056 25208
rect 26050 25168 26056 25180
rect 26108 25168 26114 25220
rect 26268 25214 26295 25245
rect 26283 25211 26295 25214
rect 26329 25211 26341 25245
rect 26970 25236 26976 25288
rect 27028 25276 27034 25288
rect 27065 25279 27123 25285
rect 27065 25276 27077 25279
rect 27028 25248 27077 25276
rect 27028 25236 27034 25248
rect 27065 25245 27077 25248
rect 27111 25276 27123 25279
rect 27801 25279 27859 25285
rect 27801 25276 27813 25279
rect 27111 25248 27813 25276
rect 27111 25245 27123 25248
rect 27065 25239 27123 25245
rect 27801 25245 27813 25248
rect 27847 25276 27859 25279
rect 28534 25276 28540 25288
rect 27847 25248 28540 25276
rect 27847 25245 27859 25248
rect 27801 25239 27859 25245
rect 28534 25236 28540 25248
rect 28592 25236 28598 25288
rect 28718 25276 28724 25288
rect 28631 25248 28724 25276
rect 28718 25236 28724 25248
rect 28776 25236 28782 25288
rect 28810 25236 28816 25288
rect 28868 25276 28874 25288
rect 29564 25285 29592 25316
rect 31110 25304 31116 25356
rect 31168 25344 31174 25356
rect 31757 25347 31815 25353
rect 31757 25344 31769 25347
rect 31168 25316 31769 25344
rect 31168 25304 31174 25316
rect 31757 25313 31769 25316
rect 31803 25313 31815 25347
rect 31757 25307 31815 25313
rect 31846 25304 31852 25356
rect 31904 25344 31910 25356
rect 32309 25347 32367 25353
rect 31904 25316 31949 25344
rect 31904 25304 31910 25316
rect 32309 25313 32321 25347
rect 32355 25344 32367 25347
rect 34514 25344 34520 25356
rect 32355 25316 34520 25344
rect 32355 25313 32367 25316
rect 32309 25307 32367 25313
rect 34514 25304 34520 25316
rect 34572 25304 34578 25356
rect 29549 25279 29607 25285
rect 28868 25248 28961 25276
rect 28868 25236 28874 25248
rect 29549 25245 29561 25279
rect 29595 25276 29607 25279
rect 30190 25276 30196 25288
rect 29595 25248 30196 25276
rect 29595 25245 29607 25248
rect 29549 25239 29607 25245
rect 30190 25236 30196 25248
rect 30248 25236 30254 25288
rect 31478 25236 31484 25288
rect 31536 25276 31542 25288
rect 31573 25279 31631 25285
rect 31573 25276 31585 25279
rect 31536 25248 31585 25276
rect 31536 25236 31542 25248
rect 31573 25245 31585 25248
rect 31619 25245 31631 25279
rect 34146 25276 34152 25288
rect 34107 25248 34152 25276
rect 31573 25239 31631 25245
rect 34146 25236 34152 25248
rect 34204 25236 34210 25288
rect 26283 25205 26341 25211
rect 28258 25140 28264 25152
rect 25424 25112 28264 25140
rect 28258 25100 28264 25112
rect 28316 25100 28322 25152
rect 28736 25140 28764 25236
rect 28828 25208 28856 25236
rect 29638 25208 29644 25220
rect 28828 25180 29644 25208
rect 29638 25168 29644 25180
rect 29696 25168 29702 25220
rect 29816 25211 29874 25217
rect 29816 25177 29828 25211
rect 29862 25208 29874 25211
rect 30650 25208 30656 25220
rect 29862 25180 30656 25208
rect 29862 25177 29874 25180
rect 29816 25171 29874 25177
rect 30650 25168 30656 25180
rect 30708 25168 30714 25220
rect 32306 25208 32312 25220
rect 30760 25180 32312 25208
rect 30760 25140 30788 25180
rect 32306 25168 32312 25180
rect 32364 25168 32370 25220
rect 32493 25211 32551 25217
rect 32493 25177 32505 25211
rect 32539 25208 32551 25211
rect 33962 25208 33968 25220
rect 32539 25180 33968 25208
rect 32539 25177 32551 25180
rect 32493 25171 32551 25177
rect 33962 25168 33968 25180
rect 34020 25168 34026 25220
rect 30926 25140 30932 25152
rect 28736 25112 30788 25140
rect 30887 25112 30932 25140
rect 30926 25100 30932 25112
rect 30984 25100 30990 25152
rect 31386 25140 31392 25152
rect 31347 25112 31392 25140
rect 31386 25100 31392 25112
rect 31444 25100 31450 25152
rect 1104 25050 34868 25072
rect 1104 24998 12214 25050
rect 12266 24998 12278 25050
rect 12330 24998 12342 25050
rect 12394 24998 12406 25050
rect 12458 24998 12470 25050
rect 12522 24998 23478 25050
rect 23530 24998 23542 25050
rect 23594 24998 23606 25050
rect 23658 24998 23670 25050
rect 23722 24998 23734 25050
rect 23786 24998 34868 25050
rect 1104 24976 34868 24998
rect 1578 24896 1584 24948
rect 1636 24936 1642 24948
rect 2685 24939 2743 24945
rect 2685 24936 2697 24939
rect 1636 24908 2697 24936
rect 1636 24896 1642 24908
rect 2685 24905 2697 24908
rect 2731 24905 2743 24939
rect 2685 24899 2743 24905
rect 13725 24939 13783 24945
rect 13725 24905 13737 24939
rect 13771 24905 13783 24939
rect 13725 24899 13783 24905
rect 13740 24868 13768 24899
rect 14550 24896 14556 24948
rect 14608 24936 14614 24948
rect 16117 24939 16175 24945
rect 16117 24936 16129 24939
rect 14608 24908 16129 24936
rect 14608 24896 14614 24908
rect 16117 24905 16129 24908
rect 16163 24905 16175 24939
rect 16117 24899 16175 24905
rect 16298 24896 16304 24948
rect 16356 24936 16362 24948
rect 19334 24936 19340 24948
rect 16356 24908 19340 24936
rect 16356 24896 16362 24908
rect 19334 24896 19340 24908
rect 19392 24896 19398 24948
rect 21910 24896 21916 24948
rect 21968 24936 21974 24948
rect 26418 24936 26424 24948
rect 21968 24908 26424 24936
rect 21968 24896 21974 24908
rect 26418 24896 26424 24908
rect 26476 24896 26482 24948
rect 28813 24939 28871 24945
rect 28813 24936 28825 24939
rect 27632 24908 28825 24936
rect 16482 24868 16488 24880
rect 13740 24840 16488 24868
rect 1394 24760 1400 24812
rect 1452 24800 1458 24812
rect 2041 24803 2099 24809
rect 2041 24800 2053 24803
rect 1452 24772 2053 24800
rect 1452 24760 1458 24772
rect 2041 24769 2053 24772
rect 2087 24769 2099 24803
rect 2041 24763 2099 24769
rect 2593 24803 2651 24809
rect 2593 24769 2605 24803
rect 2639 24800 2651 24803
rect 4430 24800 4436 24812
rect 2639 24772 4436 24800
rect 2639 24769 2651 24772
rect 2593 24763 2651 24769
rect 4430 24760 4436 24772
rect 4488 24760 4494 24812
rect 13909 24803 13967 24809
rect 13909 24769 13921 24803
rect 13955 24800 13967 24803
rect 14553 24803 14611 24809
rect 13955 24772 14504 24800
rect 13955 24769 13967 24772
rect 13909 24763 13967 24769
rect 14476 24664 14504 24772
rect 14553 24769 14565 24803
rect 14599 24769 14611 24803
rect 14553 24763 14611 24769
rect 15105 24803 15163 24809
rect 15105 24769 15117 24803
rect 15151 24800 15163 24803
rect 15838 24800 15844 24812
rect 15151 24772 15844 24800
rect 15151 24769 15163 24772
rect 15105 24763 15163 24769
rect 14568 24732 14596 24763
rect 15838 24760 15844 24772
rect 15896 24760 15902 24812
rect 15948 24809 15976 24840
rect 16482 24828 16488 24840
rect 16540 24828 16546 24880
rect 16850 24828 16856 24880
rect 16908 24868 16914 24880
rect 16908 24840 18092 24868
rect 16908 24828 16914 24840
rect 18064 24812 18092 24840
rect 18138 24828 18144 24880
rect 18196 24868 18202 24880
rect 27632 24868 27660 24908
rect 28813 24905 28825 24908
rect 28859 24936 28871 24939
rect 31846 24936 31852 24948
rect 28859 24908 28994 24936
rect 28859 24905 28871 24908
rect 28813 24899 28871 24905
rect 18196 24840 27660 24868
rect 18196 24828 18202 24840
rect 27706 24828 27712 24880
rect 27764 24868 27770 24880
rect 27801 24871 27859 24877
rect 27801 24868 27813 24871
rect 27764 24840 27813 24868
rect 27764 24828 27770 24840
rect 27801 24837 27813 24840
rect 27847 24837 27859 24871
rect 27801 24831 27859 24837
rect 28017 24871 28075 24877
rect 28017 24837 28029 24871
rect 28063 24868 28075 24871
rect 28966 24868 28994 24908
rect 29380 24908 31852 24936
rect 29380 24877 29408 24908
rect 31846 24896 31852 24908
rect 31904 24896 31910 24948
rect 29365 24871 29423 24877
rect 28063 24840 28212 24868
rect 28966 24840 29224 24868
rect 28063 24837 28075 24840
rect 28017 24831 28075 24837
rect 15933 24803 15991 24809
rect 15933 24769 15945 24803
rect 15979 24769 15991 24803
rect 15933 24763 15991 24769
rect 16206 24760 16212 24812
rect 16264 24800 16270 24812
rect 17221 24803 17279 24809
rect 17221 24800 17233 24803
rect 16264 24772 17233 24800
rect 16264 24760 16270 24772
rect 17221 24769 17233 24772
rect 17267 24769 17279 24803
rect 17221 24763 17279 24769
rect 17405 24803 17463 24809
rect 17405 24769 17417 24803
rect 17451 24800 17463 24803
rect 17494 24800 17500 24812
rect 17451 24772 17500 24800
rect 17451 24769 17463 24772
rect 17405 24763 17463 24769
rect 17494 24760 17500 24772
rect 17552 24760 17558 24812
rect 18046 24800 18052 24812
rect 18007 24772 18052 24800
rect 18046 24760 18052 24772
rect 18104 24760 18110 24812
rect 18305 24803 18363 24809
rect 18305 24800 18317 24803
rect 18156 24772 18317 24800
rect 15746 24732 15752 24744
rect 14568 24704 15424 24732
rect 15707 24704 15752 24732
rect 15102 24664 15108 24676
rect 14476 24636 15108 24664
rect 15102 24624 15108 24636
rect 15160 24624 15166 24676
rect 15286 24664 15292 24676
rect 15247 24636 15292 24664
rect 15286 24624 15292 24636
rect 15344 24624 15350 24676
rect 15396 24664 15424 24704
rect 15746 24692 15752 24704
rect 15804 24692 15810 24744
rect 17862 24692 17868 24744
rect 17920 24732 17926 24744
rect 18156 24732 18184 24772
rect 18305 24769 18317 24772
rect 18351 24769 18363 24803
rect 18305 24763 18363 24769
rect 20346 24760 20352 24812
rect 20404 24800 20410 24812
rect 20441 24803 20499 24809
rect 20441 24800 20453 24803
rect 20404 24772 20453 24800
rect 20404 24760 20410 24772
rect 20441 24769 20453 24772
rect 20487 24769 20499 24803
rect 20714 24800 20720 24812
rect 20675 24772 20720 24800
rect 20441 24763 20499 24769
rect 20714 24760 20720 24772
rect 20772 24760 20778 24812
rect 21634 24760 21640 24812
rect 21692 24800 21698 24812
rect 21821 24803 21879 24809
rect 21821 24800 21833 24803
rect 21692 24772 21833 24800
rect 21692 24760 21698 24772
rect 21821 24769 21833 24772
rect 21867 24769 21879 24803
rect 21821 24763 21879 24769
rect 22005 24803 22063 24809
rect 22005 24769 22017 24803
rect 22051 24769 22063 24803
rect 22005 24763 22063 24769
rect 17920 24704 18184 24732
rect 17920 24692 17926 24704
rect 17589 24667 17647 24673
rect 17589 24664 17601 24667
rect 15396 24636 17601 24664
rect 17589 24633 17601 24636
rect 17635 24633 17647 24667
rect 19426 24664 19432 24676
rect 19387 24636 19432 24664
rect 17589 24627 17647 24633
rect 19426 24624 19432 24636
rect 19484 24624 19490 24676
rect 19518 24624 19524 24676
rect 19576 24664 19582 24676
rect 21818 24664 21824 24676
rect 19576 24636 21824 24664
rect 19576 24624 19582 24636
rect 21818 24624 21824 24636
rect 21876 24664 21882 24676
rect 22020 24664 22048 24763
rect 22094 24760 22100 24812
rect 22152 24800 22158 24812
rect 22833 24803 22891 24809
rect 22833 24800 22845 24803
rect 22152 24772 22845 24800
rect 22152 24760 22158 24772
rect 22833 24769 22845 24772
rect 22879 24769 22891 24803
rect 23934 24800 23940 24812
rect 23847 24772 23940 24800
rect 22833 24763 22891 24769
rect 23934 24760 23940 24772
rect 23992 24800 23998 24812
rect 25406 24800 25412 24812
rect 23992 24772 25412 24800
rect 23992 24760 23998 24772
rect 25406 24760 25412 24772
rect 25464 24760 25470 24812
rect 25501 24803 25559 24809
rect 25501 24769 25513 24803
rect 25547 24800 25559 24803
rect 25590 24800 25596 24812
rect 25547 24772 25596 24800
rect 25547 24769 25559 24772
rect 25501 24763 25559 24769
rect 25590 24760 25596 24772
rect 25648 24760 25654 24812
rect 25685 24803 25743 24809
rect 25685 24769 25697 24803
rect 25731 24769 25743 24803
rect 25685 24763 25743 24769
rect 22649 24735 22707 24741
rect 22649 24701 22661 24735
rect 22695 24732 22707 24735
rect 23014 24732 23020 24744
rect 22695 24704 23020 24732
rect 22695 24701 22707 24704
rect 22649 24695 22707 24701
rect 23014 24692 23020 24704
rect 23072 24692 23078 24744
rect 23658 24732 23664 24744
rect 23619 24704 23664 24732
rect 23658 24692 23664 24704
rect 23716 24692 23722 24744
rect 25700 24732 25728 24763
rect 25774 24760 25780 24812
rect 25832 24800 25838 24812
rect 26237 24803 26295 24809
rect 25832 24772 25877 24800
rect 25832 24760 25838 24772
rect 26237 24769 26249 24803
rect 26283 24769 26295 24803
rect 27062 24800 27068 24812
rect 27023 24772 27068 24800
rect 26237 24763 26295 24769
rect 25958 24732 25964 24744
rect 25700 24704 25964 24732
rect 25958 24692 25964 24704
rect 26016 24692 26022 24744
rect 26252 24732 26280 24763
rect 27062 24760 27068 24772
rect 27120 24760 27126 24812
rect 28184 24800 28212 24840
rect 28626 24800 28632 24812
rect 27264 24772 28120 24800
rect 28184 24772 28632 24800
rect 27264 24732 27292 24772
rect 26252 24704 27292 24732
rect 27341 24735 27399 24741
rect 27341 24701 27353 24735
rect 27387 24732 27399 24735
rect 28092 24732 28120 24772
rect 28626 24760 28632 24772
rect 28684 24760 28690 24812
rect 28718 24760 28724 24812
rect 28776 24800 28782 24812
rect 28776 24772 28821 24800
rect 28776 24760 28782 24772
rect 28994 24732 29000 24744
rect 27387 24704 28028 24732
rect 28092 24704 29000 24732
rect 27387 24701 27399 24704
rect 27341 24695 27399 24701
rect 21876 24636 22048 24664
rect 21876 24624 21882 24636
rect 22094 24624 22100 24676
rect 22152 24664 22158 24676
rect 26329 24667 26387 24673
rect 22152 24636 25452 24664
rect 22152 24624 22158 24636
rect 14369 24599 14427 24605
rect 14369 24565 14381 24599
rect 14415 24596 14427 24599
rect 17770 24596 17776 24608
rect 14415 24568 17776 24596
rect 14415 24565 14427 24568
rect 14369 24559 14427 24565
rect 17770 24556 17776 24568
rect 17828 24556 17834 24608
rect 18414 24556 18420 24608
rect 18472 24596 18478 24608
rect 22189 24599 22247 24605
rect 22189 24596 22201 24599
rect 18472 24568 22201 24596
rect 18472 24556 18478 24568
rect 22189 24565 22201 24568
rect 22235 24565 22247 24599
rect 22189 24559 22247 24565
rect 22738 24556 22744 24608
rect 22796 24596 22802 24608
rect 23017 24599 23075 24605
rect 23017 24596 23029 24599
rect 22796 24568 23029 24596
rect 22796 24556 22802 24568
rect 23017 24565 23029 24568
rect 23063 24565 23075 24599
rect 23017 24559 23075 24565
rect 23106 24556 23112 24608
rect 23164 24596 23170 24608
rect 25317 24599 25375 24605
rect 25317 24596 25329 24599
rect 23164 24568 25329 24596
rect 23164 24556 23170 24568
rect 25317 24565 25329 24568
rect 25363 24565 25375 24599
rect 25424 24596 25452 24636
rect 26329 24633 26341 24667
rect 26375 24664 26387 24667
rect 27798 24664 27804 24676
rect 26375 24636 27804 24664
rect 26375 24633 26387 24636
rect 26329 24627 26387 24633
rect 27798 24624 27804 24636
rect 27856 24624 27862 24676
rect 26694 24596 26700 24608
rect 25424 24568 26700 24596
rect 25317 24559 25375 24565
rect 26694 24556 26700 24568
rect 26752 24556 26758 24608
rect 27154 24596 27160 24608
rect 27115 24568 27160 24596
rect 27154 24556 27160 24568
rect 27212 24556 27218 24608
rect 27249 24599 27307 24605
rect 27249 24565 27261 24599
rect 27295 24596 27307 24599
rect 27890 24596 27896 24608
rect 27295 24568 27896 24596
rect 27295 24565 27307 24568
rect 27249 24559 27307 24565
rect 27890 24556 27896 24568
rect 27948 24556 27954 24608
rect 28000 24605 28028 24704
rect 28994 24692 29000 24704
rect 29052 24692 29058 24744
rect 29196 24732 29224 24840
rect 29365 24837 29377 24871
rect 29411 24837 29423 24871
rect 29565 24871 29623 24877
rect 29565 24868 29577 24871
rect 29365 24831 29423 24837
rect 29564 24837 29577 24868
rect 29611 24837 29623 24871
rect 31018 24868 31024 24880
rect 29564 24831 29623 24837
rect 30392 24840 31024 24868
rect 29564 24800 29592 24831
rect 30392 24800 30420 24840
rect 31018 24828 31024 24840
rect 31076 24828 31082 24880
rect 32030 24828 32036 24880
rect 32088 24868 32094 24880
rect 32370 24871 32428 24877
rect 32370 24868 32382 24871
rect 32088 24840 32382 24868
rect 32088 24828 32094 24840
rect 32370 24837 32382 24840
rect 32416 24837 32428 24871
rect 32370 24831 32428 24837
rect 29564 24772 30420 24800
rect 30460 24803 30518 24809
rect 30460 24769 30472 24803
rect 30506 24800 30518 24803
rect 30742 24800 30748 24812
rect 30506 24772 30748 24800
rect 30506 24769 30518 24772
rect 30460 24763 30518 24769
rect 30742 24760 30748 24772
rect 30800 24760 30806 24812
rect 31294 24760 31300 24812
rect 31352 24800 31358 24812
rect 31352 24772 33180 24800
rect 31352 24760 31358 24772
rect 30190 24732 30196 24744
rect 29196 24704 30052 24732
rect 30151 24704 30196 24732
rect 28169 24667 28227 24673
rect 28169 24633 28181 24667
rect 28215 24664 28227 24667
rect 29914 24664 29920 24676
rect 28215 24636 29920 24664
rect 28215 24633 28227 24636
rect 28169 24627 28227 24633
rect 29914 24624 29920 24636
rect 29972 24624 29978 24676
rect 27985 24599 28043 24605
rect 27985 24565 27997 24599
rect 28031 24596 28043 24599
rect 28074 24596 28080 24608
rect 28031 24568 28080 24596
rect 28031 24565 28043 24568
rect 27985 24559 28043 24565
rect 28074 24556 28080 24568
rect 28132 24556 28138 24608
rect 29454 24556 29460 24608
rect 29512 24596 29518 24608
rect 29549 24599 29607 24605
rect 29549 24596 29561 24599
rect 29512 24568 29561 24596
rect 29512 24556 29518 24568
rect 29549 24565 29561 24568
rect 29595 24565 29607 24599
rect 29730 24596 29736 24608
rect 29691 24568 29736 24596
rect 29549 24559 29607 24565
rect 29730 24556 29736 24568
rect 29788 24556 29794 24608
rect 30024 24596 30052 24704
rect 30190 24692 30196 24704
rect 30248 24692 30254 24744
rect 32122 24732 32128 24744
rect 32083 24704 32128 24732
rect 32122 24692 32128 24704
rect 32180 24692 32186 24744
rect 33152 24732 33180 24772
rect 33502 24760 33508 24812
rect 33560 24800 33566 24812
rect 33965 24803 34023 24809
rect 33965 24800 33977 24803
rect 33560 24772 33977 24800
rect 33560 24760 33566 24772
rect 33965 24769 33977 24772
rect 34011 24769 34023 24803
rect 33965 24763 34023 24769
rect 34054 24760 34060 24812
rect 34112 24800 34118 24812
rect 34112 24772 34157 24800
rect 34112 24760 34118 24772
rect 33152 24704 34100 24732
rect 34072 24676 34100 24704
rect 34054 24624 34060 24676
rect 34112 24624 34118 24676
rect 31294 24596 31300 24608
rect 30024 24568 31300 24596
rect 31294 24556 31300 24568
rect 31352 24556 31358 24608
rect 31573 24599 31631 24605
rect 31573 24565 31585 24599
rect 31619 24596 31631 24599
rect 31662 24596 31668 24608
rect 31619 24568 31668 24596
rect 31619 24565 31631 24568
rect 31573 24559 31631 24565
rect 31662 24556 31668 24568
rect 31720 24556 31726 24608
rect 32306 24556 32312 24608
rect 32364 24596 32370 24608
rect 33505 24599 33563 24605
rect 33505 24596 33517 24599
rect 32364 24568 33517 24596
rect 32364 24556 32370 24568
rect 33505 24565 33517 24568
rect 33551 24565 33563 24599
rect 33505 24559 33563 24565
rect 1104 24506 34868 24528
rect 1104 24454 6582 24506
rect 6634 24454 6646 24506
rect 6698 24454 6710 24506
rect 6762 24454 6774 24506
rect 6826 24454 6838 24506
rect 6890 24454 17846 24506
rect 17898 24454 17910 24506
rect 17962 24454 17974 24506
rect 18026 24454 18038 24506
rect 18090 24454 18102 24506
rect 18154 24454 29110 24506
rect 29162 24454 29174 24506
rect 29226 24454 29238 24506
rect 29290 24454 29302 24506
rect 29354 24454 29366 24506
rect 29418 24454 34868 24506
rect 1104 24432 34868 24454
rect 15746 24352 15752 24404
rect 15804 24392 15810 24404
rect 17497 24395 17555 24401
rect 17497 24392 17509 24395
rect 15804 24364 17509 24392
rect 15804 24352 15810 24364
rect 17497 24361 17509 24364
rect 17543 24392 17555 24395
rect 18233 24395 18291 24401
rect 17543 24364 17816 24392
rect 17543 24361 17555 24364
rect 17497 24355 17555 24361
rect 15102 24216 15108 24268
rect 15160 24256 15166 24268
rect 15838 24256 15844 24268
rect 15160 24228 15844 24256
rect 15160 24216 15166 24228
rect 15838 24216 15844 24228
rect 15896 24216 15902 24268
rect 14918 24188 14924 24200
rect 14879 24160 14924 24188
rect 14918 24148 14924 24160
rect 14976 24148 14982 24200
rect 15473 24191 15531 24197
rect 15473 24157 15485 24191
rect 15519 24188 15531 24191
rect 15562 24188 15568 24200
rect 15519 24160 15568 24188
rect 15519 24157 15531 24160
rect 15473 24151 15531 24157
rect 15562 24148 15568 24160
rect 15620 24148 15626 24200
rect 15657 24191 15715 24197
rect 15657 24157 15669 24191
rect 15703 24188 15715 24191
rect 16117 24191 16175 24197
rect 16117 24188 16129 24191
rect 15703 24160 16129 24188
rect 15703 24157 15715 24160
rect 15657 24151 15715 24157
rect 16117 24157 16129 24160
rect 16163 24188 16175 24191
rect 16163 24160 16620 24188
rect 16163 24157 16175 24160
rect 16117 24151 16175 24157
rect 16592 24132 16620 24160
rect 17402 24148 17408 24200
rect 17460 24188 17466 24200
rect 17788 24188 17816 24364
rect 18233 24361 18245 24395
rect 18279 24392 18291 24395
rect 18322 24392 18328 24404
rect 18279 24364 18328 24392
rect 18279 24361 18291 24364
rect 18233 24355 18291 24361
rect 18322 24352 18328 24364
rect 18380 24352 18386 24404
rect 18506 24352 18512 24404
rect 18564 24392 18570 24404
rect 25590 24392 25596 24404
rect 18564 24364 25596 24392
rect 18564 24352 18570 24364
rect 25590 24352 25596 24364
rect 25648 24392 25654 24404
rect 31757 24395 31815 24401
rect 25648 24364 31340 24392
rect 25648 24352 25654 24364
rect 18417 24327 18475 24333
rect 18417 24293 18429 24327
rect 18463 24293 18475 24327
rect 18417 24287 18475 24293
rect 17862 24216 17868 24268
rect 17920 24256 17926 24268
rect 18432 24256 18460 24287
rect 19794 24284 19800 24336
rect 19852 24324 19858 24336
rect 20530 24324 20536 24336
rect 19852 24296 20536 24324
rect 19852 24284 19858 24296
rect 20530 24284 20536 24296
rect 20588 24324 20594 24336
rect 21269 24327 21327 24333
rect 21269 24324 21281 24327
rect 20588 24296 21281 24324
rect 20588 24284 20594 24296
rect 21269 24293 21281 24296
rect 21315 24324 21327 24327
rect 22278 24324 22284 24336
rect 21315 24296 22284 24324
rect 21315 24293 21327 24296
rect 21269 24287 21327 24293
rect 22278 24284 22284 24296
rect 22336 24284 22342 24336
rect 23106 24324 23112 24336
rect 22388 24296 23112 24324
rect 17920 24228 18348 24256
rect 18432 24228 19840 24256
rect 17920 24216 17926 24228
rect 17957 24191 18015 24197
rect 17957 24188 17969 24191
rect 17460 24160 17969 24188
rect 17460 24148 17466 24160
rect 17957 24157 17969 24160
rect 18003 24157 18015 24191
rect 18138 24188 18144 24200
rect 18099 24160 18144 24188
rect 17957 24151 18015 24157
rect 18138 24148 18144 24160
rect 18196 24148 18202 24200
rect 18233 24191 18291 24197
rect 18233 24157 18245 24191
rect 18279 24157 18291 24191
rect 18320 24188 18348 24228
rect 19518 24188 19524 24200
rect 18320 24160 19524 24188
rect 18233 24151 18291 24157
rect 14274 24080 14280 24132
rect 14332 24120 14338 24132
rect 15102 24120 15108 24132
rect 14332 24092 15108 24120
rect 14332 24080 14338 24092
rect 15102 24080 15108 24092
rect 15160 24080 15166 24132
rect 16390 24129 16396 24132
rect 16384 24083 16396 24129
rect 16448 24120 16454 24132
rect 16448 24092 16484 24120
rect 16390 24080 16396 24083
rect 16448 24080 16454 24092
rect 16574 24080 16580 24132
rect 16632 24080 16638 24132
rect 17034 24080 17040 24132
rect 17092 24120 17098 24132
rect 18248 24120 18276 24151
rect 19518 24148 19524 24160
rect 19576 24148 19582 24200
rect 19702 24188 19708 24200
rect 19663 24160 19708 24188
rect 19702 24148 19708 24160
rect 19760 24148 19766 24200
rect 19812 24197 19840 24228
rect 21542 24216 21548 24268
rect 21600 24256 21606 24268
rect 22388 24256 22416 24296
rect 23106 24284 23112 24296
rect 23164 24284 23170 24336
rect 29546 24324 29552 24336
rect 29507 24296 29552 24324
rect 29546 24284 29552 24296
rect 29604 24284 29610 24336
rect 31312 24324 31340 24364
rect 31757 24361 31769 24395
rect 31803 24392 31815 24395
rect 31846 24392 31852 24404
rect 31803 24364 31852 24392
rect 31803 24361 31815 24364
rect 31757 24355 31815 24361
rect 31846 24352 31852 24364
rect 31904 24352 31910 24404
rect 32490 24352 32496 24404
rect 32548 24352 32554 24404
rect 32508 24324 32536 24352
rect 31312 24296 32536 24324
rect 21600 24228 22416 24256
rect 21600 24216 21606 24228
rect 22554 24216 22560 24268
rect 22612 24256 22618 24268
rect 32493 24259 32551 24265
rect 22612 24228 23520 24256
rect 22612 24216 22618 24228
rect 19797 24191 19855 24197
rect 19797 24157 19809 24191
rect 19843 24157 19855 24191
rect 19797 24151 19855 24157
rect 19889 24191 19947 24197
rect 19889 24157 19901 24191
rect 19935 24157 19947 24191
rect 20070 24188 20076 24200
rect 20031 24160 20076 24188
rect 19889 24151 19947 24157
rect 17092 24092 18276 24120
rect 17092 24080 17098 24092
rect 18414 24080 18420 24132
rect 18472 24120 18478 24132
rect 19904 24120 19932 24151
rect 20070 24148 20076 24160
rect 20128 24148 20134 24200
rect 21082 24148 21088 24200
rect 21140 24188 21146 24200
rect 21140 24160 22094 24188
rect 21140 24148 21146 24160
rect 20622 24120 20628 24132
rect 18472 24092 19840 24120
rect 19904 24092 20628 24120
rect 18472 24080 18478 24092
rect 14734 24052 14740 24064
rect 14695 24024 14740 24052
rect 14734 24012 14740 24024
rect 14792 24012 14798 24064
rect 16666 24012 16672 24064
rect 16724 24052 16730 24064
rect 17862 24052 17868 24064
rect 16724 24024 17868 24052
rect 16724 24012 16730 24024
rect 17862 24012 17868 24024
rect 17920 24012 17926 24064
rect 17954 24012 17960 24064
rect 18012 24052 18018 24064
rect 18322 24052 18328 24064
rect 18012 24024 18328 24052
rect 18012 24012 18018 24024
rect 18322 24012 18328 24024
rect 18380 24012 18386 24064
rect 19429 24055 19487 24061
rect 19429 24021 19441 24055
rect 19475 24052 19487 24055
rect 19518 24052 19524 24064
rect 19475 24024 19524 24052
rect 19475 24021 19487 24024
rect 19429 24015 19487 24021
rect 19518 24012 19524 24024
rect 19576 24012 19582 24064
rect 19812 24052 19840 24092
rect 20622 24080 20628 24092
rect 20680 24120 20686 24132
rect 20993 24123 21051 24129
rect 20993 24120 21005 24123
rect 20680 24092 21005 24120
rect 20680 24080 20686 24092
rect 20993 24089 21005 24092
rect 21039 24120 21051 24123
rect 21726 24120 21732 24132
rect 21039 24092 21732 24120
rect 21039 24089 21051 24092
rect 20993 24083 21051 24089
rect 21726 24080 21732 24092
rect 21784 24080 21790 24132
rect 22066 24120 22094 24160
rect 22186 24148 22192 24200
rect 22244 24188 22250 24200
rect 22462 24188 22468 24200
rect 22244 24160 22289 24188
rect 22423 24160 22468 24188
rect 22244 24148 22250 24160
rect 22462 24148 22468 24160
rect 22520 24148 22526 24200
rect 22830 24148 22836 24200
rect 22888 24188 22894 24200
rect 23201 24191 23259 24197
rect 23201 24188 23213 24191
rect 22888 24160 23213 24188
rect 22888 24148 22894 24160
rect 23201 24157 23213 24160
rect 23247 24157 23259 24191
rect 23382 24188 23388 24200
rect 23343 24160 23388 24188
rect 23201 24151 23259 24157
rect 23382 24148 23388 24160
rect 23440 24148 23446 24200
rect 23492 24197 23520 24228
rect 32493 24225 32505 24259
rect 32539 24256 32551 24259
rect 33134 24256 33140 24268
rect 32539 24228 33140 24256
rect 32539 24225 32551 24228
rect 32493 24219 32551 24225
rect 33134 24216 33140 24228
rect 33192 24216 33198 24268
rect 34146 24256 34152 24268
rect 34107 24228 34152 24256
rect 34146 24216 34152 24228
rect 34204 24216 34210 24268
rect 23477 24191 23535 24197
rect 23477 24157 23489 24191
rect 23523 24157 23535 24191
rect 23477 24151 23535 24157
rect 24673 24191 24731 24197
rect 24673 24157 24685 24191
rect 24719 24188 24731 24191
rect 26050 24188 26056 24200
rect 24719 24160 26056 24188
rect 24719 24157 24731 24160
rect 24673 24151 24731 24157
rect 26050 24148 26056 24160
rect 26108 24148 26114 24200
rect 26142 24148 26148 24200
rect 26200 24188 26206 24200
rect 26697 24191 26755 24197
rect 26697 24188 26709 24191
rect 26200 24160 26709 24188
rect 26200 24148 26206 24160
rect 26697 24157 26709 24160
rect 26743 24157 26755 24191
rect 26697 24151 26755 24157
rect 27617 24191 27675 24197
rect 27617 24157 27629 24191
rect 27663 24188 27675 24191
rect 28350 24188 28356 24200
rect 27663 24160 28356 24188
rect 27663 24157 27675 24160
rect 27617 24151 27675 24157
rect 28350 24148 28356 24160
rect 28408 24148 28414 24200
rect 28442 24148 28448 24200
rect 28500 24188 28506 24200
rect 28500 24160 28672 24188
rect 28500 24148 28506 24160
rect 24918 24123 24976 24129
rect 24918 24120 24930 24123
rect 22066 24092 24930 24120
rect 24918 24089 24930 24092
rect 24964 24089 24976 24123
rect 24918 24083 24976 24089
rect 25866 24080 25872 24132
rect 25924 24120 25930 24132
rect 26513 24123 26571 24129
rect 26513 24120 26525 24123
rect 25924 24092 26525 24120
rect 25924 24080 25930 24092
rect 26513 24089 26525 24092
rect 26559 24089 26571 24123
rect 26513 24083 26571 24089
rect 27884 24123 27942 24129
rect 27884 24089 27896 24123
rect 27930 24120 27942 24123
rect 28534 24120 28540 24132
rect 27930 24092 28540 24120
rect 27930 24089 27942 24092
rect 27884 24083 27942 24089
rect 28534 24080 28540 24092
rect 28592 24080 28598 24132
rect 28644 24120 28672 24160
rect 29638 24148 29644 24200
rect 29696 24188 29702 24200
rect 29825 24191 29883 24197
rect 29825 24188 29837 24191
rect 29696 24160 29837 24188
rect 29696 24148 29702 24160
rect 29825 24157 29837 24160
rect 29871 24157 29883 24191
rect 29825 24151 29883 24157
rect 30190 24148 30196 24200
rect 30248 24188 30254 24200
rect 30377 24191 30435 24197
rect 30377 24188 30389 24191
rect 30248 24160 30389 24188
rect 30248 24148 30254 24160
rect 30377 24157 30389 24160
rect 30423 24188 30435 24191
rect 32122 24188 32128 24200
rect 30423 24160 32128 24188
rect 30423 24157 30435 24160
rect 30377 24151 30435 24157
rect 32122 24148 32128 24160
rect 32180 24148 32186 24200
rect 32309 24191 32367 24197
rect 32309 24157 32321 24191
rect 32355 24157 32367 24191
rect 32309 24151 32367 24157
rect 28810 24120 28816 24132
rect 28644 24092 28816 24120
rect 28810 24080 28816 24092
rect 28868 24120 28874 24132
rect 29549 24123 29607 24129
rect 29549 24120 29561 24123
rect 28868 24092 29561 24120
rect 28868 24080 28874 24092
rect 29549 24089 29561 24092
rect 29595 24089 29607 24123
rect 29549 24083 29607 24089
rect 30644 24123 30702 24129
rect 30644 24089 30656 24123
rect 30690 24120 30702 24123
rect 31386 24120 31392 24132
rect 30690 24092 31392 24120
rect 30690 24089 30702 24092
rect 30644 24083 30702 24089
rect 31386 24080 31392 24092
rect 31444 24080 31450 24132
rect 32324 24120 32352 24151
rect 34422 24120 34428 24132
rect 32324 24092 34428 24120
rect 34422 24080 34428 24092
rect 34480 24080 34486 24132
rect 20714 24052 20720 24064
rect 19812 24024 20720 24052
rect 20714 24012 20720 24024
rect 20772 24012 20778 24064
rect 21358 24012 21364 24064
rect 21416 24052 21422 24064
rect 21453 24055 21511 24061
rect 21453 24052 21465 24055
rect 21416 24024 21465 24052
rect 21416 24012 21422 24024
rect 21453 24021 21465 24024
rect 21499 24021 21511 24055
rect 21453 24015 21511 24021
rect 21634 24012 21640 24064
rect 21692 24052 21698 24064
rect 22005 24055 22063 24061
rect 22005 24052 22017 24055
rect 21692 24024 22017 24052
rect 21692 24012 21698 24024
rect 22005 24021 22017 24024
rect 22051 24021 22063 24055
rect 22370 24052 22376 24064
rect 22331 24024 22376 24052
rect 22005 24015 22063 24021
rect 22370 24012 22376 24024
rect 22428 24052 22434 24064
rect 22922 24052 22928 24064
rect 22428 24024 22928 24052
rect 22428 24012 22434 24024
rect 22922 24012 22928 24024
rect 22980 24012 22986 24064
rect 23017 24055 23075 24061
rect 23017 24021 23029 24055
rect 23063 24052 23075 24055
rect 23382 24052 23388 24064
rect 23063 24024 23388 24052
rect 23063 24021 23075 24024
rect 23017 24015 23075 24021
rect 23382 24012 23388 24024
rect 23440 24012 23446 24064
rect 23934 24012 23940 24064
rect 23992 24052 23998 24064
rect 24118 24052 24124 24064
rect 23992 24024 24124 24052
rect 23992 24012 23998 24024
rect 24118 24012 24124 24024
rect 24176 24052 24182 24064
rect 25958 24052 25964 24064
rect 24176 24024 25964 24052
rect 24176 24012 24182 24024
rect 25958 24012 25964 24024
rect 26016 24052 26022 24064
rect 26053 24055 26111 24061
rect 26053 24052 26065 24055
rect 26016 24024 26065 24052
rect 26016 24012 26022 24024
rect 26053 24021 26065 24024
rect 26099 24021 26111 24055
rect 26878 24052 26884 24064
rect 26839 24024 26884 24052
rect 26053 24015 26111 24021
rect 26878 24012 26884 24024
rect 26936 24012 26942 24064
rect 27154 24012 27160 24064
rect 27212 24052 27218 24064
rect 28997 24055 29055 24061
rect 28997 24052 29009 24055
rect 27212 24024 29009 24052
rect 27212 24012 27218 24024
rect 28997 24021 29009 24024
rect 29043 24052 29055 24055
rect 29178 24052 29184 24064
rect 29043 24024 29184 24052
rect 29043 24021 29055 24024
rect 28997 24015 29055 24021
rect 29178 24012 29184 24024
rect 29236 24052 29242 24064
rect 29454 24052 29460 24064
rect 29236 24024 29460 24052
rect 29236 24012 29242 24024
rect 29454 24012 29460 24024
rect 29512 24012 29518 24064
rect 29730 24052 29736 24064
rect 29691 24024 29736 24052
rect 29730 24012 29736 24024
rect 29788 24012 29794 24064
rect 29914 24012 29920 24064
rect 29972 24052 29978 24064
rect 33042 24052 33048 24064
rect 29972 24024 33048 24052
rect 29972 24012 29978 24024
rect 33042 24012 33048 24024
rect 33100 24012 33106 24064
rect 1104 23962 34868 23984
rect 1104 23910 12214 23962
rect 12266 23910 12278 23962
rect 12330 23910 12342 23962
rect 12394 23910 12406 23962
rect 12458 23910 12470 23962
rect 12522 23910 23478 23962
rect 23530 23910 23542 23962
rect 23594 23910 23606 23962
rect 23658 23910 23670 23962
rect 23722 23910 23734 23962
rect 23786 23910 34868 23962
rect 1104 23888 34868 23910
rect 16666 23848 16672 23860
rect 14660 23820 16672 23848
rect 14660 23712 14688 23820
rect 16666 23808 16672 23820
rect 16724 23808 16730 23860
rect 17313 23851 17371 23857
rect 17313 23817 17325 23851
rect 17359 23848 17371 23851
rect 18138 23848 18144 23860
rect 17359 23820 18144 23848
rect 17359 23817 17371 23820
rect 17313 23811 17371 23817
rect 18138 23808 18144 23820
rect 18196 23808 18202 23860
rect 18414 23848 18420 23860
rect 18331 23820 18420 23848
rect 18331 23789 18359 23820
rect 18414 23808 18420 23820
rect 18472 23808 18478 23860
rect 18506 23808 18512 23860
rect 18564 23848 18570 23860
rect 21450 23848 21456 23860
rect 18564 23820 21456 23848
rect 18564 23808 18570 23820
rect 21450 23808 21456 23820
rect 21508 23808 21514 23860
rect 22186 23808 22192 23860
rect 22244 23848 22250 23860
rect 22465 23851 22523 23857
rect 22465 23848 22477 23851
rect 22244 23820 22477 23848
rect 22244 23808 22250 23820
rect 22465 23817 22477 23820
rect 22511 23848 22523 23851
rect 27433 23851 27491 23857
rect 22511 23820 23428 23848
rect 22511 23817 22523 23820
rect 22465 23811 22523 23817
rect 18294 23783 18359 23789
rect 18294 23780 18306 23783
rect 15672 23752 18306 23780
rect 15013 23715 15071 23721
rect 15013 23712 15025 23715
rect 14660 23684 15025 23712
rect 15013 23681 15025 23684
rect 15059 23681 15071 23715
rect 15013 23675 15071 23681
rect 14829 23579 14887 23585
rect 14829 23545 14841 23579
rect 14875 23576 14887 23579
rect 15672 23576 15700 23752
rect 18294 23749 18306 23752
rect 18340 23752 18359 23783
rect 18340 23749 18352 23752
rect 18294 23743 18352 23749
rect 18690 23740 18696 23792
rect 18748 23780 18754 23792
rect 20134 23783 20192 23789
rect 20134 23780 20146 23783
rect 18748 23752 20146 23780
rect 18748 23740 18754 23752
rect 20134 23749 20146 23752
rect 20180 23749 20192 23783
rect 20134 23743 20192 23749
rect 21174 23740 21180 23792
rect 21232 23780 21238 23792
rect 21232 23752 21956 23780
rect 21232 23740 21238 23752
rect 15933 23715 15991 23721
rect 15933 23681 15945 23715
rect 15979 23712 15991 23715
rect 16482 23712 16488 23724
rect 15979 23684 16488 23712
rect 15979 23681 15991 23684
rect 15933 23675 15991 23681
rect 16482 23672 16488 23684
rect 16540 23672 16546 23724
rect 17034 23712 17040 23724
rect 16995 23684 17040 23712
rect 17034 23672 17040 23684
rect 17092 23672 17098 23724
rect 17221 23715 17279 23721
rect 17221 23681 17233 23715
rect 17267 23681 17279 23715
rect 17402 23712 17408 23724
rect 17363 23684 17408 23712
rect 17221 23675 17279 23681
rect 15749 23647 15807 23653
rect 15749 23613 15761 23647
rect 15795 23644 15807 23647
rect 17236 23644 17264 23675
rect 17402 23672 17408 23684
rect 17460 23672 17466 23724
rect 17589 23715 17647 23721
rect 17589 23681 17601 23715
rect 17635 23712 17647 23715
rect 19610 23712 19616 23724
rect 17635 23684 19616 23712
rect 17635 23681 17647 23684
rect 17589 23675 17647 23681
rect 19610 23672 19616 23684
rect 19668 23672 19674 23724
rect 19886 23712 19892 23724
rect 19847 23684 19892 23712
rect 19886 23672 19892 23684
rect 19944 23672 19950 23724
rect 21726 23672 21732 23724
rect 21784 23712 21790 23724
rect 21821 23715 21879 23721
rect 21821 23712 21833 23715
rect 21784 23684 21833 23712
rect 21784 23672 21790 23684
rect 21821 23681 21833 23684
rect 21867 23681 21879 23715
rect 21928 23712 21956 23752
rect 22922 23740 22928 23792
rect 22980 23780 22986 23792
rect 22980 23752 23290 23780
rect 22980 23740 22986 23752
rect 22002 23712 22008 23724
rect 21928 23684 22008 23712
rect 21821 23675 21879 23681
rect 22002 23672 22008 23684
rect 22060 23712 22066 23724
rect 22189 23715 22247 23721
rect 22189 23712 22201 23715
rect 22060 23684 22201 23712
rect 22060 23672 22066 23684
rect 22189 23681 22201 23684
rect 22235 23681 22247 23715
rect 22189 23675 22247 23681
rect 22278 23672 22284 23724
rect 22336 23721 22342 23724
rect 22336 23715 22364 23721
rect 22352 23681 22364 23715
rect 22336 23675 22364 23681
rect 22336 23672 22342 23675
rect 22462 23672 22468 23724
rect 22520 23712 22526 23724
rect 23262 23721 23290 23752
rect 23400 23721 23428 23820
rect 27433 23817 27445 23851
rect 27479 23848 27491 23851
rect 27982 23848 27988 23860
rect 27479 23820 27988 23848
rect 27479 23817 27491 23820
rect 27433 23811 27491 23817
rect 27982 23808 27988 23820
rect 28040 23808 28046 23860
rect 28166 23808 28172 23860
rect 28224 23848 28230 23860
rect 28442 23848 28448 23860
rect 28224 23820 28448 23848
rect 28224 23808 28230 23820
rect 28442 23808 28448 23820
rect 28500 23808 28506 23860
rect 29730 23848 29736 23860
rect 28649 23820 29736 23848
rect 23934 23740 23940 23792
rect 23992 23780 23998 23792
rect 24305 23783 24363 23789
rect 24305 23780 24317 23783
rect 23992 23752 24317 23780
rect 23992 23740 23998 23752
rect 24305 23749 24317 23752
rect 24351 23749 24363 23783
rect 25682 23780 25688 23792
rect 24305 23743 24363 23749
rect 25240 23752 25688 23780
rect 25240 23724 25268 23752
rect 25682 23740 25688 23752
rect 25740 23740 25746 23792
rect 23101 23715 23159 23721
rect 23101 23712 23113 23715
rect 22520 23684 23113 23712
rect 22520 23672 22526 23684
rect 23101 23681 23113 23684
rect 23147 23681 23159 23715
rect 23262 23715 23332 23721
rect 23262 23684 23286 23715
rect 23101 23675 23159 23681
rect 23274 23681 23286 23684
rect 23320 23681 23332 23715
rect 23274 23675 23332 23681
rect 23385 23715 23443 23721
rect 23385 23681 23397 23715
rect 23431 23681 23443 23715
rect 23385 23675 23443 23681
rect 23474 23672 23480 23724
rect 23532 23712 23538 23724
rect 24118 23712 24124 23724
rect 23532 23684 23577 23712
rect 24079 23684 24124 23712
rect 23532 23672 23538 23684
rect 24118 23672 24124 23684
rect 24176 23672 24182 23724
rect 24397 23715 24455 23721
rect 24397 23681 24409 23715
rect 24443 23681 24455 23715
rect 25222 23712 25228 23724
rect 25135 23684 25228 23712
rect 24397 23675 24455 23681
rect 17954 23644 17960 23656
rect 15795 23616 17960 23644
rect 15795 23613 15807 23616
rect 15749 23607 15807 23613
rect 17954 23604 17960 23616
rect 18012 23604 18018 23656
rect 18049 23647 18107 23653
rect 18049 23613 18061 23647
rect 18095 23613 18107 23647
rect 22097 23647 22155 23653
rect 22097 23644 22109 23647
rect 18049 23607 18107 23613
rect 21284 23616 22109 23644
rect 14875 23548 15700 23576
rect 14875 23545 14887 23548
rect 14829 23539 14887 23545
rect 16574 23536 16580 23588
rect 16632 23576 16638 23588
rect 18064 23576 18092 23607
rect 16632 23548 18092 23576
rect 16632 23536 16638 23548
rect 15194 23468 15200 23520
rect 15252 23508 15258 23520
rect 16117 23511 16175 23517
rect 16117 23508 16129 23511
rect 15252 23480 16129 23508
rect 15252 23468 15258 23480
rect 16117 23477 16129 23480
rect 16163 23477 16175 23511
rect 18064 23508 18092 23548
rect 21284 23520 21312 23616
rect 22097 23613 22109 23616
rect 22143 23644 22155 23647
rect 22925 23647 22983 23653
rect 22143 23616 22877 23644
rect 22143 23613 22155 23616
rect 22097 23607 22155 23613
rect 22002 23536 22008 23588
rect 22060 23576 22066 23588
rect 22462 23576 22468 23588
rect 22060 23548 22468 23576
rect 22060 23536 22066 23548
rect 22462 23536 22468 23548
rect 22520 23536 22526 23588
rect 22849 23576 22877 23616
rect 22925 23613 22937 23647
rect 22971 23644 22983 23647
rect 24412 23644 24440 23675
rect 25222 23672 25228 23684
rect 25280 23672 25286 23724
rect 25409 23715 25467 23721
rect 25409 23712 25421 23715
rect 25332 23684 25421 23712
rect 22971 23616 24440 23644
rect 22971 23613 22983 23616
rect 22925 23607 22983 23613
rect 24486 23604 24492 23656
rect 24544 23644 24550 23656
rect 25332 23644 25360 23684
rect 25409 23681 25421 23684
rect 25455 23681 25467 23715
rect 25409 23675 25467 23681
rect 25777 23715 25835 23721
rect 25777 23681 25789 23715
rect 25823 23681 25835 23715
rect 25777 23675 25835 23681
rect 27249 23715 27307 23721
rect 27249 23681 27261 23715
rect 27295 23681 27307 23715
rect 27522 23712 27528 23724
rect 27483 23684 27528 23712
rect 27249 23675 27307 23681
rect 25498 23644 25504 23656
rect 24544 23616 25360 23644
rect 25459 23616 25504 23644
rect 24544 23604 24550 23616
rect 25498 23604 25504 23616
rect 25556 23604 25562 23656
rect 25593 23647 25651 23653
rect 25593 23613 25605 23647
rect 25639 23644 25651 23647
rect 25682 23644 25688 23656
rect 25639 23616 25688 23644
rect 25639 23613 25651 23616
rect 25593 23607 25651 23613
rect 25682 23604 25688 23616
rect 25740 23604 25746 23656
rect 23014 23576 23020 23588
rect 22849 23548 23020 23576
rect 23014 23536 23020 23548
rect 23072 23536 23078 23588
rect 25792 23520 25820 23675
rect 27264 23644 27292 23675
rect 27522 23672 27528 23684
rect 27580 23672 27586 23724
rect 28261 23715 28319 23721
rect 28261 23681 28273 23715
rect 28307 23681 28319 23715
rect 28261 23675 28319 23681
rect 28537 23715 28595 23721
rect 28537 23681 28549 23715
rect 28583 23712 28595 23715
rect 28649 23712 28677 23820
rect 29730 23808 29736 23820
rect 29788 23848 29794 23860
rect 29914 23848 29920 23860
rect 29788 23820 29920 23848
rect 29788 23808 29794 23820
rect 29914 23808 29920 23820
rect 29972 23808 29978 23860
rect 31110 23848 31116 23860
rect 31071 23820 31116 23848
rect 31110 23808 31116 23820
rect 31168 23808 31174 23860
rect 31294 23808 31300 23860
rect 31352 23848 31358 23860
rect 31846 23848 31852 23860
rect 31352 23820 31852 23848
rect 31352 23808 31358 23820
rect 31846 23808 31852 23820
rect 31904 23808 31910 23860
rect 28718 23740 28724 23792
rect 28776 23780 28782 23792
rect 28994 23780 29000 23792
rect 28776 23752 29000 23780
rect 28776 23740 28782 23752
rect 28994 23740 29000 23752
rect 29052 23740 29058 23792
rect 34146 23780 34152 23792
rect 34107 23752 34152 23780
rect 34146 23740 34152 23752
rect 34204 23740 34210 23792
rect 28583 23684 28677 23712
rect 30929 23715 30987 23721
rect 28583 23681 28595 23684
rect 28537 23675 28595 23681
rect 30929 23681 30941 23715
rect 30975 23712 30987 23715
rect 31018 23712 31024 23724
rect 30975 23684 31024 23712
rect 30975 23681 30987 23684
rect 30929 23675 30987 23681
rect 27706 23644 27712 23656
rect 27264 23616 27712 23644
rect 27706 23604 27712 23616
rect 27764 23604 27770 23656
rect 28077 23579 28135 23585
rect 28077 23545 28089 23579
rect 28123 23576 28135 23579
rect 28166 23576 28172 23588
rect 28123 23548 28172 23576
rect 28123 23545 28135 23548
rect 28077 23539 28135 23545
rect 28166 23536 28172 23548
rect 28224 23536 28230 23588
rect 28276 23576 28304 23675
rect 31018 23672 31024 23684
rect 31076 23672 31082 23724
rect 28445 23647 28503 23653
rect 28445 23613 28457 23647
rect 28491 23644 28503 23647
rect 29043 23647 29101 23653
rect 28491 23616 28994 23644
rect 28491 23613 28503 23616
rect 28445 23607 28503 23613
rect 28966 23576 28994 23616
rect 29043 23613 29055 23647
rect 29089 23644 29101 23647
rect 29178 23644 29184 23656
rect 29089 23616 29184 23644
rect 29089 23613 29101 23616
rect 29043 23607 29101 23613
rect 29178 23604 29184 23616
rect 29236 23604 29242 23656
rect 29273 23647 29331 23653
rect 29273 23613 29285 23647
rect 29319 23644 29331 23647
rect 29638 23644 29644 23656
rect 29319 23616 29644 23644
rect 29319 23613 29331 23616
rect 29273 23607 29331 23613
rect 29288 23576 29316 23607
rect 29638 23604 29644 23616
rect 29696 23604 29702 23656
rect 30745 23647 30803 23653
rect 30745 23613 30757 23647
rect 30791 23644 30803 23647
rect 31386 23644 31392 23656
rect 30791 23616 31392 23644
rect 30791 23613 30803 23616
rect 30745 23607 30803 23613
rect 31386 23604 31392 23616
rect 31444 23644 31450 23656
rect 31662 23644 31668 23656
rect 31444 23616 31668 23644
rect 31444 23604 31450 23616
rect 31662 23604 31668 23616
rect 31720 23604 31726 23656
rect 32306 23644 32312 23656
rect 32267 23616 32312 23644
rect 32306 23604 32312 23616
rect 32364 23604 32370 23656
rect 32490 23644 32496 23656
rect 32451 23616 32496 23644
rect 32490 23604 32496 23616
rect 32548 23604 32554 23656
rect 28276 23548 28856 23576
rect 28966 23548 29316 23576
rect 19242 23508 19248 23520
rect 18064 23480 19248 23508
rect 16117 23471 16175 23477
rect 19242 23468 19248 23480
rect 19300 23468 19306 23520
rect 19334 23468 19340 23520
rect 19392 23508 19398 23520
rect 19429 23511 19487 23517
rect 19429 23508 19441 23511
rect 19392 23480 19441 23508
rect 19392 23468 19398 23480
rect 19429 23477 19441 23480
rect 19475 23477 19487 23511
rect 21266 23508 21272 23520
rect 21227 23480 21272 23508
rect 19429 23471 19487 23477
rect 21266 23468 21272 23480
rect 21324 23468 21330 23520
rect 23937 23511 23995 23517
rect 23937 23477 23949 23511
rect 23983 23508 23995 23511
rect 24670 23508 24676 23520
rect 23983 23480 24676 23508
rect 23983 23477 23995 23480
rect 23937 23471 23995 23477
rect 24670 23468 24676 23480
rect 24728 23468 24734 23520
rect 25774 23468 25780 23520
rect 25832 23468 25838 23520
rect 25961 23511 26019 23517
rect 25961 23477 25973 23511
rect 26007 23508 26019 23511
rect 26326 23508 26332 23520
rect 26007 23480 26332 23508
rect 26007 23477 26019 23480
rect 25961 23471 26019 23477
rect 26326 23468 26332 23480
rect 26384 23468 26390 23520
rect 27065 23511 27123 23517
rect 27065 23477 27077 23511
rect 27111 23508 27123 23511
rect 28718 23508 28724 23520
rect 27111 23480 28724 23508
rect 27111 23477 27123 23480
rect 27065 23471 27123 23477
rect 28718 23468 28724 23480
rect 28776 23468 28782 23520
rect 28828 23508 28856 23548
rect 29546 23508 29552 23520
rect 28828 23480 29552 23508
rect 29546 23468 29552 23480
rect 29604 23468 29610 23520
rect 30558 23468 30564 23520
rect 30616 23508 30622 23520
rect 31662 23508 31668 23520
rect 30616 23480 31668 23508
rect 30616 23468 30622 23480
rect 31662 23468 31668 23480
rect 31720 23468 31726 23520
rect 1104 23418 34868 23440
rect 1104 23366 6582 23418
rect 6634 23366 6646 23418
rect 6698 23366 6710 23418
rect 6762 23366 6774 23418
rect 6826 23366 6838 23418
rect 6890 23366 17846 23418
rect 17898 23366 17910 23418
rect 17962 23366 17974 23418
rect 18026 23366 18038 23418
rect 18090 23366 18102 23418
rect 18154 23366 29110 23418
rect 29162 23366 29174 23418
rect 29226 23366 29238 23418
rect 29290 23366 29302 23418
rect 29354 23366 29366 23418
rect 29418 23366 34868 23418
rect 1104 23344 34868 23366
rect 14461 23307 14519 23313
rect 14461 23273 14473 23307
rect 14507 23304 14519 23307
rect 16390 23304 16396 23316
rect 14507 23276 16396 23304
rect 14507 23273 14519 23276
rect 14461 23267 14519 23273
rect 16390 23264 16396 23276
rect 16448 23264 16454 23316
rect 17957 23307 18015 23313
rect 16592 23276 17908 23304
rect 16025 23239 16083 23245
rect 16025 23205 16037 23239
rect 16071 23236 16083 23239
rect 16592 23236 16620 23276
rect 16071 23208 16620 23236
rect 17880 23236 17908 23276
rect 17957 23273 17969 23307
rect 18003 23304 18015 23307
rect 18230 23304 18236 23316
rect 18003 23276 18236 23304
rect 18003 23273 18015 23276
rect 17957 23267 18015 23273
rect 18230 23264 18236 23276
rect 18288 23264 18294 23316
rect 23474 23304 23480 23316
rect 19260 23276 20208 23304
rect 19260 23236 19288 23276
rect 17880 23208 19288 23236
rect 20180 23236 20208 23276
rect 23124 23276 23480 23304
rect 22278 23236 22284 23248
rect 20180 23208 22284 23236
rect 16071 23205 16083 23208
rect 16025 23199 16083 23205
rect 22278 23196 22284 23208
rect 22336 23196 22342 23248
rect 23124 23180 23152 23276
rect 23474 23264 23480 23276
rect 23532 23264 23538 23316
rect 24857 23307 24915 23313
rect 24857 23273 24869 23307
rect 24903 23304 24915 23307
rect 25498 23304 25504 23316
rect 24903 23276 25504 23304
rect 24903 23273 24915 23276
rect 24857 23267 24915 23273
rect 25498 23264 25504 23276
rect 25556 23264 25562 23316
rect 27522 23264 27528 23316
rect 27580 23304 27586 23316
rect 28445 23307 28503 23313
rect 28445 23304 28457 23307
rect 27580 23276 28457 23304
rect 27580 23264 27586 23276
rect 28445 23273 28457 23276
rect 28491 23273 28503 23307
rect 28445 23267 28503 23273
rect 28902 23264 28908 23316
rect 28960 23304 28966 23316
rect 29730 23304 29736 23316
rect 28960 23276 29736 23304
rect 28960 23264 28966 23276
rect 29730 23264 29736 23276
rect 29788 23264 29794 23316
rect 29914 23264 29920 23316
rect 29972 23304 29978 23316
rect 30929 23307 30987 23313
rect 30929 23304 30941 23307
rect 29972 23276 30941 23304
rect 29972 23264 29978 23276
rect 30929 23273 30941 23276
rect 30975 23273 30987 23307
rect 30929 23267 30987 23273
rect 31294 23264 31300 23316
rect 31352 23304 31358 23316
rect 31481 23307 31539 23313
rect 31481 23304 31493 23307
rect 31352 23276 31493 23304
rect 31352 23264 31358 23276
rect 31481 23273 31493 23276
rect 31527 23273 31539 23307
rect 31481 23267 31539 23273
rect 23308 23208 25719 23236
rect 16574 23168 16580 23180
rect 16535 23140 16580 23168
rect 16574 23128 16580 23140
rect 16632 23128 16638 23180
rect 17696 23140 19380 23168
rect 14645 23103 14703 23109
rect 14645 23069 14657 23103
rect 14691 23100 14703 23103
rect 15194 23100 15200 23112
rect 14691 23072 15200 23100
rect 14691 23069 14703 23072
rect 14645 23063 14703 23069
rect 15194 23060 15200 23072
rect 15252 23060 15258 23112
rect 15289 23103 15347 23109
rect 15289 23069 15301 23103
rect 15335 23100 15347 23103
rect 15838 23100 15844 23112
rect 15335 23072 15844 23100
rect 15335 23069 15347 23072
rect 15289 23063 15347 23069
rect 15838 23060 15844 23072
rect 15896 23060 15902 23112
rect 15933 23103 15991 23109
rect 15933 23069 15945 23103
rect 15979 23069 15991 23103
rect 15933 23063 15991 23069
rect 16117 23103 16175 23109
rect 16117 23069 16129 23103
rect 16163 23100 16175 23103
rect 17696 23100 17724 23140
rect 16163 23072 17724 23100
rect 16163 23069 16175 23072
rect 16117 23063 16175 23069
rect 15948 23032 15976 23063
rect 17770 23060 17776 23112
rect 17828 23100 17834 23112
rect 18417 23103 18475 23109
rect 18417 23100 18429 23103
rect 17828 23072 18429 23100
rect 17828 23060 17834 23072
rect 18417 23069 18429 23072
rect 18463 23069 18475 23103
rect 19242 23100 19248 23112
rect 19203 23072 19248 23100
rect 18417 23063 18475 23069
rect 19242 23060 19248 23072
rect 19300 23060 19306 23112
rect 19352 23100 19380 23140
rect 20714 23128 20720 23180
rect 20772 23168 20778 23180
rect 20772 23140 21220 23168
rect 20772 23128 20778 23140
rect 20990 23100 20996 23112
rect 19352 23072 20996 23100
rect 20990 23060 20996 23072
rect 21048 23060 21054 23112
rect 16390 23032 16396 23044
rect 15948 23004 16396 23032
rect 16390 22992 16396 23004
rect 16448 22992 16454 23044
rect 16844 23035 16902 23041
rect 16844 23001 16856 23035
rect 16890 23032 16902 23035
rect 16942 23032 16948 23044
rect 16890 23004 16948 23032
rect 16890 23001 16902 23004
rect 16844 22995 16902 23001
rect 16942 22992 16948 23004
rect 17000 22992 17006 23044
rect 19058 22992 19064 23044
rect 19116 23032 19122 23044
rect 21192 23041 21220 23140
rect 21358 23128 21364 23180
rect 21416 23168 21422 23180
rect 22097 23171 22155 23177
rect 22097 23168 22109 23171
rect 21416 23140 22109 23168
rect 21416 23128 21422 23140
rect 22097 23137 22109 23140
rect 22143 23137 22155 23171
rect 22097 23131 22155 23137
rect 22189 23171 22247 23177
rect 22189 23137 22201 23171
rect 22235 23168 22247 23171
rect 22738 23168 22744 23180
rect 22235 23140 22744 23168
rect 22235 23137 22247 23140
rect 22189 23131 22247 23137
rect 22738 23128 22744 23140
rect 22796 23128 22802 23180
rect 23017 23171 23075 23177
rect 23017 23137 23029 23171
rect 23063 23168 23075 23171
rect 23106 23168 23112 23180
rect 23063 23140 23112 23168
rect 23063 23137 23075 23140
rect 23017 23131 23075 23137
rect 23106 23128 23112 23140
rect 23164 23128 23170 23180
rect 23198 23128 23204 23180
rect 23256 23168 23262 23180
rect 23308 23177 23336 23208
rect 23293 23171 23351 23177
rect 23293 23168 23305 23171
rect 23256 23140 23305 23168
rect 23256 23128 23262 23140
rect 23293 23137 23305 23140
rect 23339 23137 23351 23171
rect 25130 23168 25136 23180
rect 23293 23131 23351 23137
rect 24035 23140 25136 23168
rect 21818 23100 21824 23112
rect 21779 23072 21824 23100
rect 21818 23060 21824 23072
rect 21876 23060 21882 23112
rect 22002 23100 22008 23112
rect 21963 23072 22008 23100
rect 22002 23060 22008 23072
rect 22060 23060 22066 23112
rect 22384 23103 22442 23109
rect 22384 23069 22396 23103
rect 22430 23069 22442 23103
rect 22384 23063 22442 23069
rect 19490 23035 19548 23041
rect 19490 23032 19502 23035
rect 19116 23004 19502 23032
rect 19116 22992 19122 23004
rect 19490 23001 19502 23004
rect 19536 23001 19548 23035
rect 19490 22995 19548 23001
rect 21177 23035 21235 23041
rect 21177 23001 21189 23035
rect 21223 23001 21235 23035
rect 21177 22995 21235 23001
rect 21361 23035 21419 23041
rect 21361 23001 21373 23035
rect 21407 23032 21419 23035
rect 21542 23032 21548 23044
rect 21407 23004 21548 23032
rect 21407 23001 21419 23004
rect 21361 22995 21419 23001
rect 21542 22992 21548 23004
rect 21600 22992 21606 23044
rect 22186 22992 22192 23044
rect 22244 23032 22250 23044
rect 22388 23032 22416 23063
rect 22922 23060 22928 23112
rect 22980 23100 22986 23112
rect 24035 23100 24063 23140
rect 25130 23128 25136 23140
rect 25188 23128 25194 23180
rect 25225 23171 25283 23177
rect 25225 23137 25237 23171
rect 25271 23168 25283 23171
rect 25406 23168 25412 23180
rect 25271 23140 25412 23168
rect 25271 23137 25283 23140
rect 25225 23131 25283 23137
rect 22980 23072 24063 23100
rect 22980 23060 22986 23072
rect 24946 23060 24952 23112
rect 25004 23100 25010 23112
rect 25041 23103 25099 23109
rect 25041 23100 25053 23103
rect 25004 23072 25053 23100
rect 25004 23060 25010 23072
rect 25041 23069 25053 23072
rect 25087 23069 25099 23103
rect 25041 23063 25099 23069
rect 22244 23004 22416 23032
rect 22244 22992 22250 23004
rect 23014 22992 23020 23044
rect 23072 23032 23078 23044
rect 25240 23032 25268 23131
rect 25406 23128 25412 23140
rect 25464 23128 25470 23180
rect 25317 23103 25375 23109
rect 25317 23069 25329 23103
rect 25363 23100 25375 23103
rect 25590 23100 25596 23112
rect 25363 23072 25596 23100
rect 25363 23069 25375 23072
rect 25317 23063 25375 23069
rect 25590 23060 25596 23072
rect 25648 23060 25654 23112
rect 23072 23004 25268 23032
rect 25691 23032 25719 23208
rect 28166 23196 28172 23248
rect 28224 23236 28230 23248
rect 29362 23236 29368 23248
rect 28224 23208 28396 23236
rect 28224 23196 28230 23208
rect 27798 23128 27804 23180
rect 27856 23168 27862 23180
rect 27856 23140 28304 23168
rect 27856 23128 27862 23140
rect 26050 23100 26056 23112
rect 26011 23072 26056 23100
rect 26050 23060 26056 23072
rect 26108 23060 26114 23112
rect 26326 23109 26332 23112
rect 26320 23100 26332 23109
rect 26287 23072 26332 23100
rect 26320 23063 26332 23072
rect 26326 23060 26332 23063
rect 26384 23060 26390 23112
rect 27890 23100 27896 23112
rect 27851 23072 27896 23100
rect 27890 23060 27896 23072
rect 27948 23060 27954 23112
rect 28276 23109 28304 23140
rect 28261 23103 28319 23109
rect 28000 23072 28212 23100
rect 28000 23032 28028 23072
rect 28184 23044 28212 23072
rect 28261 23069 28273 23103
rect 28307 23069 28319 23103
rect 28261 23063 28319 23069
rect 25691 23004 28028 23032
rect 28077 23035 28135 23041
rect 23072 22992 23078 23004
rect 28077 23001 28089 23035
rect 28123 23001 28135 23035
rect 28077 22995 28135 23001
rect 15105 22967 15163 22973
rect 15105 22933 15117 22967
rect 15151 22964 15163 22967
rect 16482 22964 16488 22976
rect 15151 22936 16488 22964
rect 15151 22933 15163 22936
rect 15105 22927 15163 22933
rect 16482 22924 16488 22936
rect 16540 22924 16546 22976
rect 18601 22967 18659 22973
rect 18601 22933 18613 22967
rect 18647 22964 18659 22967
rect 20438 22964 20444 22976
rect 18647 22936 20444 22964
rect 18647 22933 18659 22936
rect 18601 22927 18659 22933
rect 20438 22924 20444 22936
rect 20496 22924 20502 22976
rect 20622 22964 20628 22976
rect 20583 22936 20628 22964
rect 20622 22924 20628 22936
rect 20680 22924 20686 22976
rect 20806 22924 20812 22976
rect 20864 22964 20870 22976
rect 22557 22967 22615 22973
rect 22557 22964 22569 22967
rect 20864 22936 22569 22964
rect 20864 22924 20870 22936
rect 22557 22933 22569 22936
rect 22603 22964 22615 22967
rect 24118 22964 24124 22976
rect 22603 22936 24124 22964
rect 22603 22933 22615 22936
rect 22557 22927 22615 22933
rect 24118 22924 24124 22936
rect 24176 22924 24182 22976
rect 27433 22967 27491 22973
rect 27433 22933 27445 22967
rect 27479 22964 27491 22967
rect 27522 22964 27528 22976
rect 27479 22936 27528 22964
rect 27479 22933 27491 22936
rect 27433 22927 27491 22933
rect 27522 22924 27528 22936
rect 27580 22924 27586 22976
rect 28092 22964 28120 22995
rect 28166 22992 28172 23044
rect 28224 23032 28230 23044
rect 28368 23032 28396 23208
rect 28828 23208 29368 23236
rect 28828 23032 28856 23208
rect 29362 23196 29368 23208
rect 29420 23196 29426 23248
rect 28902 23128 28908 23180
rect 28960 23168 28966 23180
rect 28960 23140 29684 23168
rect 28960 23128 28966 23140
rect 28994 23060 29000 23112
rect 29052 23100 29058 23112
rect 29549 23103 29607 23109
rect 29549 23100 29561 23103
rect 29052 23072 29561 23100
rect 29052 23060 29058 23072
rect 29549 23069 29561 23072
rect 29595 23069 29607 23103
rect 29656 23100 29684 23140
rect 31294 23128 31300 23180
rect 31352 23168 31358 23180
rect 31665 23171 31723 23177
rect 31665 23168 31677 23171
rect 31352 23140 31677 23168
rect 31352 23128 31358 23140
rect 31665 23137 31677 23140
rect 31711 23168 31723 23171
rect 32030 23168 32036 23180
rect 31711 23140 32036 23168
rect 31711 23137 31723 23140
rect 31665 23131 31723 23137
rect 32030 23128 32036 23140
rect 32088 23168 32094 23180
rect 33318 23168 33324 23180
rect 32088 23140 33324 23168
rect 32088 23128 32094 23140
rect 33318 23128 33324 23140
rect 33376 23128 33382 23180
rect 34146 23168 34152 23180
rect 34107 23140 34152 23168
rect 34146 23128 34152 23140
rect 34204 23128 34210 23180
rect 31389 23103 31447 23109
rect 31389 23100 31401 23103
rect 29656 23072 31401 23100
rect 29549 23063 29607 23069
rect 31389 23069 31401 23072
rect 31435 23069 31447 23103
rect 31389 23063 31447 23069
rect 32309 23103 32367 23109
rect 32309 23069 32321 23103
rect 32355 23069 32367 23103
rect 32309 23063 32367 23069
rect 28224 23004 28317 23032
rect 28368 23004 28856 23032
rect 28224 22992 28230 23004
rect 29362 22992 29368 23044
rect 29420 23032 29426 23044
rect 29794 23035 29852 23041
rect 29794 23032 29806 23035
rect 29420 23004 29806 23032
rect 29420 22992 29426 23004
rect 29794 23001 29806 23004
rect 29840 23001 29852 23035
rect 29794 22995 29852 23001
rect 30558 22992 30564 23044
rect 30616 23032 30622 23044
rect 32324 23032 32352 23063
rect 30616 23004 32352 23032
rect 32493 23035 32551 23041
rect 30616 22992 30622 23004
rect 32493 23001 32505 23035
rect 32539 23032 32551 23035
rect 33686 23032 33692 23044
rect 32539 23004 33692 23032
rect 32539 23001 32551 23004
rect 32493 22995 32551 23001
rect 33686 22992 33692 23004
rect 33744 22992 33750 23044
rect 30190 22964 30196 22976
rect 28092 22936 30196 22964
rect 30190 22924 30196 22936
rect 30248 22924 30254 22976
rect 30374 22924 30380 22976
rect 30432 22964 30438 22976
rect 31665 22967 31723 22973
rect 31665 22964 31677 22967
rect 30432 22936 31677 22964
rect 30432 22924 30438 22936
rect 31665 22933 31677 22936
rect 31711 22933 31723 22967
rect 31665 22927 31723 22933
rect 1104 22874 34868 22896
rect 1104 22822 12214 22874
rect 12266 22822 12278 22874
rect 12330 22822 12342 22874
rect 12394 22822 12406 22874
rect 12458 22822 12470 22874
rect 12522 22822 23478 22874
rect 23530 22822 23542 22874
rect 23594 22822 23606 22874
rect 23658 22822 23670 22874
rect 23722 22822 23734 22874
rect 23786 22822 34868 22874
rect 1104 22800 34868 22822
rect 14366 22720 14372 22772
rect 14424 22760 14430 22772
rect 17770 22760 17776 22772
rect 14424 22732 17776 22760
rect 14424 22720 14430 22732
rect 17770 22720 17776 22732
rect 17828 22720 17834 22772
rect 18049 22763 18107 22769
rect 18049 22729 18061 22763
rect 18095 22760 18107 22763
rect 18322 22760 18328 22772
rect 18095 22732 18328 22760
rect 18095 22729 18107 22732
rect 18049 22723 18107 22729
rect 18322 22720 18328 22732
rect 18380 22720 18386 22772
rect 19058 22760 19064 22772
rect 19019 22732 19064 22760
rect 19058 22720 19064 22732
rect 19116 22720 19122 22772
rect 20257 22763 20315 22769
rect 20257 22729 20269 22763
rect 20303 22760 20315 22763
rect 21910 22760 21916 22772
rect 20303 22732 21916 22760
rect 20303 22729 20315 22732
rect 20257 22723 20315 22729
rect 21910 22720 21916 22732
rect 21968 22720 21974 22772
rect 23106 22720 23112 22772
rect 23164 22760 23170 22772
rect 23569 22763 23627 22769
rect 23569 22760 23581 22763
rect 23164 22732 23581 22760
rect 23164 22720 23170 22732
rect 23569 22729 23581 22732
rect 23615 22729 23627 22763
rect 23569 22723 23627 22729
rect 24854 22720 24860 22772
rect 24912 22760 24918 22772
rect 24912 22732 25176 22760
rect 24912 22720 24918 22732
rect 16117 22695 16175 22701
rect 16117 22692 16129 22695
rect 15304 22664 16129 22692
rect 15304 22633 15332 22664
rect 16117 22661 16129 22664
rect 16163 22661 16175 22695
rect 16117 22655 16175 22661
rect 16390 22652 16396 22704
rect 16448 22692 16454 22704
rect 16574 22692 16580 22704
rect 16448 22664 16580 22692
rect 16448 22652 16454 22664
rect 16574 22652 16580 22664
rect 16632 22652 16638 22704
rect 16758 22692 16764 22704
rect 16684 22664 16764 22692
rect 15289 22627 15347 22633
rect 15289 22593 15301 22627
rect 15335 22593 15347 22627
rect 15289 22587 15347 22593
rect 15933 22627 15991 22633
rect 15933 22593 15945 22627
rect 15979 22624 15991 22627
rect 16482 22624 16488 22636
rect 15979 22596 16488 22624
rect 15979 22593 15991 22596
rect 15933 22587 15991 22593
rect 16482 22584 16488 22596
rect 16540 22584 16546 22636
rect 16684 22633 16712 22664
rect 16758 22652 16764 22664
rect 16816 22652 16822 22704
rect 19242 22652 19248 22704
rect 19300 22692 19306 22704
rect 23934 22692 23940 22704
rect 19300 22664 22094 22692
rect 19300 22652 19306 22664
rect 16669 22627 16727 22633
rect 16669 22593 16681 22627
rect 16715 22593 16727 22627
rect 16925 22627 16983 22633
rect 16925 22624 16937 22627
rect 16669 22587 16727 22593
rect 16776 22596 16937 22624
rect 15749 22559 15807 22565
rect 15749 22525 15761 22559
rect 15795 22556 15807 22559
rect 16574 22556 16580 22568
rect 15795 22528 16580 22556
rect 15795 22525 15807 22528
rect 15749 22519 15807 22525
rect 16574 22516 16580 22528
rect 16632 22516 16638 22568
rect 16776 22556 16804 22596
rect 16925 22593 16937 22596
rect 16971 22593 16983 22627
rect 16925 22587 16983 22593
rect 18414 22584 18420 22636
rect 18472 22624 18478 22636
rect 19337 22627 19395 22633
rect 19337 22624 19349 22627
rect 18472 22596 19349 22624
rect 18472 22584 18478 22596
rect 19337 22593 19349 22596
rect 19383 22593 19395 22627
rect 19518 22624 19524 22636
rect 19479 22596 19524 22624
rect 19337 22587 19395 22593
rect 19518 22584 19524 22596
rect 19576 22584 19582 22636
rect 20070 22624 20076 22636
rect 20031 22596 20076 22624
rect 20070 22584 20076 22596
rect 20128 22584 20134 22636
rect 20346 22624 20352 22636
rect 20307 22596 20352 22624
rect 20346 22584 20352 22596
rect 20404 22584 20410 22636
rect 22066 22624 22094 22664
rect 22278 22664 23940 22692
rect 22189 22627 22247 22633
rect 22189 22624 22201 22627
rect 22066 22596 22201 22624
rect 22189 22593 22201 22596
rect 22235 22593 22247 22627
rect 22189 22587 22247 22593
rect 16684 22528 16804 22556
rect 15105 22491 15163 22497
rect 15105 22457 15117 22491
rect 15151 22488 15163 22491
rect 16684 22488 16712 22528
rect 19150 22516 19156 22568
rect 19208 22556 19214 22568
rect 19245 22559 19303 22565
rect 19245 22556 19257 22559
rect 19208 22528 19257 22556
rect 19208 22516 19214 22528
rect 19245 22525 19257 22528
rect 19291 22525 19303 22559
rect 19245 22519 19303 22525
rect 19429 22559 19487 22565
rect 19429 22525 19441 22559
rect 19475 22556 19487 22559
rect 19794 22556 19800 22568
rect 19475 22528 19800 22556
rect 19475 22525 19487 22528
rect 19429 22519 19487 22525
rect 19794 22516 19800 22528
rect 19852 22516 19858 22568
rect 20530 22516 20536 22568
rect 20588 22556 20594 22568
rect 20809 22559 20867 22565
rect 20809 22556 20821 22559
rect 20588 22528 20821 22556
rect 20588 22516 20594 22528
rect 20809 22525 20821 22528
rect 20855 22525 20867 22559
rect 20809 22519 20867 22525
rect 20990 22516 20996 22568
rect 21048 22556 21054 22568
rect 22278 22556 22306 22664
rect 23934 22652 23940 22664
rect 23992 22652 23998 22704
rect 22456 22627 22514 22633
rect 22456 22593 22468 22627
rect 22502 22624 22514 22627
rect 22922 22624 22928 22636
rect 22502 22596 22928 22624
rect 22502 22593 22514 22596
rect 22456 22587 22514 22593
rect 22922 22584 22928 22596
rect 22980 22584 22986 22636
rect 24029 22627 24087 22633
rect 24029 22593 24041 22627
rect 24075 22593 24087 22627
rect 24029 22587 24087 22593
rect 24121 22627 24179 22633
rect 24121 22593 24133 22627
rect 24167 22624 24179 22627
rect 24394 22624 24400 22636
rect 24167 22596 24400 22624
rect 24167 22593 24179 22596
rect 24121 22587 24179 22593
rect 21048 22528 22306 22556
rect 24044 22556 24072 22587
rect 24394 22584 24400 22596
rect 24452 22584 24458 22636
rect 24578 22584 24584 22636
rect 24636 22624 24642 22636
rect 24903 22627 24961 22633
rect 24903 22624 24915 22627
rect 24636 22596 24915 22624
rect 24636 22584 24642 22596
rect 24903 22593 24915 22596
rect 24949 22593 24961 22627
rect 25038 22624 25044 22636
rect 24999 22596 25044 22624
rect 24903 22587 24961 22593
rect 25038 22584 25044 22596
rect 25096 22584 25102 22636
rect 25148 22633 25176 22732
rect 28258 22720 28264 22772
rect 28316 22760 28322 22772
rect 28629 22763 28687 22769
rect 28629 22760 28641 22763
rect 28316 22732 28641 22760
rect 28316 22720 28322 22732
rect 28629 22729 28641 22732
rect 28675 22729 28687 22763
rect 28629 22723 28687 22729
rect 28902 22720 28908 22772
rect 28960 22760 28966 22772
rect 30558 22760 30564 22772
rect 28960 22732 30564 22760
rect 28960 22720 28966 22732
rect 30558 22720 30564 22732
rect 30616 22720 30622 22772
rect 31021 22763 31079 22769
rect 31021 22729 31033 22763
rect 31067 22729 31079 22763
rect 31021 22723 31079 22729
rect 25222 22652 25228 22704
rect 25280 22692 25286 22704
rect 25590 22692 25596 22704
rect 25280 22664 25596 22692
rect 25280 22652 25286 22664
rect 25590 22652 25596 22664
rect 25648 22652 25654 22704
rect 25866 22652 25872 22704
rect 25924 22692 25930 22704
rect 29448 22695 29506 22701
rect 25924 22664 26096 22692
rect 25924 22652 25930 22664
rect 25133 22627 25191 22633
rect 25133 22593 25145 22627
rect 25179 22593 25191 22627
rect 25133 22587 25191 22593
rect 25317 22627 25375 22633
rect 25317 22593 25329 22627
rect 25363 22624 25375 22627
rect 25498 22624 25504 22636
rect 25363 22596 25504 22624
rect 25363 22593 25375 22596
rect 25317 22587 25375 22593
rect 25498 22584 25504 22596
rect 25556 22584 25562 22636
rect 25958 22624 25964 22636
rect 25919 22596 25964 22624
rect 25958 22584 25964 22596
rect 26016 22584 26022 22636
rect 26068 22633 26096 22664
rect 29448 22661 29460 22695
rect 29494 22692 29506 22695
rect 31036 22692 31064 22723
rect 31662 22720 31668 22772
rect 31720 22760 31726 22772
rect 32309 22763 32367 22769
rect 32309 22760 32321 22763
rect 31720 22732 32321 22760
rect 31720 22720 31726 22732
rect 32309 22729 32321 22732
rect 32355 22729 32367 22763
rect 32309 22723 32367 22729
rect 29494 22664 31064 22692
rect 29494 22661 29506 22664
rect 29448 22655 29506 22661
rect 31294 22652 31300 22704
rect 31352 22692 31358 22704
rect 33137 22695 33195 22701
rect 33137 22692 33149 22695
rect 31352 22664 33149 22692
rect 31352 22652 31358 22664
rect 33137 22661 33149 22664
rect 33183 22661 33195 22695
rect 33137 22655 33195 22661
rect 26053 22627 26111 22633
rect 26053 22593 26065 22627
rect 26099 22593 26111 22627
rect 26053 22587 26111 22593
rect 28442 22584 28448 22636
rect 28500 22624 28506 22636
rect 28537 22627 28595 22633
rect 28537 22624 28549 22627
rect 28500 22596 28549 22624
rect 28500 22584 28506 22596
rect 28537 22593 28549 22596
rect 28583 22593 28595 22627
rect 30374 22624 30380 22636
rect 28537 22587 28595 22593
rect 28635 22596 30380 22624
rect 26142 22556 26148 22568
rect 24044 22528 25912 22556
rect 26103 22528 26148 22556
rect 21048 22516 21054 22528
rect 15151 22460 16712 22488
rect 15151 22457 15163 22460
rect 15105 22451 15163 22457
rect 20622 22448 20628 22500
rect 20680 22488 20686 22500
rect 21085 22491 21143 22497
rect 21085 22488 21097 22491
rect 20680 22460 21097 22488
rect 20680 22448 20686 22460
rect 21085 22457 21097 22460
rect 21131 22457 21143 22491
rect 21085 22451 21143 22457
rect 21192 22460 22232 22488
rect 16574 22380 16580 22432
rect 16632 22420 16638 22432
rect 17034 22420 17040 22432
rect 16632 22392 17040 22420
rect 16632 22380 16638 22392
rect 17034 22380 17040 22392
rect 17092 22380 17098 22432
rect 17770 22380 17776 22432
rect 17828 22420 17834 22432
rect 19978 22420 19984 22432
rect 17828 22392 19984 22420
rect 17828 22380 17834 22392
rect 19978 22380 19984 22392
rect 20036 22380 20042 22432
rect 20073 22423 20131 22429
rect 20073 22389 20085 22423
rect 20119 22420 20131 22423
rect 21192 22420 21220 22460
rect 20119 22392 21220 22420
rect 21269 22423 21327 22429
rect 20119 22389 20131 22392
rect 20073 22383 20131 22389
rect 21269 22389 21281 22423
rect 21315 22420 21327 22423
rect 22094 22420 22100 22432
rect 21315 22392 22100 22420
rect 21315 22389 21327 22392
rect 21269 22383 21327 22389
rect 22094 22380 22100 22392
rect 22152 22380 22158 22432
rect 22204 22420 22232 22460
rect 24302 22448 24308 22500
rect 24360 22488 24366 22500
rect 25777 22491 25835 22497
rect 25777 22488 25789 22491
rect 24360 22460 25789 22488
rect 24360 22448 24366 22460
rect 25777 22457 25789 22460
rect 25823 22457 25835 22491
rect 25884 22488 25912 22528
rect 26142 22516 26148 22528
rect 26200 22516 26206 22568
rect 26234 22516 26240 22568
rect 26292 22556 26298 22568
rect 27246 22556 27252 22568
rect 26292 22528 26337 22556
rect 27207 22528 27252 22556
rect 26292 22516 26298 22528
rect 27246 22516 27252 22528
rect 27304 22516 27310 22568
rect 27338 22516 27344 22568
rect 27396 22556 27402 22568
rect 27525 22559 27583 22565
rect 27525 22556 27537 22559
rect 27396 22528 27537 22556
rect 27396 22516 27402 22528
rect 27525 22525 27537 22528
rect 27571 22525 27583 22559
rect 27525 22519 27583 22525
rect 27982 22516 27988 22568
rect 28040 22556 28046 22568
rect 28635 22556 28663 22596
rect 30374 22584 30380 22596
rect 30432 22584 30438 22636
rect 30466 22584 30472 22636
rect 30524 22624 30530 22636
rect 31021 22627 31079 22633
rect 31021 22624 31033 22627
rect 30524 22596 31033 22624
rect 30524 22584 30530 22596
rect 31021 22593 31033 22596
rect 31067 22593 31079 22627
rect 32125 22627 32183 22633
rect 32125 22624 32137 22627
rect 31021 22587 31079 22593
rect 31128 22596 32137 22624
rect 28040 22528 28663 22556
rect 28040 22516 28046 22528
rect 28994 22516 29000 22568
rect 29052 22556 29058 22568
rect 29181 22559 29239 22565
rect 29181 22556 29193 22559
rect 29052 22528 29193 22556
rect 29052 22516 29058 22528
rect 29181 22525 29193 22528
rect 29227 22525 29239 22559
rect 29181 22519 29239 22525
rect 30926 22516 30932 22568
rect 30984 22556 30990 22568
rect 31128 22556 31156 22596
rect 32125 22593 32137 22596
rect 32171 22593 32183 22627
rect 32401 22627 32459 22633
rect 32401 22624 32413 22627
rect 32125 22587 32183 22593
rect 32324 22596 32413 22624
rect 30984 22528 31156 22556
rect 31297 22559 31355 22565
rect 30984 22516 30990 22528
rect 31297 22525 31309 22559
rect 31343 22556 31355 22559
rect 31846 22556 31852 22568
rect 31343 22528 31852 22556
rect 31343 22525 31355 22528
rect 31297 22519 31355 22525
rect 31846 22516 31852 22528
rect 31904 22516 31910 22568
rect 25884 22460 27614 22488
rect 25777 22451 25835 22457
rect 24486 22420 24492 22432
rect 22204 22392 24492 22420
rect 24486 22380 24492 22392
rect 24544 22380 24550 22432
rect 24673 22423 24731 22429
rect 24673 22389 24685 22423
rect 24719 22420 24731 22423
rect 26326 22420 26332 22432
rect 24719 22392 26332 22420
rect 24719 22389 24731 22392
rect 24673 22383 24731 22389
rect 26326 22380 26332 22392
rect 26384 22380 26390 22432
rect 27586 22420 27614 22460
rect 30374 22448 30380 22500
rect 30432 22488 30438 22500
rect 31113 22491 31171 22497
rect 31113 22488 31125 22491
rect 30432 22460 31125 22488
rect 30432 22448 30438 22460
rect 31113 22457 31125 22460
rect 31159 22457 31171 22491
rect 32324 22488 32352 22596
rect 32401 22593 32413 22596
rect 32447 22593 32459 22627
rect 32401 22587 32459 22593
rect 32766 22584 32772 22636
rect 32824 22624 32830 22636
rect 32861 22627 32919 22633
rect 32861 22624 32873 22627
rect 32824 22596 32873 22624
rect 32824 22584 32830 22596
rect 32861 22593 32873 22596
rect 32907 22593 32919 22627
rect 32861 22587 32919 22593
rect 32950 22584 32956 22636
rect 33008 22624 33014 22636
rect 33781 22627 33839 22633
rect 33008 22596 33053 22624
rect 33008 22584 33014 22596
rect 33781 22593 33793 22627
rect 33827 22624 33839 22627
rect 33870 22624 33876 22636
rect 33827 22596 33876 22624
rect 33827 22593 33839 22596
rect 33781 22587 33839 22593
rect 33870 22584 33876 22596
rect 33928 22584 33934 22636
rect 33137 22559 33195 22565
rect 33137 22525 33149 22559
rect 33183 22556 33195 22559
rect 33318 22556 33324 22568
rect 33183 22528 33324 22556
rect 33183 22525 33195 22528
rect 33137 22519 33195 22525
rect 33318 22516 33324 22528
rect 33376 22516 33382 22568
rect 31113 22451 31171 22457
rect 31772 22460 32352 22488
rect 31772 22432 31800 22460
rect 32766 22448 32772 22500
rect 32824 22488 32830 22500
rect 33597 22491 33655 22497
rect 33597 22488 33609 22491
rect 32824 22460 33609 22488
rect 32824 22448 32830 22460
rect 33597 22457 33609 22460
rect 33643 22457 33655 22491
rect 33597 22451 33655 22457
rect 30098 22420 30104 22432
rect 27586 22392 30104 22420
rect 30098 22380 30104 22392
rect 30156 22420 30162 22432
rect 30561 22423 30619 22429
rect 30561 22420 30573 22423
rect 30156 22392 30573 22420
rect 30156 22380 30162 22392
rect 30561 22389 30573 22392
rect 30607 22389 30619 22423
rect 30561 22383 30619 22389
rect 31754 22380 31760 22432
rect 31812 22380 31818 22432
rect 31846 22380 31852 22432
rect 31904 22420 31910 22432
rect 32125 22423 32183 22429
rect 32125 22420 32137 22423
rect 31904 22392 32137 22420
rect 31904 22380 31910 22392
rect 32125 22389 32137 22392
rect 32171 22389 32183 22423
rect 32125 22383 32183 22389
rect 32674 22380 32680 22432
rect 32732 22420 32738 22432
rect 32858 22420 32864 22432
rect 32732 22392 32864 22420
rect 32732 22380 32738 22392
rect 32858 22380 32864 22392
rect 32916 22380 32922 22432
rect 1104 22330 34868 22352
rect 1104 22278 6582 22330
rect 6634 22278 6646 22330
rect 6698 22278 6710 22330
rect 6762 22278 6774 22330
rect 6826 22278 6838 22330
rect 6890 22278 17846 22330
rect 17898 22278 17910 22330
rect 17962 22278 17974 22330
rect 18026 22278 18038 22330
rect 18090 22278 18102 22330
rect 18154 22278 29110 22330
rect 29162 22278 29174 22330
rect 29226 22278 29238 22330
rect 29290 22278 29302 22330
rect 29354 22278 29366 22330
rect 29418 22278 34868 22330
rect 1104 22256 34868 22278
rect 16758 22216 16764 22228
rect 16408 22188 16764 22216
rect 16408 22089 16436 22188
rect 16758 22176 16764 22188
rect 16816 22176 16822 22228
rect 17034 22176 17040 22228
rect 17092 22216 17098 22228
rect 17773 22219 17831 22225
rect 17773 22216 17785 22219
rect 17092 22188 17785 22216
rect 17092 22176 17098 22188
rect 17773 22185 17785 22188
rect 17819 22185 17831 22219
rect 19334 22216 19340 22228
rect 19295 22188 19340 22216
rect 17773 22179 17831 22185
rect 19334 22176 19340 22188
rect 19392 22176 19398 22228
rect 19426 22176 19432 22228
rect 19484 22216 19490 22228
rect 20349 22219 20407 22225
rect 20349 22216 20361 22219
rect 19484 22188 20361 22216
rect 19484 22176 19490 22188
rect 20349 22185 20361 22188
rect 20395 22185 20407 22219
rect 20349 22179 20407 22185
rect 20993 22219 21051 22225
rect 20993 22185 21005 22219
rect 21039 22216 21051 22219
rect 21082 22216 21088 22228
rect 21039 22188 21088 22216
rect 21039 22185 21051 22188
rect 20993 22179 21051 22185
rect 21082 22176 21088 22188
rect 21140 22176 21146 22228
rect 21358 22176 21364 22228
rect 21416 22216 21422 22228
rect 22189 22219 22247 22225
rect 22189 22216 22201 22219
rect 21416 22188 22201 22216
rect 21416 22176 21422 22188
rect 22189 22185 22201 22188
rect 22235 22185 22247 22219
rect 22922 22216 22928 22228
rect 22883 22188 22928 22216
rect 22189 22179 22247 22185
rect 22922 22176 22928 22188
rect 22980 22176 22986 22228
rect 23106 22176 23112 22228
rect 23164 22216 23170 22228
rect 27982 22216 27988 22228
rect 23164 22188 27988 22216
rect 23164 22176 23170 22188
rect 27982 22176 27988 22188
rect 28040 22176 28046 22228
rect 28258 22176 28264 22228
rect 28316 22216 28322 22228
rect 29733 22219 29791 22225
rect 29733 22216 29745 22219
rect 28316 22188 28994 22216
rect 28316 22176 28322 22188
rect 19150 22108 19156 22160
rect 19208 22148 19214 22160
rect 20533 22151 20591 22157
rect 20533 22148 20545 22151
rect 19208 22120 20545 22148
rect 19208 22108 19214 22120
rect 20533 22117 20545 22120
rect 20579 22117 20591 22151
rect 20533 22111 20591 22117
rect 23290 22108 23296 22160
rect 23348 22108 23354 22160
rect 25866 22148 25872 22160
rect 24964 22120 25872 22148
rect 16393 22083 16451 22089
rect 16393 22049 16405 22083
rect 16439 22049 16451 22083
rect 16393 22043 16451 22049
rect 18233 22083 18291 22089
rect 18233 22049 18245 22083
rect 18279 22080 18291 22083
rect 19334 22080 19340 22092
rect 18279 22052 19340 22080
rect 18279 22049 18291 22052
rect 18233 22043 18291 22049
rect 19334 22040 19340 22052
rect 19392 22040 19398 22092
rect 19610 22040 19616 22092
rect 19668 22080 19674 22092
rect 21450 22080 21456 22092
rect 19668 22052 20300 22080
rect 19668 22040 19674 22052
rect 16022 21972 16028 22024
rect 16080 22012 16086 22024
rect 16482 22012 16488 22024
rect 16080 21984 16488 22012
rect 16080 21972 16086 21984
rect 16482 21972 16488 21984
rect 16540 21972 16546 22024
rect 17402 21972 17408 22024
rect 17460 22012 17466 22024
rect 18417 22015 18475 22021
rect 18417 22012 18429 22015
rect 17460 21984 18429 22012
rect 17460 21972 17466 21984
rect 18417 21981 18429 21984
rect 18463 21981 18475 22015
rect 19426 22012 19432 22024
rect 19387 21984 19432 22012
rect 18417 21975 18475 21981
rect 19426 21972 19432 21984
rect 19484 21972 19490 22024
rect 19518 21972 19524 22024
rect 19576 22012 19582 22024
rect 19576 21984 19621 22012
rect 19576 21972 19582 21984
rect 16660 21947 16718 21953
rect 16660 21913 16672 21947
rect 16706 21944 16718 21947
rect 17034 21944 17040 21956
rect 16706 21916 17040 21944
rect 16706 21913 16718 21916
rect 16660 21907 16718 21913
rect 17034 21904 17040 21916
rect 17092 21904 17098 21956
rect 19245 21947 19303 21953
rect 19245 21913 19257 21947
rect 19291 21913 19303 21947
rect 19245 21907 19303 21913
rect 18506 21836 18512 21888
rect 18564 21876 18570 21888
rect 18601 21879 18659 21885
rect 18601 21876 18613 21879
rect 18564 21848 18613 21876
rect 18564 21836 18570 21848
rect 18601 21845 18613 21848
rect 18647 21845 18659 21879
rect 19260 21876 19288 21907
rect 19334 21904 19340 21956
rect 19392 21944 19398 21956
rect 20165 21947 20223 21953
rect 20165 21944 20177 21947
rect 19392 21916 20177 21944
rect 19392 21904 19398 21916
rect 20165 21913 20177 21916
rect 20211 21913 20223 21947
rect 20272 21944 20300 22052
rect 21008 22052 21456 22080
rect 21008 22021 21036 22052
rect 21450 22040 21456 22052
rect 21508 22040 21514 22092
rect 22738 22080 22744 22092
rect 21928 22052 22744 22080
rect 20993 22015 21051 22021
rect 20993 21981 21005 22015
rect 21039 21981 21051 22015
rect 20993 21975 21051 21981
rect 21269 22015 21327 22021
rect 21269 21981 21281 22015
rect 21315 22012 21327 22015
rect 21358 22012 21364 22024
rect 21315 21984 21364 22012
rect 21315 21981 21327 21984
rect 21269 21975 21327 21981
rect 21358 21972 21364 21984
rect 21416 21972 21422 22024
rect 21729 22015 21787 22021
rect 21729 21981 21741 22015
rect 21775 22012 21787 22015
rect 21818 22012 21824 22024
rect 21775 21984 21824 22012
rect 21775 21981 21787 21984
rect 21729 21975 21787 21981
rect 21818 21972 21824 21984
rect 21876 21972 21882 22024
rect 21928 22021 21956 22052
rect 22738 22040 22744 22052
rect 22796 22040 22802 22092
rect 23308 22080 23336 22108
rect 24964 22092 24992 22120
rect 25866 22108 25872 22120
rect 25924 22108 25930 22160
rect 27246 22108 27252 22160
rect 27304 22148 27310 22160
rect 27433 22151 27491 22157
rect 27433 22148 27445 22151
rect 27304 22120 27445 22148
rect 27304 22108 27310 22120
rect 27433 22117 27445 22120
rect 27479 22148 27491 22151
rect 28966 22148 28994 22188
rect 29488 22188 29745 22216
rect 29178 22148 29184 22160
rect 27479 22120 28580 22148
rect 28966 22120 29184 22148
rect 27479 22117 27491 22120
rect 27433 22111 27491 22117
rect 23308 22052 23612 22080
rect 21913 22015 21971 22021
rect 21913 21981 21925 22015
rect 21959 21981 21971 22015
rect 21913 21975 21971 21981
rect 22002 21972 22008 22024
rect 22060 22012 22066 22024
rect 22060 21984 22105 22012
rect 22060 21972 22066 21984
rect 22186 21972 22192 22024
rect 22244 22012 22250 22024
rect 22281 22015 22339 22021
rect 22281 22012 22293 22015
rect 22244 21984 22293 22012
rect 22244 21972 22250 21984
rect 22281 21981 22293 21984
rect 22327 21981 22339 22015
rect 23198 22012 23204 22024
rect 23159 21984 23204 22012
rect 22281 21975 22339 21981
rect 23198 21972 23204 21984
rect 23256 21972 23262 22024
rect 23293 22015 23351 22021
rect 23293 21981 23305 22015
rect 23339 21981 23351 22015
rect 23293 21975 23351 21981
rect 20365 21947 20423 21953
rect 20365 21944 20377 21947
rect 20272 21916 20377 21944
rect 20165 21907 20223 21913
rect 20365 21913 20377 21916
rect 20411 21913 20423 21947
rect 20365 21907 20423 21913
rect 21177 21947 21235 21953
rect 21177 21913 21189 21947
rect 21223 21944 21235 21947
rect 23014 21944 23020 21956
rect 21223 21916 23020 21944
rect 21223 21913 21235 21916
rect 21177 21907 21235 21913
rect 23014 21904 23020 21916
rect 23072 21904 23078 21956
rect 23308 21944 23336 21975
rect 23382 21972 23388 22024
rect 23440 22012 23446 22024
rect 23584 22021 23612 22052
rect 23934 22040 23940 22092
rect 23992 22080 23998 22092
rect 24489 22083 24547 22089
rect 24489 22080 24501 22083
rect 23992 22052 24501 22080
rect 23992 22040 23998 22052
rect 24489 22049 24501 22052
rect 24535 22080 24547 22083
rect 24946 22080 24952 22092
rect 24535 22052 24808 22080
rect 24907 22052 24952 22080
rect 24535 22049 24547 22052
rect 24489 22043 24547 22049
rect 23569 22015 23627 22021
rect 23440 21984 23485 22012
rect 23440 21972 23446 21984
rect 23569 21981 23581 22015
rect 23615 21981 23627 22015
rect 23569 21975 23627 21981
rect 24118 21972 24124 22024
rect 24176 22012 24182 22024
rect 24302 22012 24308 22024
rect 24176 21984 24308 22012
rect 24176 21972 24182 21984
rect 24302 21972 24308 21984
rect 24360 21972 24366 22024
rect 24578 22012 24584 22024
rect 24539 21984 24584 22012
rect 24578 21972 24584 21984
rect 24636 21972 24642 22024
rect 24780 22012 24808 22052
rect 24946 22040 24952 22052
rect 25004 22040 25010 22092
rect 25590 22080 25596 22092
rect 25424 22052 25596 22080
rect 25314 22012 25320 22024
rect 24780 21984 25320 22012
rect 25314 21972 25320 21984
rect 25372 21972 25378 22024
rect 25424 22021 25452 22052
rect 25590 22040 25596 22052
rect 25648 22040 25654 22092
rect 27890 22080 27896 22092
rect 27851 22052 27896 22080
rect 27890 22040 27896 22052
rect 27948 22040 27954 22092
rect 28353 22083 28411 22089
rect 28353 22080 28365 22083
rect 28000 22052 28365 22080
rect 25409 22015 25467 22021
rect 25409 21981 25421 22015
rect 25455 21981 25467 22015
rect 25409 21975 25467 21981
rect 25498 21972 25504 22024
rect 25556 22012 25562 22024
rect 26050 22012 26056 22024
rect 25556 21984 26056 22012
rect 25556 21972 25562 21984
rect 26050 21972 26056 21984
rect 26108 21972 26114 22024
rect 26326 22021 26332 22024
rect 26320 22012 26332 22021
rect 26287 21984 26332 22012
rect 26320 21975 26332 21984
rect 26326 21972 26332 21975
rect 26384 21972 26390 22024
rect 28000 22012 28028 22052
rect 28353 22049 28365 22052
rect 28399 22049 28411 22083
rect 28552 22080 28580 22120
rect 29178 22108 29184 22120
rect 29236 22108 29242 22160
rect 28353 22043 28411 22049
rect 28460 22052 28580 22080
rect 27816 21984 28028 22012
rect 28060 22015 28118 22021
rect 25038 21944 25044 21956
rect 23308 21916 25044 21944
rect 25038 21904 25044 21916
rect 25096 21904 25102 21956
rect 27154 21944 27160 21956
rect 25424 21916 27160 21944
rect 19518 21876 19524 21888
rect 19260 21848 19524 21876
rect 18601 21839 18659 21845
rect 19518 21836 19524 21848
rect 19576 21836 19582 21888
rect 19702 21876 19708 21888
rect 19663 21848 19708 21876
rect 19702 21836 19708 21848
rect 19760 21836 19766 21888
rect 24394 21836 24400 21888
rect 24452 21876 24458 21888
rect 25424 21876 25452 21916
rect 27154 21904 27160 21916
rect 27212 21944 27218 21956
rect 27816 21944 27844 21984
rect 28060 21981 28072 22015
rect 28106 22012 28118 22015
rect 28106 21981 28120 22012
rect 28060 21975 28120 21981
rect 27212 21916 27844 21944
rect 27212 21904 27218 21916
rect 27890 21904 27896 21956
rect 27948 21944 27954 21956
rect 28092 21944 28120 21975
rect 28166 21972 28172 22024
rect 28224 22012 28230 22024
rect 28460 22021 28488 22052
rect 28445 22015 28503 22021
rect 28224 21984 28269 22012
rect 28224 21972 28230 21984
rect 28445 21981 28457 22015
rect 28491 21981 28503 22015
rect 28445 21975 28503 21981
rect 29488 22012 29516 22188
rect 29733 22185 29745 22188
rect 29779 22216 29791 22219
rect 29914 22216 29920 22228
rect 29779 22188 29920 22216
rect 29779 22185 29791 22188
rect 29733 22179 29791 22185
rect 29914 22176 29920 22188
rect 29972 22176 29978 22228
rect 31662 22216 31668 22228
rect 31128 22188 31668 22216
rect 31128 22157 31156 22188
rect 31662 22176 31668 22188
rect 31720 22176 31726 22228
rect 32030 22176 32036 22228
rect 32088 22176 32094 22228
rect 32950 22176 32956 22228
rect 33008 22216 33014 22228
rect 33318 22216 33324 22228
rect 33008 22188 33324 22216
rect 33008 22176 33014 22188
rect 33318 22176 33324 22188
rect 33376 22176 33382 22228
rect 31113 22151 31171 22157
rect 29932 22120 30696 22148
rect 29932 22092 29960 22120
rect 29914 22040 29920 22092
rect 29972 22040 29978 22092
rect 30006 22040 30012 22092
rect 30064 22080 30070 22092
rect 30449 22088 30507 22089
rect 30208 22083 30507 22088
rect 30208 22080 30461 22083
rect 30064 22060 30461 22080
rect 30064 22052 30236 22060
rect 30064 22040 30070 22052
rect 30449 22049 30461 22060
rect 30495 22049 30507 22083
rect 30449 22043 30507 22049
rect 30668 22021 30696 22120
rect 31113 22117 31125 22151
rect 31159 22117 31171 22151
rect 31113 22111 31171 22117
rect 31386 22108 31392 22160
rect 31444 22148 31450 22160
rect 31444 22120 31892 22148
rect 31444 22108 31450 22120
rect 31662 22080 31668 22092
rect 30944 22052 31668 22080
rect 30561 22015 30619 22021
rect 30561 22012 30573 22015
rect 29488 21984 30573 22012
rect 27948 21916 28120 21944
rect 27948 21904 27954 21916
rect 28258 21904 28264 21956
rect 28316 21944 28322 21956
rect 29270 21944 29276 21956
rect 28316 21916 29276 21944
rect 28316 21904 28322 21916
rect 29270 21904 29276 21916
rect 29328 21904 29334 21956
rect 24452 21848 25452 21876
rect 25501 21879 25559 21885
rect 24452 21836 24458 21848
rect 25501 21845 25513 21879
rect 25547 21876 25559 21879
rect 27246 21876 27252 21888
rect 25547 21848 27252 21876
rect 25547 21845 25559 21848
rect 25501 21839 25559 21845
rect 27246 21836 27252 21848
rect 27304 21836 27310 21888
rect 28074 21836 28080 21888
rect 28132 21876 28138 21888
rect 29488 21876 29516 21984
rect 30561 21981 30573 21984
rect 30607 21981 30619 22015
rect 30561 21975 30619 21981
rect 30653 22015 30711 22021
rect 30653 21981 30665 22015
rect 30699 21981 30711 22015
rect 30653 21975 30711 21981
rect 29549 21947 29607 21953
rect 29549 21913 29561 21947
rect 29595 21944 29607 21947
rect 30282 21944 30288 21956
rect 29595 21916 30288 21944
rect 29595 21913 29607 21916
rect 29549 21907 29607 21913
rect 30282 21904 30288 21916
rect 30340 21944 30346 21956
rect 30377 21947 30435 21953
rect 30377 21944 30389 21947
rect 30340 21916 30389 21944
rect 30340 21904 30346 21916
rect 30377 21913 30389 21916
rect 30423 21913 30435 21947
rect 30944 21944 30972 22052
rect 31662 22040 31668 22052
rect 31720 22040 31726 22092
rect 31018 21972 31024 22024
rect 31076 22012 31082 22024
rect 31389 22015 31447 22021
rect 31076 21984 31248 22012
rect 31076 21972 31082 21984
rect 31113 21947 31171 21953
rect 31113 21944 31125 21947
rect 30944 21916 31125 21944
rect 30377 21907 30435 21913
rect 31113 21913 31125 21916
rect 31159 21913 31171 21947
rect 31220 21944 31248 21984
rect 31389 21981 31401 22015
rect 31435 22012 31447 22015
rect 31754 22012 31760 22024
rect 31435 21984 31760 22012
rect 31435 21981 31447 21984
rect 31389 21975 31447 21981
rect 31754 21972 31760 21984
rect 31812 21972 31818 22024
rect 31864 22021 31892 22120
rect 32048 22080 32076 22176
rect 32125 22083 32183 22089
rect 32125 22080 32137 22083
rect 32048 22052 32137 22080
rect 32125 22049 32137 22052
rect 32171 22049 32183 22083
rect 32858 22080 32864 22092
rect 32819 22052 32864 22080
rect 32125 22043 32183 22049
rect 32858 22040 32864 22052
rect 32916 22040 32922 22092
rect 33686 22080 33692 22092
rect 33647 22052 33692 22080
rect 33686 22040 33692 22052
rect 33744 22040 33750 22092
rect 31849 22015 31907 22021
rect 31849 21981 31861 22015
rect 31895 21981 31907 22015
rect 31849 21975 31907 21981
rect 31941 22015 31999 22021
rect 31941 21981 31953 22015
rect 31987 21981 31999 22015
rect 31941 21975 31999 21981
rect 31956 21944 31984 21975
rect 32398 21972 32404 22024
rect 32456 22012 32462 22024
rect 32677 22015 32735 22021
rect 32677 22012 32689 22015
rect 32456 21984 32689 22012
rect 32456 21972 32462 21984
rect 32677 21981 32689 21984
rect 32723 21981 32735 22015
rect 33594 22012 33600 22024
rect 33555 21984 33600 22012
rect 32677 21975 32735 21981
rect 33594 21972 33600 21984
rect 33652 21972 33658 22024
rect 31220 21916 31984 21944
rect 31113 21907 31171 21913
rect 32858 21904 32864 21956
rect 32916 21944 32922 21956
rect 33318 21944 33324 21956
rect 32916 21916 33324 21944
rect 32916 21904 32922 21916
rect 33318 21904 33324 21916
rect 33376 21904 33382 21956
rect 28132 21848 29516 21876
rect 28132 21836 28138 21848
rect 29638 21836 29644 21888
rect 29696 21876 29702 21888
rect 29749 21879 29807 21885
rect 29749 21876 29761 21879
rect 29696 21848 29761 21876
rect 29696 21836 29702 21848
rect 29749 21845 29761 21848
rect 29795 21845 29807 21879
rect 29749 21839 29807 21845
rect 29917 21879 29975 21885
rect 29917 21845 29929 21879
rect 29963 21876 29975 21879
rect 30466 21876 30472 21888
rect 29963 21848 30472 21876
rect 29963 21845 29975 21848
rect 29917 21839 29975 21845
rect 30466 21836 30472 21848
rect 30524 21836 30530 21888
rect 30926 21836 30932 21888
rect 30984 21876 30990 21888
rect 31297 21879 31355 21885
rect 31297 21876 31309 21879
rect 30984 21848 31309 21876
rect 30984 21836 30990 21848
rect 31297 21845 31309 21848
rect 31343 21845 31355 21879
rect 31297 21839 31355 21845
rect 31570 21836 31576 21888
rect 31628 21876 31634 21888
rect 32125 21879 32183 21885
rect 32125 21876 32137 21879
rect 31628 21848 32137 21876
rect 31628 21836 31634 21848
rect 32125 21845 32137 21848
rect 32171 21845 32183 21879
rect 32125 21839 32183 21845
rect 1104 21786 34868 21808
rect 1104 21734 12214 21786
rect 12266 21734 12278 21786
rect 12330 21734 12342 21786
rect 12394 21734 12406 21786
rect 12458 21734 12470 21786
rect 12522 21734 23478 21786
rect 23530 21734 23542 21786
rect 23594 21734 23606 21786
rect 23658 21734 23670 21786
rect 23722 21734 23734 21786
rect 23786 21734 34868 21786
rect 1104 21712 34868 21734
rect 19518 21672 19524 21684
rect 17972 21644 19524 21672
rect 16574 21496 16580 21548
rect 16632 21536 16638 21548
rect 17402 21536 17408 21548
rect 16632 21508 17408 21536
rect 16632 21496 16638 21508
rect 17402 21496 17408 21508
rect 17460 21496 17466 21548
rect 17221 21471 17279 21477
rect 17221 21437 17233 21471
rect 17267 21468 17279 21471
rect 17972 21468 18000 21644
rect 19518 21632 19524 21644
rect 19576 21672 19582 21684
rect 19794 21672 19800 21684
rect 19576 21644 19800 21672
rect 19576 21632 19582 21644
rect 19794 21632 19800 21644
rect 19852 21672 19858 21684
rect 21269 21675 21327 21681
rect 21269 21672 21281 21675
rect 19852 21644 21281 21672
rect 19852 21632 19858 21644
rect 21269 21641 21281 21644
rect 21315 21641 21327 21675
rect 21269 21635 21327 21641
rect 23017 21675 23075 21681
rect 23017 21641 23029 21675
rect 23063 21672 23075 21675
rect 24394 21672 24400 21684
rect 23063 21644 24400 21672
rect 23063 21641 23075 21644
rect 23017 21635 23075 21641
rect 24394 21632 24400 21644
rect 24452 21632 24458 21684
rect 24762 21632 24768 21684
rect 24820 21672 24826 21684
rect 24820 21644 25176 21672
rect 24820 21632 24826 21644
rect 21082 21604 21088 21616
rect 18064 21576 21088 21604
rect 18064 21477 18092 21576
rect 18322 21545 18328 21548
rect 18316 21499 18328 21545
rect 18380 21536 18386 21548
rect 18380 21508 18416 21536
rect 18322 21496 18328 21499
rect 18380 21496 18386 21508
rect 19904 21477 19932 21576
rect 21082 21564 21088 21576
rect 21140 21564 21146 21616
rect 21358 21564 21364 21616
rect 21416 21604 21422 21616
rect 22649 21607 22707 21613
rect 21416 21576 22499 21604
rect 21416 21564 21422 21576
rect 19978 21496 19984 21548
rect 20036 21536 20042 21548
rect 20145 21539 20203 21545
rect 20145 21536 20157 21539
rect 20036 21508 20157 21536
rect 20036 21496 20042 21508
rect 20145 21505 20157 21508
rect 20191 21505 20203 21539
rect 21818 21536 21824 21548
rect 21779 21508 21824 21536
rect 20145 21499 20203 21505
rect 21818 21496 21824 21508
rect 21876 21496 21882 21548
rect 22005 21539 22063 21545
rect 22005 21505 22017 21539
rect 22051 21536 22063 21539
rect 22370 21536 22376 21548
rect 22051 21508 22376 21536
rect 22051 21505 22063 21508
rect 22005 21499 22063 21505
rect 22370 21496 22376 21508
rect 22428 21496 22434 21548
rect 22471 21536 22499 21576
rect 22649 21573 22661 21607
rect 22695 21604 22707 21607
rect 22695 21576 24992 21604
rect 22695 21573 22707 21576
rect 22649 21567 22707 21573
rect 22830 21536 22836 21548
rect 22471 21508 22836 21536
rect 22830 21496 22836 21508
rect 22888 21496 22894 21548
rect 23106 21536 23112 21548
rect 23067 21508 23112 21536
rect 23106 21496 23112 21508
rect 23164 21496 23170 21548
rect 23566 21536 23572 21548
rect 23527 21508 23572 21536
rect 23566 21496 23572 21508
rect 23624 21496 23630 21548
rect 23753 21539 23811 21545
rect 23753 21505 23765 21539
rect 23799 21536 23811 21539
rect 23934 21536 23940 21548
rect 23799 21508 23940 21536
rect 23799 21505 23811 21508
rect 23753 21499 23811 21505
rect 17267 21440 18000 21468
rect 18049 21471 18107 21477
rect 17267 21437 17279 21440
rect 17221 21431 17279 21437
rect 18049 21437 18061 21471
rect 18095 21437 18107 21471
rect 18049 21431 18107 21437
rect 19889 21471 19947 21477
rect 19889 21437 19901 21471
rect 19935 21437 19947 21471
rect 19889 21431 19947 21437
rect 16942 21360 16948 21412
rect 17000 21400 17006 21412
rect 18064 21400 18092 21431
rect 21634 21428 21640 21480
rect 21692 21468 21698 21480
rect 23768 21468 23796 21499
rect 23934 21496 23940 21508
rect 23992 21496 23998 21548
rect 24029 21539 24087 21545
rect 24029 21505 24041 21539
rect 24075 21536 24087 21539
rect 24302 21536 24308 21548
rect 24075 21508 24308 21536
rect 24075 21505 24087 21508
rect 24029 21499 24087 21505
rect 24302 21496 24308 21508
rect 24360 21496 24366 21548
rect 24486 21496 24492 21548
rect 24544 21536 24550 21548
rect 24964 21545 24992 21576
rect 25148 21545 25176 21644
rect 27246 21632 27252 21684
rect 27304 21672 27310 21684
rect 27304 21644 27660 21672
rect 27304 21632 27310 21644
rect 27154 21564 27160 21616
rect 27212 21604 27218 21616
rect 27525 21607 27583 21613
rect 27525 21604 27537 21607
rect 27212 21576 27537 21604
rect 27212 21564 27218 21576
rect 27525 21573 27537 21576
rect 27571 21573 27583 21607
rect 27632 21604 27660 21644
rect 27706 21632 27712 21684
rect 27764 21672 27770 21684
rect 27893 21675 27951 21681
rect 27893 21672 27905 21675
rect 27764 21644 27905 21672
rect 27764 21632 27770 21644
rect 27893 21641 27905 21644
rect 27939 21641 27951 21675
rect 27893 21635 27951 21641
rect 29638 21632 29644 21684
rect 29696 21672 29702 21684
rect 30006 21672 30012 21684
rect 29696 21644 30012 21672
rect 29696 21632 29702 21644
rect 30006 21632 30012 21644
rect 30064 21632 30070 21684
rect 31386 21632 31392 21684
rect 31444 21672 31450 21684
rect 31570 21672 31576 21684
rect 31444 21644 31576 21672
rect 31444 21632 31450 21644
rect 31570 21632 31576 21644
rect 31628 21632 31634 21684
rect 32122 21632 32128 21684
rect 32180 21672 32186 21684
rect 32309 21675 32367 21681
rect 32309 21672 32321 21675
rect 32180 21644 32321 21672
rect 32180 21632 32186 21644
rect 32309 21641 32321 21644
rect 32355 21641 32367 21675
rect 32309 21635 32367 21641
rect 32490 21632 32496 21684
rect 32548 21672 32554 21684
rect 33413 21675 33471 21681
rect 33413 21672 33425 21675
rect 32548 21644 33425 21672
rect 32548 21632 32554 21644
rect 33413 21641 33425 21644
rect 33459 21641 33471 21675
rect 33413 21635 33471 21641
rect 33962 21632 33968 21684
rect 34020 21672 34026 21684
rect 34057 21675 34115 21681
rect 34057 21672 34069 21675
rect 34020 21644 34069 21672
rect 34020 21632 34026 21644
rect 34057 21641 34069 21644
rect 34103 21641 34115 21675
rect 34057 21635 34115 21641
rect 31113 21607 31171 21613
rect 27632 21576 27752 21604
rect 27525 21567 27583 21573
rect 24765 21539 24823 21545
rect 24765 21536 24777 21539
rect 24544 21508 24777 21536
rect 24544 21496 24550 21508
rect 24765 21505 24777 21508
rect 24811 21505 24823 21539
rect 24765 21499 24823 21505
rect 24857 21539 24915 21545
rect 24857 21505 24869 21539
rect 24903 21505 24915 21539
rect 24857 21499 24915 21505
rect 24949 21539 25007 21545
rect 24949 21505 24961 21539
rect 24995 21505 25007 21539
rect 24949 21499 25007 21505
rect 25133 21539 25191 21545
rect 25133 21505 25145 21539
rect 25179 21505 25191 21539
rect 25774 21536 25780 21548
rect 25735 21508 25780 21536
rect 25133 21499 25191 21505
rect 24578 21468 24584 21480
rect 21692 21440 23796 21468
rect 23952 21440 24584 21468
rect 21692 21428 21698 21440
rect 17000 21372 18092 21400
rect 22189 21403 22247 21409
rect 17000 21360 17006 21372
rect 22189 21369 22201 21403
rect 22235 21400 22247 21403
rect 23382 21400 23388 21412
rect 22235 21372 23388 21400
rect 22235 21369 22247 21372
rect 22189 21363 22247 21369
rect 23382 21360 23388 21372
rect 23440 21360 23446 21412
rect 17218 21292 17224 21344
rect 17276 21332 17282 21344
rect 17589 21335 17647 21341
rect 17589 21332 17601 21335
rect 17276 21304 17601 21332
rect 17276 21292 17282 21304
rect 17589 21301 17601 21304
rect 17635 21301 17647 21335
rect 17589 21295 17647 21301
rect 18230 21292 18236 21344
rect 18288 21332 18294 21344
rect 19426 21332 19432 21344
rect 18288 21304 19432 21332
rect 18288 21292 18294 21304
rect 19426 21292 19432 21304
rect 19484 21292 19490 21344
rect 23952 21341 23980 21440
rect 24578 21428 24584 21440
rect 24636 21428 24642 21480
rect 24872 21468 24900 21499
rect 25774 21496 25780 21508
rect 25832 21536 25838 21548
rect 25832 21508 27292 21536
rect 25832 21496 25838 21508
rect 24872 21440 25176 21468
rect 25148 21412 25176 21440
rect 25314 21428 25320 21480
rect 25372 21468 25378 21480
rect 25685 21471 25743 21477
rect 25685 21468 25697 21471
rect 25372 21440 25697 21468
rect 25372 21428 25378 21440
rect 25685 21437 25697 21440
rect 25731 21437 25743 21471
rect 25685 21431 25743 21437
rect 25958 21428 25964 21480
rect 26016 21468 26022 21480
rect 26145 21471 26203 21477
rect 26145 21468 26157 21471
rect 26016 21440 26157 21468
rect 26016 21428 26022 21440
rect 26145 21437 26157 21440
rect 26191 21437 26203 21471
rect 27264 21468 27292 21508
rect 27338 21496 27344 21548
rect 27396 21536 27402 21548
rect 27724 21545 27752 21576
rect 29472 21576 30236 21604
rect 27617 21539 27675 21545
rect 27396 21508 27441 21536
rect 27396 21496 27402 21508
rect 27617 21505 27629 21539
rect 27663 21505 27675 21539
rect 27724 21539 27791 21545
rect 27724 21508 27745 21539
rect 27617 21499 27675 21505
rect 27733 21505 27745 21508
rect 27779 21505 27791 21539
rect 27733 21499 27791 21505
rect 27522 21468 27528 21480
rect 27264 21440 27528 21468
rect 26145 21431 26203 21437
rect 27522 21428 27528 21440
rect 27580 21468 27586 21480
rect 27632 21468 27660 21499
rect 28166 21496 28172 21548
rect 28224 21536 28230 21548
rect 29472 21545 29500 21576
rect 30208 21545 30236 21576
rect 31113 21573 31125 21607
rect 31159 21604 31171 21607
rect 33226 21604 33232 21616
rect 31159 21576 33232 21604
rect 31159 21573 31171 21576
rect 31113 21567 31171 21573
rect 33226 21564 33232 21576
rect 33284 21564 33290 21616
rect 28445 21539 28503 21545
rect 28445 21536 28457 21539
rect 28224 21508 28457 21536
rect 28224 21496 28230 21508
rect 28445 21505 28457 21508
rect 28491 21505 28503 21539
rect 28445 21499 28503 21505
rect 29457 21539 29515 21545
rect 29457 21505 29469 21539
rect 29503 21505 29515 21539
rect 29457 21499 29515 21505
rect 30101 21539 30159 21545
rect 30101 21505 30113 21539
rect 30147 21505 30159 21539
rect 30101 21499 30159 21505
rect 30193 21539 30251 21545
rect 30193 21505 30205 21539
rect 30239 21536 30251 21539
rect 30466 21536 30472 21548
rect 30239 21508 30472 21536
rect 30239 21505 30251 21508
rect 30193 21499 30251 21505
rect 27580 21440 27660 21468
rect 29273 21471 29331 21477
rect 27580 21428 27586 21440
rect 29273 21437 29285 21471
rect 29319 21468 29331 21471
rect 30116 21468 30144 21499
rect 30466 21496 30472 21508
rect 30524 21496 30530 21548
rect 30650 21496 30656 21548
rect 30708 21496 30714 21548
rect 30837 21539 30895 21545
rect 30837 21505 30849 21539
rect 30883 21536 30895 21539
rect 31018 21536 31024 21548
rect 30883 21508 31024 21536
rect 30883 21505 30895 21508
rect 30837 21499 30895 21505
rect 31018 21496 31024 21508
rect 31076 21496 31082 21548
rect 32217 21539 32275 21545
rect 32217 21505 32229 21539
rect 32263 21505 32275 21539
rect 32217 21499 32275 21505
rect 33321 21539 33379 21545
rect 33321 21505 33333 21539
rect 33367 21536 33379 21539
rect 33778 21536 33784 21548
rect 33367 21508 33784 21536
rect 33367 21505 33379 21508
rect 33321 21499 33379 21505
rect 29319 21440 30144 21468
rect 30377 21471 30435 21477
rect 29319 21437 29331 21440
rect 29273 21431 29331 21437
rect 25130 21360 25136 21412
rect 25188 21360 25194 21412
rect 27062 21360 27068 21412
rect 27120 21400 27126 21412
rect 29288 21400 29316 21431
rect 27120 21372 29316 21400
rect 27120 21360 27126 21372
rect 23937 21335 23995 21341
rect 23937 21301 23949 21335
rect 23983 21301 23995 21335
rect 23937 21295 23995 21301
rect 24489 21335 24547 21341
rect 24489 21301 24501 21335
rect 24535 21332 24547 21335
rect 25682 21332 25688 21344
rect 24535 21304 25688 21332
rect 24535 21301 24547 21304
rect 24489 21295 24547 21301
rect 25682 21292 25688 21304
rect 25740 21292 25746 21344
rect 26326 21292 26332 21344
rect 26384 21332 26390 21344
rect 28537 21335 28595 21341
rect 28537 21332 28549 21335
rect 26384 21304 28549 21332
rect 26384 21292 26390 21304
rect 28537 21301 28549 21304
rect 28583 21301 28595 21335
rect 28537 21295 28595 21301
rect 29546 21292 29552 21344
rect 29604 21332 29610 21344
rect 29641 21335 29699 21341
rect 29641 21332 29653 21335
rect 29604 21304 29653 21332
rect 29604 21292 29610 21304
rect 29641 21301 29653 21304
rect 29687 21301 29699 21335
rect 29840 21332 29868 21440
rect 30377 21437 30389 21471
rect 30423 21468 30435 21471
rect 30423 21440 30512 21468
rect 30423 21437 30435 21440
rect 30377 21431 30435 21437
rect 30484 21412 30512 21440
rect 29914 21360 29920 21412
rect 29972 21400 29978 21412
rect 30285 21403 30343 21409
rect 30285 21400 30297 21403
rect 29972 21372 30297 21400
rect 29972 21360 29978 21372
rect 30285 21369 30297 21372
rect 30331 21369 30343 21403
rect 30285 21363 30343 21369
rect 30466 21360 30472 21412
rect 30524 21360 30530 21412
rect 30668 21400 30696 21496
rect 30837 21403 30895 21409
rect 30837 21400 30849 21403
rect 30668 21372 30849 21400
rect 30837 21369 30849 21372
rect 30883 21369 30895 21403
rect 30837 21363 30895 21369
rect 30929 21403 30987 21409
rect 30929 21369 30941 21403
rect 30975 21400 30987 21403
rect 31846 21400 31852 21412
rect 30975 21372 31852 21400
rect 30975 21369 30987 21372
rect 30929 21363 30987 21369
rect 31846 21360 31852 21372
rect 31904 21360 31910 21412
rect 30650 21332 30656 21344
rect 29840 21304 30656 21332
rect 29641 21295 29699 21301
rect 30650 21292 30656 21304
rect 30708 21292 30714 21344
rect 31570 21292 31576 21344
rect 31628 21332 31634 21344
rect 32232 21332 32260 21499
rect 33778 21496 33784 21508
rect 33836 21496 33842 21548
rect 33870 21496 33876 21548
rect 33928 21536 33934 21548
rect 33965 21539 34023 21545
rect 33965 21536 33977 21539
rect 33928 21508 33977 21536
rect 33928 21496 33934 21508
rect 33965 21505 33977 21508
rect 34011 21505 34023 21539
rect 33965 21499 34023 21505
rect 31628 21304 32260 21332
rect 31628 21292 31634 21304
rect 1104 21242 34868 21264
rect 1104 21190 6582 21242
rect 6634 21190 6646 21242
rect 6698 21190 6710 21242
rect 6762 21190 6774 21242
rect 6826 21190 6838 21242
rect 6890 21190 17846 21242
rect 17898 21190 17910 21242
rect 17962 21190 17974 21242
rect 18026 21190 18038 21242
rect 18090 21190 18102 21242
rect 18154 21190 29110 21242
rect 29162 21190 29174 21242
rect 29226 21190 29238 21242
rect 29290 21190 29302 21242
rect 29354 21190 29366 21242
rect 29418 21190 34868 21242
rect 1104 21168 34868 21190
rect 17034 21128 17040 21140
rect 16995 21100 17040 21128
rect 17034 21088 17040 21100
rect 17092 21088 17098 21140
rect 17681 21131 17739 21137
rect 17681 21097 17693 21131
rect 17727 21128 17739 21131
rect 19978 21128 19984 21140
rect 17727 21100 19984 21128
rect 17727 21097 17739 21100
rect 17681 21091 17739 21097
rect 19978 21088 19984 21100
rect 20036 21088 20042 21140
rect 20530 21128 20536 21140
rect 20491 21100 20536 21128
rect 20530 21088 20536 21100
rect 20588 21088 20594 21140
rect 22370 21088 22376 21140
rect 22428 21128 22434 21140
rect 22465 21131 22523 21137
rect 22465 21128 22477 21131
rect 22428 21100 22477 21128
rect 22428 21088 22434 21100
rect 22465 21097 22477 21100
rect 22511 21128 22523 21131
rect 22738 21128 22744 21140
rect 22511 21100 22744 21128
rect 22511 21097 22523 21100
rect 22465 21091 22523 21097
rect 22738 21088 22744 21100
rect 22796 21128 22802 21140
rect 24302 21128 24308 21140
rect 22796 21100 24308 21128
rect 22796 21088 22802 21100
rect 24302 21088 24308 21100
rect 24360 21088 24366 21140
rect 24489 21131 24547 21137
rect 24489 21097 24501 21131
rect 24535 21128 24547 21131
rect 24854 21128 24860 21140
rect 24535 21100 24860 21128
rect 24535 21097 24547 21100
rect 24489 21091 24547 21097
rect 24854 21088 24860 21100
rect 24912 21088 24918 21140
rect 26142 21128 26148 21140
rect 25332 21100 26148 21128
rect 17402 21020 17408 21072
rect 17460 21060 17466 21072
rect 17460 21032 18828 21060
rect 17460 21020 17466 21032
rect 18693 20995 18751 21001
rect 18693 20992 18705 20995
rect 17880 20964 18705 20992
rect 17218 20924 17224 20936
rect 17179 20896 17224 20924
rect 17218 20884 17224 20896
rect 17276 20884 17282 20936
rect 17880 20933 17908 20964
rect 18693 20961 18705 20964
rect 18739 20961 18751 20995
rect 18693 20955 18751 20961
rect 17865 20927 17923 20933
rect 17865 20893 17877 20927
rect 17911 20893 17923 20927
rect 17865 20887 17923 20893
rect 18230 20884 18236 20936
rect 18288 20924 18294 20936
rect 18325 20927 18383 20933
rect 18325 20924 18337 20927
rect 18288 20896 18337 20924
rect 18288 20884 18294 20896
rect 18325 20893 18337 20896
rect 18371 20893 18383 20927
rect 18325 20887 18383 20893
rect 18509 20927 18567 20933
rect 18509 20893 18521 20927
rect 18555 20924 18567 20927
rect 18800 20924 18828 21032
rect 23290 21020 23296 21072
rect 23348 21060 23354 21072
rect 23348 21032 23612 21060
rect 23348 21020 23354 21032
rect 20806 20992 20812 21004
rect 19812 20964 20812 20992
rect 19812 20933 19840 20964
rect 20806 20952 20812 20964
rect 20864 20952 20870 21004
rect 21082 20992 21088 21004
rect 21043 20964 21088 20992
rect 21082 20952 21088 20964
rect 21140 20952 21146 21004
rect 22925 20995 22983 21001
rect 22925 20961 22937 20995
rect 22971 20961 22983 20995
rect 22925 20955 22983 20961
rect 18555 20896 18828 20924
rect 19797 20927 19855 20933
rect 18555 20893 18567 20896
rect 18509 20887 18567 20893
rect 19797 20893 19809 20927
rect 19843 20893 19855 20927
rect 19978 20924 19984 20936
rect 19939 20896 19984 20924
rect 19797 20887 19855 20893
rect 19978 20884 19984 20896
rect 20036 20884 20042 20936
rect 20438 20924 20444 20936
rect 20399 20896 20444 20924
rect 20438 20884 20444 20896
rect 20496 20884 20502 20936
rect 21352 20927 21410 20933
rect 21352 20893 21364 20927
rect 21398 20924 21410 20927
rect 22940 20924 22968 20955
rect 23014 20952 23020 21004
rect 23072 20992 23078 21004
rect 23584 20992 23612 21032
rect 24670 21020 24676 21072
rect 24728 21060 24734 21072
rect 25332 21060 25360 21100
rect 26142 21088 26148 21100
rect 26200 21088 26206 21140
rect 26694 21088 26700 21140
rect 26752 21128 26758 21140
rect 28261 21131 28319 21137
rect 28261 21128 28273 21131
rect 26752 21100 28273 21128
rect 26752 21088 26758 21100
rect 28261 21097 28273 21100
rect 28307 21097 28319 21131
rect 28261 21091 28319 21097
rect 29454 21088 29460 21140
rect 29512 21128 29518 21140
rect 29512 21100 30503 21128
rect 29512 21088 29518 21100
rect 24728 21032 25360 21060
rect 24728 21020 24734 21032
rect 25406 21020 25412 21072
rect 25464 21020 25470 21072
rect 26789 21063 26847 21069
rect 26789 21029 26801 21063
rect 26835 21060 26847 21063
rect 30475 21060 30503 21100
rect 30650 21088 30656 21140
rect 30708 21128 30714 21140
rect 30929 21131 30987 21137
rect 30929 21128 30941 21131
rect 30708 21100 30941 21128
rect 30708 21088 30714 21100
rect 30929 21097 30941 21100
rect 30975 21097 30987 21131
rect 31570 21128 31576 21140
rect 31531 21100 31576 21128
rect 30929 21091 30987 21097
rect 31570 21088 31576 21100
rect 31628 21088 31634 21140
rect 32306 21088 32312 21140
rect 32364 21128 32370 21140
rect 33873 21131 33931 21137
rect 33873 21128 33885 21131
rect 32364 21100 33885 21128
rect 32364 21088 32370 21100
rect 33873 21097 33885 21100
rect 33919 21097 33931 21131
rect 33873 21091 33931 21097
rect 26835 21032 27844 21060
rect 30475 21032 32168 21060
rect 26835 21029 26847 21032
rect 26789 21023 26847 21029
rect 24762 20992 24768 21004
rect 23072 20964 23336 20992
rect 23072 20952 23078 20964
rect 23198 20924 23204 20936
rect 21398 20896 22968 20924
rect 23159 20896 23204 20924
rect 21398 20893 21410 20896
rect 21352 20887 21410 20893
rect 23198 20884 23204 20896
rect 23256 20884 23262 20936
rect 23308 20933 23336 20964
rect 23584 20964 24768 20992
rect 23293 20927 23351 20933
rect 23293 20893 23305 20927
rect 23339 20893 23351 20927
rect 23293 20887 23351 20893
rect 23382 20884 23388 20936
rect 23440 20924 23446 20936
rect 23584 20933 23612 20964
rect 24762 20952 24768 20964
rect 24820 20952 24826 21004
rect 25424 20992 25452 21020
rect 27706 20992 27712 21004
rect 24964 20964 25452 20992
rect 27667 20964 27712 20992
rect 23569 20927 23627 20933
rect 23440 20896 23485 20924
rect 23440 20884 23446 20896
rect 23569 20893 23581 20927
rect 23615 20893 23627 20927
rect 23569 20887 23627 20893
rect 24673 20927 24731 20933
rect 24673 20893 24685 20927
rect 24719 20924 24731 20927
rect 24854 20924 24860 20936
rect 24719 20896 24860 20924
rect 24719 20893 24731 20896
rect 24673 20887 24731 20893
rect 24854 20884 24860 20896
rect 24912 20884 24918 20936
rect 24964 20933 24992 20964
rect 27706 20952 27712 20964
rect 27764 20952 27770 21004
rect 27816 20992 27844 21032
rect 28166 20992 28172 21004
rect 27816 20964 28172 20992
rect 24949 20927 25007 20933
rect 24949 20893 24961 20927
rect 24995 20893 25007 20927
rect 24949 20887 25007 20893
rect 25038 20884 25044 20936
rect 25096 20924 25102 20936
rect 25409 20927 25467 20933
rect 25409 20924 25421 20927
rect 25096 20896 25421 20924
rect 25096 20884 25102 20896
rect 25409 20893 25421 20896
rect 25455 20924 25467 20927
rect 25498 20924 25504 20936
rect 25455 20896 25504 20924
rect 25455 20893 25467 20896
rect 25409 20887 25467 20893
rect 25498 20884 25504 20896
rect 25556 20884 25562 20936
rect 25608 20896 25912 20924
rect 15286 20816 15292 20868
rect 15344 20856 15350 20868
rect 25608 20856 25636 20896
rect 25682 20865 25688 20868
rect 15344 20828 25636 20856
rect 15344 20816 15350 20828
rect 25676 20819 25688 20865
rect 25740 20856 25746 20868
rect 25884 20856 25912 20896
rect 27246 20884 27252 20936
rect 27304 20924 27310 20936
rect 27433 20927 27491 20933
rect 27433 20924 27445 20927
rect 27304 20896 27445 20924
rect 27304 20884 27310 20896
rect 27433 20893 27445 20896
rect 27479 20893 27491 20927
rect 27433 20887 27491 20893
rect 27522 20884 27528 20936
rect 27580 20924 27586 20936
rect 27816 20933 27844 20964
rect 28166 20952 28172 20964
rect 28224 20952 28230 21004
rect 27801 20927 27859 20933
rect 27580 20896 27625 20924
rect 27580 20884 27586 20896
rect 27801 20893 27813 20927
rect 27847 20893 27859 20927
rect 27801 20887 27859 20893
rect 27890 20884 27896 20936
rect 27948 20924 27954 20936
rect 28445 20927 28503 20933
rect 28445 20924 28457 20927
rect 27948 20896 28457 20924
rect 27948 20884 27954 20896
rect 28445 20893 28457 20896
rect 28491 20893 28503 20927
rect 28718 20924 28724 20936
rect 28679 20896 28724 20924
rect 28445 20887 28503 20893
rect 28718 20884 28724 20896
rect 28776 20884 28782 20936
rect 28994 20884 29000 20936
rect 29052 20924 29058 20936
rect 29454 20924 29460 20936
rect 29052 20896 29460 20924
rect 29052 20884 29058 20896
rect 29454 20884 29460 20896
rect 29512 20924 29518 20936
rect 32140 20933 32168 21032
rect 33042 20952 33048 21004
rect 33100 20992 33106 21004
rect 33100 20964 34100 20992
rect 33100 20952 33106 20964
rect 29549 20927 29607 20933
rect 29549 20924 29561 20927
rect 29512 20896 29561 20924
rect 29512 20884 29518 20896
rect 29549 20893 29561 20896
rect 29595 20893 29607 20927
rect 31481 20927 31539 20933
rect 31481 20924 31493 20927
rect 29549 20887 29607 20893
rect 29656 20896 31493 20924
rect 29656 20856 29684 20896
rect 31481 20893 31493 20896
rect 31527 20893 31539 20927
rect 31481 20887 31539 20893
rect 32125 20927 32183 20933
rect 32125 20893 32137 20927
rect 32171 20893 32183 20927
rect 32125 20887 32183 20893
rect 32309 20927 32367 20933
rect 32309 20893 32321 20927
rect 32355 20893 32367 20927
rect 32309 20887 32367 20893
rect 25740 20828 25776 20856
rect 25884 20828 29684 20856
rect 29816 20859 29874 20865
rect 25682 20816 25688 20819
rect 25740 20816 25746 20828
rect 29816 20825 29828 20859
rect 29862 20825 29874 20859
rect 29816 20819 29874 20825
rect 16850 20748 16856 20800
rect 16908 20788 16914 20800
rect 19889 20791 19947 20797
rect 19889 20788 19901 20791
rect 16908 20760 19901 20788
rect 16908 20748 16914 20760
rect 19889 20757 19901 20760
rect 19935 20788 19947 20791
rect 22370 20788 22376 20800
rect 19935 20760 22376 20788
rect 19935 20757 19947 20760
rect 19889 20751 19947 20757
rect 22370 20748 22376 20760
rect 22428 20748 22434 20800
rect 23842 20748 23848 20800
rect 23900 20788 23906 20800
rect 24578 20788 24584 20800
rect 23900 20760 24584 20788
rect 23900 20748 23906 20760
rect 24578 20748 24584 20760
rect 24636 20748 24642 20800
rect 24857 20791 24915 20797
rect 24857 20757 24869 20791
rect 24903 20788 24915 20791
rect 26878 20788 26884 20800
rect 24903 20760 26884 20788
rect 24903 20757 24915 20760
rect 24857 20751 24915 20757
rect 26878 20748 26884 20760
rect 26936 20748 26942 20800
rect 27249 20791 27307 20797
rect 27249 20757 27261 20791
rect 27295 20788 27307 20791
rect 28629 20791 28687 20797
rect 28629 20788 28641 20791
rect 27295 20760 28641 20788
rect 27295 20757 27307 20760
rect 27249 20751 27307 20757
rect 28629 20757 28641 20760
rect 28675 20757 28687 20791
rect 28629 20751 28687 20757
rect 29638 20748 29644 20800
rect 29696 20788 29702 20800
rect 29840 20788 29868 20819
rect 30190 20816 30196 20868
rect 30248 20856 30254 20868
rect 32217 20859 32275 20865
rect 32217 20856 32229 20859
rect 30248 20828 32229 20856
rect 30248 20816 30254 20828
rect 32217 20825 32229 20828
rect 32263 20825 32275 20859
rect 32217 20819 32275 20825
rect 29696 20760 29868 20788
rect 29696 20748 29702 20760
rect 31018 20748 31024 20800
rect 31076 20788 31082 20800
rect 32324 20788 32352 20887
rect 33134 20884 33140 20936
rect 33192 20924 33198 20936
rect 34072 20933 34100 20964
rect 33229 20927 33287 20933
rect 33229 20924 33241 20927
rect 33192 20896 33241 20924
rect 33192 20884 33198 20896
rect 33229 20893 33241 20896
rect 33275 20893 33287 20927
rect 33229 20887 33287 20893
rect 34057 20927 34115 20933
rect 34057 20893 34069 20927
rect 34103 20893 34115 20927
rect 34057 20887 34115 20893
rect 33244 20856 33272 20887
rect 34330 20856 34336 20868
rect 33244 20828 34336 20856
rect 34330 20816 34336 20828
rect 34388 20816 34394 20868
rect 33318 20788 33324 20800
rect 31076 20760 32352 20788
rect 33279 20760 33324 20788
rect 31076 20748 31082 20760
rect 33318 20748 33324 20760
rect 33376 20748 33382 20800
rect 1104 20698 34868 20720
rect 1104 20646 12214 20698
rect 12266 20646 12278 20698
rect 12330 20646 12342 20698
rect 12394 20646 12406 20698
rect 12458 20646 12470 20698
rect 12522 20646 23478 20698
rect 23530 20646 23542 20698
rect 23594 20646 23606 20698
rect 23658 20646 23670 20698
rect 23722 20646 23734 20698
rect 23786 20646 34868 20698
rect 1104 20624 34868 20646
rect 16114 20544 16120 20596
rect 16172 20584 16178 20596
rect 22370 20584 22376 20596
rect 16172 20556 22376 20584
rect 16172 20544 16178 20556
rect 22370 20544 22376 20556
rect 22428 20544 22434 20596
rect 22462 20544 22468 20596
rect 22520 20584 22526 20596
rect 23106 20584 23112 20596
rect 22520 20556 23112 20584
rect 22520 20544 22526 20556
rect 23106 20544 23112 20556
rect 23164 20584 23170 20596
rect 23569 20587 23627 20593
rect 23569 20584 23581 20587
rect 23164 20556 23581 20584
rect 23164 20544 23170 20556
rect 23569 20553 23581 20556
rect 23615 20553 23627 20587
rect 23934 20584 23940 20596
rect 23569 20547 23627 20553
rect 23676 20556 23940 20584
rect 21177 20519 21235 20525
rect 21177 20485 21189 20519
rect 21223 20516 21235 20519
rect 22002 20516 22008 20528
rect 21223 20488 22008 20516
rect 21223 20485 21235 20488
rect 21177 20479 21235 20485
rect 22002 20476 22008 20488
rect 22060 20476 22066 20528
rect 23474 20516 23480 20528
rect 22848 20488 23480 20516
rect 18506 20448 18512 20460
rect 18467 20420 18512 20448
rect 18506 20408 18512 20420
rect 18564 20408 18570 20460
rect 20441 20451 20499 20457
rect 20441 20417 20453 20451
rect 20487 20417 20499 20451
rect 21082 20448 21088 20460
rect 21043 20420 21088 20448
rect 20441 20411 20499 20417
rect 20456 20380 20484 20411
rect 21082 20408 21088 20420
rect 21140 20408 21146 20460
rect 21266 20448 21272 20460
rect 21227 20420 21272 20448
rect 21266 20408 21272 20420
rect 21324 20408 21330 20460
rect 21634 20408 21640 20460
rect 21692 20448 21698 20460
rect 22848 20457 22876 20488
rect 23474 20476 23480 20488
rect 23532 20476 23538 20528
rect 21913 20451 21971 20457
rect 21913 20448 21925 20451
rect 21692 20420 21925 20448
rect 21692 20408 21698 20420
rect 21913 20417 21925 20420
rect 21959 20417 21971 20451
rect 21913 20411 21971 20417
rect 22833 20451 22891 20457
rect 22833 20417 22845 20451
rect 22879 20417 22891 20451
rect 22833 20411 22891 20417
rect 23017 20451 23075 20457
rect 23017 20417 23029 20451
rect 23063 20448 23075 20451
rect 23106 20448 23112 20460
rect 23063 20420 23112 20448
rect 23063 20417 23075 20420
rect 23017 20411 23075 20417
rect 23106 20408 23112 20420
rect 23164 20408 23170 20460
rect 23676 20448 23704 20556
rect 23934 20544 23940 20556
rect 23992 20584 23998 20596
rect 24118 20584 24124 20596
rect 23992 20556 24124 20584
rect 23992 20544 23998 20556
rect 24118 20544 24124 20556
rect 24176 20544 24182 20596
rect 24302 20544 24308 20596
rect 24360 20584 24366 20596
rect 24360 20556 27568 20584
rect 24360 20544 24366 20556
rect 24486 20516 24492 20528
rect 23492 20420 23704 20448
rect 23952 20488 24492 20516
rect 21818 20380 21824 20392
rect 20456 20352 21824 20380
rect 21818 20340 21824 20352
rect 21876 20340 21882 20392
rect 22097 20383 22155 20389
rect 22097 20349 22109 20383
rect 22143 20380 22155 20383
rect 22554 20380 22560 20392
rect 22143 20352 22560 20380
rect 22143 20349 22155 20352
rect 22097 20343 22155 20349
rect 22554 20340 22560 20352
rect 22612 20340 22618 20392
rect 22741 20383 22799 20389
rect 22741 20349 22753 20383
rect 22787 20349 22799 20383
rect 22741 20343 22799 20349
rect 22925 20383 22983 20389
rect 22925 20349 22937 20383
rect 22971 20380 22983 20383
rect 23492 20380 23520 20420
rect 22971 20352 23520 20380
rect 22971 20349 22983 20352
rect 22925 20343 22983 20349
rect 18322 20312 18328 20324
rect 18283 20284 18328 20312
rect 18322 20272 18328 20284
rect 18380 20272 18386 20324
rect 20533 20315 20591 20321
rect 20533 20281 20545 20315
rect 20579 20312 20591 20315
rect 22646 20312 22652 20324
rect 20579 20284 22652 20312
rect 20579 20281 20591 20284
rect 20533 20275 20591 20281
rect 22646 20272 22652 20284
rect 22704 20272 22710 20324
rect 22756 20312 22784 20343
rect 23566 20340 23572 20392
rect 23624 20380 23630 20392
rect 23952 20389 23980 20488
rect 24486 20476 24492 20488
rect 24544 20516 24550 20528
rect 27540 20516 27568 20556
rect 28166 20544 28172 20596
rect 28224 20584 28230 20596
rect 28224 20556 28580 20584
rect 28224 20544 28230 20556
rect 28552 20525 28580 20556
rect 28626 20544 28632 20596
rect 28684 20584 28690 20596
rect 28813 20587 28871 20593
rect 28813 20584 28825 20587
rect 28684 20556 28825 20584
rect 28684 20544 28690 20556
rect 28813 20553 28825 20556
rect 28859 20553 28871 20587
rect 28813 20547 28871 20553
rect 29362 20544 29368 20596
rect 29420 20584 29426 20596
rect 29473 20587 29531 20593
rect 29473 20584 29485 20587
rect 29420 20556 29485 20584
rect 29420 20544 29426 20556
rect 29473 20553 29485 20556
rect 29519 20553 29531 20587
rect 31021 20587 31079 20593
rect 31021 20584 31033 20587
rect 29473 20547 29531 20553
rect 29580 20556 31033 20584
rect 28445 20519 28503 20525
rect 24544 20488 26372 20516
rect 24544 20476 24550 20488
rect 26344 20460 26372 20488
rect 27540 20488 28305 20516
rect 24946 20448 24952 20460
rect 24859 20420 24952 20448
rect 24946 20408 24952 20420
rect 25004 20448 25010 20460
rect 25774 20448 25780 20460
rect 25004 20420 25780 20448
rect 25004 20408 25010 20420
rect 25774 20408 25780 20420
rect 25832 20408 25838 20460
rect 25958 20448 25964 20460
rect 25919 20420 25964 20448
rect 25958 20408 25964 20420
rect 26016 20408 26022 20460
rect 26142 20448 26148 20460
rect 26103 20420 26148 20448
rect 26142 20408 26148 20420
rect 26200 20408 26206 20460
rect 26326 20448 26332 20460
rect 26287 20420 26332 20448
rect 26326 20408 26332 20420
rect 26384 20408 26390 20460
rect 26694 20408 26700 20460
rect 26752 20448 26758 20460
rect 26973 20451 27031 20457
rect 26973 20448 26985 20451
rect 26752 20420 26985 20448
rect 26752 20408 26758 20420
rect 26973 20417 26985 20420
rect 27019 20417 27031 20451
rect 27154 20448 27160 20460
rect 27115 20420 27160 20448
rect 26973 20411 27031 20417
rect 27154 20408 27160 20420
rect 27212 20408 27218 20460
rect 27338 20448 27344 20460
rect 27299 20420 27344 20448
rect 27338 20408 27344 20420
rect 27396 20408 27402 20460
rect 27540 20457 27568 20488
rect 28277 20457 28305 20488
rect 28445 20485 28457 20519
rect 28491 20485 28503 20519
rect 28445 20479 28503 20485
rect 28537 20519 28595 20525
rect 28537 20485 28549 20519
rect 28583 20485 28595 20519
rect 28537 20479 28595 20485
rect 29273 20519 29331 20525
rect 29273 20485 29285 20519
rect 29319 20485 29331 20519
rect 29580 20516 29608 20556
rect 31021 20553 31033 20556
rect 31067 20553 31079 20587
rect 31021 20547 31079 20553
rect 30466 20516 30472 20528
rect 29273 20479 29331 20485
rect 29472 20488 29608 20516
rect 29656 20488 30472 20516
rect 27525 20451 27583 20457
rect 27525 20417 27537 20451
rect 27571 20417 27583 20451
rect 27525 20411 27583 20417
rect 27709 20451 27767 20457
rect 27709 20417 27721 20451
rect 27755 20448 27767 20451
rect 28169 20451 28227 20457
rect 28169 20448 28181 20451
rect 27755 20420 28181 20448
rect 27755 20417 27767 20420
rect 27709 20411 27767 20417
rect 28169 20417 28181 20420
rect 28215 20417 28227 20451
rect 28169 20411 28227 20417
rect 28262 20451 28320 20457
rect 28262 20417 28274 20451
rect 28308 20417 28320 20451
rect 28262 20411 28320 20417
rect 23937 20383 23995 20389
rect 23937 20380 23949 20383
rect 23624 20352 23949 20380
rect 23624 20340 23630 20352
rect 23937 20349 23949 20352
rect 23983 20349 23995 20383
rect 23937 20343 23995 20349
rect 24029 20383 24087 20389
rect 24029 20349 24041 20383
rect 24075 20349 24087 20383
rect 24029 20343 24087 20349
rect 23842 20312 23848 20324
rect 22756 20284 23848 20312
rect 23842 20272 23848 20284
rect 23900 20272 23906 20324
rect 22278 20204 22284 20256
rect 22336 20244 22342 20256
rect 22557 20247 22615 20253
rect 22557 20244 22569 20247
rect 22336 20216 22569 20244
rect 22336 20204 22342 20216
rect 22557 20213 22569 20216
rect 22603 20213 22615 20247
rect 22557 20207 22615 20213
rect 22922 20204 22928 20256
rect 22980 20244 22986 20256
rect 24044 20244 24072 20343
rect 24118 20340 24124 20392
rect 24176 20380 24182 20392
rect 24673 20383 24731 20389
rect 24673 20380 24685 20383
rect 24176 20352 24685 20380
rect 24176 20340 24182 20352
rect 24673 20349 24685 20352
rect 24719 20349 24731 20383
rect 24673 20343 24731 20349
rect 26421 20383 26479 20389
rect 26421 20349 26433 20383
rect 26467 20380 26479 20383
rect 26510 20380 26516 20392
rect 26467 20352 26516 20380
rect 26467 20349 26479 20352
rect 26421 20343 26479 20349
rect 26510 20340 26516 20352
rect 26568 20380 26574 20392
rect 27249 20383 27307 20389
rect 27249 20380 27261 20383
rect 26568 20352 27261 20380
rect 26568 20340 26574 20352
rect 27249 20349 27261 20352
rect 27295 20349 27307 20383
rect 27356 20380 27384 20408
rect 28460 20380 28488 20479
rect 28634 20451 28692 20457
rect 28634 20417 28646 20451
rect 28680 20417 28692 20451
rect 28634 20411 28692 20417
rect 27356 20352 28488 20380
rect 27249 20343 27307 20349
rect 26234 20272 26240 20324
rect 26292 20312 26298 20324
rect 28649 20312 28677 20411
rect 29288 20380 29316 20479
rect 29472 20460 29500 20488
rect 29454 20408 29460 20460
rect 29512 20408 29518 20460
rect 29656 20380 29684 20488
rect 30466 20476 30472 20488
rect 30524 20476 30530 20528
rect 30929 20519 30987 20525
rect 30929 20485 30941 20519
rect 30975 20516 30987 20519
rect 31570 20516 31576 20528
rect 30975 20488 31576 20516
rect 30975 20485 30987 20488
rect 30929 20479 30987 20485
rect 31570 20476 31576 20488
rect 31628 20476 31634 20528
rect 32493 20519 32551 20525
rect 32493 20485 32505 20519
rect 32539 20516 32551 20519
rect 33318 20516 33324 20528
rect 32539 20488 33324 20516
rect 32539 20485 32551 20488
rect 32493 20479 32551 20485
rect 33318 20476 33324 20488
rect 33376 20476 33382 20528
rect 30101 20451 30159 20457
rect 30101 20448 30113 20451
rect 29288 20352 29684 20380
rect 29748 20420 30113 20448
rect 26292 20284 28677 20312
rect 26292 20272 26298 20284
rect 28718 20272 28724 20324
rect 28776 20312 28782 20324
rect 29641 20315 29699 20321
rect 29641 20312 29653 20315
rect 28776 20284 29653 20312
rect 28776 20272 28782 20284
rect 29641 20281 29653 20284
rect 29687 20312 29699 20315
rect 29748 20312 29776 20420
rect 30101 20417 30113 20420
rect 30147 20417 30159 20451
rect 30101 20411 30159 20417
rect 30377 20451 30435 20457
rect 30377 20417 30389 20451
rect 30423 20448 30435 20451
rect 31846 20448 31852 20460
rect 30423 20420 31852 20448
rect 30423 20417 30435 20420
rect 30377 20411 30435 20417
rect 31846 20408 31852 20420
rect 31904 20408 31910 20460
rect 34146 20448 34152 20460
rect 34107 20420 34152 20448
rect 34146 20408 34152 20420
rect 34204 20408 34210 20460
rect 31018 20340 31024 20392
rect 31076 20380 31082 20392
rect 32309 20383 32367 20389
rect 32309 20380 32321 20383
rect 31076 20352 32321 20380
rect 31076 20340 31082 20352
rect 32309 20349 32321 20352
rect 32355 20349 32367 20383
rect 32309 20343 32367 20349
rect 30190 20312 30196 20324
rect 29687 20284 29776 20312
rect 30151 20284 30196 20312
rect 29687 20281 29699 20284
rect 29641 20275 29699 20281
rect 30190 20272 30196 20284
rect 30248 20272 30254 20324
rect 22980 20216 24072 20244
rect 24213 20247 24271 20253
rect 22980 20204 22986 20216
rect 24213 20213 24225 20247
rect 24259 20244 24271 20247
rect 24486 20244 24492 20256
rect 24259 20216 24492 20244
rect 24259 20213 24271 20216
rect 24213 20207 24271 20213
rect 24486 20204 24492 20216
rect 24544 20204 24550 20256
rect 28626 20204 28632 20256
rect 28684 20244 28690 20256
rect 29454 20244 29460 20256
rect 28684 20216 29460 20244
rect 28684 20204 28690 20216
rect 29454 20204 29460 20216
rect 29512 20204 29518 20256
rect 30098 20244 30104 20256
rect 30059 20216 30104 20244
rect 30098 20204 30104 20216
rect 30156 20204 30162 20256
rect 30926 20204 30932 20256
rect 30984 20244 30990 20256
rect 31754 20244 31760 20256
rect 30984 20216 31760 20244
rect 30984 20204 30990 20216
rect 31754 20204 31760 20216
rect 31812 20204 31818 20256
rect 1104 20154 34868 20176
rect 1104 20102 6582 20154
rect 6634 20102 6646 20154
rect 6698 20102 6710 20154
rect 6762 20102 6774 20154
rect 6826 20102 6838 20154
rect 6890 20102 17846 20154
rect 17898 20102 17910 20154
rect 17962 20102 17974 20154
rect 18026 20102 18038 20154
rect 18090 20102 18102 20154
rect 18154 20102 29110 20154
rect 29162 20102 29174 20154
rect 29226 20102 29238 20154
rect 29290 20102 29302 20154
rect 29354 20102 29366 20154
rect 29418 20102 34868 20154
rect 1104 20080 34868 20102
rect 19978 20000 19984 20052
rect 20036 20040 20042 20052
rect 20441 20043 20499 20049
rect 20441 20040 20453 20043
rect 20036 20012 20453 20040
rect 20036 20000 20042 20012
rect 20441 20009 20453 20012
rect 20487 20009 20499 20043
rect 20441 20003 20499 20009
rect 22557 20043 22615 20049
rect 22557 20009 22569 20043
rect 22603 20040 22615 20043
rect 22830 20040 22836 20052
rect 22603 20012 22836 20040
rect 22603 20009 22615 20012
rect 22557 20003 22615 20009
rect 22830 20000 22836 20012
rect 22888 20000 22894 20052
rect 26234 20040 26240 20052
rect 26195 20012 26240 20040
rect 26234 20000 26240 20012
rect 26292 20000 26298 20052
rect 27341 20043 27399 20049
rect 27341 20009 27353 20043
rect 27387 20040 27399 20043
rect 27890 20040 27896 20052
rect 27387 20012 27896 20040
rect 27387 20009 27399 20012
rect 27341 20003 27399 20009
rect 27890 20000 27896 20012
rect 27948 20000 27954 20052
rect 27985 20043 28043 20049
rect 27985 20009 27997 20043
rect 28031 20009 28043 20043
rect 27985 20003 28043 20009
rect 23474 19932 23480 19984
rect 23532 19972 23538 19984
rect 23753 19975 23811 19981
rect 23753 19972 23765 19975
rect 23532 19944 23765 19972
rect 23532 19932 23538 19944
rect 23753 19941 23765 19944
rect 23799 19941 23811 19975
rect 26142 19972 26148 19984
rect 23753 19935 23811 19941
rect 24320 19944 26148 19972
rect 22278 19904 22284 19916
rect 22239 19876 22284 19904
rect 22278 19864 22284 19876
rect 22336 19864 22342 19916
rect 23290 19904 23296 19916
rect 23203 19876 23296 19904
rect 23290 19864 23296 19876
rect 23348 19904 23354 19916
rect 24320 19904 24348 19944
rect 26142 19932 26148 19944
rect 26200 19932 26206 19984
rect 24486 19904 24492 19916
rect 23348 19876 24348 19904
rect 24447 19876 24492 19904
rect 23348 19864 23354 19876
rect 24486 19864 24492 19876
rect 24544 19864 24550 19916
rect 24762 19864 24768 19916
rect 24820 19904 24826 19916
rect 25685 19907 25743 19913
rect 25685 19904 25697 19907
rect 24820 19876 25697 19904
rect 24820 19864 24826 19876
rect 25685 19873 25697 19876
rect 25731 19873 25743 19907
rect 25685 19867 25743 19873
rect 26160 19876 27292 19904
rect 1762 19796 1768 19848
rect 1820 19836 1826 19848
rect 1949 19839 2007 19845
rect 1949 19836 1961 19839
rect 1820 19808 1961 19836
rect 1820 19796 1826 19808
rect 1949 19805 1961 19808
rect 1995 19805 2007 19839
rect 1949 19799 2007 19805
rect 20441 19839 20499 19845
rect 20441 19805 20453 19839
rect 20487 19805 20499 19839
rect 20441 19799 20499 19805
rect 20625 19839 20683 19845
rect 20625 19805 20637 19839
rect 20671 19836 20683 19839
rect 21726 19836 21732 19848
rect 20671 19808 21732 19836
rect 20671 19805 20683 19808
rect 20625 19799 20683 19805
rect 20456 19700 20484 19799
rect 21726 19796 21732 19808
rect 21784 19796 21790 19848
rect 22186 19836 22192 19848
rect 22147 19808 22192 19836
rect 22186 19796 22192 19808
rect 22244 19796 22250 19848
rect 23385 19839 23443 19845
rect 23385 19805 23397 19839
rect 23431 19836 23443 19839
rect 23566 19836 23572 19848
rect 23431 19808 23572 19836
rect 23431 19805 23443 19808
rect 23385 19799 23443 19805
rect 23566 19796 23572 19808
rect 23624 19796 23630 19848
rect 23842 19796 23848 19848
rect 23900 19836 23906 19848
rect 24581 19839 24639 19845
rect 24581 19836 24593 19839
rect 23900 19808 24593 19836
rect 23900 19796 23906 19808
rect 24581 19805 24593 19808
rect 24627 19805 24639 19839
rect 24581 19799 24639 19805
rect 25222 19796 25228 19848
rect 25280 19796 25286 19848
rect 26160 19845 26188 19876
rect 26145 19839 26203 19845
rect 26145 19805 26157 19839
rect 26191 19805 26203 19839
rect 26145 19799 26203 19805
rect 26326 19796 26332 19848
rect 26384 19836 26390 19848
rect 26789 19839 26847 19845
rect 26789 19836 26801 19839
rect 26384 19808 26801 19836
rect 26384 19796 26390 19808
rect 26789 19805 26801 19808
rect 26835 19805 26847 19839
rect 27154 19836 27160 19848
rect 27067 19808 27160 19836
rect 26789 19799 26847 19805
rect 27154 19796 27160 19808
rect 27212 19796 27218 19848
rect 27264 19836 27292 19876
rect 28000 19848 28028 20003
rect 28074 20000 28080 20052
rect 28132 20040 28138 20052
rect 28261 20043 28319 20049
rect 28261 20040 28273 20043
rect 28132 20012 28273 20040
rect 28132 20000 28138 20012
rect 28261 20009 28273 20012
rect 28307 20009 28319 20043
rect 28261 20003 28319 20009
rect 28350 20000 28356 20052
rect 28408 20040 28414 20052
rect 28408 20012 30144 20040
rect 28408 20000 28414 20012
rect 28721 19975 28779 19981
rect 28721 19941 28733 19975
rect 28767 19941 28779 19975
rect 28721 19935 28779 19941
rect 28626 19864 28632 19916
rect 28684 19864 28690 19916
rect 28736 19904 28764 19935
rect 29454 19932 29460 19984
rect 29512 19972 29518 19984
rect 29917 19975 29975 19981
rect 29512 19944 29868 19972
rect 29512 19932 29518 19944
rect 28736 19876 29776 19904
rect 27522 19836 27528 19848
rect 27264 19808 27528 19836
rect 27522 19796 27528 19808
rect 27580 19836 27586 19848
rect 27801 19839 27859 19845
rect 27801 19836 27813 19839
rect 27580 19808 27813 19836
rect 27580 19796 27586 19808
rect 27801 19805 27813 19808
rect 27847 19805 27859 19839
rect 27801 19799 27859 19805
rect 27982 19796 27988 19848
rect 28040 19796 28046 19848
rect 28644 19836 28672 19864
rect 28905 19839 28963 19845
rect 28905 19836 28917 19839
rect 28644 19808 28917 19836
rect 28905 19805 28917 19808
rect 28951 19805 28963 19839
rect 28905 19799 28963 19805
rect 28997 19839 29055 19845
rect 28997 19805 29009 19839
rect 29043 19836 29055 19839
rect 29454 19836 29460 19848
rect 29043 19808 29460 19836
rect 29043 19805 29055 19808
rect 28997 19799 29055 19805
rect 29454 19796 29460 19808
rect 29512 19796 29518 19848
rect 29748 19845 29776 19876
rect 29733 19839 29791 19845
rect 29733 19805 29745 19839
rect 29779 19805 29791 19839
rect 29840 19836 29868 19944
rect 29917 19941 29929 19975
rect 29963 19972 29975 19975
rect 30006 19972 30012 19984
rect 29963 19944 30012 19972
rect 29963 19941 29975 19944
rect 29917 19935 29975 19941
rect 30006 19932 30012 19944
rect 30064 19932 30070 19984
rect 30116 19972 30144 20012
rect 30190 20000 30196 20052
rect 30248 20040 30254 20052
rect 30469 20043 30527 20049
rect 30469 20040 30481 20043
rect 30248 20012 30481 20040
rect 30248 20000 30254 20012
rect 30469 20009 30481 20012
rect 30515 20009 30527 20043
rect 30469 20003 30527 20009
rect 32122 19972 32128 19984
rect 30116 19944 32128 19972
rect 32122 19932 32128 19944
rect 32180 19932 32186 19984
rect 30024 19904 30052 19932
rect 30024 19876 30788 19904
rect 30009 19839 30067 19845
rect 30009 19836 30021 19839
rect 29840 19808 30021 19836
rect 29733 19799 29791 19805
rect 30009 19805 30021 19808
rect 30055 19836 30067 19839
rect 30650 19836 30656 19848
rect 30055 19808 30656 19836
rect 30055 19805 30067 19808
rect 30009 19799 30067 19805
rect 30650 19796 30656 19808
rect 30708 19796 30714 19848
rect 30760 19845 30788 19876
rect 30745 19839 30803 19845
rect 30745 19805 30757 19839
rect 30791 19805 30803 19839
rect 30745 19799 30803 19805
rect 31205 19839 31263 19845
rect 31205 19805 31217 19839
rect 31251 19805 31263 19839
rect 31205 19799 31263 19805
rect 21361 19771 21419 19777
rect 21361 19737 21373 19771
rect 21407 19768 21419 19771
rect 22554 19768 22560 19780
rect 21407 19740 22560 19768
rect 21407 19737 21419 19740
rect 21361 19731 21419 19737
rect 22554 19728 22560 19740
rect 22612 19728 22618 19780
rect 22646 19728 22652 19780
rect 22704 19768 22710 19780
rect 25240 19768 25268 19796
rect 25501 19771 25559 19777
rect 25501 19768 25513 19771
rect 22704 19740 25513 19768
rect 22704 19728 22710 19740
rect 25501 19737 25513 19740
rect 25547 19737 25559 19771
rect 26970 19768 26976 19780
rect 26931 19740 26976 19768
rect 25501 19731 25559 19737
rect 26970 19728 26976 19740
rect 27028 19728 27034 19780
rect 27065 19771 27123 19777
rect 27065 19737 27077 19771
rect 27111 19737 27123 19771
rect 27065 19731 27123 19737
rect 21453 19703 21511 19709
rect 21453 19700 21465 19703
rect 20456 19672 21465 19700
rect 21453 19669 21465 19672
rect 21499 19700 21511 19703
rect 22922 19700 22928 19712
rect 21499 19672 22928 19700
rect 21499 19669 21511 19672
rect 21453 19663 21511 19669
rect 22922 19660 22928 19672
rect 22980 19660 22986 19712
rect 24949 19703 25007 19709
rect 24949 19669 24961 19703
rect 24995 19700 25007 19703
rect 25222 19700 25228 19712
rect 24995 19672 25228 19700
rect 24995 19669 25007 19672
rect 24949 19663 25007 19669
rect 25222 19660 25228 19672
rect 25280 19660 25286 19712
rect 26510 19660 26516 19712
rect 26568 19700 26574 19712
rect 27080 19700 27108 19731
rect 26568 19672 27108 19700
rect 27172 19700 27200 19796
rect 28442 19728 28448 19780
rect 28500 19768 28506 19780
rect 28721 19771 28779 19777
rect 28721 19768 28733 19771
rect 28500 19740 28733 19768
rect 28500 19728 28506 19740
rect 28721 19737 28733 19740
rect 28767 19768 28779 19771
rect 28810 19768 28816 19780
rect 28767 19740 28816 19768
rect 28767 19737 28779 19740
rect 28721 19731 28779 19737
rect 28810 19728 28816 19740
rect 28868 19728 28874 19780
rect 30466 19768 30472 19780
rect 28966 19740 29684 19768
rect 30427 19740 30472 19768
rect 28966 19700 28994 19740
rect 27172 19672 28994 19700
rect 26568 19660 26574 19672
rect 29362 19660 29368 19712
rect 29420 19700 29426 19712
rect 29549 19703 29607 19709
rect 29549 19700 29561 19703
rect 29420 19672 29561 19700
rect 29420 19660 29426 19672
rect 29549 19669 29561 19672
rect 29595 19669 29607 19703
rect 29656 19700 29684 19740
rect 30466 19728 30472 19740
rect 30524 19768 30530 19780
rect 30926 19768 30932 19780
rect 30524 19740 30932 19768
rect 30524 19728 30530 19740
rect 30926 19728 30932 19740
rect 30984 19768 30990 19780
rect 31220 19768 31248 19799
rect 31846 19796 31852 19848
rect 31904 19836 31910 19848
rect 32309 19839 32367 19845
rect 32309 19836 32321 19839
rect 31904 19808 32321 19836
rect 31904 19796 31910 19808
rect 32309 19805 32321 19808
rect 32355 19805 32367 19839
rect 32309 19799 32367 19805
rect 30984 19740 31248 19768
rect 32493 19771 32551 19777
rect 30984 19728 30990 19740
rect 32493 19737 32505 19771
rect 32539 19768 32551 19771
rect 33226 19768 33232 19780
rect 32539 19740 33232 19768
rect 32539 19737 32551 19740
rect 32493 19731 32551 19737
rect 33226 19728 33232 19740
rect 33284 19728 33290 19780
rect 34146 19768 34152 19780
rect 34107 19740 34152 19768
rect 34146 19728 34152 19740
rect 34204 19728 34210 19780
rect 31297 19703 31355 19709
rect 31297 19700 31309 19703
rect 29656 19672 31309 19700
rect 29549 19663 29607 19669
rect 31297 19669 31309 19672
rect 31343 19669 31355 19703
rect 31297 19663 31355 19669
rect 1104 19610 34868 19632
rect 1104 19558 12214 19610
rect 12266 19558 12278 19610
rect 12330 19558 12342 19610
rect 12394 19558 12406 19610
rect 12458 19558 12470 19610
rect 12522 19558 23478 19610
rect 23530 19558 23542 19610
rect 23594 19558 23606 19610
rect 23658 19558 23670 19610
rect 23722 19558 23734 19610
rect 23786 19558 34868 19610
rect 1104 19536 34868 19558
rect 21358 19496 21364 19508
rect 20640 19468 21364 19496
rect 1762 19360 1768 19372
rect 1723 19332 1768 19360
rect 1762 19320 1768 19332
rect 1820 19320 1826 19372
rect 20640 19369 20668 19468
rect 21358 19456 21364 19468
rect 21416 19456 21422 19508
rect 22020 19468 22212 19496
rect 20717 19431 20775 19437
rect 20717 19397 20729 19431
rect 20763 19428 20775 19431
rect 22020 19428 22048 19468
rect 20763 19400 22048 19428
rect 22184 19428 22212 19468
rect 22370 19456 22376 19508
rect 22428 19496 22434 19508
rect 22557 19499 22615 19505
rect 22557 19496 22569 19499
rect 22428 19468 22569 19496
rect 22428 19456 22434 19468
rect 22557 19465 22569 19468
rect 22603 19465 22615 19499
rect 22557 19459 22615 19465
rect 23934 19456 23940 19508
rect 23992 19496 23998 19508
rect 26329 19499 26387 19505
rect 23992 19468 24348 19496
rect 23992 19456 23998 19468
rect 22184 19400 22232 19428
rect 20763 19397 20775 19400
rect 20717 19391 20775 19397
rect 20625 19363 20683 19369
rect 20625 19329 20637 19363
rect 20671 19329 20683 19363
rect 20806 19360 20812 19372
rect 20767 19332 20812 19360
rect 20625 19323 20683 19329
rect 20806 19320 20812 19332
rect 20864 19320 20870 19372
rect 21358 19320 21364 19372
rect 21416 19360 21422 19372
rect 21416 19332 22140 19360
rect 21416 19320 21422 19332
rect 1946 19292 1952 19304
rect 1907 19264 1952 19292
rect 1946 19252 1952 19264
rect 2004 19252 2010 19304
rect 2222 19292 2228 19304
rect 2183 19264 2228 19292
rect 2222 19252 2228 19264
rect 2280 19252 2286 19304
rect 22112 19224 22140 19332
rect 22204 19292 22232 19400
rect 22278 19388 22284 19440
rect 22336 19428 22342 19440
rect 23382 19428 23388 19440
rect 22336 19400 22692 19428
rect 22336 19388 22342 19400
rect 22370 19360 22376 19372
rect 22331 19332 22376 19360
rect 22370 19320 22376 19332
rect 22428 19320 22434 19372
rect 22462 19320 22468 19372
rect 22520 19320 22526 19372
rect 22664 19369 22692 19400
rect 22756 19400 23388 19428
rect 22649 19363 22707 19369
rect 22649 19329 22661 19363
rect 22695 19329 22707 19363
rect 22649 19323 22707 19329
rect 22756 19334 22784 19400
rect 23382 19388 23388 19400
rect 23440 19428 23446 19440
rect 24320 19437 24348 19468
rect 26329 19465 26341 19499
rect 26375 19496 26387 19499
rect 27246 19496 27252 19508
rect 26375 19468 27252 19496
rect 26375 19465 26387 19468
rect 26329 19459 26387 19465
rect 27246 19456 27252 19468
rect 27304 19456 27310 19508
rect 27798 19496 27804 19508
rect 27356 19468 27804 19496
rect 24121 19431 24179 19437
rect 24121 19428 24133 19431
rect 23440 19400 24133 19428
rect 23440 19388 23446 19400
rect 24121 19397 24133 19400
rect 24167 19397 24179 19431
rect 24121 19391 24179 19397
rect 24305 19431 24363 19437
rect 24305 19397 24317 19431
rect 24351 19397 24363 19431
rect 24305 19391 24363 19397
rect 26970 19388 26976 19440
rect 27028 19428 27034 19440
rect 27356 19428 27384 19468
rect 27798 19456 27804 19468
rect 27856 19496 27862 19508
rect 29270 19496 29276 19508
rect 27856 19468 29276 19496
rect 27856 19456 27862 19468
rect 29270 19456 29276 19468
rect 29328 19456 29334 19508
rect 30650 19496 30656 19508
rect 30611 19468 30656 19496
rect 30650 19456 30656 19468
rect 30708 19456 30714 19508
rect 31205 19499 31263 19505
rect 31205 19465 31217 19499
rect 31251 19496 31263 19499
rect 31570 19496 31576 19508
rect 31251 19468 31576 19496
rect 31251 19465 31263 19468
rect 31205 19459 31263 19465
rect 31570 19456 31576 19468
rect 31628 19456 31634 19508
rect 32122 19496 32128 19508
rect 32083 19468 32128 19496
rect 32122 19456 32128 19468
rect 32180 19456 32186 19508
rect 33226 19496 33232 19508
rect 33187 19468 33232 19496
rect 33226 19456 33232 19468
rect 33284 19456 33290 19508
rect 33410 19456 33416 19508
rect 33468 19496 33474 19508
rect 33965 19499 34023 19505
rect 33965 19496 33977 19499
rect 33468 19468 33977 19496
rect 33468 19456 33474 19468
rect 33965 19465 33977 19468
rect 34011 19465 34023 19499
rect 33965 19459 34023 19465
rect 27706 19428 27712 19440
rect 27028 19400 27384 19428
rect 27448 19400 27712 19428
rect 27028 19388 27034 19400
rect 23293 19363 23351 19369
rect 22480 19292 22508 19320
rect 22756 19306 22876 19334
rect 23293 19329 23305 19363
rect 23339 19360 23351 19363
rect 24210 19360 24216 19372
rect 23339 19332 24216 19360
rect 23339 19329 23351 19332
rect 23293 19323 23351 19329
rect 24210 19320 24216 19332
rect 24268 19320 24274 19372
rect 24946 19360 24952 19372
rect 24907 19332 24952 19360
rect 24946 19320 24952 19332
rect 25004 19320 25010 19372
rect 26237 19363 26295 19369
rect 26237 19329 26249 19363
rect 26283 19360 26295 19363
rect 27246 19360 27252 19372
rect 26283 19332 27108 19360
rect 27207 19332 27252 19360
rect 26283 19329 26295 19332
rect 26237 19323 26295 19329
rect 22204 19264 22508 19292
rect 22848 19224 22876 19306
rect 23198 19292 23204 19304
rect 23159 19264 23204 19292
rect 23198 19252 23204 19264
rect 23256 19252 23262 19304
rect 23661 19295 23719 19301
rect 23661 19261 23673 19295
rect 23707 19292 23719 19295
rect 23842 19292 23848 19304
rect 23707 19264 23848 19292
rect 23707 19261 23719 19264
rect 23661 19255 23719 19261
rect 23842 19252 23848 19264
rect 23900 19252 23906 19304
rect 24394 19252 24400 19304
rect 24452 19292 24458 19304
rect 24489 19295 24547 19301
rect 24489 19292 24501 19295
rect 24452 19264 24501 19292
rect 24452 19252 24458 19264
rect 24489 19261 24501 19264
rect 24535 19261 24547 19295
rect 24489 19255 24547 19261
rect 25130 19252 25136 19304
rect 25188 19292 25194 19304
rect 25225 19295 25283 19301
rect 25225 19292 25237 19295
rect 25188 19264 25237 19292
rect 25188 19252 25194 19264
rect 25225 19261 25237 19264
rect 25271 19292 25283 19295
rect 25406 19292 25412 19304
rect 25271 19264 25412 19292
rect 25271 19261 25283 19264
rect 25225 19255 25283 19261
rect 25406 19252 25412 19264
rect 25464 19252 25470 19304
rect 22112 19196 22876 19224
rect 27080 19224 27108 19332
rect 27246 19320 27252 19332
rect 27304 19320 27310 19372
rect 27448 19369 27476 19400
rect 27706 19388 27712 19400
rect 27764 19428 27770 19440
rect 28353 19431 28411 19437
rect 28353 19428 28365 19431
rect 27764 19400 28365 19428
rect 27764 19388 27770 19400
rect 28353 19397 28365 19400
rect 28399 19397 28411 19431
rect 28353 19391 28411 19397
rect 29362 19388 29368 19440
rect 29420 19428 29426 19440
rect 29518 19431 29576 19437
rect 29518 19428 29530 19431
rect 29420 19400 29530 19428
rect 29420 19388 29426 19400
rect 29518 19397 29530 19400
rect 29564 19397 29576 19431
rect 29518 19391 29576 19397
rect 27433 19363 27491 19369
rect 27433 19329 27445 19363
rect 27479 19329 27491 19363
rect 27433 19323 27491 19329
rect 28169 19363 28227 19369
rect 28169 19329 28181 19363
rect 28215 19329 28227 19363
rect 28169 19323 28227 19329
rect 27522 19292 27528 19304
rect 27483 19264 27528 19292
rect 27522 19252 27528 19264
rect 27580 19252 27586 19304
rect 27985 19295 28043 19301
rect 27985 19261 27997 19295
rect 28031 19261 28043 19295
rect 28184 19292 28212 19323
rect 28718 19320 28724 19372
rect 28776 19320 28782 19372
rect 28994 19320 29000 19372
rect 29052 19360 29058 19372
rect 29273 19363 29331 19369
rect 29052 19350 29224 19360
rect 29273 19350 29285 19363
rect 29052 19332 29285 19350
rect 29052 19320 29058 19332
rect 29196 19329 29285 19332
rect 29319 19329 29331 19363
rect 30668 19360 30696 19456
rect 31113 19363 31171 19369
rect 31113 19360 31125 19363
rect 30668 19332 31125 19360
rect 29196 19323 29331 19329
rect 31113 19329 31125 19332
rect 31159 19329 31171 19363
rect 31113 19323 31171 19329
rect 29196 19322 29316 19323
rect 31570 19320 31576 19372
rect 31628 19360 31634 19372
rect 31754 19360 31760 19372
rect 31628 19332 31760 19360
rect 31628 19320 31634 19332
rect 31754 19320 31760 19332
rect 31812 19360 31818 19372
rect 32309 19363 32367 19369
rect 32309 19360 32321 19363
rect 31812 19332 32321 19360
rect 31812 19320 31818 19332
rect 32309 19329 32321 19332
rect 32355 19329 32367 19363
rect 32309 19323 32367 19329
rect 33137 19363 33195 19369
rect 33137 19329 33149 19363
rect 33183 19329 33195 19363
rect 33137 19323 33195 19329
rect 33873 19363 33931 19369
rect 33873 19329 33885 19363
rect 33919 19360 33931 19363
rect 34054 19360 34060 19372
rect 33919 19332 34060 19360
rect 33919 19329 33931 19332
rect 33873 19323 33931 19329
rect 28736 19292 28764 19320
rect 33152 19292 33180 19323
rect 34054 19320 34060 19332
rect 34112 19320 34118 19372
rect 28184 19264 28764 19292
rect 30300 19264 33180 19292
rect 27985 19255 28043 19261
rect 28000 19224 28028 19255
rect 28718 19224 28724 19236
rect 27080 19196 28724 19224
rect 28718 19184 28724 19196
rect 28776 19184 28782 19236
rect 22189 19159 22247 19165
rect 22189 19125 22201 19159
rect 22235 19156 22247 19159
rect 23382 19156 23388 19168
rect 22235 19128 23388 19156
rect 22235 19125 22247 19128
rect 22189 19119 22247 19125
rect 23382 19116 23388 19128
rect 23440 19116 23446 19168
rect 25130 19116 25136 19168
rect 25188 19156 25194 19168
rect 26418 19156 26424 19168
rect 25188 19128 26424 19156
rect 25188 19116 25194 19128
rect 26418 19116 26424 19128
rect 26476 19116 26482 19168
rect 27062 19156 27068 19168
rect 27023 19128 27068 19156
rect 27062 19116 27068 19128
rect 27120 19116 27126 19168
rect 28626 19116 28632 19168
rect 28684 19156 28690 19168
rect 30300 19156 30328 19264
rect 30374 19184 30380 19236
rect 30432 19224 30438 19236
rect 30432 19196 31754 19224
rect 30432 19184 30438 19196
rect 28684 19128 30328 19156
rect 31726 19156 31754 19196
rect 31938 19156 31944 19168
rect 31726 19128 31944 19156
rect 28684 19116 28690 19128
rect 31938 19116 31944 19128
rect 31996 19116 32002 19168
rect 1104 19066 34868 19088
rect 1104 19014 6582 19066
rect 6634 19014 6646 19066
rect 6698 19014 6710 19066
rect 6762 19014 6774 19066
rect 6826 19014 6838 19066
rect 6890 19014 17846 19066
rect 17898 19014 17910 19066
rect 17962 19014 17974 19066
rect 18026 19014 18038 19066
rect 18090 19014 18102 19066
rect 18154 19014 29110 19066
rect 29162 19014 29174 19066
rect 29226 19014 29238 19066
rect 29290 19014 29302 19066
rect 29354 19014 29366 19066
rect 29418 19014 34868 19066
rect 1104 18992 34868 19014
rect 1946 18912 1952 18964
rect 2004 18952 2010 18964
rect 2501 18955 2559 18961
rect 2501 18952 2513 18955
rect 2004 18924 2513 18952
rect 2004 18912 2010 18924
rect 2501 18921 2513 18924
rect 2547 18921 2559 18955
rect 2501 18915 2559 18921
rect 21729 18955 21787 18961
rect 21729 18921 21741 18955
rect 21775 18952 21787 18955
rect 22186 18952 22192 18964
rect 21775 18924 22192 18952
rect 21775 18921 21787 18924
rect 21729 18915 21787 18921
rect 22186 18912 22192 18924
rect 22244 18912 22250 18964
rect 22370 18912 22376 18964
rect 22428 18952 22434 18964
rect 22741 18955 22799 18961
rect 22741 18952 22753 18955
rect 22428 18924 22753 18952
rect 22428 18912 22434 18924
rect 22741 18921 22753 18924
rect 22787 18921 22799 18955
rect 22741 18915 22799 18921
rect 24581 18955 24639 18961
rect 24581 18921 24593 18955
rect 24627 18952 24639 18955
rect 24946 18952 24952 18964
rect 24627 18924 24952 18952
rect 24627 18921 24639 18924
rect 24581 18915 24639 18921
rect 24946 18912 24952 18924
rect 25004 18952 25010 18964
rect 25866 18952 25872 18964
rect 25004 18924 25872 18952
rect 25004 18912 25010 18924
rect 25866 18912 25872 18924
rect 25924 18912 25930 18964
rect 28718 18952 28724 18964
rect 28679 18924 28724 18952
rect 28718 18912 28724 18924
rect 28776 18912 28782 18964
rect 30926 18952 30932 18964
rect 30887 18924 30932 18952
rect 30926 18912 30932 18924
rect 30984 18912 30990 18964
rect 31202 18912 31208 18964
rect 31260 18952 31266 18964
rect 31481 18955 31539 18961
rect 31481 18952 31493 18955
rect 31260 18924 31493 18952
rect 31260 18912 31266 18924
rect 31481 18921 31493 18924
rect 31527 18921 31539 18955
rect 31481 18915 31539 18921
rect 22388 18816 22416 18912
rect 25130 18884 25136 18896
rect 24136 18856 25136 18884
rect 21744 18788 22416 18816
rect 1486 18708 1492 18760
rect 1544 18748 1550 18760
rect 1673 18751 1731 18757
rect 1673 18748 1685 18751
rect 1544 18720 1685 18748
rect 1544 18708 1550 18720
rect 1673 18717 1685 18720
rect 1719 18717 1731 18751
rect 1673 18711 1731 18717
rect 2409 18751 2467 18757
rect 2409 18717 2421 18751
rect 2455 18748 2467 18751
rect 16482 18748 16488 18760
rect 2455 18720 16488 18748
rect 2455 18717 2467 18720
rect 2409 18711 2467 18717
rect 16482 18708 16488 18720
rect 16540 18708 16546 18760
rect 21744 18757 21772 18788
rect 22922 18776 22928 18828
rect 22980 18816 22986 18828
rect 23290 18816 23296 18828
rect 22980 18788 23296 18816
rect 22980 18776 22986 18788
rect 23290 18776 23296 18788
rect 23348 18776 23354 18828
rect 23753 18819 23811 18825
rect 23753 18785 23765 18819
rect 23799 18816 23811 18819
rect 23842 18816 23848 18828
rect 23799 18788 23848 18816
rect 23799 18785 23811 18788
rect 23753 18779 23811 18785
rect 23842 18776 23848 18788
rect 23900 18776 23906 18828
rect 21729 18751 21787 18757
rect 21729 18717 21741 18751
rect 21775 18717 21787 18751
rect 21910 18748 21916 18760
rect 21871 18720 21916 18748
rect 21729 18711 21787 18717
rect 21910 18708 21916 18720
rect 21968 18708 21974 18760
rect 22373 18751 22431 18757
rect 22373 18717 22385 18751
rect 22419 18717 22431 18751
rect 22373 18711 22431 18717
rect 22388 18680 22416 18711
rect 22554 18708 22560 18760
rect 22612 18748 22618 18760
rect 23198 18748 23204 18760
rect 22612 18720 23204 18748
rect 22612 18708 22618 18720
rect 23198 18708 23204 18720
rect 23256 18708 23262 18760
rect 23385 18751 23443 18757
rect 23385 18717 23397 18751
rect 23431 18748 23443 18751
rect 24136 18748 24164 18856
rect 25130 18844 25136 18856
rect 25188 18844 25194 18896
rect 34238 18884 34244 18896
rect 31726 18856 34244 18884
rect 24302 18776 24308 18828
rect 24360 18816 24366 18828
rect 24762 18816 24768 18828
rect 24360 18788 24768 18816
rect 24360 18776 24366 18788
rect 24762 18776 24768 18788
rect 24820 18776 24826 18828
rect 23431 18720 24164 18748
rect 23431 18717 23443 18720
rect 23385 18711 23443 18717
rect 24210 18708 24216 18760
rect 24268 18748 24274 18760
rect 24489 18751 24547 18757
rect 24489 18748 24501 18751
rect 24268 18720 24501 18748
rect 24268 18708 24274 18720
rect 24489 18717 24501 18720
rect 24535 18717 24547 18751
rect 24489 18711 24547 18717
rect 22738 18680 22744 18692
rect 22388 18652 22744 18680
rect 22738 18640 22744 18652
rect 22796 18640 22802 18692
rect 24504 18680 24532 18711
rect 25038 18708 25044 18760
rect 25096 18748 25102 18760
rect 25225 18751 25283 18757
rect 25225 18748 25237 18751
rect 25096 18720 25237 18748
rect 25096 18708 25102 18720
rect 25225 18717 25237 18720
rect 25271 18748 25283 18751
rect 27341 18751 27399 18757
rect 27341 18748 27353 18751
rect 25271 18720 27353 18748
rect 25271 18717 25283 18720
rect 25225 18711 25283 18717
rect 27341 18717 27353 18720
rect 27387 18748 27399 18751
rect 28994 18748 29000 18760
rect 27387 18720 29000 18748
rect 27387 18717 27399 18720
rect 27341 18711 27399 18717
rect 28994 18708 29000 18720
rect 29052 18748 29058 18760
rect 29549 18751 29607 18757
rect 29549 18748 29561 18751
rect 29052 18720 29561 18748
rect 29052 18708 29058 18720
rect 29549 18717 29561 18720
rect 29595 18717 29607 18751
rect 29549 18711 29607 18717
rect 29816 18751 29874 18757
rect 29816 18717 29828 18751
rect 29862 18748 29874 18751
rect 30098 18748 30104 18760
rect 29862 18720 30104 18748
rect 29862 18717 29874 18720
rect 29816 18711 29874 18717
rect 30098 18708 30104 18720
rect 30156 18708 30162 18760
rect 31389 18751 31447 18757
rect 31389 18717 31401 18751
rect 31435 18748 31447 18751
rect 31726 18748 31754 18856
rect 34238 18844 34244 18856
rect 34296 18844 34302 18896
rect 34146 18816 34152 18828
rect 34107 18788 34152 18816
rect 34146 18776 34152 18788
rect 34204 18776 34210 18828
rect 32306 18748 32312 18760
rect 31435 18720 31754 18748
rect 32267 18720 32312 18748
rect 31435 18717 31447 18720
rect 31389 18711 31447 18717
rect 32306 18708 32312 18720
rect 32364 18708 32370 18760
rect 25498 18689 25504 18692
rect 25492 18680 25504 18689
rect 24504 18652 25360 18680
rect 25459 18652 25504 18680
rect 24765 18615 24823 18621
rect 24765 18581 24777 18615
rect 24811 18612 24823 18615
rect 24946 18612 24952 18624
rect 24811 18584 24952 18612
rect 24811 18581 24823 18584
rect 24765 18575 24823 18581
rect 24946 18572 24952 18584
rect 25004 18572 25010 18624
rect 25332 18612 25360 18652
rect 25492 18643 25504 18652
rect 25498 18640 25504 18643
rect 25556 18640 25562 18692
rect 27608 18683 27666 18689
rect 27608 18649 27620 18683
rect 27654 18680 27666 18683
rect 27890 18680 27896 18692
rect 27654 18652 27896 18680
rect 27654 18649 27666 18652
rect 27608 18643 27666 18649
rect 27890 18640 27896 18652
rect 27948 18640 27954 18692
rect 32493 18683 32551 18689
rect 32493 18649 32505 18683
rect 32539 18680 32551 18683
rect 33686 18680 33692 18692
rect 32539 18652 33692 18680
rect 32539 18649 32551 18652
rect 32493 18643 32551 18649
rect 33686 18640 33692 18652
rect 33744 18640 33750 18692
rect 26510 18612 26516 18624
rect 25332 18584 26516 18612
rect 26510 18572 26516 18584
rect 26568 18612 26574 18624
rect 26605 18615 26663 18621
rect 26605 18612 26617 18615
rect 26568 18584 26617 18612
rect 26568 18572 26574 18584
rect 26605 18581 26617 18584
rect 26651 18581 26663 18615
rect 26605 18575 26663 18581
rect 1104 18522 34868 18544
rect 1104 18470 12214 18522
rect 12266 18470 12278 18522
rect 12330 18470 12342 18522
rect 12394 18470 12406 18522
rect 12458 18470 12470 18522
rect 12522 18470 23478 18522
rect 23530 18470 23542 18522
rect 23594 18470 23606 18522
rect 23658 18470 23670 18522
rect 23722 18470 23734 18522
rect 23786 18470 34868 18522
rect 1104 18448 34868 18470
rect 21910 18368 21916 18420
rect 21968 18408 21974 18420
rect 22465 18411 22523 18417
rect 22465 18408 22477 18411
rect 21968 18380 22477 18408
rect 21968 18368 21974 18380
rect 22465 18377 22477 18380
rect 22511 18377 22523 18411
rect 22465 18371 22523 18377
rect 24581 18411 24639 18417
rect 24581 18377 24593 18411
rect 24627 18408 24639 18411
rect 25590 18408 25596 18420
rect 24627 18380 25596 18408
rect 24627 18377 24639 18380
rect 24581 18371 24639 18377
rect 25590 18368 25596 18380
rect 25648 18368 25654 18420
rect 25774 18368 25780 18420
rect 25832 18408 25838 18420
rect 26418 18408 26424 18420
rect 25832 18380 26424 18408
rect 25832 18368 25838 18380
rect 26418 18368 26424 18380
rect 26476 18368 26482 18420
rect 27522 18368 27528 18420
rect 27580 18408 27586 18420
rect 28353 18411 28411 18417
rect 28353 18408 28365 18411
rect 27580 18380 28365 18408
rect 27580 18368 27586 18380
rect 28353 18377 28365 18380
rect 28399 18377 28411 18411
rect 29638 18408 29644 18420
rect 29599 18380 29644 18408
rect 28353 18371 28411 18377
rect 29638 18368 29644 18380
rect 29696 18368 29702 18420
rect 29730 18368 29736 18420
rect 29788 18408 29794 18420
rect 30285 18411 30343 18417
rect 30285 18408 30297 18411
rect 29788 18380 30297 18408
rect 29788 18368 29794 18380
rect 30285 18377 30297 18380
rect 30331 18377 30343 18411
rect 30285 18371 30343 18377
rect 30742 18368 30748 18420
rect 30800 18408 30806 18420
rect 31481 18411 31539 18417
rect 31481 18408 31493 18411
rect 30800 18380 31493 18408
rect 30800 18368 30806 18380
rect 31481 18377 31493 18380
rect 31527 18377 31539 18411
rect 32582 18408 32588 18420
rect 32543 18380 32588 18408
rect 31481 18371 31539 18377
rect 32582 18368 32588 18380
rect 32640 18368 32646 18420
rect 33686 18408 33692 18420
rect 33647 18380 33692 18408
rect 33686 18368 33692 18380
rect 33744 18368 33750 18420
rect 23290 18340 23296 18352
rect 22388 18312 23296 18340
rect 1486 18272 1492 18284
rect 1447 18244 1492 18272
rect 1486 18232 1492 18244
rect 1544 18232 1550 18284
rect 22388 18281 22416 18312
rect 23290 18300 23296 18312
rect 23348 18300 23354 18352
rect 24854 18340 24860 18352
rect 24412 18312 24860 18340
rect 22373 18275 22431 18281
rect 22373 18241 22385 18275
rect 22419 18241 22431 18275
rect 22373 18235 22431 18241
rect 22557 18275 22615 18281
rect 22557 18241 22569 18275
rect 22603 18272 22615 18275
rect 22738 18272 22744 18284
rect 22603 18244 22744 18272
rect 22603 18241 22615 18244
rect 22557 18235 22615 18241
rect 22738 18232 22744 18244
rect 22796 18232 22802 18284
rect 23382 18232 23388 18284
rect 23440 18272 23446 18284
rect 24412 18281 24440 18312
rect 24854 18300 24860 18312
rect 24912 18300 24918 18352
rect 25056 18312 27016 18340
rect 25056 18284 25084 18312
rect 23569 18275 23627 18281
rect 23569 18272 23581 18275
rect 23440 18244 23581 18272
rect 23440 18232 23446 18244
rect 23569 18241 23581 18244
rect 23615 18241 23627 18275
rect 23569 18235 23627 18241
rect 24397 18275 24455 18281
rect 24397 18241 24409 18275
rect 24443 18241 24455 18275
rect 24397 18235 24455 18241
rect 24581 18275 24639 18281
rect 24581 18241 24593 18275
rect 24627 18272 24639 18275
rect 24670 18272 24676 18284
rect 24627 18244 24676 18272
rect 24627 18241 24639 18244
rect 24581 18235 24639 18241
rect 24670 18232 24676 18244
rect 24728 18232 24734 18284
rect 25038 18272 25044 18284
rect 24999 18244 25044 18272
rect 25038 18232 25044 18244
rect 25096 18232 25102 18284
rect 25130 18232 25136 18284
rect 25188 18272 25194 18284
rect 26988 18281 27016 18312
rect 27062 18300 27068 18352
rect 27120 18340 27126 18352
rect 27218 18343 27276 18349
rect 27218 18340 27230 18343
rect 27120 18312 27230 18340
rect 27120 18300 27126 18312
rect 27218 18309 27230 18312
rect 27264 18309 27276 18343
rect 29914 18340 29920 18352
rect 27218 18303 27276 18309
rect 29564 18312 29920 18340
rect 25297 18275 25355 18281
rect 25297 18272 25309 18275
rect 25188 18244 25309 18272
rect 25188 18232 25194 18244
rect 25297 18241 25309 18244
rect 25343 18241 25355 18275
rect 25297 18235 25355 18241
rect 26973 18275 27031 18281
rect 26973 18241 26985 18275
rect 27019 18241 27031 18275
rect 26973 18235 27031 18241
rect 28718 18232 28724 18284
rect 28776 18272 28782 18284
rect 29564 18281 29592 18312
rect 29914 18300 29920 18312
rect 29972 18300 29978 18352
rect 31110 18300 31116 18352
rect 31168 18340 31174 18352
rect 32950 18340 32956 18352
rect 31168 18312 31616 18340
rect 31168 18300 31174 18312
rect 28813 18275 28871 18281
rect 28813 18272 28825 18275
rect 28776 18244 28825 18272
rect 28776 18232 28782 18244
rect 28813 18241 28825 18244
rect 28859 18241 28871 18275
rect 28813 18235 28871 18241
rect 29549 18275 29607 18281
rect 29549 18241 29561 18275
rect 29595 18241 29607 18275
rect 29549 18235 29607 18241
rect 29733 18275 29791 18281
rect 29733 18241 29745 18275
rect 29779 18272 29791 18275
rect 30006 18272 30012 18284
rect 29779 18244 30012 18272
rect 29779 18241 29791 18244
rect 29733 18235 29791 18241
rect 30006 18232 30012 18244
rect 30064 18232 30070 18284
rect 30193 18275 30251 18281
rect 30193 18241 30205 18275
rect 30239 18241 30251 18275
rect 30374 18272 30380 18284
rect 30335 18244 30380 18272
rect 30193 18235 30251 18241
rect 1670 18204 1676 18216
rect 1631 18176 1676 18204
rect 1670 18164 1676 18176
rect 1728 18164 1734 18216
rect 2866 18204 2872 18216
rect 2827 18176 2872 18204
rect 2866 18164 2872 18176
rect 2924 18164 2930 18216
rect 23661 18207 23719 18213
rect 23661 18173 23673 18207
rect 23707 18204 23719 18207
rect 23842 18204 23848 18216
rect 23707 18176 23848 18204
rect 23707 18173 23719 18176
rect 23661 18167 23719 18173
rect 23842 18164 23848 18176
rect 23900 18164 23906 18216
rect 29089 18207 29147 18213
rect 29089 18173 29101 18207
rect 29135 18173 29147 18207
rect 30208 18204 30236 18235
rect 30374 18232 30380 18244
rect 30432 18232 30438 18284
rect 31386 18272 31392 18284
rect 31347 18244 31392 18272
rect 31386 18232 31392 18244
rect 31444 18232 31450 18284
rect 31588 18281 31616 18312
rect 32508 18312 32956 18340
rect 32508 18284 32536 18312
rect 32950 18300 32956 18312
rect 33008 18300 33014 18352
rect 31573 18275 31631 18281
rect 31573 18241 31585 18275
rect 31619 18241 31631 18275
rect 32490 18272 32496 18284
rect 32403 18244 32496 18272
rect 31573 18235 31631 18241
rect 32490 18232 32496 18244
rect 32548 18232 32554 18284
rect 32674 18232 32680 18284
rect 32732 18272 32738 18284
rect 33594 18272 33600 18284
rect 32732 18244 33600 18272
rect 32732 18232 32738 18244
rect 33594 18232 33600 18244
rect 33652 18232 33658 18284
rect 31662 18204 31668 18216
rect 30208 18176 31668 18204
rect 29089 18167 29147 18173
rect 23937 18139 23995 18145
rect 23937 18105 23949 18139
rect 23983 18136 23995 18139
rect 24854 18136 24860 18148
rect 23983 18108 24860 18136
rect 23983 18105 23995 18108
rect 23937 18099 23995 18105
rect 24854 18096 24860 18108
rect 24912 18096 24918 18148
rect 29104 18136 29132 18167
rect 31662 18164 31668 18176
rect 31720 18164 31726 18216
rect 30650 18136 30656 18148
rect 29104 18108 30656 18136
rect 30650 18096 30656 18108
rect 30708 18096 30714 18148
rect 28810 18028 28816 18080
rect 28868 18068 28874 18080
rect 28905 18071 28963 18077
rect 28905 18068 28917 18071
rect 28868 18040 28917 18068
rect 28868 18028 28874 18040
rect 28905 18037 28917 18040
rect 28951 18037 28963 18071
rect 28905 18031 28963 18037
rect 28994 18028 29000 18080
rect 29052 18068 29058 18080
rect 29052 18040 29097 18068
rect 29052 18028 29058 18040
rect 1104 17978 34868 18000
rect 1104 17926 6582 17978
rect 6634 17926 6646 17978
rect 6698 17926 6710 17978
rect 6762 17926 6774 17978
rect 6826 17926 6838 17978
rect 6890 17926 17846 17978
rect 17898 17926 17910 17978
rect 17962 17926 17974 17978
rect 18026 17926 18038 17978
rect 18090 17926 18102 17978
rect 18154 17926 29110 17978
rect 29162 17926 29174 17978
rect 29226 17926 29238 17978
rect 29290 17926 29302 17978
rect 29354 17926 29366 17978
rect 29418 17926 34868 17978
rect 1104 17904 34868 17926
rect 1670 17824 1676 17876
rect 1728 17864 1734 17876
rect 1857 17867 1915 17873
rect 1857 17864 1869 17867
rect 1728 17836 1869 17864
rect 1728 17824 1734 17836
rect 1857 17833 1869 17836
rect 1903 17833 1915 17867
rect 1857 17827 1915 17833
rect 24949 17867 25007 17873
rect 24949 17833 24961 17867
rect 24995 17864 25007 17867
rect 25498 17864 25504 17876
rect 24995 17836 25504 17864
rect 24995 17833 25007 17836
rect 24949 17827 25007 17833
rect 25498 17824 25504 17836
rect 25556 17824 25562 17876
rect 25777 17867 25835 17873
rect 25777 17833 25789 17867
rect 25823 17864 25835 17867
rect 25866 17864 25872 17876
rect 25823 17836 25872 17864
rect 25823 17833 25835 17836
rect 25777 17827 25835 17833
rect 25866 17824 25872 17836
rect 25924 17824 25930 17876
rect 26513 17867 26571 17873
rect 26513 17833 26525 17867
rect 26559 17864 26571 17867
rect 26878 17864 26884 17876
rect 26559 17836 26884 17864
rect 26559 17833 26571 17836
rect 26513 17827 26571 17833
rect 26878 17824 26884 17836
rect 26936 17824 26942 17876
rect 27246 17824 27252 17876
rect 27304 17864 27310 17876
rect 27341 17867 27399 17873
rect 27341 17864 27353 17867
rect 27304 17836 27353 17864
rect 27304 17824 27310 17836
rect 27341 17833 27353 17836
rect 27387 17833 27399 17867
rect 28534 17864 28540 17876
rect 28495 17836 28540 17864
rect 27341 17827 27399 17833
rect 28534 17824 28540 17836
rect 28592 17824 28598 17876
rect 28902 17824 28908 17876
rect 28960 17864 28966 17876
rect 30101 17867 30159 17873
rect 30101 17864 30113 17867
rect 28960 17836 30113 17864
rect 28960 17824 28966 17836
rect 30101 17833 30113 17836
rect 30147 17833 30159 17867
rect 30101 17827 30159 17833
rect 31205 17867 31263 17873
rect 31205 17833 31217 17867
rect 31251 17864 31263 17867
rect 31478 17864 31484 17876
rect 31251 17836 31484 17864
rect 31251 17833 31263 17836
rect 31205 17827 31263 17833
rect 31478 17824 31484 17836
rect 31536 17824 31542 17876
rect 24486 17756 24492 17808
rect 24544 17796 24550 17808
rect 30561 17799 30619 17805
rect 30561 17796 30573 17799
rect 24544 17768 30573 17796
rect 24544 17756 24550 17768
rect 30561 17765 30573 17768
rect 30607 17765 30619 17799
rect 30561 17759 30619 17765
rect 1854 17688 1860 17740
rect 1912 17728 1918 17740
rect 4798 17728 4804 17740
rect 1912 17700 4804 17728
rect 1912 17688 1918 17700
rect 4798 17688 4804 17700
rect 4856 17688 4862 17740
rect 24762 17688 24768 17740
rect 24820 17728 24826 17740
rect 25961 17731 26019 17737
rect 25961 17728 25973 17731
rect 24820 17700 25973 17728
rect 24820 17688 24826 17700
rect 25961 17697 25973 17700
rect 26007 17697 26019 17731
rect 30374 17728 30380 17740
rect 25961 17691 26019 17697
rect 28736 17700 30380 17728
rect 1762 17660 1768 17672
rect 1723 17632 1768 17660
rect 1762 17620 1768 17632
rect 1820 17620 1826 17672
rect 24946 17660 24952 17672
rect 24907 17632 24952 17660
rect 24946 17620 24952 17632
rect 25004 17620 25010 17672
rect 25222 17660 25228 17672
rect 25183 17632 25228 17660
rect 25222 17620 25228 17632
rect 25280 17620 25286 17672
rect 25685 17663 25743 17669
rect 25685 17629 25697 17663
rect 25731 17660 25743 17663
rect 25774 17660 25780 17672
rect 25731 17632 25780 17660
rect 25731 17629 25743 17632
rect 25685 17623 25743 17629
rect 25774 17620 25780 17632
rect 25832 17620 25838 17672
rect 26421 17663 26479 17669
rect 26421 17629 26433 17663
rect 26467 17629 26479 17663
rect 27522 17660 27528 17672
rect 27483 17632 27528 17660
rect 26421 17623 26479 17629
rect 25038 17552 25044 17604
rect 25096 17592 25102 17604
rect 25133 17595 25191 17601
rect 25133 17592 25145 17595
rect 25096 17564 25145 17592
rect 25096 17552 25102 17564
rect 25133 17561 25145 17564
rect 25179 17592 25191 17595
rect 25406 17592 25412 17604
rect 25179 17564 25412 17592
rect 25179 17561 25191 17564
rect 25133 17555 25191 17561
rect 25406 17552 25412 17564
rect 25464 17552 25470 17604
rect 26436 17592 26464 17623
rect 27522 17620 27528 17632
rect 27580 17620 27586 17672
rect 27617 17663 27675 17669
rect 27617 17629 27629 17663
rect 27663 17660 27675 17663
rect 27706 17660 27712 17672
rect 27663 17632 27712 17660
rect 27663 17629 27675 17632
rect 27617 17623 27675 17629
rect 27706 17620 27712 17632
rect 27764 17620 27770 17672
rect 28736 17669 28764 17700
rect 30374 17688 30380 17700
rect 30432 17688 30438 17740
rect 32490 17728 32496 17740
rect 30760 17700 32496 17728
rect 28537 17663 28595 17669
rect 28537 17629 28549 17663
rect 28583 17629 28595 17663
rect 28537 17623 28595 17629
rect 28721 17663 28779 17669
rect 28721 17629 28733 17663
rect 28767 17629 28779 17663
rect 30190 17660 30196 17672
rect 28721 17623 28779 17629
rect 29380 17632 30196 17660
rect 25516 17564 26464 17592
rect 27341 17595 27399 17601
rect 24578 17484 24584 17536
rect 24636 17524 24642 17536
rect 25516 17524 25544 17564
rect 27341 17561 27353 17595
rect 27387 17592 27399 17595
rect 28442 17592 28448 17604
rect 27387 17564 28448 17592
rect 27387 17561 27399 17564
rect 27341 17555 27399 17561
rect 28442 17552 28448 17564
rect 28500 17552 28506 17604
rect 28552 17592 28580 17623
rect 29380 17592 29408 17632
rect 30190 17620 30196 17632
rect 30248 17620 30254 17672
rect 30558 17660 30564 17672
rect 30519 17632 30564 17660
rect 30558 17620 30564 17632
rect 30616 17620 30622 17672
rect 30760 17669 30788 17700
rect 32490 17688 32496 17700
rect 32548 17688 32554 17740
rect 34146 17728 34152 17740
rect 34107 17700 34152 17728
rect 34146 17688 34152 17700
rect 34204 17688 34210 17740
rect 30745 17663 30803 17669
rect 30745 17629 30757 17663
rect 30791 17629 30803 17663
rect 30745 17623 30803 17629
rect 31205 17663 31263 17669
rect 31205 17629 31217 17663
rect 31251 17629 31263 17663
rect 31205 17623 31263 17629
rect 31389 17663 31447 17669
rect 31389 17629 31401 17663
rect 31435 17660 31447 17663
rect 31435 17632 31754 17660
rect 31435 17629 31447 17632
rect 31389 17623 31447 17629
rect 28552 17564 29408 17592
rect 29454 17552 29460 17604
rect 29512 17592 29518 17604
rect 31220 17592 31248 17623
rect 29512 17564 31248 17592
rect 29512 17552 29518 17564
rect 25958 17524 25964 17536
rect 24636 17496 25544 17524
rect 25919 17496 25964 17524
rect 24636 17484 24642 17496
rect 25958 17484 25964 17496
rect 26016 17484 26022 17536
rect 29546 17484 29552 17536
rect 29604 17524 29610 17536
rect 31478 17524 31484 17536
rect 29604 17496 31484 17524
rect 29604 17484 29610 17496
rect 31478 17484 31484 17496
rect 31536 17484 31542 17536
rect 31726 17524 31754 17632
rect 31938 17620 31944 17672
rect 31996 17660 32002 17672
rect 32309 17663 32367 17669
rect 32309 17660 32321 17663
rect 31996 17632 32321 17660
rect 31996 17620 32002 17632
rect 32309 17629 32321 17632
rect 32355 17629 32367 17663
rect 32309 17623 32367 17629
rect 32493 17595 32551 17601
rect 32493 17561 32505 17595
rect 32539 17592 32551 17595
rect 33778 17592 33784 17604
rect 32539 17564 33784 17592
rect 32539 17561 32551 17564
rect 32493 17555 32551 17561
rect 33778 17552 33784 17564
rect 33836 17552 33842 17604
rect 32398 17524 32404 17536
rect 31726 17496 32404 17524
rect 32398 17484 32404 17496
rect 32456 17484 32462 17536
rect 1104 17434 34868 17456
rect 1104 17382 12214 17434
rect 12266 17382 12278 17434
rect 12330 17382 12342 17434
rect 12394 17382 12406 17434
rect 12458 17382 12470 17434
rect 12522 17382 23478 17434
rect 23530 17382 23542 17434
rect 23594 17382 23606 17434
rect 23658 17382 23670 17434
rect 23722 17382 23734 17434
rect 23786 17382 34868 17434
rect 1104 17360 34868 17382
rect 5074 17280 5080 17332
rect 5132 17320 5138 17332
rect 24857 17323 24915 17329
rect 5132 17292 24624 17320
rect 5132 17280 5138 17292
rect 1489 17119 1547 17125
rect 1489 17085 1501 17119
rect 1535 17085 1547 17119
rect 1670 17116 1676 17128
rect 1631 17088 1676 17116
rect 1489 17079 1547 17085
rect 1504 17048 1532 17079
rect 1670 17076 1676 17088
rect 1728 17076 1734 17128
rect 1946 17116 1952 17128
rect 1907 17088 1952 17116
rect 1946 17076 1952 17088
rect 2004 17076 2010 17128
rect 12894 17076 12900 17128
rect 12952 17116 12958 17128
rect 24486 17116 24492 17128
rect 12952 17088 24492 17116
rect 12952 17076 12958 17088
rect 24486 17076 24492 17088
rect 24544 17076 24550 17128
rect 24596 17116 24624 17292
rect 24857 17289 24869 17323
rect 24903 17320 24915 17323
rect 25038 17320 25044 17332
rect 24903 17292 25044 17320
rect 24903 17289 24915 17292
rect 24857 17283 24915 17289
rect 25038 17280 25044 17292
rect 25096 17280 25102 17332
rect 25314 17280 25320 17332
rect 25372 17320 25378 17332
rect 25501 17323 25559 17329
rect 25501 17320 25513 17323
rect 25372 17292 25513 17320
rect 25372 17280 25378 17292
rect 25501 17289 25513 17292
rect 25547 17289 25559 17323
rect 27890 17320 27896 17332
rect 27851 17292 27896 17320
rect 25501 17283 25559 17289
rect 27890 17280 27896 17292
rect 27948 17280 27954 17332
rect 30466 17280 30472 17332
rect 30524 17320 30530 17332
rect 31481 17323 31539 17329
rect 31481 17320 31493 17323
rect 30524 17292 31493 17320
rect 30524 17280 30530 17292
rect 31481 17289 31493 17292
rect 31527 17289 31539 17323
rect 31481 17283 31539 17289
rect 24673 17255 24731 17261
rect 24673 17221 24685 17255
rect 24719 17252 24731 17255
rect 25958 17252 25964 17264
rect 24719 17224 25964 17252
rect 24719 17221 24731 17224
rect 24673 17215 24731 17221
rect 25958 17212 25964 17224
rect 26016 17212 26022 17264
rect 28994 17252 29000 17264
rect 27816 17224 29000 17252
rect 24946 17144 24952 17196
rect 25004 17184 25010 17196
rect 25004 17156 25049 17184
rect 25004 17144 25010 17156
rect 25406 17144 25412 17196
rect 25464 17184 25470 17196
rect 25593 17187 25651 17193
rect 25464 17156 25509 17184
rect 25464 17144 25470 17156
rect 25593 17153 25605 17187
rect 25639 17184 25651 17187
rect 25682 17184 25688 17196
rect 25639 17156 25688 17184
rect 25639 17153 25651 17156
rect 25593 17147 25651 17153
rect 25682 17144 25688 17156
rect 25740 17144 25746 17196
rect 27816 17193 27844 17224
rect 28994 17212 29000 17224
rect 29052 17212 29058 17264
rect 32306 17252 32312 17264
rect 30944 17224 32312 17252
rect 27801 17187 27859 17193
rect 27801 17153 27813 17187
rect 27847 17153 27859 17187
rect 27801 17147 27859 17153
rect 27985 17187 28043 17193
rect 27985 17153 27997 17187
rect 28031 17153 28043 17187
rect 30282 17184 30288 17196
rect 30243 17156 30288 17184
rect 27985 17147 28043 17153
rect 24596 17088 25268 17116
rect 2590 17048 2596 17060
rect 1504 17020 2596 17048
rect 2590 17008 2596 17020
rect 2648 17008 2654 17060
rect 24673 17051 24731 17057
rect 24673 17017 24685 17051
rect 24719 17048 24731 17051
rect 25130 17048 25136 17060
rect 24719 17020 25136 17048
rect 24719 17017 24731 17020
rect 24673 17011 24731 17017
rect 25130 17008 25136 17020
rect 25188 17008 25194 17060
rect 25240 17048 25268 17088
rect 27706 17076 27712 17128
rect 27764 17116 27770 17128
rect 28000 17116 28028 17147
rect 30282 17144 30288 17156
rect 30340 17144 30346 17196
rect 30944 17193 30972 17224
rect 32306 17212 32312 17224
rect 32364 17212 32370 17264
rect 30929 17187 30987 17193
rect 30929 17153 30941 17187
rect 30975 17153 30987 17187
rect 30929 17147 30987 17153
rect 31294 17144 31300 17196
rect 31352 17184 31358 17196
rect 31389 17187 31447 17193
rect 31389 17184 31401 17187
rect 31352 17156 31401 17184
rect 31352 17144 31358 17156
rect 31389 17153 31401 17156
rect 31435 17153 31447 17187
rect 31389 17147 31447 17153
rect 31478 17144 31484 17196
rect 31536 17184 31542 17196
rect 31573 17187 31631 17193
rect 31573 17184 31585 17187
rect 31536 17156 31585 17184
rect 31536 17144 31542 17156
rect 31573 17153 31585 17156
rect 31619 17153 31631 17187
rect 31846 17184 31852 17196
rect 31573 17147 31631 17153
rect 31726 17156 31852 17184
rect 27764 17088 28028 17116
rect 29641 17119 29699 17125
rect 27764 17076 27770 17088
rect 29641 17085 29653 17119
rect 29687 17116 29699 17119
rect 31726 17116 31754 17156
rect 31846 17144 31852 17156
rect 31904 17144 31910 17196
rect 29687 17088 31754 17116
rect 29687 17085 29699 17088
rect 29641 17079 29699 17085
rect 32030 17076 32036 17128
rect 32088 17116 32094 17128
rect 32309 17119 32367 17125
rect 32309 17116 32321 17119
rect 32088 17088 32321 17116
rect 32088 17076 32094 17088
rect 32309 17085 32321 17088
rect 32355 17085 32367 17119
rect 32309 17079 32367 17085
rect 32493 17119 32551 17125
rect 32493 17085 32505 17119
rect 32539 17116 32551 17119
rect 33134 17116 33140 17128
rect 32539 17088 33140 17116
rect 32539 17085 32551 17088
rect 32493 17079 32551 17085
rect 33134 17076 33140 17088
rect 33192 17076 33198 17128
rect 34146 17116 34152 17128
rect 34107 17088 34152 17116
rect 34146 17076 34152 17088
rect 34204 17076 34210 17128
rect 32950 17048 32956 17060
rect 25240 17020 32956 17048
rect 32950 17008 32956 17020
rect 33008 17008 33014 17060
rect 31662 16940 31668 16992
rect 31720 16980 31726 16992
rect 33410 16980 33416 16992
rect 31720 16952 33416 16980
rect 31720 16940 31726 16952
rect 33410 16940 33416 16952
rect 33468 16940 33474 16992
rect 1104 16890 34868 16912
rect 1104 16838 6582 16890
rect 6634 16838 6646 16890
rect 6698 16838 6710 16890
rect 6762 16838 6774 16890
rect 6826 16838 6838 16890
rect 6890 16838 17846 16890
rect 17898 16838 17910 16890
rect 17962 16838 17974 16890
rect 18026 16838 18038 16890
rect 18090 16838 18102 16890
rect 18154 16838 29110 16890
rect 29162 16838 29174 16890
rect 29226 16838 29238 16890
rect 29290 16838 29302 16890
rect 29354 16838 29366 16890
rect 29418 16838 34868 16890
rect 1104 16816 34868 16838
rect 1670 16736 1676 16788
rect 1728 16776 1734 16788
rect 1857 16779 1915 16785
rect 1857 16776 1869 16779
rect 1728 16748 1869 16776
rect 1728 16736 1734 16748
rect 1857 16745 1869 16748
rect 1903 16745 1915 16779
rect 2590 16776 2596 16788
rect 2551 16748 2596 16776
rect 1857 16739 1915 16745
rect 2590 16736 2596 16748
rect 2648 16736 2654 16788
rect 31018 16776 31024 16788
rect 30979 16748 31024 16776
rect 31018 16736 31024 16748
rect 31076 16736 31082 16788
rect 31665 16779 31723 16785
rect 31665 16745 31677 16779
rect 31711 16776 31723 16779
rect 32306 16776 32312 16788
rect 31711 16748 32312 16776
rect 31711 16745 31723 16748
rect 31665 16739 31723 16745
rect 32306 16736 32312 16748
rect 32364 16736 32370 16788
rect 30377 16711 30435 16717
rect 30377 16677 30389 16711
rect 30423 16708 30435 16711
rect 34514 16708 34520 16720
rect 30423 16680 34520 16708
rect 30423 16677 30435 16680
rect 30377 16671 30435 16677
rect 34514 16668 34520 16680
rect 34572 16668 34578 16720
rect 1670 16600 1676 16652
rect 1728 16640 1734 16652
rect 1854 16640 1860 16652
rect 1728 16612 1860 16640
rect 1728 16600 1734 16612
rect 1780 16581 1808 16612
rect 1854 16600 1860 16612
rect 1912 16600 1918 16652
rect 30098 16600 30104 16652
rect 30156 16640 30162 16652
rect 31662 16640 31668 16652
rect 30156 16612 31668 16640
rect 30156 16600 30162 16612
rect 31662 16600 31668 16612
rect 31720 16600 31726 16652
rect 32858 16640 32864 16652
rect 32140 16612 32864 16640
rect 32140 16581 32168 16612
rect 32858 16600 32864 16612
rect 32916 16600 32922 16652
rect 32950 16600 32956 16652
rect 33008 16640 33014 16652
rect 33008 16612 33088 16640
rect 33008 16600 33014 16612
rect 1765 16575 1823 16581
rect 1765 16541 1777 16575
rect 1811 16541 1823 16575
rect 1765 16535 1823 16541
rect 32125 16575 32183 16581
rect 32125 16541 32137 16575
rect 32171 16541 32183 16575
rect 32125 16535 32183 16541
rect 32309 16575 32367 16581
rect 32309 16541 32321 16575
rect 32355 16572 32367 16575
rect 32398 16572 32404 16584
rect 32355 16544 32404 16572
rect 32355 16541 32367 16544
rect 32309 16535 32367 16541
rect 32398 16532 32404 16544
rect 32456 16532 32462 16584
rect 33060 16581 33088 16612
rect 33410 16600 33416 16652
rect 33468 16640 33474 16652
rect 33468 16612 33732 16640
rect 33468 16600 33474 16612
rect 33045 16575 33103 16581
rect 33045 16541 33057 16575
rect 33091 16541 33103 16575
rect 33045 16535 33103 16541
rect 33134 16532 33140 16584
rect 33192 16572 33198 16584
rect 33704 16581 33732 16612
rect 33689 16575 33747 16581
rect 33192 16544 33237 16572
rect 33192 16532 33198 16544
rect 33689 16541 33701 16575
rect 33735 16541 33747 16575
rect 33689 16535 33747 16541
rect 33778 16532 33784 16584
rect 33836 16572 33842 16584
rect 33836 16544 33881 16572
rect 33836 16532 33842 16544
rect 32122 16396 32128 16448
rect 32180 16436 32186 16448
rect 32217 16439 32275 16445
rect 32217 16436 32229 16439
rect 32180 16408 32229 16436
rect 32180 16396 32186 16408
rect 32217 16405 32229 16408
rect 32263 16405 32275 16439
rect 32217 16399 32275 16405
rect 1104 16346 34868 16368
rect 1104 16294 12214 16346
rect 12266 16294 12278 16346
rect 12330 16294 12342 16346
rect 12394 16294 12406 16346
rect 12458 16294 12470 16346
rect 12522 16294 23478 16346
rect 23530 16294 23542 16346
rect 23594 16294 23606 16346
rect 23658 16294 23670 16346
rect 23722 16294 23734 16346
rect 23786 16294 34868 16346
rect 1104 16272 34868 16294
rect 34146 16164 34152 16176
rect 34107 16136 34152 16164
rect 34146 16124 34152 16136
rect 34204 16124 34210 16176
rect 31573 16099 31631 16105
rect 31573 16065 31585 16099
rect 31619 16096 31631 16099
rect 31938 16096 31944 16108
rect 31619 16068 31944 16096
rect 31619 16065 31631 16068
rect 31573 16059 31631 16065
rect 31938 16056 31944 16068
rect 31996 16056 32002 16108
rect 32306 16096 32312 16108
rect 32267 16068 32312 16096
rect 32306 16056 32312 16068
rect 32364 16056 32370 16108
rect 30929 16031 30987 16037
rect 30929 15997 30941 16031
rect 30975 16028 30987 16031
rect 32030 16028 32036 16040
rect 30975 16000 32036 16028
rect 30975 15997 30987 16000
rect 30929 15991 30987 15997
rect 32030 15988 32036 16000
rect 32088 15988 32094 16040
rect 32493 16031 32551 16037
rect 32493 15997 32505 16031
rect 32539 16028 32551 16031
rect 33686 16028 33692 16040
rect 32539 16000 33692 16028
rect 32539 15997 32551 16000
rect 32493 15991 32551 15997
rect 33686 15988 33692 16000
rect 33744 15988 33750 16040
rect 1394 15852 1400 15904
rect 1452 15892 1458 15904
rect 1857 15895 1915 15901
rect 1857 15892 1869 15895
rect 1452 15864 1869 15892
rect 1452 15852 1458 15864
rect 1857 15861 1869 15864
rect 1903 15861 1915 15895
rect 1857 15855 1915 15861
rect 1104 15802 34868 15824
rect 1104 15750 6582 15802
rect 6634 15750 6646 15802
rect 6698 15750 6710 15802
rect 6762 15750 6774 15802
rect 6826 15750 6838 15802
rect 6890 15750 17846 15802
rect 17898 15750 17910 15802
rect 17962 15750 17974 15802
rect 18026 15750 18038 15802
rect 18090 15750 18102 15802
rect 18154 15750 29110 15802
rect 29162 15750 29174 15802
rect 29226 15750 29238 15802
rect 29290 15750 29302 15802
rect 29354 15750 29366 15802
rect 29418 15750 34868 15802
rect 1104 15728 34868 15750
rect 33686 15688 33692 15700
rect 33647 15660 33692 15688
rect 33686 15648 33692 15660
rect 33744 15648 33750 15700
rect 33137 15623 33195 15629
rect 33137 15589 33149 15623
rect 33183 15620 33195 15623
rect 34422 15620 34428 15632
rect 33183 15592 34428 15620
rect 33183 15589 33195 15592
rect 33137 15583 33195 15589
rect 34422 15580 34428 15592
rect 34480 15580 34486 15632
rect 1394 15552 1400 15564
rect 1355 15524 1400 15552
rect 1394 15512 1400 15524
rect 1452 15512 1458 15564
rect 2774 15552 2780 15564
rect 2735 15524 2780 15552
rect 2774 15512 2780 15524
rect 2832 15512 2838 15564
rect 33594 15484 33600 15496
rect 33555 15456 33600 15484
rect 33594 15444 33600 15456
rect 33652 15444 33658 15496
rect 1578 15416 1584 15428
rect 1539 15388 1584 15416
rect 1578 15376 1584 15388
rect 1636 15376 1642 15428
rect 1104 15258 34868 15280
rect 1104 15206 12214 15258
rect 12266 15206 12278 15258
rect 12330 15206 12342 15258
rect 12394 15206 12406 15258
rect 12458 15206 12470 15258
rect 12522 15206 23478 15258
rect 23530 15206 23542 15258
rect 23594 15206 23606 15258
rect 23658 15206 23670 15258
rect 23722 15206 23734 15258
rect 23786 15206 34868 15258
rect 1104 15184 34868 15206
rect 1578 15104 1584 15156
rect 1636 15144 1642 15156
rect 2041 15147 2099 15153
rect 2041 15144 2053 15147
rect 1636 15116 2053 15144
rect 1636 15104 1642 15116
rect 2041 15113 2053 15116
rect 2087 15113 2099 15147
rect 2041 15107 2099 15113
rect 1949 15011 2007 15017
rect 1949 14977 1961 15011
rect 1995 15008 2007 15011
rect 2222 15008 2228 15020
rect 1995 14980 2228 15008
rect 1995 14977 2007 14980
rect 1949 14971 2007 14977
rect 2222 14968 2228 14980
rect 2280 14968 2286 15020
rect 32950 14968 32956 15020
rect 33008 15008 33014 15020
rect 33045 15011 33103 15017
rect 33045 15008 33057 15011
rect 33008 14980 33057 15008
rect 33008 14968 33014 14980
rect 33045 14977 33057 14980
rect 33091 15008 33103 15011
rect 33689 15011 33747 15017
rect 33689 15008 33701 15011
rect 33091 14980 33701 15008
rect 33091 14977 33103 14980
rect 33045 14971 33103 14977
rect 33689 14977 33701 14980
rect 33735 14977 33747 15011
rect 33689 14971 33747 14977
rect 1394 14764 1400 14816
rect 1452 14804 1458 14816
rect 2777 14807 2835 14813
rect 2777 14804 2789 14807
rect 1452 14776 2789 14804
rect 1452 14764 1458 14776
rect 2777 14773 2789 14776
rect 2823 14773 2835 14807
rect 2777 14767 2835 14773
rect 32306 14764 32312 14816
rect 32364 14804 32370 14816
rect 32585 14807 32643 14813
rect 32585 14804 32597 14807
rect 32364 14776 32597 14804
rect 32364 14764 32370 14776
rect 32585 14773 32597 14776
rect 32631 14773 32643 14807
rect 33134 14804 33140 14816
rect 33095 14776 33140 14804
rect 32585 14767 32643 14773
rect 33134 14764 33140 14776
rect 33192 14764 33198 14816
rect 33778 14804 33784 14816
rect 33739 14776 33784 14804
rect 33778 14764 33784 14776
rect 33836 14764 33842 14816
rect 1104 14714 34868 14736
rect 1104 14662 6582 14714
rect 6634 14662 6646 14714
rect 6698 14662 6710 14714
rect 6762 14662 6774 14714
rect 6826 14662 6838 14714
rect 6890 14662 17846 14714
rect 17898 14662 17910 14714
rect 17962 14662 17974 14714
rect 18026 14662 18038 14714
rect 18090 14662 18102 14714
rect 18154 14662 29110 14714
rect 29162 14662 29174 14714
rect 29226 14662 29238 14714
rect 29290 14662 29302 14714
rect 29354 14662 29366 14714
rect 29418 14662 34868 14714
rect 1104 14640 34868 14662
rect 1394 14464 1400 14476
rect 1355 14436 1400 14464
rect 1394 14424 1400 14436
rect 1452 14424 1458 14476
rect 1946 14464 1952 14476
rect 1907 14436 1952 14464
rect 1946 14424 1952 14436
rect 2004 14424 2010 14476
rect 32306 14464 32312 14476
rect 32267 14436 32312 14464
rect 32306 14424 32312 14436
rect 32364 14424 32370 14476
rect 32493 14467 32551 14473
rect 32493 14433 32505 14467
rect 32539 14464 32551 14467
rect 33134 14464 33140 14476
rect 32539 14436 33140 14464
rect 32539 14433 32551 14436
rect 32493 14427 32551 14433
rect 33134 14424 33140 14436
rect 33192 14424 33198 14476
rect 1581 14331 1639 14337
rect 1581 14297 1593 14331
rect 1627 14328 1639 14331
rect 1854 14328 1860 14340
rect 1627 14300 1860 14328
rect 1627 14297 1639 14300
rect 1581 14291 1639 14297
rect 1854 14288 1860 14300
rect 1912 14288 1918 14340
rect 34146 14328 34152 14340
rect 34107 14300 34152 14328
rect 34146 14288 34152 14300
rect 34204 14288 34210 14340
rect 1104 14170 34868 14192
rect 1104 14118 12214 14170
rect 12266 14118 12278 14170
rect 12330 14118 12342 14170
rect 12394 14118 12406 14170
rect 12458 14118 12470 14170
rect 12522 14118 23478 14170
rect 23530 14118 23542 14170
rect 23594 14118 23606 14170
rect 23658 14118 23670 14170
rect 23722 14118 23734 14170
rect 23786 14118 34868 14170
rect 1104 14096 34868 14118
rect 1854 14056 1860 14068
rect 1815 14028 1860 14056
rect 1854 14016 1860 14028
rect 1912 14016 1918 14068
rect 32493 13991 32551 13997
rect 32493 13957 32505 13991
rect 32539 13988 32551 13991
rect 33778 13988 33784 14000
rect 32539 13960 33784 13988
rect 32539 13957 32551 13960
rect 32493 13951 32551 13957
rect 33778 13948 33784 13960
rect 33836 13948 33842 14000
rect 1670 13880 1676 13932
rect 1728 13920 1734 13932
rect 1765 13923 1823 13929
rect 1765 13920 1777 13923
rect 1728 13892 1777 13920
rect 1728 13880 1734 13892
rect 1765 13889 1777 13892
rect 1811 13920 1823 13923
rect 1854 13920 1860 13932
rect 1811 13892 1860 13920
rect 1811 13889 1823 13892
rect 1765 13883 1823 13889
rect 1854 13880 1860 13892
rect 1912 13880 1918 13932
rect 2593 13923 2651 13929
rect 2593 13889 2605 13923
rect 2639 13920 2651 13923
rect 3050 13920 3056 13932
rect 2639 13892 3056 13920
rect 2639 13889 2651 13892
rect 2593 13883 2651 13889
rect 3050 13880 3056 13892
rect 3108 13920 3114 13932
rect 7926 13920 7932 13932
rect 3108 13892 7932 13920
rect 3108 13880 3114 13892
rect 7926 13880 7932 13892
rect 7984 13880 7990 13932
rect 31573 13855 31631 13861
rect 31573 13821 31585 13855
rect 31619 13852 31631 13855
rect 32309 13855 32367 13861
rect 32309 13852 32321 13855
rect 31619 13824 32321 13852
rect 31619 13821 31631 13824
rect 31573 13815 31631 13821
rect 32309 13821 32321 13824
rect 32355 13821 32367 13855
rect 34146 13852 34152 13864
rect 34107 13824 34152 13852
rect 32309 13815 32367 13821
rect 34146 13812 34152 13824
rect 34204 13812 34210 13864
rect 1578 13676 1584 13728
rect 1636 13716 1642 13728
rect 2685 13719 2743 13725
rect 2685 13716 2697 13719
rect 1636 13688 2697 13716
rect 1636 13676 1642 13688
rect 2685 13685 2697 13688
rect 2731 13685 2743 13719
rect 3418 13716 3424 13728
rect 3379 13688 3424 13716
rect 2685 13679 2743 13685
rect 3418 13676 3424 13688
rect 3476 13676 3482 13728
rect 1104 13626 34868 13648
rect 1104 13574 6582 13626
rect 6634 13574 6646 13626
rect 6698 13574 6710 13626
rect 6762 13574 6774 13626
rect 6826 13574 6838 13626
rect 6890 13574 17846 13626
rect 17898 13574 17910 13626
rect 17962 13574 17974 13626
rect 18026 13574 18038 13626
rect 18090 13574 18102 13626
rect 18154 13574 29110 13626
rect 29162 13574 29174 13626
rect 29226 13574 29238 13626
rect 29290 13574 29302 13626
rect 29354 13574 29366 13626
rect 29418 13574 34868 13626
rect 1104 13552 34868 13574
rect 3418 13444 3424 13456
rect 1412 13416 3424 13444
rect 1412 13385 1440 13416
rect 3418 13404 3424 13416
rect 3476 13404 3482 13456
rect 1397 13379 1455 13385
rect 1397 13345 1409 13379
rect 1443 13345 1455 13379
rect 1578 13376 1584 13388
rect 1539 13348 1584 13376
rect 1397 13339 1455 13345
rect 1578 13336 1584 13348
rect 1636 13336 1642 13388
rect 2774 13376 2780 13388
rect 2735 13348 2780 13376
rect 2774 13336 2780 13348
rect 2832 13336 2838 13388
rect 32306 13268 32312 13320
rect 32364 13308 32370 13320
rect 32493 13311 32551 13317
rect 32493 13308 32505 13311
rect 32364 13280 32505 13308
rect 32364 13268 32370 13280
rect 32493 13277 32505 13280
rect 32539 13277 32551 13311
rect 33134 13308 33140 13320
rect 33095 13280 33140 13308
rect 32493 13271 32551 13277
rect 33134 13268 33140 13280
rect 33192 13268 33198 13320
rect 33410 13268 33416 13320
rect 33468 13308 33474 13320
rect 33597 13311 33655 13317
rect 33597 13308 33609 13311
rect 33468 13280 33609 13308
rect 33468 13268 33474 13280
rect 33597 13277 33609 13280
rect 33643 13277 33655 13311
rect 33597 13271 33655 13277
rect 32490 13132 32496 13184
rect 32548 13172 32554 13184
rect 33689 13175 33747 13181
rect 33689 13172 33701 13175
rect 32548 13144 33701 13172
rect 32548 13132 32554 13144
rect 33689 13141 33701 13144
rect 33735 13141 33747 13175
rect 33689 13135 33747 13141
rect 1104 13082 34868 13104
rect 1104 13030 12214 13082
rect 12266 13030 12278 13082
rect 12330 13030 12342 13082
rect 12394 13030 12406 13082
rect 12458 13030 12470 13082
rect 12522 13030 23478 13082
rect 23530 13030 23542 13082
rect 23594 13030 23606 13082
rect 23658 13030 23670 13082
rect 23722 13030 23734 13082
rect 23786 13030 34868 13082
rect 1104 13008 34868 13030
rect 32490 12900 32496 12912
rect 32451 12872 32496 12900
rect 32490 12860 32496 12872
rect 32548 12860 32554 12912
rect 34146 12900 34152 12912
rect 34107 12872 34152 12900
rect 34146 12860 34152 12872
rect 34204 12860 34210 12912
rect 32306 12832 32312 12844
rect 32267 12804 32312 12832
rect 32306 12792 32312 12804
rect 32364 12792 32370 12844
rect 1578 12588 1584 12640
rect 1636 12628 1642 12640
rect 1857 12631 1915 12637
rect 1857 12628 1869 12631
rect 1636 12600 1869 12628
rect 1636 12588 1642 12600
rect 1857 12597 1869 12600
rect 1903 12597 1915 12631
rect 1857 12591 1915 12597
rect 1104 12538 34868 12560
rect 1104 12486 6582 12538
rect 6634 12486 6646 12538
rect 6698 12486 6710 12538
rect 6762 12486 6774 12538
rect 6826 12486 6838 12538
rect 6890 12486 17846 12538
rect 17898 12486 17910 12538
rect 17962 12486 17974 12538
rect 18026 12486 18038 12538
rect 18090 12486 18102 12538
rect 18154 12486 29110 12538
rect 29162 12486 29174 12538
rect 29226 12486 29238 12538
rect 29290 12486 29302 12538
rect 29354 12486 29366 12538
rect 29418 12486 34868 12538
rect 1104 12464 34868 12486
rect 32309 12291 32367 12297
rect 32309 12257 32321 12291
rect 32355 12288 32367 12291
rect 33134 12288 33140 12300
rect 32355 12260 33140 12288
rect 32355 12257 32367 12260
rect 32309 12251 32367 12257
rect 33134 12248 33140 12260
rect 33192 12248 33198 12300
rect 34146 12288 34152 12300
rect 34107 12260 34152 12288
rect 34146 12248 34152 12260
rect 34204 12248 34210 12300
rect 1949 12223 2007 12229
rect 1949 12189 1961 12223
rect 1995 12220 2007 12223
rect 2222 12220 2228 12232
rect 1995 12192 2228 12220
rect 1995 12189 2007 12192
rect 1949 12183 2007 12189
rect 2222 12180 2228 12192
rect 2280 12220 2286 12232
rect 14366 12220 14372 12232
rect 2280 12192 14372 12220
rect 2280 12180 2286 12192
rect 14366 12180 14372 12192
rect 14424 12220 14430 12232
rect 20898 12220 20904 12232
rect 14424 12192 20904 12220
rect 14424 12180 14430 12192
rect 20898 12180 20904 12192
rect 20956 12180 20962 12232
rect 32493 12155 32551 12161
rect 32493 12121 32505 12155
rect 32539 12152 32551 12155
rect 33686 12152 33692 12164
rect 32539 12124 33692 12152
rect 32539 12121 32551 12124
rect 32493 12115 32551 12121
rect 33686 12112 33692 12124
rect 33744 12112 33750 12164
rect 1762 12044 1768 12096
rect 1820 12084 1826 12096
rect 2041 12087 2099 12093
rect 2041 12084 2053 12087
rect 1820 12056 2053 12084
rect 1820 12044 1826 12056
rect 2041 12053 2053 12056
rect 2087 12053 2099 12087
rect 2041 12047 2099 12053
rect 1104 11994 34868 12016
rect 1104 11942 12214 11994
rect 12266 11942 12278 11994
rect 12330 11942 12342 11994
rect 12394 11942 12406 11994
rect 12458 11942 12470 11994
rect 12522 11942 23478 11994
rect 23530 11942 23542 11994
rect 23594 11942 23606 11994
rect 23658 11942 23670 11994
rect 23722 11942 23734 11994
rect 23786 11942 34868 11994
rect 1104 11920 34868 11942
rect 1762 11812 1768 11824
rect 1723 11784 1768 11812
rect 1762 11772 1768 11784
rect 1820 11772 1826 11824
rect 32493 11815 32551 11821
rect 32493 11781 32505 11815
rect 32539 11812 32551 11815
rect 32766 11812 32772 11824
rect 32539 11784 32772 11812
rect 32539 11781 32551 11784
rect 32493 11775 32551 11781
rect 32766 11772 32772 11784
rect 32824 11772 32830 11824
rect 1578 11744 1584 11756
rect 1539 11716 1584 11744
rect 1578 11704 1584 11716
rect 1636 11704 1642 11756
rect 2774 11676 2780 11688
rect 2735 11648 2780 11676
rect 2774 11636 2780 11648
rect 2832 11636 2838 11688
rect 32309 11679 32367 11685
rect 32309 11645 32321 11679
rect 32355 11645 32367 11679
rect 32309 11639 32367 11645
rect 32324 11608 32352 11639
rect 32674 11636 32680 11688
rect 32732 11676 32738 11688
rect 32769 11679 32827 11685
rect 32769 11676 32781 11679
rect 32732 11648 32781 11676
rect 32732 11636 32738 11648
rect 32769 11645 32781 11648
rect 32815 11645 32827 11679
rect 32769 11639 32827 11645
rect 33962 11608 33968 11620
rect 32324 11580 33968 11608
rect 33962 11568 33968 11580
rect 34020 11568 34026 11620
rect 1104 11450 34868 11472
rect 1104 11398 6582 11450
rect 6634 11398 6646 11450
rect 6698 11398 6710 11450
rect 6762 11398 6774 11450
rect 6826 11398 6838 11450
rect 6890 11398 17846 11450
rect 17898 11398 17910 11450
rect 17962 11398 17974 11450
rect 18026 11398 18038 11450
rect 18090 11398 18102 11450
rect 18154 11398 29110 11450
rect 29162 11398 29174 11450
rect 29226 11398 29238 11450
rect 29290 11398 29302 11450
rect 29354 11398 29366 11450
rect 29418 11398 34868 11450
rect 1104 11376 34868 11398
rect 33686 11336 33692 11348
rect 33647 11308 33692 11336
rect 33686 11296 33692 11308
rect 33744 11296 33750 11348
rect 1854 11200 1860 11212
rect 1815 11172 1860 11200
rect 1854 11160 1860 11172
rect 1912 11160 1918 11212
rect 1394 11132 1400 11144
rect 1355 11104 1400 11132
rect 1394 11092 1400 11104
rect 1452 11092 1458 11144
rect 33594 11132 33600 11144
rect 33555 11104 33600 11132
rect 33594 11092 33600 11104
rect 33652 11092 33658 11144
rect 1578 11064 1584 11076
rect 1539 11036 1584 11064
rect 1578 11024 1584 11036
rect 1636 11024 1642 11076
rect 1104 10906 34868 10928
rect 1104 10854 12214 10906
rect 12266 10854 12278 10906
rect 12330 10854 12342 10906
rect 12394 10854 12406 10906
rect 12458 10854 12470 10906
rect 12522 10854 23478 10906
rect 23530 10854 23542 10906
rect 23594 10854 23606 10906
rect 23658 10854 23670 10906
rect 23722 10854 23734 10906
rect 23786 10854 34868 10906
rect 1104 10832 34868 10854
rect 1578 10752 1584 10804
rect 1636 10792 1642 10804
rect 1949 10795 2007 10801
rect 1949 10792 1961 10795
rect 1636 10764 1961 10792
rect 1636 10752 1642 10764
rect 1949 10761 1961 10764
rect 1995 10761 2007 10795
rect 1949 10755 2007 10761
rect 1857 10659 1915 10665
rect 1857 10625 1869 10659
rect 1903 10656 1915 10659
rect 2130 10656 2136 10668
rect 1903 10628 2136 10656
rect 1903 10625 1915 10628
rect 1857 10619 1915 10625
rect 2130 10616 2136 10628
rect 2188 10616 2194 10668
rect 33962 10656 33968 10668
rect 33923 10628 33968 10656
rect 33962 10616 33968 10628
rect 34020 10616 34026 10668
rect 1394 10548 1400 10600
rect 1452 10588 1458 10600
rect 2685 10591 2743 10597
rect 2685 10588 2697 10591
rect 1452 10560 2697 10588
rect 1452 10548 1458 10560
rect 2685 10557 2697 10560
rect 2731 10557 2743 10591
rect 2685 10551 2743 10557
rect 1104 10362 34868 10384
rect 1104 10310 6582 10362
rect 6634 10310 6646 10362
rect 6698 10310 6710 10362
rect 6762 10310 6774 10362
rect 6826 10310 6838 10362
rect 6890 10310 17846 10362
rect 17898 10310 17910 10362
rect 17962 10310 17974 10362
rect 18026 10310 18038 10362
rect 18090 10310 18102 10362
rect 18154 10310 29110 10362
rect 29162 10310 29174 10362
rect 29226 10310 29238 10362
rect 29290 10310 29302 10362
rect 29354 10310 29366 10362
rect 29418 10310 34868 10362
rect 1104 10288 34868 10310
rect 31570 10208 31576 10260
rect 31628 10248 31634 10260
rect 34057 10251 34115 10257
rect 34057 10248 34069 10251
rect 31628 10220 34069 10248
rect 31628 10208 31634 10220
rect 34057 10217 34069 10220
rect 34103 10217 34115 10251
rect 34057 10211 34115 10217
rect 1762 10044 1768 10056
rect 1723 10016 1768 10044
rect 1762 10004 1768 10016
rect 1820 10004 1826 10056
rect 2590 10044 2596 10056
rect 2551 10016 2596 10044
rect 2590 10004 2596 10016
rect 2648 10004 2654 10056
rect 32122 10004 32128 10056
rect 32180 10044 32186 10056
rect 33229 10047 33287 10053
rect 33229 10044 33241 10047
rect 32180 10016 33241 10044
rect 32180 10004 32186 10016
rect 33229 10013 33241 10016
rect 33275 10013 33287 10047
rect 33229 10007 33287 10013
rect 33962 9976 33968 9988
rect 33923 9948 33968 9976
rect 33962 9936 33968 9948
rect 34020 9936 34026 9988
rect 1670 9868 1676 9920
rect 1728 9908 1734 9920
rect 1857 9911 1915 9917
rect 1857 9908 1869 9911
rect 1728 9880 1869 9908
rect 1728 9868 1734 9880
rect 1857 9877 1869 9880
rect 1903 9877 1915 9911
rect 33318 9908 33324 9920
rect 33279 9880 33324 9908
rect 1857 9871 1915 9877
rect 33318 9868 33324 9880
rect 33376 9868 33382 9920
rect 1104 9818 34868 9840
rect 1104 9766 12214 9818
rect 12266 9766 12278 9818
rect 12330 9766 12342 9818
rect 12394 9766 12406 9818
rect 12458 9766 12470 9818
rect 12522 9766 23478 9818
rect 23530 9766 23542 9818
rect 23594 9766 23606 9818
rect 23658 9766 23670 9818
rect 23722 9766 23734 9818
rect 23786 9766 34868 9818
rect 1104 9744 34868 9766
rect 1670 9636 1676 9648
rect 1631 9608 1676 9636
rect 1670 9596 1676 9608
rect 1728 9596 1734 9648
rect 32493 9639 32551 9645
rect 32493 9605 32505 9639
rect 32539 9636 32551 9639
rect 33318 9636 33324 9648
rect 32539 9608 33324 9636
rect 32539 9605 32551 9608
rect 32493 9599 32551 9605
rect 33318 9596 33324 9608
rect 33376 9596 33382 9648
rect 1489 9503 1547 9509
rect 1489 9469 1501 9503
rect 1535 9500 1547 9503
rect 2590 9500 2596 9512
rect 1535 9472 2596 9500
rect 1535 9469 1547 9472
rect 1489 9463 1547 9469
rect 2590 9460 2596 9472
rect 2648 9460 2654 9512
rect 2866 9500 2872 9512
rect 2827 9472 2872 9500
rect 2866 9460 2872 9472
rect 2924 9460 2930 9512
rect 32309 9503 32367 9509
rect 32309 9469 32321 9503
rect 32355 9500 32367 9503
rect 33962 9500 33968 9512
rect 32355 9472 33968 9500
rect 32355 9469 32367 9472
rect 32309 9463 32367 9469
rect 33962 9460 33968 9472
rect 34020 9460 34026 9512
rect 34146 9500 34152 9512
rect 34107 9472 34152 9500
rect 34146 9460 34152 9472
rect 34204 9460 34210 9512
rect 1104 9274 34868 9296
rect 1104 9222 6582 9274
rect 6634 9222 6646 9274
rect 6698 9222 6710 9274
rect 6762 9222 6774 9274
rect 6826 9222 6838 9274
rect 6890 9222 17846 9274
rect 17898 9222 17910 9274
rect 17962 9222 17974 9274
rect 18026 9222 18038 9274
rect 18090 9222 18102 9274
rect 18154 9222 29110 9274
rect 29162 9222 29174 9274
rect 29226 9222 29238 9274
rect 29290 9222 29302 9274
rect 29354 9222 29366 9274
rect 29418 9222 34868 9274
rect 1104 9200 34868 9222
rect 33962 9160 33968 9172
rect 33923 9132 33968 9160
rect 33962 9120 33968 9132
rect 34020 9120 34026 9172
rect 2774 9024 2780 9036
rect 2735 8996 2780 9024
rect 2774 8984 2780 8996
rect 2832 8984 2838 9036
rect 1394 8956 1400 8968
rect 1355 8928 1400 8956
rect 1394 8916 1400 8928
rect 1452 8916 1458 8968
rect 1581 8891 1639 8897
rect 1581 8857 1593 8891
rect 1627 8888 1639 8891
rect 1946 8888 1952 8900
rect 1627 8860 1952 8888
rect 1627 8857 1639 8860
rect 1581 8851 1639 8857
rect 1946 8848 1952 8860
rect 2004 8848 2010 8900
rect 1104 8730 34868 8752
rect 1104 8678 12214 8730
rect 12266 8678 12278 8730
rect 12330 8678 12342 8730
rect 12394 8678 12406 8730
rect 12458 8678 12470 8730
rect 12522 8678 23478 8730
rect 23530 8678 23542 8730
rect 23594 8678 23606 8730
rect 23658 8678 23670 8730
rect 23722 8678 23734 8730
rect 23786 8678 34868 8730
rect 1104 8656 34868 8678
rect 1946 8616 1952 8628
rect 1907 8588 1952 8616
rect 1946 8576 1952 8588
rect 2004 8576 2010 8628
rect 1394 8508 1400 8560
rect 1452 8548 1458 8560
rect 1452 8520 2728 8548
rect 1452 8508 1458 8520
rect 1857 8483 1915 8489
rect 1857 8449 1869 8483
rect 1903 8480 1915 8483
rect 2314 8480 2320 8492
rect 1903 8452 2320 8480
rect 1903 8449 1915 8452
rect 1857 8443 1915 8449
rect 2314 8440 2320 8452
rect 2372 8440 2378 8492
rect 2700 8489 2728 8520
rect 2685 8483 2743 8489
rect 2685 8449 2697 8483
rect 2731 8449 2743 8483
rect 2685 8443 2743 8449
rect 1104 8186 34868 8208
rect 1104 8134 6582 8186
rect 6634 8134 6646 8186
rect 6698 8134 6710 8186
rect 6762 8134 6774 8186
rect 6826 8134 6838 8186
rect 6890 8134 17846 8186
rect 17898 8134 17910 8186
rect 17962 8134 17974 8186
rect 18026 8134 18038 8186
rect 18090 8134 18102 8186
rect 18154 8134 29110 8186
rect 29162 8134 29174 8186
rect 29226 8134 29238 8186
rect 29290 8134 29302 8186
rect 29354 8134 29366 8186
rect 29418 8134 34868 8186
rect 1104 8112 34868 8134
rect 2038 8072 2044 8084
rect 1999 8044 2044 8072
rect 2038 8032 2044 8044
rect 2096 8032 2102 8084
rect 1946 7868 1952 7880
rect 1907 7840 1952 7868
rect 1946 7828 1952 7840
rect 2004 7828 2010 7880
rect 2777 7871 2835 7877
rect 2777 7837 2789 7871
rect 2823 7837 2835 7871
rect 2777 7831 2835 7837
rect 1578 7760 1584 7812
rect 1636 7800 1642 7812
rect 2792 7800 2820 7831
rect 32582 7828 32588 7880
rect 32640 7868 32646 7880
rect 33965 7871 34023 7877
rect 33965 7868 33977 7871
rect 32640 7840 33977 7868
rect 32640 7828 32646 7840
rect 33965 7837 33977 7840
rect 34011 7837 34023 7871
rect 33965 7831 34023 7837
rect 1636 7772 2820 7800
rect 1636 7760 1642 7772
rect 1104 7642 34868 7664
rect 1104 7590 12214 7642
rect 12266 7590 12278 7642
rect 12330 7590 12342 7642
rect 12394 7590 12406 7642
rect 12458 7590 12470 7642
rect 12522 7590 23478 7642
rect 23530 7590 23542 7642
rect 23594 7590 23606 7642
rect 23658 7590 23670 7642
rect 23722 7590 23734 7642
rect 23786 7590 34868 7642
rect 1104 7568 34868 7590
rect 1578 7392 1584 7404
rect 1539 7364 1584 7392
rect 1578 7352 1584 7364
rect 1636 7352 1642 7404
rect 1762 7324 1768 7336
rect 1723 7296 1768 7324
rect 1762 7284 1768 7296
rect 1820 7284 1826 7336
rect 2774 7324 2780 7336
rect 2735 7296 2780 7324
rect 2774 7284 2780 7296
rect 2832 7284 2838 7336
rect 3878 7148 3884 7200
rect 3936 7188 3942 7200
rect 4065 7191 4123 7197
rect 4065 7188 4077 7191
rect 3936 7160 4077 7188
rect 3936 7148 3942 7160
rect 4065 7157 4077 7160
rect 4111 7157 4123 7191
rect 4065 7151 4123 7157
rect 29730 7148 29736 7200
rect 29788 7188 29794 7200
rect 33321 7191 33379 7197
rect 33321 7188 33333 7191
rect 29788 7160 33333 7188
rect 29788 7148 29794 7160
rect 33321 7157 33333 7160
rect 33367 7157 33379 7191
rect 33962 7188 33968 7200
rect 33923 7160 33968 7188
rect 33321 7151 33379 7157
rect 33962 7148 33968 7160
rect 34020 7148 34026 7200
rect 1104 7098 34868 7120
rect 1104 7046 6582 7098
rect 6634 7046 6646 7098
rect 6698 7046 6710 7098
rect 6762 7046 6774 7098
rect 6826 7046 6838 7098
rect 6890 7046 17846 7098
rect 17898 7046 17910 7098
rect 17962 7046 17974 7098
rect 18026 7046 18038 7098
rect 18090 7046 18102 7098
rect 18154 7046 29110 7098
rect 29162 7046 29174 7098
rect 29226 7046 29238 7098
rect 29290 7046 29302 7098
rect 29354 7046 29366 7098
rect 29418 7046 34868 7098
rect 1104 7024 34868 7046
rect 1762 6944 1768 6996
rect 1820 6984 1826 6996
rect 2041 6987 2099 6993
rect 2041 6984 2053 6987
rect 1820 6956 2053 6984
rect 1820 6944 1826 6956
rect 2041 6953 2053 6956
rect 2087 6953 2099 6987
rect 2041 6947 2099 6953
rect 32309 6851 32367 6857
rect 32309 6817 32321 6851
rect 32355 6848 32367 6851
rect 33962 6848 33968 6860
rect 32355 6820 33968 6848
rect 32355 6817 32367 6820
rect 32309 6811 32367 6817
rect 33962 6808 33968 6820
rect 34020 6808 34026 6860
rect 34146 6848 34152 6860
rect 34107 6820 34152 6848
rect 34146 6808 34152 6820
rect 34204 6808 34210 6860
rect 1946 6780 1952 6792
rect 1907 6752 1952 6780
rect 1946 6740 1952 6752
rect 2004 6740 2010 6792
rect 2777 6783 2835 6789
rect 2777 6749 2789 6783
rect 2823 6780 2835 6783
rect 3142 6780 3148 6792
rect 2823 6752 3148 6780
rect 2823 6749 2835 6752
rect 2777 6743 2835 6749
rect 3142 6740 3148 6752
rect 3200 6740 3206 6792
rect 3786 6780 3792 6792
rect 3747 6752 3792 6780
rect 3786 6740 3792 6752
rect 3844 6740 3850 6792
rect 31662 6740 31668 6792
rect 31720 6780 31726 6792
rect 31849 6783 31907 6789
rect 31849 6780 31861 6783
rect 31720 6752 31861 6780
rect 31720 6740 31726 6752
rect 31849 6749 31861 6752
rect 31895 6749 31907 6783
rect 31849 6743 31907 6749
rect 32493 6715 32551 6721
rect 32493 6681 32505 6715
rect 32539 6712 32551 6715
rect 33686 6712 33692 6724
rect 32539 6684 33692 6712
rect 32539 6681 32551 6684
rect 32493 6675 32551 6681
rect 33686 6672 33692 6684
rect 33744 6672 33750 6724
rect 3881 6647 3939 6653
rect 3881 6613 3893 6647
rect 3927 6644 3939 6647
rect 3970 6644 3976 6656
rect 3927 6616 3976 6644
rect 3927 6613 3939 6616
rect 3881 6607 3939 6613
rect 3970 6604 3976 6616
rect 4028 6604 4034 6656
rect 1104 6554 34868 6576
rect 1104 6502 12214 6554
rect 12266 6502 12278 6554
rect 12330 6502 12342 6554
rect 12394 6502 12406 6554
rect 12458 6502 12470 6554
rect 12522 6502 23478 6554
rect 23530 6502 23542 6554
rect 23594 6502 23606 6554
rect 23658 6502 23670 6554
rect 23722 6502 23734 6554
rect 23786 6502 34868 6554
rect 1104 6480 34868 6502
rect 33686 6440 33692 6452
rect 33647 6412 33692 6440
rect 33686 6400 33692 6412
rect 33744 6400 33750 6452
rect 32950 6304 32956 6316
rect 32911 6276 32956 6304
rect 32950 6264 32956 6276
rect 33008 6264 33014 6316
rect 33410 6264 33416 6316
rect 33468 6304 33474 6316
rect 33597 6307 33655 6313
rect 33597 6304 33609 6307
rect 33468 6276 33609 6304
rect 33468 6264 33474 6276
rect 33597 6273 33609 6276
rect 33643 6273 33655 6307
rect 33597 6267 33655 6273
rect 2041 6239 2099 6245
rect 2041 6205 2053 6239
rect 2087 6205 2099 6239
rect 2041 6199 2099 6205
rect 2225 6239 2283 6245
rect 2225 6205 2237 6239
rect 2271 6236 2283 6239
rect 2866 6236 2872 6248
rect 2271 6208 2872 6236
rect 2271 6205 2283 6208
rect 2225 6199 2283 6205
rect 2056 6168 2084 6199
rect 2866 6196 2872 6208
rect 2924 6196 2930 6248
rect 3234 6236 3240 6248
rect 3195 6208 3240 6236
rect 3234 6196 3240 6208
rect 3292 6196 3298 6248
rect 6454 6168 6460 6180
rect 2056 6140 6460 6168
rect 6454 6128 6460 6140
rect 6512 6128 6518 6180
rect 1394 6060 1400 6112
rect 1452 6100 1458 6112
rect 1581 6103 1639 6109
rect 1581 6100 1593 6103
rect 1452 6072 1593 6100
rect 1452 6060 1458 6072
rect 1581 6069 1593 6072
rect 1627 6069 1639 6103
rect 4522 6100 4528 6112
rect 4483 6072 4528 6100
rect 1581 6063 1639 6069
rect 4522 6060 4528 6072
rect 4580 6060 4586 6112
rect 5166 6100 5172 6112
rect 5127 6072 5172 6100
rect 5166 6060 5172 6072
rect 5224 6060 5230 6112
rect 30466 6060 30472 6112
rect 30524 6100 30530 6112
rect 31573 6103 31631 6109
rect 31573 6100 31585 6103
rect 30524 6072 31585 6100
rect 30524 6060 30530 6072
rect 31573 6069 31585 6072
rect 31619 6069 31631 6103
rect 32490 6100 32496 6112
rect 32451 6072 32496 6100
rect 31573 6063 31631 6069
rect 32490 6060 32496 6072
rect 32548 6060 32554 6112
rect 33042 6100 33048 6112
rect 33003 6072 33048 6100
rect 33042 6060 33048 6072
rect 33100 6060 33106 6112
rect 1104 6010 34868 6032
rect 1104 5958 6582 6010
rect 6634 5958 6646 6010
rect 6698 5958 6710 6010
rect 6762 5958 6774 6010
rect 6826 5958 6838 6010
rect 6890 5958 17846 6010
rect 17898 5958 17910 6010
rect 17962 5958 17974 6010
rect 18026 5958 18038 6010
rect 18090 5958 18102 6010
rect 18154 5958 29110 6010
rect 29162 5958 29174 6010
rect 29226 5958 29238 6010
rect 29290 5958 29302 6010
rect 29354 5958 29366 6010
rect 29418 5958 34868 6010
rect 1104 5936 34868 5958
rect 31205 5899 31263 5905
rect 31205 5865 31217 5899
rect 31251 5896 31263 5899
rect 32306 5896 32312 5908
rect 31251 5868 32312 5896
rect 31251 5865 31263 5868
rect 31205 5859 31263 5865
rect 32306 5856 32312 5868
rect 32364 5856 32370 5908
rect 4522 5828 4528 5840
rect 1412 5800 4528 5828
rect 1412 5769 1440 5800
rect 4522 5788 4528 5800
rect 4580 5788 4586 5840
rect 24026 5788 24032 5840
rect 24084 5828 24090 5840
rect 24084 5800 34008 5828
rect 24084 5788 24090 5800
rect 1397 5763 1455 5769
rect 1397 5729 1409 5763
rect 1443 5729 1455 5763
rect 1854 5760 1860 5772
rect 1815 5732 1860 5760
rect 1397 5723 1455 5729
rect 1854 5720 1860 5732
rect 1912 5720 1918 5772
rect 3786 5760 3792 5772
rect 3747 5732 3792 5760
rect 3786 5720 3792 5732
rect 3844 5720 3850 5772
rect 3970 5760 3976 5772
rect 3931 5732 3976 5760
rect 3970 5720 3976 5732
rect 4028 5720 4034 5772
rect 4154 5720 4160 5772
rect 4212 5760 4218 5772
rect 4249 5763 4307 5769
rect 4249 5760 4261 5763
rect 4212 5732 4261 5760
rect 4212 5720 4218 5732
rect 4249 5729 4261 5732
rect 4295 5729 4307 5763
rect 31662 5760 31668 5772
rect 31623 5732 31668 5760
rect 4249 5723 4307 5729
rect 31662 5720 31668 5732
rect 31720 5720 31726 5772
rect 33134 5760 33140 5772
rect 33095 5732 33140 5760
rect 33134 5720 33140 5732
rect 33192 5720 33198 5772
rect 6270 5692 6276 5704
rect 6231 5664 6276 5692
rect 6270 5652 6276 5664
rect 6328 5652 6334 5704
rect 30561 5695 30619 5701
rect 30561 5661 30573 5695
rect 30607 5692 30619 5695
rect 31478 5692 31484 5704
rect 30607 5664 31484 5692
rect 30607 5661 30619 5664
rect 30561 5655 30619 5661
rect 31478 5652 31484 5664
rect 31536 5652 31542 5704
rect 33980 5701 34008 5800
rect 33965 5695 34023 5701
rect 33965 5661 33977 5695
rect 34011 5661 34023 5695
rect 33965 5655 34023 5661
rect 1578 5624 1584 5636
rect 1539 5596 1584 5624
rect 1578 5584 1584 5596
rect 1636 5584 1642 5636
rect 31846 5624 31852 5636
rect 31807 5596 31852 5624
rect 31846 5584 31852 5596
rect 31904 5584 31910 5636
rect 34054 5556 34060 5568
rect 34015 5528 34060 5556
rect 34054 5516 34060 5528
rect 34112 5516 34118 5568
rect 1104 5466 34868 5488
rect 1104 5414 12214 5466
rect 12266 5414 12278 5466
rect 12330 5414 12342 5466
rect 12394 5414 12406 5466
rect 12458 5414 12470 5466
rect 12522 5414 23478 5466
rect 23530 5414 23542 5466
rect 23594 5414 23606 5466
rect 23658 5414 23670 5466
rect 23722 5414 23734 5466
rect 23786 5414 34868 5466
rect 1104 5392 34868 5414
rect 1578 5312 1584 5364
rect 1636 5352 1642 5364
rect 1857 5355 1915 5361
rect 1857 5352 1869 5355
rect 1636 5324 1869 5352
rect 1636 5312 1642 5324
rect 1857 5321 1869 5324
rect 1903 5321 1915 5355
rect 1857 5315 1915 5321
rect 4706 5312 4712 5364
rect 4764 5352 4770 5364
rect 32950 5352 32956 5364
rect 4764 5324 32956 5352
rect 4764 5312 4770 5324
rect 32950 5312 32956 5324
rect 33008 5312 33014 5364
rect 5166 5284 5172 5296
rect 2608 5256 5172 5284
rect 1670 5176 1676 5228
rect 1728 5216 1734 5228
rect 2608 5225 2636 5256
rect 5166 5244 5172 5256
rect 5224 5244 5230 5296
rect 31481 5287 31539 5293
rect 31481 5253 31493 5287
rect 31527 5284 31539 5287
rect 32493 5287 32551 5293
rect 32493 5284 32505 5287
rect 31527 5256 32505 5284
rect 31527 5253 31539 5256
rect 31481 5247 31539 5253
rect 32493 5253 32505 5256
rect 32539 5253 32551 5287
rect 32493 5247 32551 5253
rect 1765 5219 1823 5225
rect 1765 5216 1777 5219
rect 1728 5188 1777 5216
rect 1728 5176 1734 5188
rect 1765 5185 1777 5188
rect 1811 5185 1823 5219
rect 1765 5179 1823 5185
rect 2593 5219 2651 5225
rect 2593 5185 2605 5219
rect 2639 5185 2651 5219
rect 2593 5179 2651 5185
rect 6454 5176 6460 5228
rect 6512 5216 6518 5228
rect 6549 5219 6607 5225
rect 6549 5216 6561 5219
rect 6512 5188 6561 5216
rect 6512 5176 6518 5188
rect 6549 5185 6561 5188
rect 6595 5185 6607 5219
rect 6549 5179 6607 5185
rect 27614 5176 27620 5228
rect 27672 5216 27678 5228
rect 29457 5219 29515 5225
rect 29457 5216 29469 5219
rect 27672 5188 29469 5216
rect 27672 5176 27678 5188
rect 29457 5185 29469 5188
rect 29503 5185 29515 5219
rect 29457 5179 29515 5185
rect 29638 5176 29644 5228
rect 29696 5216 29702 5228
rect 29822 5216 29828 5228
rect 29696 5188 29828 5216
rect 29696 5176 29702 5188
rect 29822 5176 29828 5188
rect 29880 5216 29886 5228
rect 30745 5219 30803 5225
rect 30745 5216 30757 5219
rect 29880 5188 30757 5216
rect 29880 5176 29886 5188
rect 30745 5185 30757 5188
rect 30791 5185 30803 5219
rect 30745 5179 30803 5185
rect 2774 5148 2780 5160
rect 2735 5120 2780 5148
rect 2774 5108 2780 5120
rect 2832 5108 2838 5160
rect 3050 5148 3056 5160
rect 3011 5120 3056 5148
rect 3050 5108 3056 5120
rect 3108 5108 3114 5160
rect 30760 5148 30788 5179
rect 31386 5176 31392 5228
rect 31444 5216 31450 5228
rect 31444 5188 31489 5216
rect 31444 5176 31450 5188
rect 32214 5148 32220 5160
rect 30760 5120 32220 5148
rect 32214 5108 32220 5120
rect 32272 5108 32278 5160
rect 32309 5151 32367 5157
rect 32309 5117 32321 5151
rect 32355 5148 32367 5151
rect 32582 5148 32588 5160
rect 32355 5120 32588 5148
rect 32355 5117 32367 5120
rect 32309 5111 32367 5117
rect 32582 5108 32588 5120
rect 32640 5108 32646 5160
rect 34146 5148 34152 5160
rect 34107 5120 34152 5148
rect 34146 5108 34152 5120
rect 34204 5108 34210 5160
rect 30374 5040 30380 5092
rect 30432 5080 30438 5092
rect 31386 5080 31392 5092
rect 30432 5052 31392 5080
rect 30432 5040 30438 5052
rect 31386 5040 31392 5052
rect 31444 5080 31450 5092
rect 33870 5080 33876 5092
rect 31444 5052 33876 5080
rect 31444 5040 31450 5052
rect 33870 5040 33876 5052
rect 33928 5040 33934 5092
rect 4430 4972 4436 5024
rect 4488 5012 4494 5024
rect 5077 5015 5135 5021
rect 5077 5012 5089 5015
rect 4488 4984 5089 5012
rect 4488 4972 4494 4984
rect 5077 4981 5089 4984
rect 5123 4981 5135 5015
rect 5077 4975 5135 4981
rect 5166 4972 5172 5024
rect 5224 5012 5230 5024
rect 5721 5015 5779 5021
rect 5721 5012 5733 5015
rect 5224 4984 5733 5012
rect 5224 4972 5230 4984
rect 5721 4981 5733 4984
rect 5767 4981 5779 5015
rect 29546 5012 29552 5024
rect 29507 4984 29552 5012
rect 5721 4975 5779 4981
rect 29546 4972 29552 4984
rect 29604 4972 29610 5024
rect 29822 4972 29828 5024
rect 29880 5012 29886 5024
rect 30285 5015 30343 5021
rect 30285 5012 30297 5015
rect 29880 4984 30297 5012
rect 29880 4972 29886 4984
rect 30285 4981 30297 4984
rect 30331 4981 30343 5015
rect 30834 5012 30840 5024
rect 30795 4984 30840 5012
rect 30285 4975 30343 4981
rect 30834 4972 30840 4984
rect 30892 4972 30898 5024
rect 1104 4922 34868 4944
rect 1104 4870 6582 4922
rect 6634 4870 6646 4922
rect 6698 4870 6710 4922
rect 6762 4870 6774 4922
rect 6826 4870 6838 4922
rect 6890 4870 17846 4922
rect 17898 4870 17910 4922
rect 17962 4870 17974 4922
rect 18026 4870 18038 4922
rect 18090 4870 18102 4922
rect 18154 4870 29110 4922
rect 29162 4870 29174 4922
rect 29226 4870 29238 4922
rect 29290 4870 29302 4922
rect 29354 4870 29366 4922
rect 29418 4870 34868 4922
rect 1104 4848 34868 4870
rect 2774 4768 2780 4820
rect 2832 4808 2838 4820
rect 3881 4811 3939 4817
rect 3881 4808 3893 4811
rect 2832 4780 3893 4808
rect 2832 4768 2838 4780
rect 3881 4777 3893 4780
rect 3927 4777 3939 4811
rect 3881 4771 3939 4777
rect 2958 4700 2964 4752
rect 3016 4740 3022 4752
rect 3016 4712 5672 4740
rect 3016 4700 3022 4712
rect 2777 4675 2835 4681
rect 2777 4641 2789 4675
rect 2823 4672 2835 4675
rect 2866 4672 2872 4684
rect 2823 4644 2872 4672
rect 2823 4641 2835 4644
rect 2777 4635 2835 4641
rect 2866 4632 2872 4644
rect 2924 4632 2930 4684
rect 4890 4672 4896 4684
rect 3712 4644 4896 4672
rect 1857 4607 1915 4613
rect 1857 4573 1869 4607
rect 1903 4573 1915 4607
rect 1857 4567 1915 4573
rect 2685 4607 2743 4613
rect 2685 4573 2697 4607
rect 2731 4604 2743 4607
rect 3712 4604 3740 4644
rect 4890 4632 4896 4644
rect 4948 4632 4954 4684
rect 5166 4672 5172 4684
rect 5127 4644 5172 4672
rect 5166 4632 5172 4644
rect 5224 4632 5230 4684
rect 5644 4681 5672 4712
rect 29546 4700 29552 4752
rect 29604 4740 29610 4752
rect 29604 4712 30052 4740
rect 29604 4700 29610 4712
rect 5629 4675 5687 4681
rect 5629 4641 5641 4675
rect 5675 4641 5687 4675
rect 29822 4672 29828 4684
rect 29783 4644 29828 4672
rect 5629 4635 5687 4641
rect 29822 4632 29828 4644
rect 29880 4632 29886 4684
rect 30024 4681 30052 4712
rect 30009 4675 30067 4681
rect 30009 4641 30021 4675
rect 30055 4641 30067 4675
rect 30926 4672 30932 4684
rect 30887 4644 30932 4672
rect 30009 4635 30067 4641
rect 30926 4632 30932 4644
rect 30984 4632 30990 4684
rect 32306 4672 32312 4684
rect 32267 4644 32312 4672
rect 32306 4632 32312 4644
rect 32364 4632 32370 4684
rect 32493 4675 32551 4681
rect 32493 4641 32505 4675
rect 32539 4672 32551 4675
rect 33042 4672 33048 4684
rect 32539 4644 33048 4672
rect 32539 4641 32551 4644
rect 32493 4635 32551 4641
rect 33042 4632 33048 4644
rect 33100 4632 33106 4684
rect 2731 4576 3740 4604
rect 3789 4607 3847 4613
rect 2731 4573 2743 4576
rect 2685 4567 2743 4573
rect 3789 4573 3801 4607
rect 3835 4573 3847 4607
rect 3789 4567 3847 4573
rect 1872 4536 1900 4567
rect 2774 4536 2780 4548
rect 1872 4508 2780 4536
rect 2774 4496 2780 4508
rect 2832 4496 2838 4548
rect 3804 4536 3832 4567
rect 4246 4564 4252 4616
rect 4304 4604 4310 4616
rect 4433 4607 4491 4613
rect 4433 4604 4445 4607
rect 4304 4576 4445 4604
rect 4304 4564 4310 4576
rect 4433 4573 4445 4576
rect 4479 4573 4491 4607
rect 4433 4567 4491 4573
rect 7742 4564 7748 4616
rect 7800 4604 7806 4616
rect 8021 4607 8079 4613
rect 8021 4604 8033 4607
rect 7800 4576 8033 4604
rect 7800 4564 7806 4576
rect 8021 4573 8033 4576
rect 8067 4573 8079 4607
rect 9858 4604 9864 4616
rect 9819 4576 9864 4604
rect 8021 4567 8079 4573
rect 9858 4564 9864 4576
rect 9916 4564 9922 4616
rect 10502 4604 10508 4616
rect 10463 4576 10508 4604
rect 10502 4564 10508 4576
rect 10560 4564 10566 4616
rect 4706 4536 4712 4548
rect 3804 4508 4712 4536
rect 4706 4496 4712 4508
rect 4764 4496 4770 4548
rect 5350 4536 5356 4548
rect 5311 4508 5356 4536
rect 5350 4496 5356 4508
rect 5408 4496 5414 4548
rect 34146 4536 34152 4548
rect 34107 4508 34152 4536
rect 34146 4496 34152 4508
rect 34204 4496 34210 4548
rect 1578 4428 1584 4480
rect 1636 4468 1642 4480
rect 1949 4471 2007 4477
rect 1949 4468 1961 4471
rect 1636 4440 1961 4468
rect 1636 4428 1642 4440
rect 1949 4437 1961 4440
rect 1995 4437 2007 4471
rect 1949 4431 2007 4437
rect 4525 4471 4583 4477
rect 4525 4437 4537 4471
rect 4571 4468 4583 4471
rect 6362 4468 6368 4480
rect 4571 4440 6368 4468
rect 4571 4437 4583 4440
rect 4525 4431 4583 4437
rect 6362 4428 6368 4440
rect 6420 4428 6426 4480
rect 1104 4378 34868 4400
rect 1104 4326 12214 4378
rect 12266 4326 12278 4378
rect 12330 4326 12342 4378
rect 12394 4326 12406 4378
rect 12458 4326 12470 4378
rect 12522 4326 23478 4378
rect 23530 4326 23542 4378
rect 23594 4326 23606 4378
rect 23658 4326 23670 4378
rect 23722 4326 23734 4378
rect 23786 4326 34868 4378
rect 1104 4304 34868 4326
rect 2498 4156 2504 4208
rect 2556 4196 2562 4208
rect 4246 4196 4252 4208
rect 2556 4168 3188 4196
rect 2556 4156 2562 4168
rect 1765 4063 1823 4069
rect 1765 4029 1777 4063
rect 1811 4029 1823 4063
rect 1765 4023 1823 4029
rect 1949 4063 2007 4069
rect 1949 4029 1961 4063
rect 1995 4029 2007 4063
rect 2866 4060 2872 4072
rect 2827 4032 2872 4060
rect 1949 4023 2007 4029
rect 1780 3924 1808 4023
rect 1964 3992 1992 4023
rect 2866 4020 2872 4032
rect 2924 4020 2930 4072
rect 3160 4060 3188 4168
rect 4080 4168 4252 4196
rect 4080 4137 4108 4168
rect 4246 4156 4252 4168
rect 4304 4156 4310 4208
rect 29917 4199 29975 4205
rect 29917 4196 29929 4199
rect 29564 4168 29929 4196
rect 4065 4131 4123 4137
rect 4065 4097 4077 4131
rect 4111 4097 4123 4131
rect 4709 4131 4767 4137
rect 4709 4128 4721 4131
rect 4065 4091 4123 4097
rect 4172 4100 4721 4128
rect 4172 4060 4200 4100
rect 4709 4097 4721 4100
rect 4755 4097 4767 4131
rect 7742 4128 7748 4140
rect 7703 4100 7748 4128
rect 4709 4091 4767 4097
rect 7742 4088 7748 4100
rect 7800 4088 7806 4140
rect 10229 4131 10287 4137
rect 10229 4097 10241 4131
rect 10275 4128 10287 4131
rect 13814 4128 13820 4140
rect 10275 4100 13820 4128
rect 10275 4097 10287 4100
rect 10229 4091 10287 4097
rect 13814 4088 13820 4100
rect 13872 4088 13878 4140
rect 20533 4131 20591 4137
rect 20533 4097 20545 4131
rect 20579 4128 20591 4131
rect 21818 4128 21824 4140
rect 20579 4100 21824 4128
rect 20579 4097 20591 4100
rect 20533 4091 20591 4097
rect 21818 4088 21824 4100
rect 21876 4088 21882 4140
rect 29089 4131 29147 4137
rect 29089 4097 29101 4131
rect 29135 4097 29147 4131
rect 29089 4091 29147 4097
rect 29181 4131 29239 4137
rect 29181 4097 29193 4131
rect 29227 4128 29239 4131
rect 29564 4128 29592 4168
rect 29917 4165 29929 4168
rect 29963 4165 29975 4199
rect 29917 4159 29975 4165
rect 29730 4128 29736 4140
rect 29227 4100 29592 4128
rect 29691 4100 29736 4128
rect 29227 4097 29239 4100
rect 29181 4091 29239 4097
rect 3160 4032 4200 4060
rect 4338 4020 4344 4072
rect 4396 4060 4402 4072
rect 6549 4063 6607 4069
rect 6549 4060 6561 4063
rect 4396 4032 6561 4060
rect 4396 4020 4402 4032
rect 6549 4029 6561 4032
rect 6595 4029 6607 4063
rect 6549 4023 6607 4029
rect 7929 4063 7987 4069
rect 7929 4029 7941 4063
rect 7975 4060 7987 4063
rect 8018 4060 8024 4072
rect 7975 4032 8024 4060
rect 7975 4029 7987 4032
rect 7929 4023 7987 4029
rect 8018 4020 8024 4032
rect 8076 4020 8082 4072
rect 8386 4060 8392 4072
rect 8347 4032 8392 4060
rect 8386 4020 8392 4032
rect 8444 4020 8450 4072
rect 27706 4020 27712 4072
rect 27764 4060 27770 4072
rect 28902 4060 28908 4072
rect 27764 4032 28908 4060
rect 27764 4020 27770 4032
rect 28902 4020 28908 4032
rect 28960 4060 28966 4072
rect 29104 4060 29132 4091
rect 29730 4088 29736 4100
rect 29788 4088 29794 4140
rect 31478 4088 31484 4140
rect 31536 4128 31542 4140
rect 32125 4131 32183 4137
rect 32125 4128 32137 4131
rect 31536 4100 32137 4128
rect 31536 4088 31542 4100
rect 32125 4097 32137 4100
rect 32171 4097 32183 4131
rect 32125 4091 32183 4097
rect 30742 4060 30748 4072
rect 28960 4032 30748 4060
rect 28960 4020 28966 4032
rect 30742 4020 30748 4032
rect 30800 4020 30806 4072
rect 31573 4063 31631 4069
rect 31573 4029 31585 4063
rect 31619 4060 31631 4063
rect 32030 4060 32036 4072
rect 31619 4032 32036 4060
rect 31619 4029 31631 4032
rect 31573 4023 31631 4029
rect 32030 4020 32036 4032
rect 32088 4020 32094 4072
rect 32306 4060 32312 4072
rect 32267 4032 32312 4060
rect 32306 4020 32312 4032
rect 32364 4020 32370 4072
rect 33042 4060 33048 4072
rect 33003 4032 33048 4060
rect 33042 4020 33048 4032
rect 33100 4020 33106 4072
rect 4157 3995 4215 4001
rect 4157 3992 4169 3995
rect 1964 3964 4169 3992
rect 4157 3961 4169 3964
rect 4203 3961 4215 3995
rect 4157 3955 4215 3961
rect 5350 3952 5356 4004
rect 5408 3992 5414 4004
rect 20349 3995 20407 4001
rect 20349 3992 20361 3995
rect 5408 3964 20361 3992
rect 5408 3952 5414 3964
rect 20349 3961 20361 3964
rect 20395 3961 20407 3995
rect 20349 3955 20407 3961
rect 28350 3952 28356 4004
rect 28408 3992 28414 4004
rect 30374 3992 30380 4004
rect 28408 3964 30380 3992
rect 28408 3952 28414 3964
rect 30374 3952 30380 3964
rect 30432 3952 30438 4004
rect 3142 3924 3148 3936
rect 1780 3896 3148 3924
rect 3142 3884 3148 3896
rect 3200 3884 3206 3936
rect 4614 3884 4620 3936
rect 4672 3924 4678 3936
rect 4801 3927 4859 3933
rect 4801 3924 4813 3927
rect 4672 3896 4813 3924
rect 4672 3884 4678 3896
rect 4801 3893 4813 3896
rect 4847 3893 4859 3927
rect 5534 3924 5540 3936
rect 5495 3896 5540 3924
rect 4801 3887 4859 3893
rect 5534 3884 5540 3896
rect 5592 3884 5598 3936
rect 6914 3884 6920 3936
rect 6972 3924 6978 3936
rect 7193 3927 7251 3933
rect 7193 3924 7205 3927
rect 6972 3896 7205 3924
rect 6972 3884 6978 3896
rect 7193 3893 7205 3896
rect 7239 3893 7251 3927
rect 7193 3887 7251 3893
rect 9766 3884 9772 3936
rect 9824 3924 9830 3936
rect 10321 3927 10379 3933
rect 10321 3924 10333 3927
rect 9824 3896 10333 3924
rect 9824 3884 9830 3896
rect 10321 3893 10333 3896
rect 10367 3893 10379 3927
rect 10321 3887 10379 3893
rect 14274 3884 14280 3936
rect 14332 3924 14338 3936
rect 14553 3927 14611 3933
rect 14553 3924 14565 3927
rect 14332 3896 14565 3924
rect 14332 3884 14338 3896
rect 14553 3893 14565 3896
rect 14599 3893 14611 3927
rect 14553 3887 14611 3893
rect 15470 3884 15476 3936
rect 15528 3924 15534 3936
rect 15749 3927 15807 3933
rect 15749 3924 15761 3927
rect 15528 3896 15761 3924
rect 15528 3884 15534 3896
rect 15749 3893 15761 3896
rect 15795 3893 15807 3927
rect 15749 3887 15807 3893
rect 19426 3884 19432 3936
rect 19484 3924 19490 3936
rect 19705 3927 19763 3933
rect 19705 3924 19717 3927
rect 19484 3896 19717 3924
rect 19484 3884 19490 3896
rect 19705 3893 19717 3896
rect 19751 3893 19763 3927
rect 19705 3887 19763 3893
rect 20806 3884 20812 3936
rect 20864 3924 20870 3936
rect 21269 3927 21327 3933
rect 21269 3924 21281 3927
rect 20864 3896 21281 3924
rect 20864 3884 20870 3896
rect 21269 3893 21281 3896
rect 21315 3893 21327 3927
rect 21269 3887 21327 3893
rect 28629 3927 28687 3933
rect 28629 3893 28641 3927
rect 28675 3924 28687 3927
rect 29638 3924 29644 3936
rect 28675 3896 29644 3924
rect 28675 3893 28687 3896
rect 28629 3887 28687 3893
rect 29638 3884 29644 3896
rect 29696 3884 29702 3936
rect 1104 3834 34868 3856
rect 1104 3782 6582 3834
rect 6634 3782 6646 3834
rect 6698 3782 6710 3834
rect 6762 3782 6774 3834
rect 6826 3782 6838 3834
rect 6890 3782 17846 3834
rect 17898 3782 17910 3834
rect 17962 3782 17974 3834
rect 18026 3782 18038 3834
rect 18090 3782 18102 3834
rect 18154 3782 29110 3834
rect 29162 3782 29174 3834
rect 29226 3782 29238 3834
rect 29290 3782 29302 3834
rect 29354 3782 29366 3834
rect 29418 3782 34868 3834
rect 1104 3760 34868 3782
rect 4246 3680 4252 3732
rect 4304 3720 4310 3732
rect 7834 3720 7840 3732
rect 4304 3692 7840 3720
rect 4304 3680 4310 3692
rect 7834 3680 7840 3692
rect 7892 3680 7898 3732
rect 8018 3720 8024 3732
rect 7979 3692 8024 3720
rect 8018 3680 8024 3692
rect 8076 3680 8082 3732
rect 28350 3720 28356 3732
rect 8772 3692 28356 3720
rect 658 3612 664 3664
rect 716 3652 722 3664
rect 716 3624 1900 3652
rect 716 3612 722 3624
rect 1394 3584 1400 3596
rect 1355 3556 1400 3584
rect 1394 3544 1400 3556
rect 1452 3544 1458 3596
rect 1578 3584 1584 3596
rect 1539 3556 1584 3584
rect 1578 3544 1584 3556
rect 1636 3544 1642 3596
rect 1872 3593 1900 3624
rect 1857 3587 1915 3593
rect 1857 3553 1869 3587
rect 1903 3553 1915 3587
rect 4430 3584 4436 3596
rect 4391 3556 4436 3584
rect 1857 3547 1915 3553
rect 4430 3544 4436 3556
rect 4488 3544 4494 3596
rect 4614 3584 4620 3596
rect 4575 3556 4620 3584
rect 4614 3544 4620 3556
rect 4672 3544 4678 3596
rect 5166 3584 5172 3596
rect 5127 3556 5172 3584
rect 5166 3544 5172 3556
rect 5224 3544 5230 3596
rect 5258 3544 5264 3596
rect 5316 3584 5322 3596
rect 6917 3587 6975 3593
rect 6917 3584 6929 3587
rect 5316 3556 6929 3584
rect 5316 3544 5322 3556
rect 6917 3553 6929 3556
rect 6963 3553 6975 3587
rect 6917 3547 6975 3553
rect 2774 3476 2780 3528
rect 2832 3516 2838 3528
rect 3789 3519 3847 3525
rect 3789 3516 3801 3519
rect 2832 3488 3801 3516
rect 2832 3476 2838 3488
rect 3789 3485 3801 3488
rect 3835 3485 3847 3519
rect 7926 3516 7932 3528
rect 7839 3488 7932 3516
rect 3789 3479 3847 3485
rect 3804 3448 3832 3479
rect 7926 3476 7932 3488
rect 7984 3516 7990 3528
rect 8772 3516 8800 3692
rect 28350 3680 28356 3692
rect 28408 3680 28414 3732
rect 28905 3723 28963 3729
rect 28905 3689 28917 3723
rect 28951 3720 28963 3723
rect 32306 3720 32312 3732
rect 28951 3692 32312 3720
rect 28951 3689 28963 3692
rect 28905 3683 28963 3689
rect 32306 3680 32312 3692
rect 32364 3680 32370 3732
rect 10502 3652 10508 3664
rect 9600 3624 10508 3652
rect 9600 3593 9628 3624
rect 10502 3612 10508 3624
rect 10560 3612 10566 3664
rect 27709 3655 27767 3661
rect 14200 3624 26924 3652
rect 9585 3587 9643 3593
rect 9585 3553 9597 3587
rect 9631 3553 9643 3587
rect 9766 3584 9772 3596
rect 9727 3556 9772 3584
rect 9585 3547 9643 3553
rect 9766 3544 9772 3556
rect 9824 3544 9830 3596
rect 9950 3544 9956 3596
rect 10008 3584 10014 3596
rect 10045 3587 10103 3593
rect 10045 3584 10057 3587
rect 10008 3556 10057 3584
rect 10008 3544 10014 3556
rect 10045 3553 10057 3556
rect 10091 3553 10103 3587
rect 10045 3547 10103 3553
rect 8938 3516 8944 3528
rect 7984 3488 8800 3516
rect 8899 3488 8944 3516
rect 7984 3476 7990 3488
rect 8938 3476 8944 3488
rect 8996 3476 9002 3528
rect 10962 3476 10968 3528
rect 11020 3516 11026 3528
rect 12069 3519 12127 3525
rect 12069 3516 12081 3519
rect 11020 3488 12081 3516
rect 11020 3476 11026 3488
rect 12069 3485 12081 3488
rect 12115 3485 12127 3519
rect 13173 3519 13231 3525
rect 13173 3516 13185 3519
rect 12069 3479 12127 3485
rect 12406 3488 13185 3516
rect 3804 3420 11744 3448
rect 2498 3340 2504 3392
rect 2556 3380 2562 3392
rect 3881 3383 3939 3389
rect 3881 3380 3893 3383
rect 2556 3352 3893 3380
rect 2556 3340 2562 3352
rect 3881 3349 3893 3352
rect 3927 3349 3939 3383
rect 3881 3343 3939 3349
rect 9033 3383 9091 3389
rect 9033 3349 9045 3383
rect 9079 3380 9091 3383
rect 9306 3380 9312 3392
rect 9079 3352 9312 3380
rect 9079 3349 9091 3352
rect 9033 3343 9091 3349
rect 9306 3340 9312 3352
rect 9364 3340 9370 3392
rect 11716 3380 11744 3420
rect 11974 3408 11980 3460
rect 12032 3448 12038 3460
rect 12406 3448 12434 3488
rect 13173 3485 13185 3488
rect 13219 3485 13231 3519
rect 13173 3479 13231 3485
rect 12032 3420 12434 3448
rect 12032 3408 12038 3420
rect 14200 3380 14228 3624
rect 15470 3584 15476 3596
rect 15431 3556 15476 3584
rect 15470 3544 15476 3556
rect 15528 3544 15534 3596
rect 16114 3584 16120 3596
rect 16075 3556 16120 3584
rect 16114 3544 16120 3556
rect 16172 3544 16178 3596
rect 20806 3584 20812 3596
rect 20767 3556 20812 3584
rect 20806 3544 20812 3556
rect 20864 3544 20870 3596
rect 22189 3587 22247 3593
rect 22189 3553 22201 3587
rect 22235 3553 22247 3587
rect 22189 3547 22247 3553
rect 14277 3519 14335 3525
rect 14277 3485 14289 3519
rect 14323 3516 14335 3519
rect 14366 3516 14372 3528
rect 14323 3488 14372 3516
rect 14323 3485 14335 3488
rect 14277 3479 14335 3485
rect 14366 3476 14372 3488
rect 14424 3476 14430 3528
rect 16850 3476 16856 3528
rect 16908 3516 16914 3528
rect 17957 3519 18015 3525
rect 17957 3516 17969 3519
rect 16908 3488 17969 3516
rect 16908 3476 16914 3488
rect 17957 3485 17969 3488
rect 18003 3485 18015 3519
rect 17957 3479 18015 3485
rect 18414 3476 18420 3528
rect 18472 3516 18478 3528
rect 19242 3516 19248 3528
rect 18472 3488 19248 3516
rect 18472 3476 18478 3488
rect 19242 3476 19248 3488
rect 19300 3516 19306 3528
rect 19429 3519 19487 3525
rect 19429 3516 19441 3519
rect 19300 3488 19441 3516
rect 19300 3476 19306 3488
rect 19429 3485 19441 3488
rect 19475 3485 19487 3519
rect 20346 3516 20352 3528
rect 20307 3488 20352 3516
rect 19429 3479 19487 3485
rect 20346 3476 20352 3488
rect 20404 3476 20410 3528
rect 15654 3448 15660 3460
rect 15615 3420 15660 3448
rect 15654 3408 15660 3420
rect 15712 3408 15718 3460
rect 20993 3451 21051 3457
rect 20993 3417 21005 3451
rect 21039 3448 21051 3451
rect 21910 3448 21916 3460
rect 21039 3420 21916 3448
rect 21039 3417 21051 3420
rect 20993 3411 21051 3417
rect 21910 3408 21916 3420
rect 21968 3408 21974 3460
rect 11716 3352 14228 3380
rect 14369 3383 14427 3389
rect 14369 3349 14381 3383
rect 14415 3380 14427 3383
rect 14458 3380 14464 3392
rect 14415 3352 14464 3380
rect 14415 3349 14427 3352
rect 14369 3343 14427 3349
rect 14458 3340 14464 3352
rect 14516 3340 14522 3392
rect 19521 3383 19579 3389
rect 19521 3349 19533 3383
rect 19567 3380 19579 3383
rect 19610 3380 19616 3392
rect 19567 3352 19616 3380
rect 19567 3349 19579 3352
rect 19521 3343 19579 3349
rect 19610 3340 19616 3352
rect 19668 3340 19674 3392
rect 21266 3340 21272 3392
rect 21324 3380 21330 3392
rect 22204 3380 22232 3547
rect 23842 3476 23848 3528
rect 23900 3516 23906 3528
rect 24581 3519 24639 3525
rect 24581 3516 24593 3519
rect 23900 3488 24593 3516
rect 23900 3476 23906 3488
rect 24581 3485 24593 3488
rect 24627 3485 24639 3519
rect 24581 3479 24639 3485
rect 21324 3352 22232 3380
rect 26896 3380 26924 3624
rect 27709 3621 27721 3655
rect 27755 3652 27767 3655
rect 30190 3652 30196 3664
rect 27755 3624 30196 3652
rect 27755 3621 27767 3624
rect 27709 3615 27767 3621
rect 30190 3612 30196 3624
rect 30248 3612 30254 3664
rect 28353 3587 28411 3593
rect 28353 3553 28365 3587
rect 28399 3584 28411 3587
rect 30469 3587 30527 3593
rect 30469 3584 30481 3587
rect 28399 3556 30481 3584
rect 28399 3553 28411 3556
rect 28353 3547 28411 3553
rect 30469 3553 30481 3556
rect 30515 3553 30527 3587
rect 30469 3547 30527 3553
rect 32309 3587 32367 3593
rect 32309 3553 32321 3587
rect 32355 3584 32367 3587
rect 35434 3584 35440 3596
rect 32355 3556 35440 3584
rect 32355 3553 32367 3556
rect 32309 3547 32367 3553
rect 35434 3544 35440 3556
rect 35492 3544 35498 3596
rect 27890 3476 27896 3528
rect 27948 3516 27954 3528
rect 28813 3519 28871 3525
rect 28813 3516 28825 3519
rect 27948 3488 28825 3516
rect 27948 3476 27954 3488
rect 28813 3485 28825 3488
rect 28859 3485 28871 3519
rect 28813 3479 28871 3485
rect 29454 3476 29460 3528
rect 29512 3518 29518 3528
rect 29549 3519 29607 3525
rect 29549 3518 29561 3519
rect 29512 3490 29561 3518
rect 29512 3476 29518 3490
rect 29549 3485 29561 3490
rect 29595 3485 29607 3519
rect 29549 3479 29607 3485
rect 32214 3476 32220 3528
rect 32272 3516 32278 3528
rect 32953 3519 33011 3525
rect 32953 3516 32965 3519
rect 32272 3488 32965 3516
rect 32272 3476 32278 3488
rect 32953 3485 32965 3488
rect 32999 3485 33011 3519
rect 32953 3479 33011 3485
rect 28994 3408 29000 3460
rect 29052 3448 29058 3460
rect 29825 3451 29883 3457
rect 29825 3448 29837 3451
rect 29052 3420 29837 3448
rect 29052 3408 29058 3420
rect 29825 3417 29837 3420
rect 29871 3417 29883 3451
rect 30650 3448 30656 3460
rect 30611 3420 30656 3448
rect 29825 3411 29883 3417
rect 30650 3408 30656 3420
rect 30708 3408 30714 3460
rect 33778 3448 33784 3460
rect 31726 3420 33784 3448
rect 31726 3380 31754 3420
rect 33778 3408 33784 3420
rect 33836 3408 33842 3460
rect 26896 3352 31754 3380
rect 21324 3340 21330 3352
rect 1104 3290 34868 3312
rect 1104 3238 12214 3290
rect 12266 3238 12278 3290
rect 12330 3238 12342 3290
rect 12394 3238 12406 3290
rect 12458 3238 12470 3290
rect 12522 3238 23478 3290
rect 23530 3238 23542 3290
rect 23594 3238 23606 3290
rect 23658 3238 23670 3290
rect 23722 3238 23734 3290
rect 23786 3238 34868 3290
rect 1104 3216 34868 3238
rect 5534 3176 5540 3188
rect 2332 3148 5540 3176
rect 2332 3049 2360 3148
rect 5534 3136 5540 3148
rect 5592 3136 5598 3188
rect 15746 3176 15752 3188
rect 5644 3148 15752 3176
rect 2498 3108 2504 3120
rect 2459 3080 2504 3108
rect 2498 3068 2504 3080
rect 2556 3068 2562 3120
rect 2590 3068 2596 3120
rect 2648 3108 2654 3120
rect 2648 3080 4660 3108
rect 2648 3068 2654 3080
rect 4632 3049 4660 3080
rect 5644 3049 5672 3148
rect 15746 3136 15752 3148
rect 15804 3176 15810 3188
rect 21910 3176 21916 3188
rect 15804 3148 20484 3176
rect 21871 3148 21916 3176
rect 15804 3136 15810 3148
rect 5721 3111 5779 3117
rect 5721 3077 5733 3111
rect 5767 3108 5779 3111
rect 6549 3111 6607 3117
rect 6549 3108 6561 3111
rect 5767 3080 6561 3108
rect 5767 3077 5779 3080
rect 5721 3071 5779 3077
rect 6549 3077 6561 3080
rect 6595 3077 6607 3111
rect 9858 3108 9864 3120
rect 6549 3071 6607 3077
rect 9140 3080 9864 3108
rect 1673 3043 1731 3049
rect 1673 3009 1685 3043
rect 1719 3009 1731 3043
rect 1673 3003 1731 3009
rect 2317 3043 2375 3049
rect 2317 3009 2329 3043
rect 2363 3009 2375 3043
rect 2317 3003 2375 3009
rect 4617 3043 4675 3049
rect 4617 3009 4629 3043
rect 4663 3009 4675 3043
rect 4617 3003 4675 3009
rect 5629 3043 5687 3049
rect 5629 3009 5641 3043
rect 5675 3009 5687 3043
rect 5629 3003 5687 3009
rect 1688 2904 1716 3003
rect 2590 2932 2596 2984
rect 2648 2972 2654 2984
rect 2777 2975 2835 2981
rect 2777 2972 2789 2975
rect 2648 2944 2789 2972
rect 2648 2932 2654 2944
rect 2777 2941 2789 2944
rect 2823 2941 2835 2975
rect 4246 2972 4252 2984
rect 2777 2935 2835 2941
rect 3160 2944 4252 2972
rect 3160 2904 3188 2944
rect 4246 2932 4252 2944
rect 4304 2932 4310 2984
rect 5644 2972 5672 3003
rect 6270 3000 6276 3052
rect 6328 3040 6334 3052
rect 9140 3049 9168 3080
rect 9858 3068 9864 3080
rect 9916 3068 9922 3120
rect 14458 3108 14464 3120
rect 14419 3080 14464 3108
rect 14458 3068 14464 3080
rect 14516 3068 14522 3120
rect 20346 3108 20352 3120
rect 19444 3080 20352 3108
rect 6365 3043 6423 3049
rect 6365 3040 6377 3043
rect 6328 3012 6377 3040
rect 6328 3000 6334 3012
rect 6365 3009 6377 3012
rect 6411 3009 6423 3043
rect 6365 3003 6423 3009
rect 9125 3043 9183 3049
rect 9125 3009 9137 3043
rect 9171 3009 9183 3043
rect 11974 3040 11980 3052
rect 11935 3012 11980 3040
rect 9125 3003 9183 3009
rect 11974 3000 11980 3012
rect 12032 3000 12038 3052
rect 14274 3040 14280 3052
rect 14235 3012 14280 3040
rect 14274 3000 14280 3012
rect 14332 3000 14338 3052
rect 16850 3040 16856 3052
rect 16811 3012 16856 3040
rect 16850 3000 16856 3012
rect 16908 3000 16914 3052
rect 19444 3049 19472 3080
rect 20346 3068 20352 3080
rect 20404 3068 20410 3120
rect 20456 3108 20484 3148
rect 21910 3136 21916 3148
rect 21968 3136 21974 3188
rect 28994 3176 29000 3188
rect 22066 3148 29000 3176
rect 22066 3108 22094 3148
rect 28994 3136 29000 3148
rect 29052 3136 29058 3188
rect 29089 3179 29147 3185
rect 29089 3145 29101 3179
rect 29135 3176 29147 3179
rect 30650 3176 30656 3188
rect 29135 3148 30656 3176
rect 29135 3145 29147 3148
rect 29089 3139 29147 3145
rect 30650 3136 30656 3148
rect 30708 3136 30714 3188
rect 20456 3080 22094 3108
rect 23293 3111 23351 3117
rect 23293 3077 23305 3111
rect 23339 3108 23351 3111
rect 24029 3111 24087 3117
rect 24029 3108 24041 3111
rect 23339 3080 24041 3108
rect 23339 3077 23351 3080
rect 23293 3071 23351 3077
rect 24029 3077 24041 3080
rect 24075 3077 24087 3111
rect 24029 3071 24087 3077
rect 25240 3080 27844 3108
rect 19429 3043 19487 3049
rect 19429 3009 19441 3043
rect 19475 3009 19487 3043
rect 21818 3040 21824 3052
rect 21779 3012 21824 3040
rect 19429 3003 19487 3009
rect 21818 3000 21824 3012
rect 21876 3040 21882 3052
rect 23201 3043 23259 3049
rect 23201 3040 23213 3043
rect 21876 3012 23213 3040
rect 21876 3000 21882 3012
rect 23201 3009 23213 3012
rect 23247 3009 23259 3043
rect 23842 3040 23848 3052
rect 23803 3012 23848 3040
rect 23201 3003 23259 3009
rect 6825 2975 6883 2981
rect 6825 2972 6837 2975
rect 4356 2944 5672 2972
rect 6472 2944 6837 2972
rect 1688 2876 3188 2904
rect 1578 2796 1584 2848
rect 1636 2836 1642 2848
rect 1765 2839 1823 2845
rect 1765 2836 1777 2839
rect 1636 2808 1777 2836
rect 1636 2796 1642 2808
rect 1765 2805 1777 2808
rect 1811 2805 1823 2839
rect 1765 2799 1823 2805
rect 1946 2796 1952 2848
rect 2004 2836 2010 2848
rect 4356 2836 4384 2944
rect 6472 2916 6500 2944
rect 6825 2941 6837 2944
rect 6871 2941 6883 2975
rect 6825 2935 6883 2941
rect 9309 2975 9367 2981
rect 9309 2941 9321 2975
rect 9355 2941 9367 2975
rect 9674 2972 9680 2984
rect 9635 2944 9680 2972
rect 9309 2935 9367 2941
rect 6454 2864 6460 2916
rect 6512 2864 6518 2916
rect 9324 2904 9352 2935
rect 9674 2932 9680 2944
rect 9732 2932 9738 2984
rect 12161 2975 12219 2981
rect 12161 2941 12173 2975
rect 12207 2972 12219 2975
rect 13170 2972 13176 2984
rect 12207 2944 13176 2972
rect 12207 2941 12219 2944
rect 12161 2935 12219 2941
rect 13170 2932 13176 2944
rect 13228 2932 13234 2984
rect 13538 2972 13544 2984
rect 13499 2944 13544 2972
rect 13538 2932 13544 2944
rect 13596 2932 13602 2984
rect 14826 2972 14832 2984
rect 14787 2944 14832 2972
rect 14826 2932 14832 2944
rect 14884 2932 14890 2984
rect 17034 2972 17040 2984
rect 16995 2944 17040 2972
rect 17034 2932 17040 2944
rect 17092 2932 17098 2984
rect 17402 2972 17408 2984
rect 17363 2944 17408 2972
rect 17402 2932 17408 2944
rect 17460 2932 17466 2984
rect 19613 2975 19671 2981
rect 19613 2941 19625 2975
rect 19659 2941 19671 2975
rect 20622 2972 20628 2984
rect 20583 2944 20628 2972
rect 19613 2935 19671 2941
rect 10870 2904 10876 2916
rect 9324 2876 10876 2904
rect 10870 2864 10876 2876
rect 10928 2864 10934 2916
rect 19628 2904 19656 2935
rect 20622 2932 20628 2944
rect 20680 2932 20686 2984
rect 21910 2904 21916 2916
rect 19628 2876 21916 2904
rect 21910 2864 21916 2876
rect 21968 2864 21974 2916
rect 23216 2904 23244 3003
rect 23842 3000 23848 3012
rect 23900 3000 23906 3052
rect 24486 2972 24492 2984
rect 24447 2944 24492 2972
rect 24486 2932 24492 2944
rect 24544 2932 24550 2984
rect 25240 2904 25268 3080
rect 27706 3040 27712 3052
rect 27667 3012 27712 3040
rect 27706 3000 27712 3012
rect 27764 3000 27770 3052
rect 23216 2876 25268 2904
rect 27816 2904 27844 3080
rect 29012 3049 29040 3136
rect 32493 3111 32551 3117
rect 32493 3077 32505 3111
rect 32539 3108 32551 3111
rect 34054 3108 34060 3120
rect 32539 3080 34060 3108
rect 32539 3077 32551 3080
rect 32493 3071 32551 3077
rect 34054 3068 34060 3080
rect 34112 3068 34118 3120
rect 28353 3043 28411 3049
rect 28353 3009 28365 3043
rect 28399 3009 28411 3043
rect 28353 3003 28411 3009
rect 28997 3043 29055 3049
rect 28997 3009 29009 3043
rect 29043 3009 29055 3043
rect 29638 3040 29644 3052
rect 29599 3012 29644 3040
rect 28997 3003 29055 3009
rect 27890 2932 27896 2984
rect 27948 2972 27954 2984
rect 28368 2972 28396 3003
rect 29638 3000 29644 3012
rect 29696 3000 29702 3052
rect 27948 2944 28396 2972
rect 28445 2975 28503 2981
rect 27948 2932 27954 2944
rect 28445 2941 28457 2975
rect 28491 2972 28503 2975
rect 29825 2975 29883 2981
rect 29825 2972 29837 2975
rect 28491 2944 29837 2972
rect 28491 2941 28503 2944
rect 28445 2935 28503 2941
rect 29825 2941 29837 2944
rect 29871 2941 29883 2975
rect 30282 2972 30288 2984
rect 30243 2944 30288 2972
rect 29825 2935 29883 2941
rect 30282 2932 30288 2944
rect 30340 2932 30346 2984
rect 32309 2975 32367 2981
rect 32309 2941 32321 2975
rect 32355 2972 32367 2975
rect 32490 2972 32496 2984
rect 32355 2944 32496 2972
rect 32355 2941 32367 2944
rect 32309 2935 32367 2941
rect 32490 2932 32496 2944
rect 32548 2932 32554 2984
rect 34149 2975 34207 2981
rect 34149 2941 34161 2975
rect 34195 2972 34207 2975
rect 34790 2972 34796 2984
rect 34195 2944 34796 2972
rect 34195 2941 34207 2944
rect 34149 2935 34207 2941
rect 34790 2932 34796 2944
rect 34848 2932 34854 2984
rect 33226 2904 33232 2916
rect 27816 2876 33232 2904
rect 33226 2864 33232 2876
rect 33284 2864 33290 2916
rect 4706 2836 4712 2848
rect 2004 2808 4384 2836
rect 4667 2808 4712 2836
rect 2004 2796 2010 2808
rect 4706 2796 4712 2808
rect 4764 2796 4770 2848
rect 7834 2796 7840 2848
rect 7892 2836 7898 2848
rect 12434 2836 12440 2848
rect 7892 2808 12440 2836
rect 7892 2796 7898 2808
rect 12434 2796 12440 2808
rect 12492 2796 12498 2848
rect 19242 2796 19248 2848
rect 19300 2836 19306 2848
rect 27706 2836 27712 2848
rect 19300 2808 27712 2836
rect 19300 2796 19306 2808
rect 27706 2796 27712 2808
rect 27764 2796 27770 2848
rect 27801 2839 27859 2845
rect 27801 2805 27813 2839
rect 27847 2836 27859 2839
rect 29914 2836 29920 2848
rect 27847 2808 29920 2836
rect 27847 2805 27859 2808
rect 27801 2799 27859 2805
rect 29914 2796 29920 2808
rect 29972 2796 29978 2848
rect 32214 2796 32220 2848
rect 32272 2836 32278 2848
rect 33134 2836 33140 2848
rect 32272 2808 33140 2836
rect 32272 2796 32278 2808
rect 33134 2796 33140 2808
rect 33192 2796 33198 2848
rect 1104 2746 34868 2768
rect 1104 2694 6582 2746
rect 6634 2694 6646 2746
rect 6698 2694 6710 2746
rect 6762 2694 6774 2746
rect 6826 2694 6838 2746
rect 6890 2694 17846 2746
rect 17898 2694 17910 2746
rect 17962 2694 17974 2746
rect 18026 2694 18038 2746
rect 18090 2694 18102 2746
rect 18154 2694 29110 2746
rect 29162 2694 29174 2746
rect 29226 2694 29238 2746
rect 29290 2694 29302 2746
rect 29354 2694 29366 2746
rect 29418 2694 34868 2746
rect 1104 2672 34868 2694
rect 3418 2592 3424 2644
rect 3476 2632 3482 2644
rect 9674 2632 9680 2644
rect 3476 2604 9680 2632
rect 3476 2592 3482 2604
rect 9674 2592 9680 2604
rect 9732 2592 9738 2644
rect 13170 2592 13176 2644
rect 13228 2632 13234 2644
rect 13265 2635 13323 2641
rect 13265 2632 13277 2635
rect 13228 2604 13277 2632
rect 13228 2592 13234 2604
rect 13265 2601 13277 2604
rect 13311 2601 13323 2635
rect 13265 2595 13323 2601
rect 15654 2592 15660 2644
rect 15712 2632 15718 2644
rect 15841 2635 15899 2641
rect 15841 2632 15853 2635
rect 15712 2604 15853 2632
rect 15712 2592 15718 2604
rect 15841 2601 15853 2604
rect 15887 2601 15899 2635
rect 15841 2595 15899 2601
rect 16945 2635 17003 2641
rect 16945 2601 16957 2635
rect 16991 2632 17003 2635
rect 17034 2632 17040 2644
rect 16991 2604 17040 2632
rect 16991 2601 17003 2604
rect 16945 2595 17003 2601
rect 17034 2592 17040 2604
rect 17092 2592 17098 2644
rect 17494 2592 17500 2644
rect 17552 2632 17558 2644
rect 18325 2635 18383 2641
rect 18325 2632 18337 2635
rect 17552 2604 18337 2632
rect 17552 2592 17558 2604
rect 18325 2601 18337 2604
rect 18371 2601 18383 2635
rect 21910 2632 21916 2644
rect 21871 2604 21916 2632
rect 18325 2595 18383 2601
rect 21910 2592 21916 2604
rect 21968 2592 21974 2644
rect 28905 2635 28963 2641
rect 28905 2601 28917 2635
rect 28951 2632 28963 2635
rect 31846 2632 31852 2644
rect 28951 2604 31852 2632
rect 28951 2601 28963 2604
rect 28905 2595 28963 2601
rect 31846 2592 31852 2604
rect 31904 2592 31910 2644
rect 4338 2564 4344 2576
rect 3896 2536 4344 2564
rect 1578 2496 1584 2508
rect 1539 2468 1584 2496
rect 1578 2456 1584 2468
rect 1636 2456 1642 2508
rect 2774 2496 2780 2508
rect 2735 2468 2780 2496
rect 2774 2456 2780 2468
rect 2832 2456 2838 2508
rect 3896 2505 3924 2536
rect 4338 2524 4344 2536
rect 4396 2524 4402 2576
rect 4522 2524 4528 2576
rect 4580 2564 4586 2576
rect 10962 2564 10968 2576
rect 4580 2536 4844 2564
rect 4580 2524 4586 2536
rect 3881 2499 3939 2505
rect 3881 2465 3893 2499
rect 3927 2465 3939 2499
rect 3881 2459 3939 2465
rect 4065 2499 4123 2505
rect 4065 2465 4077 2499
rect 4111 2496 4123 2499
rect 4706 2496 4712 2508
rect 4111 2468 4712 2496
rect 4111 2465 4123 2468
rect 4065 2459 4123 2465
rect 4706 2456 4712 2468
rect 4764 2456 4770 2508
rect 4816 2505 4844 2536
rect 5644 2536 7052 2564
rect 4801 2499 4859 2505
rect 4801 2465 4813 2499
rect 4847 2465 4859 2499
rect 4801 2459 4859 2465
rect 1397 2431 1455 2437
rect 1397 2397 1409 2431
rect 1443 2397 1455 2431
rect 1397 2391 1455 2397
rect 1412 2360 1440 2391
rect 5258 2360 5264 2372
rect 1412 2332 5264 2360
rect 5258 2320 5264 2332
rect 5316 2320 5322 2372
rect 3234 2252 3240 2304
rect 3292 2292 3298 2304
rect 5644 2292 5672 2536
rect 6365 2499 6423 2505
rect 6365 2465 6377 2499
rect 6411 2496 6423 2499
rect 6914 2496 6920 2508
rect 6411 2468 6920 2496
rect 6411 2465 6423 2468
rect 6365 2459 6423 2465
rect 6914 2456 6920 2468
rect 6972 2456 6978 2508
rect 7024 2505 7052 2536
rect 9140 2536 10968 2564
rect 9140 2505 9168 2536
rect 10962 2524 10968 2536
rect 11020 2524 11026 2576
rect 30466 2564 30472 2576
rect 16868 2536 29684 2564
rect 7009 2499 7067 2505
rect 7009 2465 7021 2499
rect 7055 2465 7067 2499
rect 7009 2459 7067 2465
rect 9125 2499 9183 2505
rect 9125 2465 9137 2499
rect 9171 2465 9183 2499
rect 9306 2496 9312 2508
rect 9267 2468 9312 2496
rect 9125 2459 9183 2465
rect 9306 2456 9312 2468
rect 9364 2456 9370 2508
rect 10318 2496 10324 2508
rect 10279 2468 10324 2496
rect 10318 2456 10324 2468
rect 10376 2456 10382 2508
rect 10870 2456 10876 2508
rect 10928 2496 10934 2508
rect 14185 2499 14243 2505
rect 14185 2496 14197 2499
rect 10928 2468 14197 2496
rect 10928 2456 10934 2468
rect 14185 2465 14197 2468
rect 14231 2465 14243 2499
rect 16868 2496 16896 2536
rect 19426 2496 19432 2508
rect 14185 2459 14243 2465
rect 14936 2468 16896 2496
rect 19387 2468 19432 2496
rect 12434 2388 12440 2440
rect 12492 2428 12498 2440
rect 13173 2431 13231 2437
rect 13173 2428 13185 2431
rect 12492 2400 13185 2428
rect 12492 2388 12498 2400
rect 13173 2397 13185 2400
rect 13219 2397 13231 2431
rect 14090 2428 14096 2440
rect 14051 2400 14096 2428
rect 13173 2391 13231 2397
rect 6362 2320 6368 2372
rect 6420 2360 6426 2372
rect 6549 2363 6607 2369
rect 6549 2360 6561 2363
rect 6420 2332 6561 2360
rect 6420 2320 6426 2332
rect 6549 2329 6561 2332
rect 6595 2329 6607 2363
rect 13188 2360 13216 2391
rect 14090 2388 14096 2400
rect 14148 2428 14154 2440
rect 14936 2428 14964 2468
rect 15746 2428 15752 2440
rect 14148 2400 14964 2428
rect 15707 2400 15752 2428
rect 14148 2388 14154 2400
rect 15746 2388 15752 2400
rect 15804 2388 15810 2440
rect 16868 2437 16896 2468
rect 19426 2456 19432 2468
rect 19484 2456 19490 2508
rect 19610 2496 19616 2508
rect 19571 2468 19616 2496
rect 19610 2456 19616 2468
rect 19668 2456 19674 2508
rect 19978 2496 19984 2508
rect 19939 2468 19984 2496
rect 19978 2456 19984 2468
rect 20036 2456 20042 2508
rect 29546 2496 29552 2508
rect 26206 2468 29552 2496
rect 16853 2431 16911 2437
rect 16853 2397 16865 2431
rect 16899 2397 16911 2431
rect 16853 2391 16911 2397
rect 21821 2431 21879 2437
rect 21821 2397 21833 2431
rect 21867 2428 21879 2431
rect 26206 2428 26234 2468
rect 29546 2456 29552 2468
rect 29604 2456 29610 2508
rect 28810 2428 28816 2440
rect 21867 2400 26234 2428
rect 28771 2400 28816 2428
rect 21867 2397 21879 2400
rect 21821 2391 21879 2397
rect 28810 2388 28816 2400
rect 28868 2388 28874 2440
rect 15378 2360 15384 2372
rect 13188 2332 15384 2360
rect 6549 2323 6607 2329
rect 15378 2320 15384 2332
rect 15436 2320 15442 2372
rect 18046 2320 18052 2372
rect 18104 2360 18110 2372
rect 18233 2363 18291 2369
rect 18233 2360 18245 2363
rect 18104 2332 18245 2360
rect 18104 2320 18110 2332
rect 18233 2329 18245 2332
rect 18279 2329 18291 2363
rect 18233 2323 18291 2329
rect 3292 2264 5672 2292
rect 29656 2292 29684 2536
rect 29748 2536 30472 2564
rect 29748 2505 29776 2536
rect 30466 2524 30472 2536
rect 30524 2524 30530 2576
rect 29733 2499 29791 2505
rect 29733 2465 29745 2499
rect 29779 2465 29791 2499
rect 29914 2496 29920 2508
rect 29875 2468 29920 2496
rect 29733 2459 29791 2465
rect 29914 2456 29920 2468
rect 29972 2456 29978 2508
rect 30190 2456 30196 2508
rect 30248 2496 30254 2508
rect 31573 2499 31631 2505
rect 30248 2468 31156 2496
rect 30248 2456 30254 2468
rect 31128 2428 31156 2468
rect 31573 2465 31585 2499
rect 31619 2496 31631 2499
rect 32858 2496 32864 2508
rect 31619 2468 32864 2496
rect 31619 2465 31631 2468
rect 31573 2459 31631 2465
rect 32858 2456 32864 2468
rect 32916 2456 32922 2508
rect 32309 2431 32367 2437
rect 32309 2428 32321 2431
rect 31128 2400 32321 2428
rect 32309 2397 32321 2400
rect 32355 2397 32367 2431
rect 32309 2391 32367 2397
rect 30834 2320 30840 2372
rect 30892 2360 30898 2372
rect 32493 2363 32551 2369
rect 32493 2360 32505 2363
rect 30892 2332 32505 2360
rect 30892 2320 30898 2332
rect 32493 2329 32505 2332
rect 32539 2329 32551 2363
rect 32493 2323 32551 2329
rect 34149 2363 34207 2369
rect 34149 2329 34161 2363
rect 34195 2360 34207 2363
rect 34422 2360 34428 2372
rect 34195 2332 34428 2360
rect 34195 2329 34207 2332
rect 34149 2323 34207 2329
rect 34422 2320 34428 2332
rect 34480 2320 34486 2372
rect 33594 2292 33600 2304
rect 29656 2264 33600 2292
rect 3292 2252 3298 2264
rect 33594 2252 33600 2264
rect 33652 2252 33658 2304
rect 1104 2202 34868 2224
rect 1104 2150 12214 2202
rect 12266 2150 12278 2202
rect 12330 2150 12342 2202
rect 12394 2150 12406 2202
rect 12458 2150 12470 2202
rect 12522 2150 23478 2202
rect 23530 2150 23542 2202
rect 23594 2150 23606 2202
rect 23658 2150 23670 2202
rect 23722 2150 23734 2202
rect 23786 2150 34868 2202
rect 1104 2128 34868 2150
<< via1 >>
rect 13636 40876 13688 40928
rect 20168 40876 20220 40928
rect 12072 40808 12124 40860
rect 30380 40808 30432 40860
rect 4436 40740 4488 40792
rect 18604 40740 18656 40792
rect 14740 40672 14792 40724
rect 19892 40672 19944 40724
rect 11704 40604 11756 40656
rect 12992 40604 13044 40656
rect 26424 40604 26476 40656
rect 12624 40536 12676 40588
rect 31852 40536 31904 40588
rect 16028 40468 16080 40520
rect 29920 40468 29972 40520
rect 15384 40400 15436 40452
rect 30104 40400 30156 40452
rect 14464 40332 14516 40384
rect 30288 40332 30340 40384
rect 30012 40264 30064 40316
rect 15844 40196 15896 40248
rect 19800 40196 19852 40248
rect 19892 40196 19944 40248
rect 27252 40196 27304 40248
rect 13544 40128 13596 40180
rect 31944 40128 31996 40180
rect 12716 40060 12768 40112
rect 15936 40060 15988 40112
rect 19616 40060 19668 40112
rect 11796 39992 11848 40044
rect 19248 39992 19300 40044
rect 22652 39992 22704 40044
rect 29644 39992 29696 40044
rect 12256 39924 12308 39976
rect 22192 39924 22244 39976
rect 23756 39924 23808 39976
rect 32496 39924 32548 39976
rect 13912 39856 13964 39908
rect 18880 39856 18932 39908
rect 18972 39856 19024 39908
rect 26700 39856 26752 39908
rect 12900 39788 12952 39840
rect 17776 39788 17828 39840
rect 20812 39788 20864 39840
rect 27896 39788 27948 39840
rect 6582 39686 6634 39738
rect 6646 39686 6698 39738
rect 6710 39686 6762 39738
rect 6774 39686 6826 39738
rect 6838 39686 6890 39738
rect 17846 39686 17898 39738
rect 17910 39686 17962 39738
rect 17974 39686 18026 39738
rect 18038 39686 18090 39738
rect 18102 39686 18154 39738
rect 29110 39686 29162 39738
rect 29174 39686 29226 39738
rect 29238 39686 29290 39738
rect 29302 39686 29354 39738
rect 29366 39686 29418 39738
rect 10324 39627 10376 39636
rect 10324 39593 10333 39627
rect 10333 39593 10367 39627
rect 10367 39593 10376 39627
rect 10324 39584 10376 39593
rect 8300 39516 8352 39568
rect 9588 39516 9640 39568
rect 12256 39559 12308 39568
rect 12256 39525 12265 39559
rect 12265 39525 12299 39559
rect 12299 39525 12308 39559
rect 12256 39516 12308 39525
rect 4988 39448 5040 39500
rect 16396 39584 16448 39636
rect 17316 39584 17368 39636
rect 19064 39584 19116 39636
rect 23756 39627 23808 39636
rect 16304 39516 16356 39568
rect 23756 39593 23765 39627
rect 23765 39593 23799 39627
rect 23799 39593 23808 39627
rect 23756 39584 23808 39593
rect 25688 39584 25740 39636
rect 26240 39584 26292 39636
rect 26424 39627 26476 39636
rect 26424 39593 26433 39627
rect 26433 39593 26467 39627
rect 26467 39593 26476 39627
rect 26424 39584 26476 39593
rect 26516 39584 26568 39636
rect 31576 39584 31628 39636
rect 13544 39491 13596 39500
rect 13544 39457 13553 39491
rect 13553 39457 13587 39491
rect 13587 39457 13596 39491
rect 16672 39491 16724 39500
rect 13544 39448 13596 39457
rect 1400 39423 1452 39432
rect 1400 39389 1409 39423
rect 1409 39389 1443 39423
rect 1443 39389 1452 39423
rect 1400 39380 1452 39389
rect 3608 39380 3660 39432
rect 4068 39380 4120 39432
rect 4620 39423 4672 39432
rect 4620 39389 4629 39423
rect 4629 39389 4663 39423
rect 4663 39389 4672 39423
rect 4620 39380 4672 39389
rect 5264 39423 5316 39432
rect 5264 39389 5273 39423
rect 5273 39389 5307 39423
rect 5307 39389 5316 39423
rect 5264 39380 5316 39389
rect 5356 39380 5408 39432
rect 7196 39380 7248 39432
rect 8576 39380 8628 39432
rect 10968 39423 11020 39432
rect 10968 39389 10977 39423
rect 10977 39389 11011 39423
rect 11011 39389 11020 39423
rect 10968 39380 11020 39389
rect 13452 39380 13504 39432
rect 13820 39380 13872 39432
rect 14464 39423 14516 39432
rect 14464 39389 14473 39423
rect 14473 39389 14507 39423
rect 14507 39389 14516 39423
rect 14464 39380 14516 39389
rect 14924 39380 14976 39432
rect 15200 39380 15252 39432
rect 16672 39457 16681 39491
rect 16681 39457 16715 39491
rect 16715 39457 16724 39491
rect 16672 39448 16724 39457
rect 17408 39491 17460 39500
rect 17408 39457 17417 39491
rect 17417 39457 17451 39491
rect 17451 39457 17460 39491
rect 17408 39448 17460 39457
rect 17500 39448 17552 39500
rect 19984 39491 20036 39500
rect 19984 39457 19993 39491
rect 19993 39457 20027 39491
rect 20027 39457 20036 39491
rect 19984 39448 20036 39457
rect 25228 39516 25280 39568
rect 26792 39516 26844 39568
rect 30196 39516 30248 39568
rect 18052 39380 18104 39432
rect 19340 39380 19392 39432
rect 21916 39423 21968 39432
rect 21916 39389 21925 39423
rect 21925 39389 21959 39423
rect 21959 39389 21968 39423
rect 21916 39380 21968 39389
rect 22008 39423 22060 39432
rect 22008 39389 22017 39423
rect 22017 39389 22051 39423
rect 22051 39389 22060 39423
rect 22652 39423 22704 39432
rect 22008 39380 22060 39389
rect 22652 39389 22661 39423
rect 22661 39389 22695 39423
rect 22695 39389 22704 39423
rect 22652 39380 22704 39389
rect 23664 39423 23716 39432
rect 23664 39389 23673 39423
rect 23673 39389 23707 39423
rect 23707 39389 23716 39423
rect 23664 39380 23716 39389
rect 24584 39423 24636 39432
rect 24584 39389 24593 39423
rect 24593 39389 24627 39423
rect 24627 39389 24636 39423
rect 24584 39380 24636 39389
rect 26148 39423 26200 39432
rect 7012 39312 7064 39364
rect 7932 39312 7984 39364
rect 12716 39312 12768 39364
rect 15660 39312 15712 39364
rect 16120 39355 16172 39364
rect 16120 39321 16129 39355
rect 16129 39321 16163 39355
rect 16163 39321 16172 39355
rect 16120 39312 16172 39321
rect 16580 39312 16632 39364
rect 17316 39312 17368 39364
rect 18788 39312 18840 39364
rect 19432 39312 19484 39364
rect 20444 39312 20496 39364
rect 22836 39312 22888 39364
rect 26148 39389 26157 39423
rect 26157 39389 26191 39423
rect 26191 39389 26200 39423
rect 26148 39380 26200 39389
rect 26240 39423 26292 39432
rect 26240 39389 26249 39423
rect 26249 39389 26283 39423
rect 26283 39389 26292 39423
rect 26240 39380 26292 39389
rect 3148 39287 3200 39296
rect 3148 39253 3157 39287
rect 3157 39253 3191 39287
rect 3191 39253 3200 39287
rect 3148 39244 3200 39253
rect 3240 39244 3292 39296
rect 15200 39287 15252 39296
rect 15200 39253 15209 39287
rect 15209 39253 15243 39287
rect 15243 39253 15252 39287
rect 15200 39244 15252 39253
rect 15568 39244 15620 39296
rect 16396 39244 16448 39296
rect 16488 39244 16540 39296
rect 18972 39244 19024 39296
rect 20720 39244 20772 39296
rect 23848 39244 23900 39296
rect 26056 39312 26108 39364
rect 27160 39448 27212 39500
rect 30472 39448 30524 39500
rect 26976 39423 27028 39432
rect 26976 39389 26985 39423
rect 26985 39389 27019 39423
rect 27019 39389 27028 39423
rect 26976 39380 27028 39389
rect 34152 39491 34204 39500
rect 34152 39457 34161 39491
rect 34161 39457 34195 39491
rect 34195 39457 34204 39491
rect 34152 39448 34204 39457
rect 29460 39312 29512 39364
rect 30840 39380 30892 39432
rect 32312 39423 32364 39432
rect 32312 39389 32321 39423
rect 32321 39389 32355 39423
rect 32355 39389 32364 39423
rect 32312 39380 32364 39389
rect 30932 39312 30984 39364
rect 28908 39244 28960 39296
rect 30840 39244 30892 39296
rect 12214 39142 12266 39194
rect 12278 39142 12330 39194
rect 12342 39142 12394 39194
rect 12406 39142 12458 39194
rect 12470 39142 12522 39194
rect 23478 39142 23530 39194
rect 23542 39142 23594 39194
rect 23606 39142 23658 39194
rect 23670 39142 23722 39194
rect 23734 39142 23786 39194
rect 4620 39040 4672 39092
rect 12900 39083 12952 39092
rect 3148 38972 3200 39024
rect 4068 38972 4120 39024
rect 7932 38947 7984 38956
rect 1676 38879 1728 38888
rect 1676 38845 1685 38879
rect 1685 38845 1719 38879
rect 1719 38845 1728 38879
rect 1676 38836 1728 38845
rect 664 38768 716 38820
rect 5356 38836 5408 38888
rect 4160 38768 4212 38820
rect 7012 38836 7064 38888
rect 7932 38913 7941 38947
rect 7941 38913 7975 38947
rect 7975 38913 7984 38947
rect 7932 38904 7984 38913
rect 8576 38947 8628 38956
rect 8576 38913 8585 38947
rect 8585 38913 8619 38947
rect 8619 38913 8628 38947
rect 8576 38904 8628 38913
rect 11796 38947 11848 38956
rect 11796 38913 11805 38947
rect 11805 38913 11839 38947
rect 11839 38913 11848 38947
rect 11796 38904 11848 38913
rect 12624 38904 12676 38956
rect 9220 38836 9272 38888
rect 9312 38879 9364 38888
rect 9312 38845 9321 38879
rect 9321 38845 9355 38879
rect 9355 38845 9364 38879
rect 12900 39049 12909 39083
rect 12909 39049 12943 39083
rect 12943 39049 12952 39083
rect 12900 39040 12952 39049
rect 13452 39040 13504 39092
rect 13728 39040 13780 39092
rect 14924 39040 14976 39092
rect 15200 39040 15252 39092
rect 16120 38972 16172 39024
rect 13820 38904 13872 38956
rect 14188 38879 14240 38888
rect 9312 38836 9364 38845
rect 14188 38845 14197 38879
rect 14197 38845 14231 38879
rect 14231 38845 14240 38879
rect 14188 38836 14240 38845
rect 14372 38879 14424 38888
rect 14372 38845 14381 38879
rect 14381 38845 14415 38879
rect 14415 38845 14424 38879
rect 14372 38836 14424 38845
rect 14832 38879 14884 38888
rect 14832 38845 14841 38879
rect 14841 38845 14875 38879
rect 14875 38845 14884 38879
rect 14832 38836 14884 38845
rect 15108 38836 15160 38888
rect 15752 38836 15804 38888
rect 16488 38836 16540 38888
rect 8300 38768 8352 38820
rect 17132 38904 17184 38956
rect 16948 38836 17000 38888
rect 18052 38972 18104 39024
rect 18788 39040 18840 39092
rect 20996 39040 21048 39092
rect 22100 39040 22152 39092
rect 26792 39040 26844 39092
rect 30380 39083 30432 39092
rect 27252 39015 27304 39024
rect 27252 38981 27261 39015
rect 27261 38981 27295 39015
rect 27295 38981 27304 39015
rect 27252 38972 27304 38981
rect 27896 39015 27948 39024
rect 27896 38981 27905 39015
rect 27905 38981 27939 39015
rect 27939 38981 27948 39015
rect 27896 38972 27948 38981
rect 30380 39049 30389 39083
rect 30389 39049 30423 39083
rect 30423 39049 30432 39083
rect 30380 39040 30432 39049
rect 29828 38972 29880 39024
rect 32496 39015 32548 39024
rect 32496 38981 32505 39015
rect 32505 38981 32539 39015
rect 32539 38981 32548 39015
rect 32496 38972 32548 38981
rect 18880 38904 18932 38956
rect 22192 38947 22244 38956
rect 18236 38879 18288 38888
rect 17224 38768 17276 38820
rect 18236 38845 18245 38879
rect 18245 38845 18279 38879
rect 18279 38845 18288 38879
rect 18236 38836 18288 38845
rect 18328 38836 18380 38888
rect 19708 38836 19760 38888
rect 19892 38879 19944 38888
rect 19892 38845 19901 38879
rect 19901 38845 19935 38879
rect 19935 38845 19944 38879
rect 19892 38836 19944 38845
rect 19340 38768 19392 38820
rect 6460 38700 6512 38752
rect 9128 38700 9180 38752
rect 9220 38700 9272 38752
rect 13728 38700 13780 38752
rect 13820 38700 13872 38752
rect 17316 38700 17368 38752
rect 22192 38913 22201 38947
rect 22201 38913 22235 38947
rect 22235 38913 22244 38947
rect 22192 38904 22244 38913
rect 24492 38947 24544 38956
rect 24492 38913 24501 38947
rect 24501 38913 24535 38947
rect 24535 38913 24544 38947
rect 24492 38904 24544 38913
rect 20996 38768 21048 38820
rect 22100 38768 22152 38820
rect 22468 38836 22520 38888
rect 22560 38836 22612 38888
rect 25136 38879 25188 38888
rect 25136 38845 25145 38879
rect 25145 38845 25179 38879
rect 25179 38845 25188 38879
rect 25136 38836 25188 38845
rect 27712 38879 27764 38888
rect 27712 38845 27721 38879
rect 27721 38845 27755 38879
rect 27755 38845 27764 38879
rect 27712 38836 27764 38845
rect 28356 38879 28408 38888
rect 28356 38845 28365 38879
rect 28365 38845 28399 38879
rect 28399 38845 28408 38879
rect 28356 38836 28408 38845
rect 28448 38836 28500 38888
rect 21088 38700 21140 38752
rect 21916 38700 21968 38752
rect 22560 38700 22612 38752
rect 23756 38700 23808 38752
rect 27528 38768 27580 38820
rect 31944 38904 31996 38956
rect 33508 38879 33560 38888
rect 33508 38845 33517 38879
rect 33517 38845 33551 38879
rect 33551 38845 33560 38879
rect 33508 38836 33560 38845
rect 31484 38768 31536 38820
rect 30656 38700 30708 38752
rect 6582 38598 6634 38650
rect 6646 38598 6698 38650
rect 6710 38598 6762 38650
rect 6774 38598 6826 38650
rect 6838 38598 6890 38650
rect 17846 38598 17898 38650
rect 17910 38598 17962 38650
rect 17974 38598 18026 38650
rect 18038 38598 18090 38650
rect 18102 38598 18154 38650
rect 29110 38598 29162 38650
rect 29174 38598 29226 38650
rect 29238 38598 29290 38650
rect 29302 38598 29354 38650
rect 29366 38598 29418 38650
rect 14188 38496 14240 38548
rect 14372 38496 14424 38548
rect 14648 38496 14700 38548
rect 18420 38496 18472 38548
rect 18788 38496 18840 38548
rect 19340 38539 19392 38548
rect 19340 38505 19349 38539
rect 19349 38505 19383 38539
rect 19383 38505 19392 38539
rect 19340 38496 19392 38505
rect 1860 38428 1912 38480
rect 1308 38360 1360 38412
rect 5632 38360 5684 38412
rect 5816 38403 5868 38412
rect 5816 38369 5825 38403
rect 5825 38369 5859 38403
rect 5859 38369 5868 38403
rect 5816 38360 5868 38369
rect 6460 38360 6512 38412
rect 7104 38403 7156 38412
rect 7104 38369 7113 38403
rect 7113 38369 7147 38403
rect 7147 38369 7156 38403
rect 7104 38360 7156 38369
rect 1584 38267 1636 38276
rect 1584 38233 1593 38267
rect 1593 38233 1627 38267
rect 1627 38233 1636 38267
rect 1584 38224 1636 38233
rect 5356 38224 5408 38276
rect 6736 38267 6788 38276
rect 6736 38233 6745 38267
rect 6745 38233 6779 38267
rect 6779 38233 6788 38267
rect 6736 38224 6788 38233
rect 8392 38428 8444 38480
rect 12256 38471 12308 38480
rect 9128 38403 9180 38412
rect 9128 38369 9137 38403
rect 9137 38369 9171 38403
rect 9171 38369 9180 38403
rect 9128 38360 9180 38369
rect 12256 38437 12265 38471
rect 12265 38437 12299 38471
rect 12299 38437 12308 38471
rect 12256 38428 12308 38437
rect 13452 38428 13504 38480
rect 17684 38428 17736 38480
rect 11336 38360 11388 38412
rect 13084 38360 13136 38412
rect 8116 38292 8168 38344
rect 12900 38335 12952 38344
rect 12900 38301 12909 38335
rect 12909 38301 12943 38335
rect 12943 38301 12952 38335
rect 12900 38292 12952 38301
rect 14648 38360 14700 38412
rect 15660 38403 15712 38412
rect 15660 38369 15669 38403
rect 15669 38369 15703 38403
rect 15703 38369 15712 38403
rect 15660 38360 15712 38369
rect 16116 38403 16168 38412
rect 16116 38369 16129 38403
rect 16129 38369 16163 38403
rect 16163 38369 16168 38403
rect 16116 38360 16168 38369
rect 17408 38360 17460 38412
rect 19708 38428 19760 38480
rect 21916 38428 21968 38480
rect 23756 38471 23808 38480
rect 23756 38437 23765 38471
rect 23765 38437 23799 38471
rect 23799 38437 23808 38471
rect 23756 38428 23808 38437
rect 24032 38428 24084 38480
rect 18144 38360 18196 38412
rect 19984 38360 20036 38412
rect 20260 38403 20312 38412
rect 20260 38369 20269 38403
rect 20269 38369 20303 38403
rect 20303 38369 20312 38403
rect 20260 38360 20312 38369
rect 20628 38360 20680 38412
rect 21732 38360 21784 38412
rect 22284 38360 22336 38412
rect 25780 38403 25832 38412
rect 25780 38369 25789 38403
rect 25789 38369 25823 38403
rect 25823 38369 25832 38403
rect 25780 38360 25832 38369
rect 28632 38403 28684 38412
rect 28632 38369 28641 38403
rect 28641 38369 28675 38403
rect 28675 38369 28684 38403
rect 28632 38360 28684 38369
rect 29000 38360 29052 38412
rect 31852 38360 31904 38412
rect 34152 38403 34204 38412
rect 34152 38369 34161 38403
rect 34161 38369 34195 38403
rect 34195 38369 34204 38403
rect 34152 38360 34204 38369
rect 14372 38335 14424 38344
rect 14372 38301 14381 38335
rect 14381 38301 14415 38335
rect 14415 38301 14424 38335
rect 14372 38292 14424 38301
rect 14464 38292 14516 38344
rect 16856 38292 16908 38344
rect 13268 38224 13320 38276
rect 5264 38156 5316 38208
rect 11612 38156 11664 38208
rect 12624 38156 12676 38208
rect 13084 38156 13136 38208
rect 16948 38224 17000 38276
rect 17132 38292 17184 38344
rect 17868 38292 17920 38344
rect 19064 38292 19116 38344
rect 19156 38292 19208 38344
rect 19340 38292 19392 38344
rect 22376 38335 22428 38344
rect 22376 38301 22385 38335
rect 22385 38301 22419 38335
rect 22419 38301 22428 38335
rect 22376 38292 22428 38301
rect 25136 38335 25188 38344
rect 25136 38301 25145 38335
rect 25145 38301 25179 38335
rect 25179 38301 25188 38335
rect 25136 38292 25188 38301
rect 26516 38292 26568 38344
rect 27528 38292 27580 38344
rect 28816 38292 28868 38344
rect 29552 38335 29604 38344
rect 29552 38301 29561 38335
rect 29561 38301 29595 38335
rect 29595 38301 29604 38335
rect 29552 38292 29604 38301
rect 13728 38156 13780 38208
rect 15016 38156 15068 38208
rect 15108 38156 15160 38208
rect 22192 38156 22244 38208
rect 22744 38224 22796 38276
rect 24768 38224 24820 38276
rect 25044 38224 25096 38276
rect 32496 38267 32548 38276
rect 32496 38233 32505 38267
rect 32505 38233 32539 38267
rect 32539 38233 32548 38267
rect 32496 38224 32548 38233
rect 24676 38156 24728 38208
rect 27804 38199 27856 38208
rect 27804 38165 27813 38199
rect 27813 38165 27847 38199
rect 27847 38165 27856 38199
rect 27804 38156 27856 38165
rect 12214 38054 12266 38106
rect 12278 38054 12330 38106
rect 12342 38054 12394 38106
rect 12406 38054 12458 38106
rect 12470 38054 12522 38106
rect 23478 38054 23530 38106
rect 23542 38054 23594 38106
rect 23606 38054 23658 38106
rect 23670 38054 23722 38106
rect 23734 38054 23786 38106
rect 1676 37952 1728 38004
rect 5356 37995 5408 38004
rect 5356 37961 5365 37995
rect 5365 37961 5399 37995
rect 5399 37961 5408 37995
rect 5356 37952 5408 37961
rect 6736 37952 6788 38004
rect 11612 37995 11664 38004
rect 11612 37961 11621 37995
rect 11621 37961 11655 37995
rect 11655 37961 11664 37995
rect 11612 37952 11664 37961
rect 12716 37952 12768 38004
rect 13912 37952 13964 38004
rect 14188 37952 14240 38004
rect 3240 37884 3292 37936
rect 10416 37884 10468 37936
rect 14464 37884 14516 37936
rect 1860 37859 1912 37868
rect 1860 37825 1869 37859
rect 1869 37825 1903 37859
rect 1903 37825 1912 37859
rect 1860 37816 1912 37825
rect 4804 37816 4856 37868
rect 5540 37816 5592 37868
rect 7196 37859 7248 37868
rect 7196 37825 7205 37859
rect 7205 37825 7239 37859
rect 7239 37825 7248 37859
rect 7196 37816 7248 37825
rect 10324 37859 10376 37868
rect 10324 37825 10333 37859
rect 10333 37825 10367 37859
rect 10367 37825 10376 37859
rect 10324 37816 10376 37825
rect 10968 37859 11020 37868
rect 10968 37825 10977 37859
rect 10977 37825 11011 37859
rect 11011 37825 11020 37859
rect 10968 37816 11020 37825
rect 12072 37816 12124 37868
rect 12440 37859 12492 37868
rect 12440 37825 12449 37859
rect 12449 37825 12483 37859
rect 12483 37825 12492 37859
rect 12440 37816 12492 37825
rect 2964 37748 3016 37800
rect 7380 37791 7432 37800
rect 7380 37757 7389 37791
rect 7389 37757 7423 37791
rect 7423 37757 7432 37791
rect 7380 37748 7432 37757
rect 7748 37791 7800 37800
rect 7748 37757 7757 37791
rect 7757 37757 7791 37791
rect 7791 37757 7800 37791
rect 7748 37748 7800 37757
rect 13820 37816 13872 37868
rect 14372 37816 14424 37868
rect 15016 37884 15068 37936
rect 18144 37884 18196 37936
rect 18236 37884 18288 37936
rect 15936 37859 15988 37868
rect 4620 37680 4672 37732
rect 9680 37723 9732 37732
rect 9680 37689 9689 37723
rect 9689 37689 9723 37723
rect 9723 37689 9732 37723
rect 9680 37680 9732 37689
rect 12716 37680 12768 37732
rect 13728 37680 13780 37732
rect 13912 37748 13964 37800
rect 15936 37825 15945 37859
rect 15945 37825 15979 37859
rect 15979 37825 15988 37859
rect 15936 37816 15988 37825
rect 16028 37859 16080 37868
rect 16028 37825 16037 37859
rect 16037 37825 16071 37859
rect 16071 37825 16080 37859
rect 16028 37816 16080 37825
rect 14924 37748 14976 37800
rect 16764 37816 16816 37868
rect 16948 37859 17000 37868
rect 16948 37825 16982 37859
rect 16982 37825 17000 37859
rect 16948 37816 17000 37825
rect 17224 37816 17276 37868
rect 18328 37816 18380 37868
rect 18788 37859 18840 37868
rect 18788 37825 18822 37859
rect 18822 37825 18840 37859
rect 19892 37884 19944 37936
rect 20996 37952 21048 38004
rect 23020 37952 23072 38004
rect 23388 37952 23440 38004
rect 24032 37995 24084 38004
rect 24032 37961 24041 37995
rect 24041 37961 24075 37995
rect 24075 37961 24084 37995
rect 24032 37952 24084 37961
rect 18788 37816 18840 37825
rect 20260 37816 20312 37868
rect 20536 37859 20588 37868
rect 20536 37825 20545 37859
rect 20545 37825 20579 37859
rect 20579 37825 20588 37859
rect 20536 37816 20588 37825
rect 22192 37884 22244 37936
rect 29920 37927 29972 37936
rect 29920 37893 29929 37927
rect 29929 37893 29963 37927
rect 29963 37893 29972 37927
rect 29920 37884 29972 37893
rect 33048 37884 33100 37936
rect 34060 37884 34112 37936
rect 22376 37816 22428 37868
rect 23020 37816 23072 37868
rect 24400 37816 24452 37868
rect 25688 37859 25740 37868
rect 25688 37825 25697 37859
rect 25697 37825 25731 37859
rect 25731 37825 25740 37859
rect 25688 37816 25740 37825
rect 27528 37816 27580 37868
rect 28908 37816 28960 37868
rect 32036 37816 32088 37868
rect 16580 37748 16632 37800
rect 17684 37748 17736 37800
rect 18236 37748 18288 37800
rect 18512 37791 18564 37800
rect 18512 37757 18521 37791
rect 18521 37757 18555 37791
rect 18555 37757 18564 37791
rect 18512 37748 18564 37757
rect 20996 37748 21048 37800
rect 25412 37748 25464 37800
rect 25872 37748 25924 37800
rect 26608 37748 26660 37800
rect 28540 37748 28592 37800
rect 29736 37791 29788 37800
rect 29736 37757 29745 37791
rect 29745 37757 29779 37791
rect 29779 37757 29788 37791
rect 29736 37748 29788 37757
rect 15568 37612 15620 37664
rect 17776 37612 17828 37664
rect 22836 37680 22888 37732
rect 22008 37612 22060 37664
rect 24584 37612 24636 37664
rect 24768 37612 24820 37664
rect 26240 37612 26292 37664
rect 6582 37510 6634 37562
rect 6646 37510 6698 37562
rect 6710 37510 6762 37562
rect 6774 37510 6826 37562
rect 6838 37510 6890 37562
rect 17846 37510 17898 37562
rect 17910 37510 17962 37562
rect 17974 37510 18026 37562
rect 18038 37510 18090 37562
rect 18102 37510 18154 37562
rect 29110 37510 29162 37562
rect 29174 37510 29226 37562
rect 29238 37510 29290 37562
rect 29302 37510 29354 37562
rect 29366 37510 29418 37562
rect 1584 37408 1636 37460
rect 7380 37451 7432 37460
rect 7380 37417 7389 37451
rect 7389 37417 7423 37451
rect 7423 37417 7432 37451
rect 7380 37408 7432 37417
rect 8116 37451 8168 37460
rect 8116 37417 8125 37451
rect 8125 37417 8159 37451
rect 8159 37417 8168 37451
rect 8116 37408 8168 37417
rect 9772 37408 9824 37460
rect 10876 37451 10928 37460
rect 10876 37417 10885 37451
rect 10885 37417 10919 37451
rect 10919 37417 10928 37451
rect 10876 37408 10928 37417
rect 12348 37408 12400 37460
rect 12440 37408 12492 37460
rect 16488 37408 16540 37460
rect 16856 37408 16908 37460
rect 17500 37408 17552 37460
rect 18236 37408 18288 37460
rect 18328 37408 18380 37460
rect 18696 37408 18748 37460
rect 19340 37451 19392 37460
rect 19340 37417 19349 37451
rect 19349 37417 19383 37451
rect 19383 37417 19392 37451
rect 19340 37408 19392 37417
rect 21456 37451 21508 37460
rect 21456 37417 21465 37451
rect 21465 37417 21499 37451
rect 21499 37417 21508 37451
rect 21456 37408 21508 37417
rect 2320 37204 2372 37256
rect 12624 37340 12676 37392
rect 15660 37340 15712 37392
rect 15752 37340 15804 37392
rect 16212 37340 16264 37392
rect 3332 37272 3384 37324
rect 5172 37272 5224 37324
rect 10232 37315 10284 37324
rect 10232 37281 10241 37315
rect 10241 37281 10275 37315
rect 10275 37281 10284 37315
rect 10232 37272 10284 37281
rect 3792 37247 3844 37256
rect 3792 37213 3801 37247
rect 3801 37213 3835 37247
rect 3835 37213 3844 37247
rect 3792 37204 3844 37213
rect 3056 37136 3108 37188
rect 4712 37136 4764 37188
rect 7012 37136 7064 37188
rect 12440 37136 12492 37188
rect 12900 37272 12952 37324
rect 17224 37340 17276 37392
rect 17684 37340 17736 37392
rect 26516 37408 26568 37460
rect 31208 37408 31260 37460
rect 26332 37340 26384 37392
rect 18328 37315 18380 37324
rect 13176 37204 13228 37256
rect 13268 37247 13320 37256
rect 13268 37213 13277 37247
rect 13277 37213 13311 37247
rect 13311 37213 13320 37247
rect 14372 37247 14424 37256
rect 13268 37204 13320 37213
rect 14372 37213 14381 37247
rect 14381 37213 14415 37247
rect 14415 37213 14424 37247
rect 14372 37204 14424 37213
rect 15844 37204 15896 37256
rect 17040 37247 17092 37256
rect 17040 37213 17049 37247
rect 17049 37213 17083 37247
rect 17083 37213 17092 37247
rect 17040 37204 17092 37213
rect 17500 37204 17552 37256
rect 18328 37281 18337 37315
rect 18337 37281 18371 37315
rect 18371 37281 18380 37315
rect 18328 37272 18380 37281
rect 19156 37272 19208 37324
rect 19800 37272 19852 37324
rect 21088 37315 21140 37324
rect 21088 37281 21097 37315
rect 21097 37281 21131 37315
rect 21131 37281 21140 37315
rect 21088 37272 21140 37281
rect 21732 37272 21784 37324
rect 22376 37315 22428 37324
rect 22376 37281 22385 37315
rect 22385 37281 22419 37315
rect 22419 37281 22428 37315
rect 22376 37272 22428 37281
rect 24124 37272 24176 37324
rect 24676 37272 24728 37324
rect 32864 37315 32916 37324
rect 18604 37204 18656 37256
rect 19248 37204 19300 37256
rect 15016 37179 15068 37188
rect 11980 37111 12032 37120
rect 11980 37077 11989 37111
rect 11989 37077 12023 37111
rect 12023 37077 12032 37111
rect 11980 37068 12032 37077
rect 12624 37111 12676 37120
rect 12624 37077 12633 37111
rect 12633 37077 12667 37111
rect 12667 37077 12676 37111
rect 12624 37068 12676 37077
rect 14372 37068 14424 37120
rect 15016 37145 15025 37179
rect 15025 37145 15059 37179
rect 15059 37145 15068 37179
rect 15016 37136 15068 37145
rect 16212 37179 16264 37188
rect 16212 37145 16221 37179
rect 16221 37145 16255 37179
rect 16255 37145 16264 37179
rect 16212 37136 16264 37145
rect 16396 37136 16448 37188
rect 16672 37068 16724 37120
rect 17316 37136 17368 37188
rect 19892 37204 19944 37256
rect 20260 37247 20312 37256
rect 20260 37213 20269 37247
rect 20269 37213 20303 37247
rect 20303 37213 20312 37247
rect 20260 37204 20312 37213
rect 20352 37204 20404 37256
rect 20812 37204 20864 37256
rect 21364 37204 21416 37256
rect 24308 37204 24360 37256
rect 32864 37281 32873 37315
rect 32873 37281 32907 37315
rect 32907 37281 32916 37315
rect 32864 37272 32916 37281
rect 27160 37204 27212 37256
rect 28908 37204 28960 37256
rect 30656 37247 30708 37256
rect 30656 37213 30665 37247
rect 30665 37213 30699 37247
rect 30699 37213 30708 37247
rect 30656 37204 30708 37213
rect 32128 37247 32180 37256
rect 32128 37213 32137 37247
rect 32137 37213 32171 37247
rect 32171 37213 32180 37247
rect 32128 37204 32180 37213
rect 17592 37068 17644 37120
rect 18328 37068 18380 37120
rect 20720 37136 20772 37188
rect 19708 37068 19760 37120
rect 20260 37068 20312 37120
rect 21548 37068 21600 37120
rect 23296 37068 23348 37120
rect 24860 37136 24912 37188
rect 26240 37136 26292 37188
rect 26332 37136 26384 37188
rect 25320 37068 25372 37120
rect 30564 37136 30616 37188
rect 31300 37179 31352 37188
rect 31300 37145 31309 37179
rect 31309 37145 31343 37179
rect 31343 37145 31352 37179
rect 31300 37136 31352 37145
rect 32312 37179 32364 37188
rect 28448 37068 28500 37120
rect 28724 37111 28776 37120
rect 28724 37077 28733 37111
rect 28733 37077 28767 37111
rect 28767 37077 28776 37111
rect 28724 37068 28776 37077
rect 31668 37111 31720 37120
rect 31668 37077 31677 37111
rect 31677 37077 31711 37111
rect 31711 37077 31720 37111
rect 31668 37068 31720 37077
rect 32312 37145 32321 37179
rect 32321 37145 32355 37179
rect 32355 37145 32364 37179
rect 32312 37136 32364 37145
rect 33416 37068 33468 37120
rect 12214 36966 12266 37018
rect 12278 36966 12330 37018
rect 12342 36966 12394 37018
rect 12406 36966 12458 37018
rect 12470 36966 12522 37018
rect 23478 36966 23530 37018
rect 23542 36966 23594 37018
rect 23606 36966 23658 37018
rect 23670 36966 23722 37018
rect 23734 36966 23786 37018
rect 4712 36864 4764 36916
rect 7932 36864 7984 36916
rect 10876 36864 10928 36916
rect 13452 36864 13504 36916
rect 3976 36839 4028 36848
rect 3976 36805 3985 36839
rect 3985 36805 4019 36839
rect 4019 36805 4028 36839
rect 3976 36796 4028 36805
rect 5080 36839 5132 36848
rect 5080 36805 5089 36839
rect 5089 36805 5123 36839
rect 5123 36805 5132 36839
rect 5080 36796 5132 36805
rect 5540 36796 5592 36848
rect 3792 36728 3844 36780
rect 5632 36728 5684 36780
rect 10416 36728 10468 36780
rect 10784 36728 10836 36780
rect 12900 36796 12952 36848
rect 12440 36771 12492 36780
rect 12440 36737 12449 36771
rect 12449 36737 12483 36771
rect 12483 36737 12492 36771
rect 12440 36728 12492 36737
rect 16396 36796 16448 36848
rect 16672 36864 16724 36916
rect 21364 36864 21416 36916
rect 22008 36864 22060 36916
rect 22928 36864 22980 36916
rect 31116 36864 31168 36916
rect 32496 36864 32548 36916
rect 17040 36796 17092 36848
rect 17224 36796 17276 36848
rect 13912 36728 13964 36780
rect 14372 36771 14424 36780
rect 14372 36737 14381 36771
rect 14381 36737 14415 36771
rect 14415 36737 14424 36771
rect 14372 36728 14424 36737
rect 3884 36660 3936 36712
rect 2688 36592 2740 36644
rect 4804 36592 4856 36644
rect 12072 36592 12124 36644
rect 12164 36524 12216 36576
rect 14556 36703 14608 36712
rect 14556 36669 14565 36703
rect 14565 36669 14599 36703
rect 14599 36669 14608 36703
rect 15200 36728 15252 36780
rect 15936 36771 15988 36780
rect 15936 36737 15945 36771
rect 15945 36737 15979 36771
rect 15979 36737 15988 36771
rect 15936 36728 15988 36737
rect 16028 36771 16080 36780
rect 16028 36737 16037 36771
rect 16037 36737 16071 36771
rect 16071 36737 16080 36771
rect 16028 36728 16080 36737
rect 16304 36728 16356 36780
rect 18236 36728 18288 36780
rect 18512 36771 18564 36780
rect 18512 36737 18521 36771
rect 18521 36737 18555 36771
rect 18555 36737 18564 36771
rect 18512 36728 18564 36737
rect 14556 36660 14608 36669
rect 16396 36660 16448 36712
rect 16672 36703 16724 36712
rect 16672 36669 16681 36703
rect 16681 36669 16715 36703
rect 16715 36669 16724 36703
rect 16672 36660 16724 36669
rect 21548 36796 21600 36848
rect 21732 36796 21784 36848
rect 18788 36771 18840 36780
rect 18788 36737 18811 36771
rect 18811 36737 18840 36771
rect 18788 36728 18840 36737
rect 19156 36728 19208 36780
rect 16488 36592 16540 36644
rect 12716 36524 12768 36576
rect 19524 36660 19576 36712
rect 19892 36660 19944 36712
rect 20628 36728 20680 36780
rect 21180 36728 21232 36780
rect 21824 36771 21876 36780
rect 21824 36737 21833 36771
rect 21833 36737 21867 36771
rect 21867 36737 21876 36771
rect 21824 36728 21876 36737
rect 22560 36728 22612 36780
rect 22836 36796 22888 36848
rect 23204 36796 23256 36848
rect 23388 36771 23440 36780
rect 23388 36737 23397 36771
rect 23397 36737 23431 36771
rect 23431 36737 23440 36771
rect 23388 36728 23440 36737
rect 23480 36728 23532 36780
rect 25780 36796 25832 36848
rect 26608 36796 26660 36848
rect 26700 36796 26752 36848
rect 17776 36592 17828 36644
rect 18420 36524 18472 36576
rect 21548 36592 21600 36644
rect 24400 36771 24452 36780
rect 24400 36737 24409 36771
rect 24409 36737 24443 36771
rect 24443 36737 24452 36771
rect 25872 36771 25924 36780
rect 24400 36728 24452 36737
rect 25872 36737 25881 36771
rect 25881 36737 25915 36771
rect 25915 36737 25924 36771
rect 25872 36728 25924 36737
rect 25964 36728 26016 36780
rect 32312 36796 32364 36848
rect 28908 36728 28960 36780
rect 30288 36771 30340 36780
rect 30288 36737 30297 36771
rect 30297 36737 30331 36771
rect 30331 36737 30340 36771
rect 30288 36728 30340 36737
rect 31392 36771 31444 36780
rect 31392 36737 31401 36771
rect 31401 36737 31435 36771
rect 31435 36737 31444 36771
rect 31392 36728 31444 36737
rect 31852 36728 31904 36780
rect 34152 36771 34204 36780
rect 34152 36737 34161 36771
rect 34161 36737 34195 36771
rect 34195 36737 34204 36771
rect 34152 36728 34204 36737
rect 24676 36660 24728 36712
rect 26516 36660 26568 36712
rect 27160 36703 27212 36712
rect 27160 36669 27169 36703
rect 27169 36669 27203 36703
rect 27203 36669 27212 36703
rect 27160 36660 27212 36669
rect 28172 36660 28224 36712
rect 30564 36703 30616 36712
rect 23572 36592 23624 36644
rect 23664 36592 23716 36644
rect 19892 36567 19944 36576
rect 19892 36533 19901 36567
rect 19901 36533 19935 36567
rect 19935 36533 19944 36567
rect 20720 36567 20772 36576
rect 19892 36524 19944 36533
rect 20720 36533 20729 36567
rect 20729 36533 20763 36567
rect 20763 36533 20772 36567
rect 20720 36524 20772 36533
rect 22744 36567 22796 36576
rect 22744 36533 22753 36567
rect 22753 36533 22787 36567
rect 22787 36533 22796 36567
rect 22744 36524 22796 36533
rect 22928 36567 22980 36576
rect 22928 36533 22937 36567
rect 22937 36533 22971 36567
rect 22971 36533 22980 36567
rect 22928 36524 22980 36533
rect 23112 36524 23164 36576
rect 23480 36524 23532 36576
rect 23756 36567 23808 36576
rect 23756 36533 23765 36567
rect 23765 36533 23799 36567
rect 23799 36533 23808 36567
rect 23756 36524 23808 36533
rect 24308 36592 24360 36644
rect 25320 36524 25372 36576
rect 25412 36524 25464 36576
rect 25688 36524 25740 36576
rect 27804 36524 27856 36576
rect 28356 36524 28408 36576
rect 30564 36669 30573 36703
rect 30573 36669 30607 36703
rect 30607 36669 30616 36703
rect 30564 36660 30616 36669
rect 31024 36660 31076 36712
rect 31944 36660 31996 36712
rect 29736 36592 29788 36644
rect 30564 36524 30616 36576
rect 30656 36524 30708 36576
rect 34336 36524 34388 36576
rect 6582 36422 6634 36474
rect 6646 36422 6698 36474
rect 6710 36422 6762 36474
rect 6774 36422 6826 36474
rect 6838 36422 6890 36474
rect 17846 36422 17898 36474
rect 17910 36422 17962 36474
rect 17974 36422 18026 36474
rect 18038 36422 18090 36474
rect 18102 36422 18154 36474
rect 29110 36422 29162 36474
rect 29174 36422 29226 36474
rect 29238 36422 29290 36474
rect 29302 36422 29354 36474
rect 29366 36422 29418 36474
rect 2320 36320 2372 36372
rect 4988 36363 5040 36372
rect 2688 36252 2740 36304
rect 4988 36329 4997 36363
rect 4997 36329 5031 36363
rect 5031 36329 5040 36363
rect 4988 36320 5040 36329
rect 10876 36320 10928 36372
rect 2412 36184 2464 36236
rect 2780 36227 2832 36236
rect 2780 36193 2789 36227
rect 2789 36193 2823 36227
rect 2823 36193 2832 36227
rect 2780 36184 2832 36193
rect 11428 36252 11480 36304
rect 11612 36295 11664 36304
rect 11612 36261 11621 36295
rect 11621 36261 11655 36295
rect 11655 36261 11664 36295
rect 11612 36252 11664 36261
rect 13636 36320 13688 36372
rect 13912 36320 13964 36372
rect 15844 36320 15896 36372
rect 16120 36320 16172 36372
rect 16212 36320 16264 36372
rect 16948 36320 17000 36372
rect 18696 36363 18748 36372
rect 12900 36252 12952 36304
rect 16396 36252 16448 36304
rect 12348 36184 12400 36236
rect 12440 36184 12492 36236
rect 17316 36252 17368 36304
rect 18696 36329 18705 36363
rect 18705 36329 18739 36363
rect 18739 36329 18748 36363
rect 18696 36320 18748 36329
rect 20720 36320 20772 36372
rect 21548 36320 21600 36372
rect 23756 36320 23808 36372
rect 24032 36320 24084 36372
rect 23296 36252 23348 36304
rect 23572 36295 23624 36304
rect 23572 36261 23581 36295
rect 23581 36261 23615 36295
rect 23615 36261 23624 36295
rect 23572 36252 23624 36261
rect 3516 36116 3568 36168
rect 3792 36116 3844 36168
rect 4436 36159 4488 36168
rect 4436 36125 4445 36159
rect 4445 36125 4479 36159
rect 4479 36125 4488 36159
rect 4436 36116 4488 36125
rect 5172 36159 5224 36168
rect 5172 36125 5181 36159
rect 5181 36125 5215 36159
rect 5215 36125 5224 36159
rect 5172 36116 5224 36125
rect 11336 36116 11388 36168
rect 12808 36116 12860 36168
rect 12900 36159 12952 36168
rect 12900 36125 12909 36159
rect 12909 36125 12943 36159
rect 12943 36125 12952 36159
rect 13544 36159 13596 36168
rect 12900 36116 12952 36125
rect 13544 36125 13553 36159
rect 13553 36125 13587 36159
rect 13587 36125 13596 36159
rect 13544 36116 13596 36125
rect 14372 36116 14424 36168
rect 14464 36116 14516 36168
rect 14924 36116 14976 36168
rect 15292 36116 15344 36168
rect 15476 36116 15528 36168
rect 16948 36184 17000 36236
rect 1584 36091 1636 36100
rect 1584 36057 1593 36091
rect 1593 36057 1627 36091
rect 1627 36057 1636 36091
rect 1584 36048 1636 36057
rect 13728 36048 13780 36100
rect 15200 36048 15252 36100
rect 15568 36048 15620 36100
rect 16764 36116 16816 36168
rect 18512 36184 18564 36236
rect 18696 36184 18748 36236
rect 16948 36048 17000 36100
rect 17132 36048 17184 36100
rect 17224 36048 17276 36100
rect 18972 36116 19024 36168
rect 20536 36184 20588 36236
rect 21272 36116 21324 36168
rect 12716 36023 12768 36032
rect 12716 35989 12725 36023
rect 12725 35989 12759 36023
rect 12759 35989 12768 36023
rect 12716 35980 12768 35989
rect 13360 36023 13412 36032
rect 13360 35989 13369 36023
rect 13369 35989 13403 36023
rect 13403 35989 13412 36023
rect 13360 35980 13412 35989
rect 13544 35980 13596 36032
rect 14372 35980 14424 36032
rect 15016 35980 15068 36032
rect 17776 36048 17828 36100
rect 22376 36116 22428 36168
rect 22744 36116 22796 36168
rect 24124 36184 24176 36236
rect 25872 36320 25924 36372
rect 25504 36252 25556 36304
rect 25688 36252 25740 36304
rect 25964 36184 26016 36236
rect 26148 36184 26200 36236
rect 28356 36320 28408 36372
rect 28448 36320 28500 36372
rect 29644 36320 29696 36372
rect 30012 36320 30064 36372
rect 27896 36252 27948 36304
rect 23480 36116 23532 36168
rect 28448 36184 28500 36236
rect 27804 36116 27856 36168
rect 29000 36184 29052 36236
rect 31116 36227 31168 36236
rect 31116 36193 31125 36227
rect 31125 36193 31159 36227
rect 31159 36193 31168 36227
rect 31116 36184 31168 36193
rect 32312 36227 32364 36236
rect 32312 36193 32321 36227
rect 32321 36193 32355 36227
rect 32355 36193 32364 36227
rect 32312 36184 32364 36193
rect 32956 36227 33008 36236
rect 32956 36193 32965 36227
rect 32965 36193 32999 36227
rect 32999 36193 33008 36227
rect 32956 36184 33008 36193
rect 17684 35980 17736 36032
rect 18512 35980 18564 36032
rect 18788 35980 18840 36032
rect 19984 35980 20036 36032
rect 25412 36048 25464 36100
rect 26608 36091 26660 36100
rect 26608 36057 26617 36091
rect 26617 36057 26651 36091
rect 26651 36057 26660 36091
rect 26608 36048 26660 36057
rect 29644 36159 29696 36168
rect 22376 35980 22428 36032
rect 22928 35980 22980 36032
rect 25964 35980 26016 36032
rect 26516 36023 26568 36032
rect 26516 35989 26525 36023
rect 26525 35989 26559 36023
rect 26559 35989 26568 36023
rect 26516 35980 26568 35989
rect 27620 35980 27672 36032
rect 28540 36091 28592 36100
rect 28540 36057 28549 36091
rect 28549 36057 28583 36091
rect 28583 36057 28592 36091
rect 28540 36048 28592 36057
rect 27896 36023 27948 36032
rect 27896 35989 27905 36023
rect 27905 35989 27939 36023
rect 27939 35989 27948 36023
rect 27896 35980 27948 35989
rect 28356 35980 28408 36032
rect 29644 36125 29653 36159
rect 29653 36125 29687 36159
rect 29687 36125 29696 36159
rect 29644 36116 29696 36125
rect 30288 36116 30340 36168
rect 30380 36048 30432 36100
rect 29552 35980 29604 36032
rect 12214 35878 12266 35930
rect 12278 35878 12330 35930
rect 12342 35878 12394 35930
rect 12406 35878 12458 35930
rect 12470 35878 12522 35930
rect 23478 35878 23530 35930
rect 23542 35878 23594 35930
rect 23606 35878 23658 35930
rect 23670 35878 23722 35930
rect 23734 35878 23786 35930
rect 1584 35776 1636 35828
rect 3516 35776 3568 35828
rect 11704 35776 11756 35828
rect 1400 35683 1452 35692
rect 1400 35649 1409 35683
rect 1409 35649 1443 35683
rect 1443 35649 1452 35683
rect 1400 35640 1452 35649
rect 2136 35683 2188 35692
rect 2136 35649 2145 35683
rect 2145 35649 2179 35683
rect 2179 35649 2188 35683
rect 2136 35640 2188 35649
rect 13268 35708 13320 35760
rect 3884 35640 3936 35692
rect 4620 35683 4672 35692
rect 4620 35649 4629 35683
rect 4629 35649 4663 35683
rect 4663 35649 4672 35683
rect 4620 35640 4672 35649
rect 13176 35640 13228 35692
rect 16764 35776 16816 35828
rect 18696 35776 18748 35828
rect 19340 35776 19392 35828
rect 17132 35708 17184 35760
rect 19708 35751 19760 35760
rect 19708 35717 19717 35751
rect 19717 35717 19751 35751
rect 19751 35717 19760 35751
rect 19708 35708 19760 35717
rect 19892 35708 19944 35760
rect 20076 35776 20128 35828
rect 20536 35776 20588 35828
rect 21364 35776 21416 35828
rect 20996 35708 21048 35760
rect 22100 35751 22152 35760
rect 22100 35717 22134 35751
rect 22134 35717 22152 35751
rect 22468 35776 22520 35828
rect 25780 35776 25832 35828
rect 29000 35776 29052 35828
rect 22100 35708 22152 35717
rect 13912 35572 13964 35624
rect 14372 35640 14424 35692
rect 15292 35640 15344 35692
rect 14924 35572 14976 35624
rect 15752 35615 15804 35624
rect 15752 35581 15761 35615
rect 15761 35581 15795 35615
rect 15795 35581 15804 35615
rect 15752 35572 15804 35581
rect 15936 35683 15988 35692
rect 15936 35649 15945 35683
rect 15945 35649 15979 35683
rect 15979 35649 15988 35683
rect 15936 35640 15988 35649
rect 16212 35640 16264 35692
rect 16396 35640 16448 35692
rect 16488 35572 16540 35624
rect 16672 35615 16724 35624
rect 16672 35581 16681 35615
rect 16681 35581 16715 35615
rect 16715 35581 16724 35615
rect 16672 35572 16724 35581
rect 17776 35640 17828 35692
rect 18420 35640 18472 35692
rect 18696 35683 18748 35692
rect 18696 35649 18705 35683
rect 18705 35649 18739 35683
rect 18739 35649 18748 35683
rect 18696 35640 18748 35649
rect 19800 35640 19852 35692
rect 12532 35547 12584 35556
rect 12532 35513 12541 35547
rect 12541 35513 12575 35547
rect 12575 35513 12584 35547
rect 12532 35504 12584 35513
rect 13176 35504 13228 35556
rect 19432 35572 19484 35624
rect 2136 35436 2188 35488
rect 13452 35436 13504 35488
rect 13820 35479 13872 35488
rect 13820 35445 13829 35479
rect 13829 35445 13863 35479
rect 13863 35445 13872 35479
rect 14464 35479 14516 35488
rect 13820 35436 13872 35445
rect 14464 35445 14473 35479
rect 14473 35445 14507 35479
rect 14507 35445 14516 35479
rect 14464 35436 14516 35445
rect 14924 35436 14976 35488
rect 17776 35436 17828 35488
rect 20076 35572 20128 35624
rect 20628 35640 20680 35692
rect 22376 35640 22428 35692
rect 22560 35640 22612 35692
rect 23572 35640 23624 35692
rect 24216 35708 24268 35760
rect 24124 35640 24176 35692
rect 21272 35572 21324 35624
rect 26240 35683 26292 35692
rect 26240 35649 26249 35683
rect 26249 35649 26283 35683
rect 26283 35649 26292 35683
rect 26240 35640 26292 35649
rect 27068 35640 27120 35692
rect 27160 35640 27212 35692
rect 25320 35572 25372 35624
rect 27896 35640 27948 35692
rect 28540 35640 28592 35692
rect 19524 35436 19576 35488
rect 20352 35436 20404 35488
rect 22928 35436 22980 35488
rect 23296 35436 23348 35488
rect 26700 35504 26752 35556
rect 29184 35708 29236 35760
rect 29920 35640 29972 35692
rect 25780 35436 25832 35488
rect 27988 35436 28040 35488
rect 31300 35708 31352 35760
rect 32496 35708 32548 35760
rect 32036 35640 32088 35692
rect 32404 35640 32456 35692
rect 33324 35683 33376 35692
rect 33324 35649 33333 35683
rect 33333 35649 33367 35683
rect 33367 35649 33376 35683
rect 33324 35640 33376 35649
rect 29460 35436 29512 35488
rect 30472 35436 30524 35488
rect 32220 35436 32272 35488
rect 6582 35334 6634 35386
rect 6646 35334 6698 35386
rect 6710 35334 6762 35386
rect 6774 35334 6826 35386
rect 6838 35334 6890 35386
rect 17846 35334 17898 35386
rect 17910 35334 17962 35386
rect 17974 35334 18026 35386
rect 18038 35334 18090 35386
rect 18102 35334 18154 35386
rect 29110 35334 29162 35386
rect 29174 35334 29226 35386
rect 29238 35334 29290 35386
rect 29302 35334 29354 35386
rect 29366 35334 29418 35386
rect 1768 35232 1820 35284
rect 2780 35139 2832 35148
rect 2780 35105 2789 35139
rect 2789 35105 2823 35139
rect 2823 35105 2832 35139
rect 2780 35096 2832 35105
rect 14096 35232 14148 35284
rect 15016 35232 15068 35284
rect 15752 35232 15804 35284
rect 16948 35275 17000 35284
rect 16948 35241 16957 35275
rect 16957 35241 16991 35275
rect 16991 35241 17000 35275
rect 16948 35232 17000 35241
rect 17132 35232 17184 35284
rect 18328 35232 18380 35284
rect 13176 35207 13228 35216
rect 13176 35173 13185 35207
rect 13185 35173 13219 35207
rect 13219 35173 13228 35207
rect 13176 35164 13228 35173
rect 14924 35207 14976 35216
rect 14924 35173 14933 35207
rect 14933 35173 14967 35207
rect 14967 35173 14976 35207
rect 14924 35164 14976 35173
rect 15200 35164 15252 35216
rect 14280 35096 14332 35148
rect 1400 35071 1452 35080
rect 1400 35037 1409 35071
rect 1409 35037 1443 35071
rect 1443 35037 1452 35071
rect 1400 35028 1452 35037
rect 2044 34960 2096 35012
rect 12808 35028 12860 35080
rect 13544 35028 13596 35080
rect 13912 35028 13964 35080
rect 15476 35096 15528 35148
rect 16580 35164 16632 35216
rect 20904 35232 20956 35284
rect 14648 35028 14700 35080
rect 15292 35028 15344 35080
rect 16672 35096 16724 35148
rect 17224 35096 17276 35148
rect 17316 35096 17368 35148
rect 19340 35164 19392 35216
rect 19616 35164 19668 35216
rect 20812 35164 20864 35216
rect 23388 35275 23440 35284
rect 23388 35241 23397 35275
rect 23397 35241 23431 35275
rect 23431 35241 23440 35275
rect 23388 35232 23440 35241
rect 23572 35232 23624 35284
rect 25320 35164 25372 35216
rect 27068 35164 27120 35216
rect 29644 35164 29696 35216
rect 18788 35096 18840 35148
rect 19156 35096 19208 35148
rect 17040 35028 17092 35080
rect 17500 35028 17552 35080
rect 17776 35028 17828 35080
rect 18420 35028 18472 35080
rect 18604 35028 18656 35080
rect 21088 35096 21140 35148
rect 21272 35096 21324 35148
rect 13820 34960 13872 35012
rect 15936 34960 15988 35012
rect 16580 34960 16632 35012
rect 17224 34960 17276 35012
rect 18972 34960 19024 35012
rect 19524 35071 19576 35080
rect 19524 35037 19533 35071
rect 19533 35037 19567 35071
rect 19567 35037 19576 35071
rect 19892 35071 19944 35080
rect 19524 35028 19576 35037
rect 19892 35037 19901 35071
rect 19901 35037 19935 35071
rect 19935 35037 19944 35071
rect 19892 35028 19944 35037
rect 19616 35003 19668 35012
rect 14372 34892 14424 34944
rect 14556 34892 14608 34944
rect 17040 34892 17092 34944
rect 17408 34892 17460 34944
rect 17776 34935 17828 34944
rect 17776 34901 17785 34935
rect 17785 34901 17819 34935
rect 17819 34901 17828 34935
rect 17776 34892 17828 34901
rect 19616 34969 19625 35003
rect 19625 34969 19659 35003
rect 19659 34969 19668 35003
rect 19616 34960 19668 34969
rect 20260 35028 20312 35080
rect 20444 35071 20496 35080
rect 20444 35037 20453 35071
rect 20453 35037 20487 35071
rect 20487 35037 20496 35071
rect 20444 35028 20496 35037
rect 20628 35028 20680 35080
rect 20812 35028 20864 35080
rect 20076 34960 20128 35012
rect 19156 34892 19208 34944
rect 19340 34892 19392 34944
rect 23296 35028 23348 35080
rect 23480 35028 23532 35080
rect 24584 35071 24636 35080
rect 23204 34960 23256 35012
rect 23020 34892 23072 34944
rect 24584 35037 24593 35071
rect 24593 35037 24627 35071
rect 24627 35037 24636 35071
rect 24584 35028 24636 35037
rect 24860 35096 24912 35148
rect 25136 35096 25188 35148
rect 26700 35096 26752 35148
rect 29368 35096 29420 35148
rect 26424 35028 26476 35080
rect 27620 35028 27672 35080
rect 27804 35071 27856 35080
rect 27804 35037 27813 35071
rect 27813 35037 27847 35071
rect 27847 35037 27856 35071
rect 27804 35028 27856 35037
rect 27988 35071 28040 35080
rect 27988 35037 28023 35071
rect 28023 35037 28040 35071
rect 27988 35028 28040 35037
rect 28172 35071 28224 35080
rect 28172 35037 28181 35071
rect 28181 35037 28215 35071
rect 28215 35037 28224 35071
rect 28172 35028 28224 35037
rect 23756 34960 23808 35012
rect 24676 35003 24728 35012
rect 23848 34935 23900 34944
rect 23848 34901 23857 34935
rect 23857 34901 23891 34935
rect 23891 34901 23900 34935
rect 23848 34892 23900 34901
rect 24400 34935 24452 34944
rect 24400 34901 24409 34935
rect 24409 34901 24443 34935
rect 24443 34901 24452 34935
rect 24400 34892 24452 34901
rect 24676 34969 24685 35003
rect 24685 34969 24719 35003
rect 24719 34969 24728 35003
rect 24676 34960 24728 34969
rect 24768 35003 24820 35012
rect 24768 34969 24777 35003
rect 24777 34969 24811 35003
rect 24811 34969 24820 35003
rect 24768 34960 24820 34969
rect 28356 34960 28408 35012
rect 28632 35003 28684 35012
rect 28632 34969 28641 35003
rect 28641 34969 28675 35003
rect 28675 34969 28684 35003
rect 28632 34960 28684 34969
rect 29644 35028 29696 35080
rect 30472 35164 30524 35216
rect 32404 35164 32456 35216
rect 33508 35164 33560 35216
rect 30472 35071 30524 35080
rect 30472 35037 30481 35071
rect 30481 35037 30515 35071
rect 30515 35037 30524 35071
rect 30472 35028 30524 35037
rect 31944 35028 31996 35080
rect 26148 34892 26200 34944
rect 27436 34892 27488 34944
rect 28540 34892 28592 34944
rect 30196 34960 30248 35012
rect 32128 34960 32180 35012
rect 34152 35003 34204 35012
rect 34152 34969 34161 35003
rect 34161 34969 34195 35003
rect 34195 34969 34204 35003
rect 34152 34960 34204 34969
rect 31300 34892 31352 34944
rect 32404 34892 32456 34944
rect 12214 34790 12266 34842
rect 12278 34790 12330 34842
rect 12342 34790 12394 34842
rect 12406 34790 12458 34842
rect 12470 34790 12522 34842
rect 23478 34790 23530 34842
rect 23542 34790 23594 34842
rect 23606 34790 23658 34842
rect 23670 34790 23722 34842
rect 23734 34790 23786 34842
rect 12716 34731 12768 34740
rect 12716 34697 12725 34731
rect 12725 34697 12759 34731
rect 12759 34697 12768 34731
rect 12716 34688 12768 34697
rect 13360 34731 13412 34740
rect 13360 34697 13369 34731
rect 13369 34697 13403 34731
rect 13403 34697 13412 34731
rect 13360 34688 13412 34697
rect 15016 34688 15068 34740
rect 15476 34688 15528 34740
rect 13636 34620 13688 34672
rect 15200 34620 15252 34672
rect 1400 34552 1452 34604
rect 12992 34552 13044 34604
rect 14188 34595 14240 34604
rect 14188 34561 14197 34595
rect 14197 34561 14231 34595
rect 14231 34561 14240 34595
rect 14188 34552 14240 34561
rect 14556 34552 14608 34604
rect 14740 34552 14792 34604
rect 15016 34552 15068 34604
rect 15752 34552 15804 34604
rect 14464 34484 14516 34536
rect 16488 34620 16540 34672
rect 16580 34620 16632 34672
rect 16764 34620 16816 34672
rect 20996 34688 21048 34740
rect 23388 34688 23440 34740
rect 23848 34688 23900 34740
rect 26148 34731 26200 34740
rect 16396 34552 16448 34604
rect 2412 34459 2464 34468
rect 2412 34425 2421 34459
rect 2421 34425 2455 34459
rect 2455 34425 2464 34459
rect 2412 34416 2464 34425
rect 12256 34459 12308 34468
rect 12256 34425 12265 34459
rect 12265 34425 12299 34459
rect 12299 34425 12308 34459
rect 12256 34416 12308 34425
rect 14004 34459 14056 34468
rect 14004 34425 14013 34459
rect 14013 34425 14047 34459
rect 14047 34425 14056 34459
rect 14004 34416 14056 34425
rect 16580 34484 16632 34536
rect 17040 34552 17092 34604
rect 18052 34620 18104 34672
rect 18236 34620 18288 34672
rect 18972 34620 19024 34672
rect 17592 34552 17644 34604
rect 17684 34527 17736 34536
rect 11888 34348 11940 34400
rect 14924 34416 14976 34468
rect 15200 34416 15252 34468
rect 15292 34416 15344 34468
rect 16304 34416 16356 34468
rect 16488 34416 16540 34468
rect 17224 34416 17276 34468
rect 17684 34493 17693 34527
rect 17693 34493 17727 34527
rect 17727 34493 17736 34527
rect 18696 34552 18748 34604
rect 19248 34552 19300 34604
rect 19708 34552 19760 34604
rect 19892 34595 19944 34604
rect 19892 34561 19926 34595
rect 19926 34561 19944 34595
rect 19892 34552 19944 34561
rect 17684 34484 17736 34493
rect 18788 34484 18840 34536
rect 18880 34484 18932 34536
rect 19524 34484 19576 34536
rect 21088 34620 21140 34672
rect 24400 34620 24452 34672
rect 26148 34697 26157 34731
rect 26157 34697 26191 34731
rect 26191 34697 26200 34731
rect 26148 34688 26200 34697
rect 31576 34688 31628 34740
rect 32128 34731 32180 34740
rect 32128 34697 32137 34731
rect 32137 34697 32171 34731
rect 32171 34697 32180 34731
rect 32128 34688 32180 34697
rect 32496 34688 32548 34740
rect 21272 34552 21324 34604
rect 22652 34552 22704 34604
rect 23756 34484 23808 34536
rect 25320 34552 25372 34604
rect 27344 34620 27396 34672
rect 28172 34620 28224 34672
rect 29368 34620 29420 34672
rect 29460 34620 29512 34672
rect 25964 34595 26016 34604
rect 25964 34561 25973 34595
rect 25973 34561 26007 34595
rect 26007 34561 26016 34595
rect 25964 34552 26016 34561
rect 27620 34552 27672 34604
rect 27896 34552 27948 34604
rect 28816 34595 28868 34604
rect 28816 34561 28825 34595
rect 28825 34561 28859 34595
rect 28859 34561 28868 34595
rect 28816 34552 28868 34561
rect 28908 34552 28960 34604
rect 30472 34620 30524 34672
rect 30748 34552 30800 34604
rect 31576 34552 31628 34604
rect 32312 34552 32364 34604
rect 32496 34595 32548 34604
rect 32496 34561 32505 34595
rect 32505 34561 32539 34595
rect 32539 34561 32548 34595
rect 32496 34552 32548 34561
rect 32680 34620 32732 34672
rect 33232 34663 33284 34672
rect 33232 34629 33241 34663
rect 33241 34629 33275 34663
rect 33275 34629 33284 34663
rect 33232 34620 33284 34629
rect 32772 34595 32824 34604
rect 32772 34561 32781 34595
rect 32781 34561 32815 34595
rect 32815 34561 32824 34595
rect 33416 34595 33468 34604
rect 32772 34552 32824 34561
rect 33416 34561 33425 34595
rect 33425 34561 33459 34595
rect 33459 34561 33468 34595
rect 33416 34552 33468 34561
rect 33692 34595 33744 34604
rect 33692 34561 33701 34595
rect 33701 34561 33735 34595
rect 33735 34561 33744 34595
rect 33692 34552 33744 34561
rect 27436 34484 27488 34536
rect 14188 34348 14240 34400
rect 17040 34348 17092 34400
rect 17408 34348 17460 34400
rect 18236 34416 18288 34468
rect 20996 34459 21048 34468
rect 19432 34348 19484 34400
rect 20996 34425 21005 34459
rect 21005 34425 21039 34459
rect 21039 34425 21048 34459
rect 20996 34416 21048 34425
rect 22100 34416 22152 34468
rect 21364 34348 21416 34400
rect 23572 34416 23624 34468
rect 23112 34348 23164 34400
rect 25320 34391 25372 34400
rect 25320 34357 25329 34391
rect 25329 34357 25363 34391
rect 25363 34357 25372 34391
rect 25320 34348 25372 34357
rect 25596 34416 25648 34468
rect 27528 34416 27580 34468
rect 29000 34416 29052 34468
rect 28540 34348 28592 34400
rect 30288 34348 30340 34400
rect 31024 34391 31076 34400
rect 31024 34357 31033 34391
rect 31033 34357 31067 34391
rect 31067 34357 31076 34391
rect 31024 34348 31076 34357
rect 6582 34246 6634 34298
rect 6646 34246 6698 34298
rect 6710 34246 6762 34298
rect 6774 34246 6826 34298
rect 6838 34246 6890 34298
rect 17846 34246 17898 34298
rect 17910 34246 17962 34298
rect 17974 34246 18026 34298
rect 18038 34246 18090 34298
rect 18102 34246 18154 34298
rect 29110 34246 29162 34298
rect 29174 34246 29226 34298
rect 29238 34246 29290 34298
rect 29302 34246 29354 34298
rect 29366 34246 29418 34298
rect 12900 34187 12952 34196
rect 12900 34153 12909 34187
rect 12909 34153 12943 34187
rect 12943 34153 12952 34187
rect 12900 34144 12952 34153
rect 13084 34144 13136 34196
rect 15752 34144 15804 34196
rect 15936 34144 15988 34196
rect 16212 34144 16264 34196
rect 16304 34144 16356 34196
rect 16580 34144 16632 34196
rect 2504 34076 2556 34128
rect 2780 34051 2832 34060
rect 2780 34017 2789 34051
rect 2789 34017 2823 34051
rect 2823 34017 2832 34051
rect 2780 34008 2832 34017
rect 13268 34008 13320 34060
rect 13452 34076 13504 34128
rect 14556 34008 14608 34060
rect 15476 34076 15528 34128
rect 18512 34076 18564 34128
rect 18972 34076 19024 34128
rect 20444 34144 20496 34196
rect 20720 34144 20772 34196
rect 23388 34144 23440 34196
rect 24676 34144 24728 34196
rect 24768 34144 24820 34196
rect 28632 34144 28684 34196
rect 30748 34187 30800 34196
rect 30748 34153 30757 34187
rect 30757 34153 30791 34187
rect 30791 34153 30800 34187
rect 30748 34144 30800 34153
rect 31392 34144 31444 34196
rect 32772 34144 32824 34196
rect 31208 34076 31260 34128
rect 1400 33983 1452 33992
rect 1400 33949 1409 33983
rect 1409 33949 1443 33983
rect 1443 33949 1452 33983
rect 1400 33940 1452 33949
rect 2596 33872 2648 33924
rect 14004 33940 14056 33992
rect 14188 33940 14240 33992
rect 14648 33940 14700 33992
rect 15476 33940 15528 33992
rect 15936 33940 15988 33992
rect 16212 34008 16264 34060
rect 13268 33872 13320 33924
rect 16304 33940 16356 33992
rect 16672 34051 16724 34060
rect 16672 34017 16681 34051
rect 16681 34017 16715 34051
rect 16715 34017 16724 34051
rect 16672 34008 16724 34017
rect 18696 34008 18748 34060
rect 18788 34008 18840 34060
rect 18880 33940 18932 33992
rect 19248 33983 19300 33992
rect 19248 33949 19257 33983
rect 19257 33949 19291 33983
rect 19291 33949 19300 33983
rect 19248 33940 19300 33949
rect 20260 34008 20312 34060
rect 23112 34008 23164 34060
rect 23572 34008 23624 34060
rect 21640 33940 21692 33992
rect 21916 33940 21968 33992
rect 22284 33940 22336 33992
rect 22928 33940 22980 33992
rect 23480 33940 23532 33992
rect 23756 33940 23808 33992
rect 24124 33940 24176 33992
rect 24584 33983 24636 33992
rect 24584 33949 24593 33983
rect 24593 33949 24627 33983
rect 24627 33949 24636 33983
rect 24584 33940 24636 33949
rect 14464 33804 14516 33856
rect 15752 33804 15804 33856
rect 16212 33872 16264 33924
rect 17316 33804 17368 33856
rect 17960 33804 18012 33856
rect 18052 33804 18104 33856
rect 19156 33804 19208 33856
rect 19340 33872 19392 33924
rect 20628 33872 20680 33924
rect 25136 34008 25188 34060
rect 24860 33940 24912 33992
rect 26516 33940 26568 33992
rect 30748 34008 30800 34060
rect 28540 33940 28592 33992
rect 29644 33983 29696 33992
rect 29644 33949 29653 33983
rect 29653 33949 29687 33983
rect 29687 33949 29696 33983
rect 29644 33940 29696 33949
rect 30104 33983 30156 33992
rect 30104 33949 30113 33983
rect 30113 33949 30147 33983
rect 30147 33949 30156 33983
rect 30104 33940 30156 33949
rect 31024 33983 31076 33992
rect 31024 33949 31033 33983
rect 31033 33949 31067 33983
rect 31067 33949 31076 33983
rect 31024 33940 31076 33949
rect 32496 34008 32548 34060
rect 34152 34051 34204 34060
rect 34152 34017 34161 34051
rect 34161 34017 34195 34051
rect 34195 34017 34204 34051
rect 34152 34008 34204 34017
rect 27344 33872 27396 33924
rect 20536 33804 20588 33856
rect 21456 33804 21508 33856
rect 22008 33847 22060 33856
rect 22008 33813 22017 33847
rect 22017 33813 22051 33847
rect 22051 33813 22060 33847
rect 22008 33804 22060 33813
rect 22744 33804 22796 33856
rect 23296 33804 23348 33856
rect 23848 33804 23900 33856
rect 26056 33804 26108 33856
rect 27252 33804 27304 33856
rect 28448 33872 28500 33924
rect 27804 33804 27856 33856
rect 30472 33872 30524 33924
rect 31208 33983 31260 33992
rect 31208 33949 31217 33983
rect 31217 33949 31251 33983
rect 31251 33949 31260 33983
rect 31208 33940 31260 33949
rect 31392 33983 31444 33992
rect 31392 33949 31401 33983
rect 31401 33949 31435 33983
rect 31435 33949 31444 33983
rect 31392 33940 31444 33949
rect 29644 33804 29696 33856
rect 32496 33915 32548 33924
rect 32496 33881 32505 33915
rect 32505 33881 32539 33915
rect 32539 33881 32548 33915
rect 32496 33872 32548 33881
rect 33232 33804 33284 33856
rect 12214 33702 12266 33754
rect 12278 33702 12330 33754
rect 12342 33702 12394 33754
rect 12406 33702 12458 33754
rect 12470 33702 12522 33754
rect 23478 33702 23530 33754
rect 23542 33702 23594 33754
rect 23606 33702 23658 33754
rect 23670 33702 23722 33754
rect 23734 33702 23786 33754
rect 2596 33643 2648 33652
rect 2596 33609 2605 33643
rect 2605 33609 2639 33643
rect 2639 33609 2648 33643
rect 2596 33600 2648 33609
rect 13176 33600 13228 33652
rect 13636 33600 13688 33652
rect 1400 33464 1452 33516
rect 2504 33507 2556 33516
rect 2504 33473 2513 33507
rect 2513 33473 2547 33507
rect 2547 33473 2556 33507
rect 2504 33464 2556 33473
rect 12716 33507 12768 33516
rect 12716 33473 12725 33507
rect 12725 33473 12759 33507
rect 12759 33473 12768 33507
rect 12716 33464 12768 33473
rect 13084 33464 13136 33516
rect 13360 33507 13412 33516
rect 13360 33473 13369 33507
rect 13369 33473 13403 33507
rect 13403 33473 13412 33507
rect 13360 33464 13412 33473
rect 13452 33464 13504 33516
rect 18052 33600 18104 33652
rect 14464 33532 14516 33584
rect 15660 33532 15712 33584
rect 16580 33532 16632 33584
rect 14556 33464 14608 33516
rect 18420 33532 18472 33584
rect 18696 33532 18748 33584
rect 18972 33532 19024 33584
rect 16856 33507 16908 33516
rect 12164 33396 12216 33448
rect 13912 33396 13964 33448
rect 16856 33473 16865 33507
rect 16865 33473 16899 33507
rect 16899 33473 16908 33507
rect 16856 33464 16908 33473
rect 18144 33507 18196 33516
rect 18144 33473 18153 33507
rect 18153 33473 18187 33507
rect 18187 33473 18196 33507
rect 18144 33464 18196 33473
rect 18236 33464 18288 33516
rect 19340 33600 19392 33652
rect 20444 33532 20496 33584
rect 21824 33643 21876 33652
rect 21824 33609 21833 33643
rect 21833 33609 21867 33643
rect 21867 33609 21876 33643
rect 21824 33600 21876 33609
rect 22100 33600 22152 33652
rect 24584 33600 24636 33652
rect 25320 33600 25372 33652
rect 25412 33600 25464 33652
rect 27804 33643 27856 33652
rect 27804 33609 27813 33643
rect 27813 33609 27847 33643
rect 27847 33609 27856 33643
rect 27804 33600 27856 33609
rect 28816 33600 28868 33652
rect 31208 33600 31260 33652
rect 32680 33600 32732 33652
rect 19616 33464 19668 33516
rect 19800 33507 19852 33516
rect 19800 33473 19809 33507
rect 19809 33473 19843 33507
rect 19843 33473 19852 33507
rect 19800 33464 19852 33473
rect 20076 33507 20128 33516
rect 14372 33328 14424 33380
rect 14556 33328 14608 33380
rect 17408 33396 17460 33448
rect 16396 33328 16448 33380
rect 17224 33328 17276 33380
rect 18052 33396 18104 33448
rect 19524 33396 19576 33448
rect 20076 33473 20085 33507
rect 20085 33473 20119 33507
rect 20119 33473 20128 33507
rect 20076 33464 20128 33473
rect 21640 33464 21692 33516
rect 22100 33507 22152 33516
rect 22100 33473 22109 33507
rect 22109 33473 22143 33507
rect 22143 33473 22152 33507
rect 22100 33464 22152 33473
rect 22376 33507 22428 33516
rect 22376 33473 22385 33507
rect 22385 33473 22419 33507
rect 22419 33473 22428 33507
rect 22376 33464 22428 33473
rect 22652 33464 22704 33516
rect 18512 33328 18564 33380
rect 19156 33328 19208 33380
rect 12808 33303 12860 33312
rect 12808 33269 12817 33303
rect 12817 33269 12851 33303
rect 12851 33269 12860 33303
rect 12808 33260 12860 33269
rect 13176 33260 13228 33312
rect 15936 33260 15988 33312
rect 16028 33260 16080 33312
rect 16212 33260 16264 33312
rect 17316 33260 17368 33312
rect 17408 33260 17460 33312
rect 18788 33303 18840 33312
rect 18788 33269 18797 33303
rect 18797 33269 18831 33303
rect 18831 33269 18840 33303
rect 18788 33260 18840 33269
rect 18880 33260 18932 33312
rect 19064 33260 19116 33312
rect 19800 33328 19852 33380
rect 22100 33328 22152 33380
rect 22744 33396 22796 33448
rect 23020 33507 23072 33516
rect 23020 33473 23029 33507
rect 23029 33473 23063 33507
rect 23063 33473 23072 33507
rect 23020 33464 23072 33473
rect 23848 33464 23900 33516
rect 24124 33507 24176 33516
rect 24124 33473 24133 33507
rect 24133 33473 24167 33507
rect 24167 33473 24176 33507
rect 24124 33464 24176 33473
rect 22652 33328 22704 33380
rect 23664 33396 23716 33448
rect 26056 33507 26108 33516
rect 26056 33473 26065 33507
rect 26065 33473 26099 33507
rect 26099 33473 26108 33507
rect 26056 33464 26108 33473
rect 27252 33532 27304 33584
rect 27528 33532 27580 33584
rect 28448 33532 28500 33584
rect 29368 33532 29420 33584
rect 29828 33532 29880 33584
rect 31852 33532 31904 33584
rect 22928 33328 22980 33380
rect 25320 33396 25372 33448
rect 27436 33439 27488 33448
rect 27436 33405 27445 33439
rect 27445 33405 27479 33439
rect 27479 33405 27488 33439
rect 27436 33396 27488 33405
rect 19524 33260 19576 33312
rect 26056 33328 26108 33380
rect 27988 33396 28040 33448
rect 28356 33396 28408 33448
rect 28908 33464 28960 33516
rect 29460 33464 29512 33516
rect 29000 33439 29052 33448
rect 29000 33405 29009 33439
rect 29009 33405 29043 33439
rect 29043 33405 29052 33439
rect 29000 33396 29052 33405
rect 29276 33396 29328 33448
rect 31300 33507 31352 33516
rect 30012 33439 30064 33448
rect 29460 33328 29512 33380
rect 30012 33405 30021 33439
rect 30021 33405 30055 33439
rect 30055 33405 30064 33439
rect 30012 33396 30064 33405
rect 31300 33473 31309 33507
rect 31309 33473 31343 33507
rect 31343 33473 31352 33507
rect 31300 33464 31352 33473
rect 32312 33507 32364 33516
rect 32312 33473 32321 33507
rect 32321 33473 32355 33507
rect 32355 33473 32364 33507
rect 32312 33464 32364 33473
rect 30748 33396 30800 33448
rect 33692 33396 33744 33448
rect 34152 33439 34204 33448
rect 34152 33405 34161 33439
rect 34161 33405 34195 33439
rect 34195 33405 34204 33439
rect 34152 33396 34204 33405
rect 31300 33328 31352 33380
rect 23112 33260 23164 33312
rect 28356 33260 28408 33312
rect 29828 33260 29880 33312
rect 30288 33260 30340 33312
rect 30748 33260 30800 33312
rect 32036 33260 32088 33312
rect 6582 33158 6634 33210
rect 6646 33158 6698 33210
rect 6710 33158 6762 33210
rect 6774 33158 6826 33210
rect 6838 33158 6890 33210
rect 17846 33158 17898 33210
rect 17910 33158 17962 33210
rect 17974 33158 18026 33210
rect 18038 33158 18090 33210
rect 18102 33158 18154 33210
rect 29110 33158 29162 33210
rect 29174 33158 29226 33210
rect 29238 33158 29290 33210
rect 29302 33158 29354 33210
rect 29366 33158 29418 33210
rect 12164 33056 12216 33108
rect 16396 33056 16448 33108
rect 16488 33056 16540 33108
rect 18512 33056 18564 33108
rect 18604 33056 18656 33108
rect 18788 33056 18840 33108
rect 19064 33056 19116 33108
rect 19432 33056 19484 33108
rect 22192 33056 22244 33108
rect 22376 33056 22428 33108
rect 13544 32988 13596 33040
rect 12900 32895 12952 32904
rect 12900 32861 12909 32895
rect 12909 32861 12943 32895
rect 12943 32861 12952 32895
rect 12900 32852 12952 32861
rect 13176 32852 13228 32904
rect 13636 32852 13688 32904
rect 12808 32784 12860 32836
rect 14740 32920 14792 32972
rect 16580 32988 16632 33040
rect 14464 32895 14516 32904
rect 14464 32861 14473 32895
rect 14473 32861 14507 32895
rect 14507 32861 14516 32895
rect 14464 32852 14516 32861
rect 14556 32852 14608 32904
rect 14924 32852 14976 32904
rect 16120 32920 16172 32972
rect 17132 32920 17184 32972
rect 15200 32784 15252 32836
rect 15660 32852 15712 32904
rect 16304 32852 16356 32904
rect 16856 32852 16908 32904
rect 16948 32852 17000 32904
rect 18972 32988 19024 33040
rect 19156 32988 19208 33040
rect 20720 32988 20772 33040
rect 21916 32988 21968 33040
rect 22560 33031 22612 33040
rect 22560 32997 22569 33031
rect 22569 32997 22603 33031
rect 22603 32997 22612 33031
rect 22560 32988 22612 32997
rect 22652 32988 22704 33040
rect 24492 32988 24544 33040
rect 25780 32988 25832 33040
rect 27436 32988 27488 33040
rect 27804 32988 27856 33040
rect 19248 32963 19300 32972
rect 17684 32784 17736 32836
rect 19248 32929 19257 32963
rect 19257 32929 19291 32963
rect 19291 32929 19300 32963
rect 19248 32920 19300 32929
rect 23112 32920 23164 32972
rect 23204 32920 23256 32972
rect 21364 32895 21416 32904
rect 21364 32861 21373 32895
rect 21373 32861 21407 32895
rect 21407 32861 21416 32895
rect 21364 32852 21416 32861
rect 21548 32895 21600 32904
rect 21548 32861 21557 32895
rect 21557 32861 21591 32895
rect 21591 32861 21600 32895
rect 21548 32852 21600 32861
rect 21640 32895 21692 32904
rect 21640 32861 21649 32895
rect 21649 32861 21683 32895
rect 21683 32861 21692 32895
rect 21640 32852 21692 32861
rect 22100 32852 22152 32904
rect 18972 32784 19024 32836
rect 15476 32716 15528 32768
rect 15568 32716 15620 32768
rect 16396 32716 16448 32768
rect 16488 32759 16540 32768
rect 16488 32725 16497 32759
rect 16497 32725 16531 32759
rect 16531 32725 16540 32759
rect 16488 32716 16540 32725
rect 17224 32716 17276 32768
rect 18604 32716 18656 32768
rect 18788 32716 18840 32768
rect 19156 32716 19208 32768
rect 19524 32827 19576 32836
rect 19524 32793 19558 32827
rect 19558 32793 19576 32827
rect 19524 32784 19576 32793
rect 19892 32784 19944 32836
rect 21088 32784 21140 32836
rect 21824 32784 21876 32836
rect 22652 32852 22704 32904
rect 22836 32852 22888 32904
rect 23020 32895 23072 32904
rect 23020 32861 23029 32895
rect 23029 32861 23063 32895
rect 23063 32861 23072 32895
rect 23020 32852 23072 32861
rect 23756 32920 23808 32972
rect 24768 32920 24820 32972
rect 20904 32716 20956 32768
rect 23572 32784 23624 32836
rect 24032 32784 24084 32836
rect 22468 32716 22520 32768
rect 23112 32716 23164 32768
rect 25688 32852 25740 32904
rect 27252 32963 27304 32972
rect 27252 32929 27261 32963
rect 27261 32929 27295 32963
rect 27295 32929 27304 32963
rect 27252 32920 27304 32929
rect 28724 32988 28776 33040
rect 29092 32988 29144 33040
rect 29000 32920 29052 32972
rect 28080 32852 28132 32904
rect 28356 32895 28408 32904
rect 28356 32861 28365 32895
rect 28365 32861 28399 32895
rect 28399 32861 28408 32895
rect 28356 32852 28408 32861
rect 27988 32784 28040 32836
rect 26148 32716 26200 32768
rect 27804 32716 27856 32768
rect 28356 32716 28408 32768
rect 29736 33056 29788 33108
rect 29276 32988 29328 33040
rect 29552 32988 29604 33040
rect 30104 33056 30156 33108
rect 31208 33056 31260 33108
rect 29552 32895 29604 32904
rect 29552 32861 29561 32895
rect 29561 32861 29595 32895
rect 29595 32861 29604 32895
rect 29920 32988 29972 33040
rect 29736 32920 29788 32972
rect 29552 32852 29604 32861
rect 29828 32852 29880 32904
rect 31484 32988 31536 33040
rect 31944 32988 31996 33040
rect 31668 32895 31720 32904
rect 31668 32861 31677 32895
rect 31677 32861 31711 32895
rect 31711 32861 31720 32895
rect 31668 32852 31720 32861
rect 32036 32895 32088 32904
rect 32036 32861 32045 32895
rect 32045 32861 32079 32895
rect 32079 32861 32088 32895
rect 32036 32852 32088 32861
rect 33324 32852 33376 32904
rect 28816 32716 28868 32768
rect 29460 32716 29512 32768
rect 29828 32716 29880 32768
rect 30012 32716 30064 32768
rect 30380 32716 30432 32768
rect 31852 32716 31904 32768
rect 33048 32716 33100 32768
rect 12214 32614 12266 32666
rect 12278 32614 12330 32666
rect 12342 32614 12394 32666
rect 12406 32614 12458 32666
rect 12470 32614 12522 32666
rect 23478 32614 23530 32666
rect 23542 32614 23594 32666
rect 23606 32614 23658 32666
rect 23670 32614 23722 32666
rect 23734 32614 23786 32666
rect 12808 32512 12860 32564
rect 12900 32512 12952 32564
rect 16212 32512 16264 32564
rect 16396 32512 16448 32564
rect 17316 32512 17368 32564
rect 17868 32555 17920 32564
rect 17868 32521 17877 32555
rect 17877 32521 17911 32555
rect 17911 32521 17920 32555
rect 17868 32512 17920 32521
rect 18328 32512 18380 32564
rect 12992 32487 13044 32496
rect 12992 32453 13001 32487
rect 13001 32453 13035 32487
rect 13035 32453 13044 32487
rect 12992 32444 13044 32453
rect 12624 32376 12676 32428
rect 12900 32419 12952 32428
rect 12900 32385 12909 32419
rect 12909 32385 12943 32419
rect 12943 32385 12952 32419
rect 12900 32376 12952 32385
rect 13084 32419 13136 32428
rect 13084 32385 13093 32419
rect 13093 32385 13127 32419
rect 13127 32385 13136 32419
rect 13084 32376 13136 32385
rect 14556 32444 14608 32496
rect 14648 32444 14700 32496
rect 14924 32444 14976 32496
rect 16120 32444 16172 32496
rect 16580 32444 16632 32496
rect 17040 32444 17092 32496
rect 11796 32351 11848 32360
rect 11796 32317 11805 32351
rect 11805 32317 11839 32351
rect 11839 32317 11848 32351
rect 11796 32308 11848 32317
rect 14464 32376 14516 32428
rect 15568 32376 15620 32428
rect 12348 32240 12400 32292
rect 16488 32376 16540 32428
rect 15844 32351 15896 32360
rect 15844 32317 15853 32351
rect 15853 32317 15887 32351
rect 15887 32317 15896 32351
rect 15844 32308 15896 32317
rect 16212 32308 16264 32360
rect 17500 32376 17552 32428
rect 17776 32376 17828 32428
rect 17040 32308 17092 32360
rect 17960 32376 18012 32428
rect 18236 32376 18288 32428
rect 19248 32444 19300 32496
rect 19064 32376 19116 32428
rect 19340 32376 19392 32428
rect 19800 32512 19852 32564
rect 20904 32555 20956 32564
rect 20904 32521 20913 32555
rect 20913 32521 20947 32555
rect 20947 32521 20956 32555
rect 20904 32512 20956 32521
rect 20996 32555 21048 32564
rect 20996 32521 21005 32555
rect 21005 32521 21039 32555
rect 21039 32521 21048 32555
rect 20996 32512 21048 32521
rect 22744 32512 22796 32564
rect 22836 32512 22888 32564
rect 30288 32512 30340 32564
rect 30656 32512 30708 32564
rect 20444 32444 20496 32496
rect 21548 32444 21600 32496
rect 20536 32376 20588 32428
rect 21824 32376 21876 32428
rect 23020 32444 23072 32496
rect 23204 32444 23256 32496
rect 22192 32376 22244 32428
rect 22468 32376 22520 32428
rect 22928 32376 22980 32428
rect 23480 32419 23532 32428
rect 23480 32385 23489 32419
rect 23489 32385 23523 32419
rect 23523 32385 23532 32419
rect 23480 32376 23532 32385
rect 25412 32376 25464 32428
rect 25780 32376 25832 32428
rect 23388 32308 23440 32360
rect 13636 32215 13688 32224
rect 13636 32181 13645 32215
rect 13645 32181 13679 32215
rect 13679 32181 13688 32215
rect 13636 32172 13688 32181
rect 14556 32172 14608 32224
rect 17960 32240 18012 32292
rect 15476 32172 15528 32224
rect 16028 32172 16080 32224
rect 17316 32172 17368 32224
rect 17684 32172 17736 32224
rect 20720 32240 20772 32292
rect 20996 32240 21048 32292
rect 22652 32240 22704 32292
rect 20168 32172 20220 32224
rect 21732 32172 21784 32224
rect 22100 32172 22152 32224
rect 22192 32172 22244 32224
rect 22376 32172 22428 32224
rect 23020 32240 23072 32292
rect 24492 32240 24544 32292
rect 25320 32283 25372 32292
rect 23296 32172 23348 32224
rect 23388 32172 23440 32224
rect 24860 32215 24912 32224
rect 24860 32181 24869 32215
rect 24869 32181 24903 32215
rect 24903 32181 24912 32215
rect 24860 32172 24912 32181
rect 25320 32249 25329 32283
rect 25329 32249 25363 32283
rect 25363 32249 25372 32283
rect 25320 32240 25372 32249
rect 27252 32308 27304 32360
rect 27896 32376 27948 32428
rect 28356 32376 28408 32428
rect 28448 32419 28500 32428
rect 28448 32385 28457 32419
rect 28457 32385 28491 32419
rect 28491 32385 28500 32419
rect 28448 32376 28500 32385
rect 27620 32308 27672 32360
rect 27804 32351 27856 32360
rect 27804 32317 27813 32351
rect 27813 32317 27847 32351
rect 27847 32317 27856 32351
rect 27804 32308 27856 32317
rect 28816 32419 28868 32428
rect 28816 32385 28825 32419
rect 28825 32385 28859 32419
rect 28859 32385 28868 32419
rect 28816 32376 28868 32385
rect 30012 32376 30064 32428
rect 26424 32283 26476 32292
rect 26424 32249 26433 32283
rect 26433 32249 26467 32283
rect 26467 32249 26476 32283
rect 26424 32240 26476 32249
rect 27988 32240 28040 32292
rect 25504 32172 25556 32224
rect 28632 32240 28684 32292
rect 28908 32240 28960 32292
rect 29000 32172 29052 32224
rect 34152 32487 34204 32496
rect 34152 32453 34161 32487
rect 34161 32453 34195 32487
rect 34195 32453 34204 32487
rect 34152 32444 34204 32453
rect 31484 32376 31536 32428
rect 32312 32419 32364 32428
rect 32312 32385 32321 32419
rect 32321 32385 32355 32419
rect 32355 32385 32364 32419
rect 32312 32376 32364 32385
rect 30748 32351 30800 32360
rect 30748 32317 30757 32351
rect 30757 32317 30791 32351
rect 30791 32317 30800 32351
rect 30748 32308 30800 32317
rect 31668 32308 31720 32360
rect 33784 32240 33836 32292
rect 30104 32172 30156 32224
rect 30748 32172 30800 32224
rect 6582 32070 6634 32122
rect 6646 32070 6698 32122
rect 6710 32070 6762 32122
rect 6774 32070 6826 32122
rect 6838 32070 6890 32122
rect 17846 32070 17898 32122
rect 17910 32070 17962 32122
rect 17974 32070 18026 32122
rect 18038 32070 18090 32122
rect 18102 32070 18154 32122
rect 29110 32070 29162 32122
rect 29174 32070 29226 32122
rect 29238 32070 29290 32122
rect 29302 32070 29354 32122
rect 29366 32070 29418 32122
rect 14740 31968 14792 32020
rect 14924 31968 14976 32020
rect 15660 31968 15712 32020
rect 16212 31968 16264 32020
rect 16396 31968 16448 32020
rect 16580 31968 16632 32020
rect 16764 31968 16816 32020
rect 18236 31968 18288 32020
rect 18512 32011 18564 32020
rect 18512 31977 18521 32011
rect 18521 31977 18555 32011
rect 18555 31977 18564 32011
rect 18512 31968 18564 31977
rect 18604 31968 18656 32020
rect 18972 31968 19024 32020
rect 19064 31968 19116 32020
rect 20720 31968 20772 32020
rect 21640 31968 21692 32020
rect 22192 31968 22244 32020
rect 22284 31968 22336 32020
rect 23204 32011 23256 32020
rect 14556 31900 14608 31952
rect 16488 31900 16540 31952
rect 1492 31764 1544 31816
rect 12348 31807 12400 31816
rect 12348 31773 12357 31807
rect 12357 31773 12391 31807
rect 12391 31773 12400 31807
rect 12348 31764 12400 31773
rect 12808 31807 12860 31816
rect 12808 31773 12817 31807
rect 12817 31773 12851 31807
rect 12851 31773 12860 31807
rect 12808 31764 12860 31773
rect 12992 31807 13044 31816
rect 12992 31773 13001 31807
rect 13001 31773 13035 31807
rect 13035 31773 13044 31807
rect 12992 31764 13044 31773
rect 14372 31764 14424 31816
rect 14464 31696 14516 31748
rect 14924 31764 14976 31816
rect 15108 31696 15160 31748
rect 16580 31832 16632 31884
rect 12716 31628 12768 31680
rect 13728 31628 13780 31680
rect 15292 31628 15344 31680
rect 16028 31764 16080 31816
rect 18144 31832 18196 31884
rect 17776 31764 17828 31816
rect 15936 31696 15988 31748
rect 16580 31696 16632 31748
rect 16856 31696 16908 31748
rect 18604 31764 18656 31816
rect 18880 31832 18932 31884
rect 19340 31900 19392 31952
rect 20444 31900 20496 31952
rect 23204 31977 23213 32011
rect 23213 31977 23247 32011
rect 23247 31977 23256 32011
rect 23204 31968 23256 31977
rect 23296 31968 23348 32020
rect 24860 31968 24912 32020
rect 19156 31832 19208 31884
rect 19708 31832 19760 31884
rect 20536 31875 20588 31884
rect 20536 31841 20545 31875
rect 20545 31841 20579 31875
rect 20579 31841 20588 31875
rect 20536 31832 20588 31841
rect 20904 31832 20956 31884
rect 21456 31832 21508 31884
rect 21824 31832 21876 31884
rect 21916 31832 21968 31884
rect 23296 31832 23348 31884
rect 25228 31900 25280 31952
rect 26332 31900 26384 31952
rect 16212 31628 16264 31680
rect 16396 31628 16448 31680
rect 19064 31696 19116 31748
rect 19616 31739 19668 31748
rect 19616 31705 19625 31739
rect 19625 31705 19659 31739
rect 19659 31705 19668 31739
rect 19616 31696 19668 31705
rect 19708 31696 19760 31748
rect 21640 31696 21692 31748
rect 22008 31764 22060 31816
rect 22836 31764 22888 31816
rect 23388 31764 23440 31816
rect 22652 31696 22704 31748
rect 18512 31628 18564 31680
rect 18604 31628 18656 31680
rect 18880 31628 18932 31680
rect 19524 31628 19576 31680
rect 20076 31628 20128 31680
rect 20628 31628 20680 31680
rect 20720 31628 20772 31680
rect 22744 31628 22796 31680
rect 26148 31832 26200 31884
rect 24584 31764 24636 31816
rect 25504 31807 25556 31816
rect 24676 31696 24728 31748
rect 25504 31773 25513 31807
rect 25513 31773 25547 31807
rect 25547 31773 25556 31807
rect 25504 31764 25556 31773
rect 25596 31764 25648 31816
rect 26056 31696 26108 31748
rect 26884 31807 26936 31816
rect 26884 31773 26893 31807
rect 26893 31773 26927 31807
rect 26927 31773 26936 31807
rect 27068 31807 27120 31816
rect 26884 31764 26936 31773
rect 27068 31773 27077 31807
rect 27077 31773 27111 31807
rect 27111 31773 27120 31807
rect 27068 31764 27120 31773
rect 27804 31875 27856 31884
rect 27804 31841 27813 31875
rect 27813 31841 27847 31875
rect 27847 31841 27856 31875
rect 27804 31832 27856 31841
rect 27896 31832 27948 31884
rect 27896 31696 27948 31748
rect 28080 31764 28132 31816
rect 30564 31968 30616 32020
rect 28632 31900 28684 31952
rect 29276 31900 29328 31952
rect 30104 31832 30156 31884
rect 30380 31832 30432 31884
rect 30932 31968 30984 32020
rect 28724 31807 28776 31816
rect 28724 31773 28733 31807
rect 28733 31773 28767 31807
rect 28767 31773 28776 31807
rect 28724 31764 28776 31773
rect 29000 31807 29052 31816
rect 29000 31773 29009 31807
rect 29009 31773 29043 31807
rect 29043 31773 29052 31807
rect 29000 31764 29052 31773
rect 30656 31764 30708 31816
rect 29828 31696 29880 31748
rect 30196 31696 30248 31748
rect 24216 31628 24268 31680
rect 25688 31628 25740 31680
rect 26608 31628 26660 31680
rect 28080 31671 28132 31680
rect 28080 31637 28089 31671
rect 28089 31637 28123 31671
rect 28123 31637 28132 31671
rect 28080 31628 28132 31637
rect 28632 31628 28684 31680
rect 29000 31628 29052 31680
rect 31668 31968 31720 32020
rect 31484 31900 31536 31952
rect 32036 31900 32088 31952
rect 33416 31900 33468 31952
rect 31944 31832 31996 31884
rect 32312 31875 32364 31884
rect 32312 31841 32321 31875
rect 32321 31841 32355 31875
rect 32355 31841 32364 31875
rect 32312 31832 32364 31841
rect 32588 31832 32640 31884
rect 34152 31875 34204 31884
rect 34152 31841 34161 31875
rect 34161 31841 34195 31875
rect 34195 31841 34204 31875
rect 34152 31832 34204 31841
rect 31484 31807 31536 31816
rect 31484 31773 31493 31807
rect 31493 31773 31527 31807
rect 31527 31773 31536 31807
rect 31484 31764 31536 31773
rect 12214 31526 12266 31578
rect 12278 31526 12330 31578
rect 12342 31526 12394 31578
rect 12406 31526 12458 31578
rect 12470 31526 12522 31578
rect 23478 31526 23530 31578
rect 23542 31526 23594 31578
rect 23606 31526 23658 31578
rect 23670 31526 23722 31578
rect 23734 31526 23786 31578
rect 12992 31424 13044 31476
rect 1492 31331 1544 31340
rect 1492 31297 1501 31331
rect 1501 31297 1535 31331
rect 1535 31297 1544 31331
rect 1492 31288 1544 31297
rect 12256 31331 12308 31340
rect 12256 31297 12265 31331
rect 12265 31297 12299 31331
rect 12299 31297 12308 31331
rect 12256 31288 12308 31297
rect 12900 31288 12952 31340
rect 14648 31356 14700 31408
rect 15108 31356 15160 31408
rect 16764 31399 16816 31408
rect 1860 31220 1912 31272
rect 1952 31263 2004 31272
rect 1952 31229 1961 31263
rect 1961 31229 1995 31263
rect 1995 31229 2004 31263
rect 13728 31288 13780 31340
rect 13820 31288 13872 31340
rect 14556 31288 14608 31340
rect 1952 31220 2004 31229
rect 14004 31220 14056 31272
rect 16488 31288 16540 31340
rect 16764 31365 16773 31399
rect 16773 31365 16807 31399
rect 16807 31365 16816 31399
rect 16764 31356 16816 31365
rect 18236 31399 18288 31408
rect 17040 31288 17092 31340
rect 17224 31288 17276 31340
rect 18236 31365 18245 31399
rect 18245 31365 18279 31399
rect 18279 31365 18288 31399
rect 18236 31356 18288 31365
rect 18512 31424 18564 31476
rect 18052 31288 18104 31340
rect 18328 31288 18380 31340
rect 15844 31220 15896 31272
rect 13544 31127 13596 31136
rect 13544 31093 13553 31127
rect 13553 31093 13587 31127
rect 13587 31093 13596 31127
rect 13544 31084 13596 31093
rect 14004 31084 14056 31136
rect 14556 31084 14608 31136
rect 15936 31152 15988 31204
rect 16488 31152 16540 31204
rect 16856 31152 16908 31204
rect 17132 31220 17184 31272
rect 17500 31220 17552 31272
rect 17684 31220 17736 31272
rect 18788 31288 18840 31340
rect 18880 31220 18932 31272
rect 16672 31084 16724 31136
rect 16948 31084 17000 31136
rect 21456 31424 21508 31476
rect 24124 31424 24176 31476
rect 24216 31424 24268 31476
rect 27068 31424 27120 31476
rect 27436 31424 27488 31476
rect 27988 31424 28040 31476
rect 28264 31424 28316 31476
rect 28540 31424 28592 31476
rect 19340 31288 19392 31340
rect 20168 31288 20220 31340
rect 21548 31288 21600 31340
rect 22100 31356 22152 31408
rect 22744 31356 22796 31408
rect 24676 31356 24728 31408
rect 29644 31424 29696 31476
rect 30196 31467 30248 31476
rect 30196 31433 30205 31467
rect 30205 31433 30239 31467
rect 30239 31433 30248 31467
rect 30196 31424 30248 31433
rect 32128 31424 32180 31476
rect 22928 31288 22980 31340
rect 23112 31288 23164 31340
rect 23480 31288 23532 31340
rect 23756 31331 23808 31340
rect 21088 31220 21140 31272
rect 20628 31152 20680 31204
rect 20720 31152 20772 31204
rect 21456 31220 21508 31272
rect 21364 31152 21416 31204
rect 21640 31152 21692 31204
rect 23572 31220 23624 31272
rect 23756 31297 23785 31331
rect 23785 31297 23808 31331
rect 23756 31288 23808 31297
rect 24400 31288 24452 31340
rect 24860 31331 24912 31340
rect 24860 31297 24869 31331
rect 24869 31297 24903 31331
rect 24903 31297 24912 31331
rect 24860 31288 24912 31297
rect 25412 31288 25464 31340
rect 30380 31331 30432 31340
rect 30380 31297 30389 31331
rect 30389 31297 30423 31331
rect 30423 31297 30432 31331
rect 30380 31288 30432 31297
rect 30564 31331 30616 31340
rect 30564 31297 30573 31331
rect 30573 31297 30607 31331
rect 30607 31297 30616 31331
rect 30564 31288 30616 31297
rect 30840 31288 30892 31340
rect 23848 31220 23900 31272
rect 25044 31220 25096 31272
rect 27528 31263 27580 31272
rect 27528 31229 27537 31263
rect 27537 31229 27571 31263
rect 27571 31229 27580 31263
rect 27528 31220 27580 31229
rect 27988 31263 28040 31272
rect 22376 31195 22428 31204
rect 22376 31161 22385 31195
rect 22385 31161 22419 31195
rect 22419 31161 22428 31195
rect 22376 31152 22428 31161
rect 27988 31229 27997 31263
rect 27997 31229 28031 31263
rect 28031 31229 28040 31263
rect 27988 31220 28040 31229
rect 18788 31084 18840 31136
rect 18880 31084 18932 31136
rect 19432 31084 19484 31136
rect 19616 31084 19668 31136
rect 21088 31127 21140 31136
rect 21088 31093 21097 31127
rect 21097 31093 21131 31127
rect 21131 31093 21140 31127
rect 21088 31084 21140 31093
rect 21272 31084 21324 31136
rect 22008 31084 22060 31136
rect 23848 31084 23900 31136
rect 24124 31084 24176 31136
rect 24216 31084 24268 31136
rect 26240 31084 26292 31136
rect 27252 31084 27304 31136
rect 29736 31220 29788 31272
rect 30288 31220 30340 31272
rect 34152 31331 34204 31340
rect 34152 31297 34161 31331
rect 34161 31297 34195 31331
rect 34195 31297 34204 31331
rect 34152 31288 34204 31297
rect 30564 31152 30616 31204
rect 32312 31263 32364 31272
rect 32312 31229 32321 31263
rect 32321 31229 32355 31263
rect 32355 31229 32364 31263
rect 32312 31220 32364 31229
rect 34060 31220 34112 31272
rect 29000 31084 29052 31136
rect 31576 31084 31628 31136
rect 6582 30982 6634 31034
rect 6646 30982 6698 31034
rect 6710 30982 6762 31034
rect 6774 30982 6826 31034
rect 6838 30982 6890 31034
rect 17846 30982 17898 31034
rect 17910 30982 17962 31034
rect 17974 30982 18026 31034
rect 18038 30982 18090 31034
rect 18102 30982 18154 31034
rect 29110 30982 29162 31034
rect 29174 30982 29226 31034
rect 29238 30982 29290 31034
rect 29302 30982 29354 31034
rect 29366 30982 29418 31034
rect 1860 30923 1912 30932
rect 1860 30889 1869 30923
rect 1869 30889 1903 30923
rect 1903 30889 1912 30923
rect 1860 30880 1912 30889
rect 12072 30923 12124 30932
rect 12072 30889 12081 30923
rect 12081 30889 12115 30923
rect 12115 30889 12124 30923
rect 12072 30880 12124 30889
rect 13084 30880 13136 30932
rect 13544 30880 13596 30932
rect 15200 30880 15252 30932
rect 15292 30880 15344 30932
rect 12256 30812 12308 30864
rect 12808 30787 12860 30796
rect 12808 30753 12817 30787
rect 12817 30753 12851 30787
rect 12851 30753 12860 30787
rect 12808 30744 12860 30753
rect 15660 30855 15712 30864
rect 15660 30821 15669 30855
rect 15669 30821 15703 30855
rect 15703 30821 15712 30855
rect 15936 30880 15988 30932
rect 15660 30812 15712 30821
rect 17132 30812 17184 30864
rect 18696 30923 18748 30932
rect 18696 30889 18705 30923
rect 18705 30889 18739 30923
rect 18739 30889 18748 30923
rect 18696 30880 18748 30889
rect 24676 30880 24728 30932
rect 25228 30880 25280 30932
rect 27896 30923 27948 30932
rect 20260 30812 20312 30864
rect 21456 30812 21508 30864
rect 1768 30719 1820 30728
rect 1768 30685 1777 30719
rect 1777 30685 1811 30719
rect 1811 30685 1820 30719
rect 1768 30676 1820 30685
rect 11980 30676 12032 30728
rect 12624 30676 12676 30728
rect 12992 30676 13044 30728
rect 13544 30719 13596 30728
rect 13176 30608 13228 30660
rect 13544 30685 13553 30719
rect 13553 30685 13587 30719
rect 13587 30685 13596 30719
rect 13544 30676 13596 30685
rect 15108 30676 15160 30728
rect 15844 30744 15896 30796
rect 16028 30744 16080 30796
rect 16396 30744 16448 30796
rect 17316 30787 17368 30796
rect 15936 30676 15988 30728
rect 16304 30719 16356 30728
rect 16304 30685 16313 30719
rect 16313 30685 16347 30719
rect 16347 30685 16356 30719
rect 16304 30676 16356 30685
rect 16672 30676 16724 30728
rect 17316 30753 17325 30787
rect 17325 30753 17359 30787
rect 17359 30753 17368 30787
rect 17316 30744 17368 30753
rect 14648 30608 14700 30660
rect 14832 30608 14884 30660
rect 15292 30608 15344 30660
rect 15476 30651 15528 30660
rect 15476 30617 15485 30651
rect 15485 30617 15519 30651
rect 15519 30617 15528 30651
rect 15476 30608 15528 30617
rect 15844 30608 15896 30660
rect 14464 30540 14516 30592
rect 18144 30676 18196 30728
rect 19616 30744 19668 30796
rect 18420 30676 18472 30728
rect 18696 30676 18748 30728
rect 18972 30676 19024 30728
rect 19340 30676 19392 30728
rect 19800 30676 19852 30728
rect 20812 30676 20864 30728
rect 20996 30744 21048 30796
rect 21180 30676 21232 30728
rect 21732 30744 21784 30796
rect 23388 30812 23440 30864
rect 25136 30855 25188 30864
rect 25136 30821 25145 30855
rect 25145 30821 25179 30855
rect 25179 30821 25188 30855
rect 25136 30812 25188 30821
rect 25412 30812 25464 30864
rect 25780 30812 25832 30864
rect 25964 30812 26016 30864
rect 27896 30889 27905 30923
rect 27905 30889 27939 30923
rect 27939 30889 27948 30923
rect 27896 30880 27948 30889
rect 28264 30880 28316 30932
rect 30840 30880 30892 30932
rect 22100 30787 22152 30796
rect 22100 30753 22109 30787
rect 22109 30753 22143 30787
rect 22143 30753 22152 30787
rect 22100 30744 22152 30753
rect 22836 30744 22888 30796
rect 23572 30744 23624 30796
rect 25596 30744 25648 30796
rect 19708 30608 19760 30660
rect 20168 30608 20220 30660
rect 22008 30608 22060 30660
rect 22928 30676 22980 30728
rect 23204 30719 23256 30728
rect 23204 30685 23213 30719
rect 23213 30685 23247 30719
rect 23247 30685 23256 30719
rect 23204 30676 23256 30685
rect 22376 30608 22428 30660
rect 24308 30676 24360 30728
rect 24952 30676 25004 30728
rect 25780 30719 25832 30728
rect 25780 30685 25789 30719
rect 25789 30685 25823 30719
rect 25823 30685 25832 30719
rect 25780 30676 25832 30685
rect 26332 30744 26384 30796
rect 28540 30787 28592 30796
rect 28540 30753 28549 30787
rect 28549 30753 28583 30787
rect 28583 30753 28592 30787
rect 28540 30744 28592 30753
rect 26516 30719 26568 30728
rect 22192 30540 22244 30592
rect 22468 30540 22520 30592
rect 25320 30608 25372 30660
rect 25412 30608 25464 30660
rect 26516 30685 26525 30719
rect 26525 30685 26559 30719
rect 26559 30685 26568 30719
rect 26516 30676 26568 30685
rect 26608 30676 26660 30728
rect 27160 30676 27212 30728
rect 29736 30744 29788 30796
rect 30012 30744 30064 30796
rect 31944 30812 31996 30864
rect 32036 30744 32088 30796
rect 32220 30787 32272 30796
rect 32220 30753 32229 30787
rect 32229 30753 32263 30787
rect 32263 30753 32272 30787
rect 32220 30744 32272 30753
rect 28724 30719 28776 30728
rect 28724 30685 28753 30719
rect 28753 30685 28776 30719
rect 28724 30676 28776 30685
rect 30104 30719 30156 30728
rect 30104 30685 30113 30719
rect 30113 30685 30147 30719
rect 30147 30685 30156 30719
rect 30104 30676 30156 30685
rect 31484 30676 31536 30728
rect 31576 30676 31628 30728
rect 31944 30676 31996 30728
rect 32312 30719 32364 30728
rect 32312 30685 32321 30719
rect 32321 30685 32355 30719
rect 32355 30685 32364 30719
rect 32312 30676 32364 30685
rect 33508 30744 33560 30796
rect 34244 30744 34296 30796
rect 33876 30719 33928 30728
rect 27804 30608 27856 30660
rect 27896 30608 27948 30660
rect 28908 30608 28960 30660
rect 29644 30608 29696 30660
rect 22836 30540 22888 30592
rect 24400 30540 24452 30592
rect 27344 30540 27396 30592
rect 27988 30540 28040 30592
rect 30656 30540 30708 30592
rect 31024 30540 31076 30592
rect 31944 30583 31996 30592
rect 31944 30549 31953 30583
rect 31953 30549 31987 30583
rect 31987 30549 31996 30583
rect 31944 30540 31996 30549
rect 33048 30608 33100 30660
rect 33876 30685 33885 30719
rect 33885 30685 33919 30719
rect 33919 30685 33928 30719
rect 33876 30676 33928 30685
rect 33968 30676 34020 30728
rect 12214 30438 12266 30490
rect 12278 30438 12330 30490
rect 12342 30438 12394 30490
rect 12406 30438 12458 30490
rect 12470 30438 12522 30490
rect 23478 30438 23530 30490
rect 23542 30438 23594 30490
rect 23606 30438 23658 30490
rect 23670 30438 23722 30490
rect 23734 30438 23786 30490
rect 13820 30336 13872 30388
rect 16948 30336 17000 30388
rect 17684 30336 17736 30388
rect 11796 30200 11848 30252
rect 12440 30200 12492 30252
rect 14832 30268 14884 30320
rect 15476 30268 15528 30320
rect 16580 30268 16632 30320
rect 20996 30336 21048 30388
rect 12624 30200 12676 30252
rect 12808 30200 12860 30252
rect 13268 30200 13320 30252
rect 13728 30200 13780 30252
rect 14280 30200 14332 30252
rect 14556 30200 14608 30252
rect 15108 30200 15160 30252
rect 15844 30200 15896 30252
rect 16028 30200 16080 30252
rect 16304 30200 16356 30252
rect 16856 30200 16908 30252
rect 17132 30243 17184 30252
rect 17132 30209 17141 30243
rect 17141 30209 17175 30243
rect 17175 30209 17184 30243
rect 17132 30200 17184 30209
rect 17316 30200 17368 30252
rect 17592 30200 17644 30252
rect 18420 30268 18472 30320
rect 21732 30336 21784 30388
rect 17960 30243 18012 30252
rect 17960 30209 17983 30243
rect 17983 30209 18012 30243
rect 17960 30200 18012 30209
rect 18328 30200 18380 30252
rect 19248 30200 19300 30252
rect 19524 30243 19576 30252
rect 19524 30209 19533 30243
rect 19533 30209 19567 30243
rect 19567 30209 19576 30243
rect 19524 30200 19576 30209
rect 20260 30200 20312 30252
rect 20536 30200 20588 30252
rect 17040 30064 17092 30116
rect 17500 30064 17552 30116
rect 13176 29996 13228 30048
rect 14188 29996 14240 30048
rect 14924 29996 14976 30048
rect 15476 29996 15528 30048
rect 16212 29996 16264 30048
rect 16304 29996 16356 30048
rect 20996 30132 21048 30184
rect 22173 30246 22225 30252
rect 22376 30336 22428 30388
rect 22560 30268 22612 30320
rect 22744 30268 22796 30320
rect 22173 30212 22198 30246
rect 22198 30212 22225 30246
rect 22173 30200 22225 30212
rect 22652 30200 22704 30252
rect 22836 30132 22888 30184
rect 23480 30200 23532 30252
rect 23940 30243 23992 30252
rect 23940 30209 23949 30243
rect 23949 30209 23983 30243
rect 23983 30209 23992 30243
rect 23940 30200 23992 30209
rect 24124 30200 24176 30252
rect 25136 30268 25188 30320
rect 25780 30268 25832 30320
rect 30012 30336 30064 30388
rect 25504 30200 25556 30252
rect 25596 30200 25648 30252
rect 29000 30268 29052 30320
rect 29644 30268 29696 30320
rect 24952 30175 25004 30184
rect 24952 30141 24961 30175
rect 24961 30141 24995 30175
rect 24995 30141 25004 30175
rect 26056 30175 26108 30184
rect 24952 30132 25004 30141
rect 26056 30141 26065 30175
rect 26065 30141 26099 30175
rect 26099 30141 26108 30175
rect 26056 30132 26108 30141
rect 18696 29996 18748 30048
rect 20536 29996 20588 30048
rect 23296 30064 23348 30116
rect 25412 30064 25464 30116
rect 25872 30064 25924 30116
rect 28264 30243 28316 30252
rect 28264 30209 28298 30243
rect 28298 30209 28316 30243
rect 28264 30200 28316 30209
rect 28540 30200 28592 30252
rect 30564 30336 30616 30388
rect 30656 30336 30708 30388
rect 26516 30132 26568 30184
rect 27160 30132 27212 30184
rect 23940 29996 23992 30048
rect 27896 30064 27948 30116
rect 29000 30064 29052 30116
rect 30748 30268 30800 30320
rect 30840 30268 30892 30320
rect 31668 30268 31720 30320
rect 33876 30268 33928 30320
rect 30656 30200 30708 30252
rect 33140 30200 33192 30252
rect 33784 30243 33836 30252
rect 33784 30209 33793 30243
rect 33793 30209 33827 30243
rect 33827 30209 33836 30243
rect 33784 30200 33836 30209
rect 31852 30132 31904 30184
rect 31944 30132 31996 30184
rect 29644 30064 29696 30116
rect 30288 30064 30340 30116
rect 31208 30107 31260 30116
rect 31208 30073 31217 30107
rect 31217 30073 31251 30107
rect 31251 30073 31260 30107
rect 31208 30064 31260 30073
rect 30380 29996 30432 30048
rect 30840 30039 30892 30048
rect 30840 30005 30849 30039
rect 30849 30005 30883 30039
rect 30883 30005 30892 30039
rect 30840 29996 30892 30005
rect 31300 29996 31352 30048
rect 31484 29996 31536 30048
rect 33140 29996 33192 30048
rect 33416 29996 33468 30048
rect 6582 29894 6634 29946
rect 6646 29894 6698 29946
rect 6710 29894 6762 29946
rect 6774 29894 6826 29946
rect 6838 29894 6890 29946
rect 17846 29894 17898 29946
rect 17910 29894 17962 29946
rect 17974 29894 18026 29946
rect 18038 29894 18090 29946
rect 18102 29894 18154 29946
rect 29110 29894 29162 29946
rect 29174 29894 29226 29946
rect 29238 29894 29290 29946
rect 29302 29894 29354 29946
rect 29366 29894 29418 29946
rect 15292 29792 15344 29844
rect 20444 29792 20496 29844
rect 22836 29835 22888 29844
rect 11796 29724 11848 29776
rect 15936 29724 15988 29776
rect 16028 29724 16080 29776
rect 17040 29724 17092 29776
rect 19432 29724 19484 29776
rect 17132 29656 17184 29708
rect 19524 29699 19576 29708
rect 11888 29588 11940 29640
rect 12716 29631 12768 29640
rect 12716 29597 12725 29631
rect 12725 29597 12759 29631
rect 12759 29597 12768 29631
rect 12716 29588 12768 29597
rect 12900 29631 12952 29640
rect 12900 29597 12909 29631
rect 12909 29597 12943 29631
rect 12943 29597 12952 29631
rect 12900 29588 12952 29597
rect 13360 29631 13412 29640
rect 13360 29597 13369 29631
rect 13369 29597 13403 29631
rect 13403 29597 13412 29631
rect 13360 29588 13412 29597
rect 14004 29588 14056 29640
rect 14188 29588 14240 29640
rect 14372 29588 14424 29640
rect 14832 29588 14884 29640
rect 15384 29631 15436 29640
rect 15384 29597 15393 29631
rect 15393 29597 15427 29631
rect 15427 29597 15436 29631
rect 15384 29588 15436 29597
rect 15476 29631 15528 29640
rect 15476 29597 15485 29631
rect 15485 29597 15519 29631
rect 15519 29597 15528 29631
rect 15476 29588 15528 29597
rect 15752 29588 15804 29640
rect 15936 29588 15988 29640
rect 17316 29588 17368 29640
rect 17776 29588 17828 29640
rect 18052 29631 18104 29640
rect 18052 29597 18061 29631
rect 18061 29597 18095 29631
rect 18095 29597 18104 29631
rect 18052 29588 18104 29597
rect 18144 29588 18196 29640
rect 16396 29520 16448 29572
rect 16672 29520 16724 29572
rect 17040 29520 17092 29572
rect 13268 29452 13320 29504
rect 14648 29452 14700 29504
rect 15752 29452 15804 29504
rect 16028 29452 16080 29504
rect 17960 29520 18012 29572
rect 18604 29588 18656 29640
rect 18972 29588 19024 29640
rect 19524 29665 19533 29699
rect 19533 29665 19567 29699
rect 19567 29665 19576 29699
rect 19524 29656 19576 29665
rect 20628 29724 20680 29776
rect 21824 29724 21876 29776
rect 22284 29724 22336 29776
rect 22468 29767 22520 29776
rect 22468 29733 22477 29767
rect 22477 29733 22511 29767
rect 22511 29733 22520 29767
rect 22468 29724 22520 29733
rect 22836 29801 22845 29835
rect 22845 29801 22879 29835
rect 22879 29801 22888 29835
rect 22836 29792 22888 29801
rect 23388 29792 23440 29844
rect 23848 29792 23900 29844
rect 24584 29792 24636 29844
rect 21916 29656 21968 29708
rect 20628 29588 20680 29640
rect 17224 29452 17276 29504
rect 17500 29452 17552 29504
rect 18236 29495 18288 29504
rect 18236 29461 18245 29495
rect 18245 29461 18279 29495
rect 18279 29461 18288 29495
rect 18236 29452 18288 29461
rect 19616 29452 19668 29504
rect 20996 29452 21048 29504
rect 21088 29452 21140 29504
rect 21456 29452 21508 29504
rect 21824 29631 21876 29640
rect 21824 29597 21833 29631
rect 21833 29597 21867 29631
rect 21867 29597 21876 29631
rect 25044 29656 25096 29708
rect 27620 29792 27672 29844
rect 27896 29792 27948 29844
rect 28264 29792 28316 29844
rect 28724 29792 28776 29844
rect 30288 29792 30340 29844
rect 32036 29792 32088 29844
rect 32496 29792 32548 29844
rect 33048 29792 33100 29844
rect 27436 29724 27488 29776
rect 29644 29724 29696 29776
rect 30196 29724 30248 29776
rect 21824 29588 21876 29597
rect 22376 29588 22428 29640
rect 22744 29588 22796 29640
rect 25412 29631 25464 29640
rect 22192 29520 22244 29572
rect 22560 29520 22612 29572
rect 23480 29520 23532 29572
rect 24124 29520 24176 29572
rect 24676 29520 24728 29572
rect 24952 29520 25004 29572
rect 25412 29597 25421 29631
rect 25421 29597 25455 29631
rect 25455 29597 25464 29631
rect 25412 29588 25464 29597
rect 25504 29631 25556 29640
rect 25504 29597 25513 29631
rect 25513 29597 25547 29631
rect 25547 29597 25556 29631
rect 25504 29588 25556 29597
rect 25872 29520 25924 29572
rect 26332 29631 26384 29640
rect 26332 29597 26341 29631
rect 26341 29597 26375 29631
rect 26375 29597 26384 29631
rect 26332 29588 26384 29597
rect 27068 29588 27120 29640
rect 27344 29631 27396 29640
rect 27344 29597 27353 29631
rect 27353 29597 27387 29631
rect 27387 29597 27396 29631
rect 27344 29588 27396 29597
rect 28448 29588 28500 29640
rect 28724 29631 28776 29640
rect 28724 29597 28733 29631
rect 28733 29597 28767 29631
rect 28767 29597 28776 29631
rect 28724 29588 28776 29597
rect 29368 29588 29420 29640
rect 30472 29656 30524 29708
rect 30840 29656 30892 29708
rect 30656 29588 30708 29640
rect 26884 29520 26936 29572
rect 29276 29520 29328 29572
rect 22744 29452 22796 29504
rect 23296 29452 23348 29504
rect 25964 29452 26016 29504
rect 27804 29452 27856 29504
rect 29368 29452 29420 29504
rect 30012 29452 30064 29504
rect 31300 29452 31352 29504
rect 32128 29631 32180 29640
rect 32128 29597 32137 29631
rect 32137 29597 32171 29631
rect 32171 29597 32180 29631
rect 32128 29588 32180 29597
rect 34152 29588 34204 29640
rect 32864 29520 32916 29572
rect 33692 29452 33744 29504
rect 12214 29350 12266 29402
rect 12278 29350 12330 29402
rect 12342 29350 12394 29402
rect 12406 29350 12458 29402
rect 12470 29350 12522 29402
rect 23478 29350 23530 29402
rect 23542 29350 23594 29402
rect 23606 29350 23658 29402
rect 23670 29350 23722 29402
rect 23734 29350 23786 29402
rect 12992 29291 13044 29300
rect 12992 29257 13001 29291
rect 13001 29257 13035 29291
rect 13035 29257 13044 29291
rect 12992 29248 13044 29257
rect 14188 29248 14240 29300
rect 13820 29180 13872 29232
rect 14648 29223 14700 29232
rect 14648 29189 14657 29223
rect 14657 29189 14691 29223
rect 14691 29189 14700 29223
rect 14648 29180 14700 29189
rect 15660 29248 15712 29300
rect 22560 29248 22612 29300
rect 16580 29180 16632 29232
rect 13268 29155 13320 29164
rect 13268 29121 13277 29155
rect 13277 29121 13311 29155
rect 13311 29121 13320 29155
rect 13268 29112 13320 29121
rect 13636 29112 13688 29164
rect 14556 29155 14608 29164
rect 13728 29044 13780 29096
rect 13820 29044 13872 29096
rect 14004 29087 14056 29096
rect 14004 29053 14013 29087
rect 14013 29053 14047 29087
rect 14047 29053 14056 29087
rect 14004 29044 14056 29053
rect 14556 29121 14565 29155
rect 14565 29121 14599 29155
rect 14599 29121 14608 29155
rect 14556 29112 14608 29121
rect 15108 29112 15160 29164
rect 15476 29112 15528 29164
rect 15660 29112 15712 29164
rect 14832 29044 14884 29096
rect 15568 29044 15620 29096
rect 16120 29155 16172 29164
rect 16120 29121 16129 29155
rect 16129 29121 16163 29155
rect 16163 29121 16172 29155
rect 16120 29112 16172 29121
rect 15292 29019 15344 29028
rect 15292 28985 15301 29019
rect 15301 28985 15335 29019
rect 15335 28985 15344 29019
rect 15292 28976 15344 28985
rect 12164 28951 12216 28960
rect 12164 28917 12173 28951
rect 12173 28917 12207 28951
rect 12207 28917 12216 28951
rect 12164 28908 12216 28917
rect 13452 28951 13504 28960
rect 13452 28917 13461 28951
rect 13461 28917 13495 28951
rect 13495 28917 13504 28951
rect 13452 28908 13504 28917
rect 13636 28908 13688 28960
rect 14004 28908 14056 28960
rect 15016 28908 15068 28960
rect 16120 28976 16172 29028
rect 16212 28976 16264 29028
rect 17408 29180 17460 29232
rect 18328 29180 18380 29232
rect 18512 29180 18564 29232
rect 20444 29180 20496 29232
rect 21824 29223 21876 29232
rect 16948 29087 17000 29096
rect 16948 29053 16957 29087
rect 16957 29053 16991 29087
rect 16991 29053 17000 29087
rect 16948 29044 17000 29053
rect 18052 29112 18104 29164
rect 18604 29112 18656 29164
rect 18972 29155 19024 29164
rect 18972 29121 18981 29155
rect 18981 29121 19015 29155
rect 19015 29121 19024 29155
rect 18972 29112 19024 29121
rect 20996 29155 21048 29164
rect 20996 29121 21005 29155
rect 21005 29121 21039 29155
rect 21039 29121 21048 29155
rect 20996 29112 21048 29121
rect 21364 29112 21416 29164
rect 21824 29189 21833 29223
rect 21833 29189 21867 29223
rect 21867 29189 21876 29223
rect 21824 29180 21876 29189
rect 22008 29223 22060 29232
rect 22008 29189 22017 29223
rect 22017 29189 22051 29223
rect 22051 29189 22060 29223
rect 24308 29248 24360 29300
rect 25412 29248 25464 29300
rect 31668 29248 31720 29300
rect 32864 29291 32916 29300
rect 32864 29257 32873 29291
rect 32873 29257 32907 29291
rect 32907 29257 32916 29291
rect 32864 29248 32916 29257
rect 33324 29248 33376 29300
rect 34060 29291 34112 29300
rect 34060 29257 34069 29291
rect 34069 29257 34103 29291
rect 34103 29257 34112 29291
rect 34060 29248 34112 29257
rect 22008 29180 22060 29189
rect 22744 29223 22796 29232
rect 22744 29189 22753 29223
rect 22753 29189 22787 29223
rect 22787 29189 22796 29223
rect 22744 29180 22796 29189
rect 22468 29112 22520 29164
rect 22836 29112 22888 29164
rect 23020 29155 23072 29164
rect 23020 29121 23043 29155
rect 23043 29121 23072 29155
rect 23020 29112 23072 29121
rect 23250 29155 23302 29164
rect 23250 29121 23268 29155
rect 23268 29121 23302 29155
rect 23250 29112 23302 29121
rect 23480 29112 23532 29164
rect 24400 29155 24452 29164
rect 24400 29121 24434 29155
rect 24434 29121 24452 29155
rect 19616 29087 19668 29096
rect 18972 28976 19024 29028
rect 19248 28976 19300 29028
rect 19616 29053 19625 29087
rect 19625 29053 19659 29087
rect 19659 29053 19668 29087
rect 19616 29044 19668 29053
rect 20168 28976 20220 29028
rect 21824 28976 21876 29028
rect 22100 29044 22152 29096
rect 24400 29112 24452 29121
rect 24676 29112 24728 29164
rect 25964 29155 26016 29164
rect 25964 29121 25973 29155
rect 25973 29121 26007 29155
rect 26007 29121 26016 29155
rect 25964 29112 26016 29121
rect 26148 29155 26200 29164
rect 26148 29121 26157 29155
rect 26157 29121 26191 29155
rect 26191 29121 26200 29155
rect 26148 29112 26200 29121
rect 26608 29112 26660 29164
rect 27068 29180 27120 29232
rect 30104 29180 30156 29232
rect 29092 29155 29144 29164
rect 29092 29121 29126 29155
rect 29126 29121 29144 29155
rect 29092 29112 29144 29121
rect 29368 29112 29420 29164
rect 30380 29112 30432 29164
rect 31300 29087 31352 29096
rect 31300 29053 31309 29087
rect 31309 29053 31343 29087
rect 31343 29053 31352 29087
rect 31300 29044 31352 29053
rect 31668 29112 31720 29164
rect 31852 29112 31904 29164
rect 33048 29112 33100 29164
rect 33600 29180 33652 29232
rect 33508 29155 33560 29164
rect 33508 29121 33517 29155
rect 33517 29121 33551 29155
rect 33551 29121 33560 29155
rect 33508 29112 33560 29121
rect 33876 29112 33928 29164
rect 22560 28976 22612 29028
rect 22652 28976 22704 29028
rect 22100 28908 22152 28960
rect 22284 28908 22336 28960
rect 23940 28908 23992 28960
rect 25688 28908 25740 28960
rect 28724 28908 28776 28960
rect 32496 28976 32548 29028
rect 30196 28951 30248 28960
rect 30196 28917 30205 28951
rect 30205 28917 30239 28951
rect 30239 28917 30248 28951
rect 30196 28908 30248 28917
rect 6582 28806 6634 28858
rect 6646 28806 6698 28858
rect 6710 28806 6762 28858
rect 6774 28806 6826 28858
rect 6838 28806 6890 28858
rect 17846 28806 17898 28858
rect 17910 28806 17962 28858
rect 17974 28806 18026 28858
rect 18038 28806 18090 28858
rect 18102 28806 18154 28858
rect 29110 28806 29162 28858
rect 29174 28806 29226 28858
rect 29238 28806 29290 28858
rect 29302 28806 29354 28858
rect 29366 28806 29418 28858
rect 16580 28704 16632 28756
rect 16672 28704 16724 28756
rect 19064 28704 19116 28756
rect 16212 28636 16264 28688
rect 17500 28636 17552 28688
rect 18512 28636 18564 28688
rect 18604 28636 18656 28688
rect 18880 28636 18932 28688
rect 12164 28568 12216 28620
rect 16120 28568 16172 28620
rect 18972 28568 19024 28620
rect 19524 28704 19576 28756
rect 19616 28704 19668 28756
rect 20260 28636 20312 28688
rect 20444 28636 20496 28688
rect 22008 28704 22060 28756
rect 22100 28704 22152 28756
rect 21088 28679 21140 28688
rect 21088 28645 21097 28679
rect 21097 28645 21131 28679
rect 21131 28645 21140 28679
rect 21088 28636 21140 28645
rect 22192 28636 22244 28688
rect 13452 28500 13504 28552
rect 13728 28500 13780 28552
rect 14648 28543 14700 28552
rect 14648 28509 14657 28543
rect 14657 28509 14691 28543
rect 14691 28509 14700 28543
rect 14648 28500 14700 28509
rect 14832 28500 14884 28552
rect 15108 28500 15160 28552
rect 15292 28543 15344 28552
rect 15292 28509 15301 28543
rect 15301 28509 15335 28543
rect 15335 28509 15344 28543
rect 15292 28500 15344 28509
rect 15476 28500 15528 28552
rect 16948 28500 17000 28552
rect 17316 28500 17368 28552
rect 13268 28432 13320 28484
rect 16856 28364 16908 28416
rect 17776 28432 17828 28484
rect 19340 28432 19392 28484
rect 19708 28432 19760 28484
rect 20260 28500 20312 28552
rect 21364 28500 21416 28552
rect 22468 28611 22520 28620
rect 22468 28577 22477 28611
rect 22477 28577 22511 28611
rect 22511 28577 22520 28611
rect 23572 28704 23624 28756
rect 28080 28704 28132 28756
rect 29000 28704 29052 28756
rect 23848 28636 23900 28688
rect 24216 28636 24268 28688
rect 27528 28636 27580 28688
rect 28632 28636 28684 28688
rect 22468 28568 22520 28577
rect 22560 28500 22612 28552
rect 22744 28543 22796 28552
rect 22744 28509 22778 28543
rect 22778 28509 22796 28543
rect 22744 28500 22796 28509
rect 27252 28543 27304 28552
rect 23020 28432 23072 28484
rect 23572 28432 23624 28484
rect 24768 28475 24820 28484
rect 24768 28441 24777 28475
rect 24777 28441 24811 28475
rect 24811 28441 24820 28475
rect 24768 28432 24820 28441
rect 18328 28407 18380 28416
rect 18328 28373 18337 28407
rect 18337 28373 18371 28407
rect 18371 28373 18380 28407
rect 18328 28364 18380 28373
rect 18512 28407 18564 28416
rect 18512 28373 18521 28407
rect 18521 28373 18555 28407
rect 18555 28373 18564 28407
rect 18512 28364 18564 28373
rect 18696 28407 18748 28416
rect 18696 28373 18705 28407
rect 18705 28373 18739 28407
rect 18739 28373 18748 28407
rect 18696 28364 18748 28373
rect 18880 28364 18932 28416
rect 19156 28364 19208 28416
rect 19616 28364 19668 28416
rect 19800 28364 19852 28416
rect 22284 28364 22336 28416
rect 22376 28364 22428 28416
rect 23112 28364 23164 28416
rect 23204 28364 23256 28416
rect 24216 28364 24268 28416
rect 24676 28364 24728 28416
rect 27252 28509 27261 28543
rect 27261 28509 27295 28543
rect 27295 28509 27304 28543
rect 27252 28500 27304 28509
rect 27436 28543 27488 28552
rect 27436 28509 27445 28543
rect 27445 28509 27479 28543
rect 27479 28509 27488 28543
rect 27436 28500 27488 28509
rect 27988 28543 28040 28552
rect 27068 28432 27120 28484
rect 27528 28432 27580 28484
rect 27988 28509 27997 28543
rect 27997 28509 28031 28543
rect 28031 28509 28040 28543
rect 27988 28500 28040 28509
rect 28264 28568 28316 28620
rect 30104 28611 30156 28620
rect 30104 28577 30113 28611
rect 30113 28577 30147 28611
rect 30147 28577 30156 28611
rect 30104 28568 30156 28577
rect 31576 28568 31628 28620
rect 29000 28543 29052 28552
rect 29000 28509 29009 28543
rect 29009 28509 29043 28543
rect 29043 28509 29052 28543
rect 29000 28500 29052 28509
rect 30196 28500 30248 28552
rect 31944 28543 31996 28552
rect 31944 28509 31953 28543
rect 31953 28509 31987 28543
rect 31987 28509 31996 28543
rect 31944 28500 31996 28509
rect 32128 28500 32180 28552
rect 32956 28568 33008 28620
rect 32588 28500 32640 28552
rect 33232 28636 33284 28688
rect 33324 28543 33376 28552
rect 29460 28432 29512 28484
rect 27988 28364 28040 28416
rect 28908 28364 28960 28416
rect 29000 28364 29052 28416
rect 29920 28364 29972 28416
rect 31392 28364 31444 28416
rect 32036 28364 32088 28416
rect 32772 28364 32824 28416
rect 33324 28509 33333 28543
rect 33333 28509 33367 28543
rect 33367 28509 33376 28543
rect 33324 28500 33376 28509
rect 33784 28543 33836 28552
rect 33784 28509 33793 28543
rect 33793 28509 33827 28543
rect 33827 28509 33836 28543
rect 33784 28500 33836 28509
rect 33692 28432 33744 28484
rect 33508 28364 33560 28416
rect 12214 28262 12266 28314
rect 12278 28262 12330 28314
rect 12342 28262 12394 28314
rect 12406 28262 12458 28314
rect 12470 28262 12522 28314
rect 23478 28262 23530 28314
rect 23542 28262 23594 28314
rect 23606 28262 23658 28314
rect 23670 28262 23722 28314
rect 23734 28262 23786 28314
rect 13268 28203 13320 28212
rect 13268 28169 13277 28203
rect 13277 28169 13311 28203
rect 13311 28169 13320 28203
rect 13268 28160 13320 28169
rect 17408 28160 17460 28212
rect 20260 28160 20312 28212
rect 21272 28203 21324 28212
rect 21272 28169 21281 28203
rect 21281 28169 21315 28203
rect 21315 28169 21324 28203
rect 21272 28160 21324 28169
rect 21916 28160 21968 28212
rect 22376 28160 22428 28212
rect 23020 28160 23072 28212
rect 23940 28203 23992 28212
rect 23940 28169 23949 28203
rect 23949 28169 23983 28203
rect 23983 28169 23992 28203
rect 23940 28160 23992 28169
rect 26148 28160 26200 28212
rect 26332 28203 26384 28212
rect 26332 28169 26341 28203
rect 26341 28169 26375 28203
rect 26375 28169 26384 28203
rect 26332 28160 26384 28169
rect 27252 28160 27304 28212
rect 27344 28160 27396 28212
rect 31392 28160 31444 28212
rect 13820 28092 13872 28144
rect 14648 28135 14700 28144
rect 14648 28101 14657 28135
rect 14657 28101 14691 28135
rect 14691 28101 14700 28135
rect 14648 28092 14700 28101
rect 15108 28092 15160 28144
rect 14004 28024 14056 28076
rect 14464 28024 14516 28076
rect 14556 28067 14608 28076
rect 14556 28033 14565 28067
rect 14565 28033 14599 28067
rect 14599 28033 14608 28067
rect 14556 28024 14608 28033
rect 14924 28024 14976 28076
rect 15200 28067 15252 28076
rect 15200 28033 15209 28067
rect 15209 28033 15243 28067
rect 15243 28033 15252 28067
rect 15200 28024 15252 28033
rect 15752 28024 15804 28076
rect 16212 28092 16264 28144
rect 16672 28092 16724 28144
rect 18512 28092 18564 28144
rect 18880 28092 18932 28144
rect 19064 28092 19116 28144
rect 16120 28067 16172 28076
rect 16120 28033 16129 28067
rect 16129 28033 16163 28067
rect 16163 28033 16172 28067
rect 16120 28024 16172 28033
rect 16304 28024 16356 28076
rect 14188 27956 14240 28008
rect 14556 27888 14608 27940
rect 16764 27956 16816 28008
rect 17132 28067 17184 28076
rect 17132 28033 17141 28067
rect 17141 28033 17175 28067
rect 17175 28033 17184 28067
rect 17132 28024 17184 28033
rect 17316 28024 17368 28076
rect 18052 28067 18104 28076
rect 18052 28033 18061 28067
rect 18061 28033 18095 28067
rect 18095 28033 18104 28067
rect 18052 28024 18104 28033
rect 17960 27956 18012 28008
rect 19524 28024 19576 28076
rect 21088 28092 21140 28144
rect 22468 28092 22520 28144
rect 22560 28092 22612 28144
rect 24124 28092 24176 28144
rect 24400 28092 24452 28144
rect 24492 28092 24544 28144
rect 16396 27888 16448 27940
rect 15752 27820 15804 27872
rect 17316 27820 17368 27872
rect 17592 27888 17644 27940
rect 19800 27956 19852 28008
rect 21180 27956 21232 28008
rect 21916 27956 21968 28008
rect 22100 28024 22152 28076
rect 22284 28067 22336 28076
rect 22284 28033 22293 28067
rect 22293 28033 22327 28067
rect 22327 28033 22336 28067
rect 22744 28067 22796 28076
rect 22284 28024 22336 28033
rect 22744 28033 22753 28067
rect 22753 28033 22787 28067
rect 22787 28033 22796 28067
rect 22744 28024 22796 28033
rect 22836 28067 22888 28076
rect 22836 28033 22846 28067
rect 22846 28033 22880 28067
rect 22880 28033 22888 28067
rect 23020 28067 23072 28076
rect 22836 28024 22888 28033
rect 23020 28033 23029 28067
rect 23029 28033 23063 28067
rect 23063 28033 23072 28067
rect 23020 28024 23072 28033
rect 23112 28067 23164 28076
rect 23112 28033 23121 28067
rect 23121 28033 23155 28067
rect 23155 28033 23164 28067
rect 23112 28024 23164 28033
rect 23480 28024 23532 28076
rect 23848 28067 23900 28076
rect 23848 28033 23857 28067
rect 23857 28033 23891 28067
rect 23891 28033 23900 28067
rect 23848 28024 23900 28033
rect 24584 28024 24636 28076
rect 24676 28024 24728 28076
rect 24952 28067 25004 28076
rect 24952 28033 24961 28067
rect 24961 28033 24995 28067
rect 24995 28033 25004 28067
rect 24952 28024 25004 28033
rect 28080 28092 28132 28144
rect 25320 28067 25372 28076
rect 25320 28033 25329 28067
rect 25329 28033 25363 28067
rect 25363 28033 25372 28067
rect 25320 28024 25372 28033
rect 24308 27956 24360 28008
rect 25136 27999 25188 28008
rect 25136 27965 25145 27999
rect 25145 27965 25179 27999
rect 25179 27965 25188 27999
rect 25136 27956 25188 27965
rect 25412 27956 25464 28008
rect 19340 27888 19392 27940
rect 21824 27888 21876 27940
rect 26332 28024 26384 28076
rect 27528 28067 27580 28076
rect 26240 27956 26292 28008
rect 27528 28033 27537 28067
rect 27537 28033 27571 28067
rect 27571 28033 27580 28067
rect 27528 28024 27580 28033
rect 28816 28024 28868 28076
rect 27712 27956 27764 28008
rect 29644 28092 29696 28144
rect 29920 28024 29972 28076
rect 30380 28067 30432 28076
rect 30380 28033 30389 28067
rect 30389 28033 30423 28067
rect 30423 28033 30432 28067
rect 30380 28024 30432 28033
rect 30748 28024 30800 28076
rect 31024 28024 31076 28076
rect 27896 27888 27948 27940
rect 29552 27888 29604 27940
rect 29920 27888 29972 27940
rect 30196 27888 30248 27940
rect 32312 28067 32364 28076
rect 32312 28033 32321 28067
rect 32321 28033 32355 28067
rect 32355 28033 32364 28067
rect 32312 28024 32364 28033
rect 34152 27999 34204 28008
rect 34152 27965 34161 27999
rect 34161 27965 34195 27999
rect 34195 27965 34204 27999
rect 34152 27956 34204 27965
rect 23388 27863 23440 27872
rect 23388 27829 23397 27863
rect 23397 27829 23431 27863
rect 23431 27829 23440 27863
rect 23388 27820 23440 27829
rect 24124 27863 24176 27872
rect 24124 27829 24133 27863
rect 24133 27829 24167 27863
rect 24167 27829 24176 27863
rect 24124 27820 24176 27829
rect 25872 27820 25924 27872
rect 27804 27820 27856 27872
rect 31300 27863 31352 27872
rect 31300 27829 31309 27863
rect 31309 27829 31343 27863
rect 31343 27829 31352 27863
rect 31300 27820 31352 27829
rect 31484 27820 31536 27872
rect 31760 27820 31812 27872
rect 32864 27820 32916 27872
rect 6582 27718 6634 27770
rect 6646 27718 6698 27770
rect 6710 27718 6762 27770
rect 6774 27718 6826 27770
rect 6838 27718 6890 27770
rect 17846 27718 17898 27770
rect 17910 27718 17962 27770
rect 17974 27718 18026 27770
rect 18038 27718 18090 27770
rect 18102 27718 18154 27770
rect 29110 27718 29162 27770
rect 29174 27718 29226 27770
rect 29238 27718 29290 27770
rect 29302 27718 29354 27770
rect 29366 27718 29418 27770
rect 14464 27616 14516 27668
rect 15016 27548 15068 27600
rect 15752 27548 15804 27600
rect 18052 27548 18104 27600
rect 18420 27616 18472 27668
rect 19892 27616 19944 27668
rect 22192 27616 22244 27668
rect 22376 27616 22428 27668
rect 26240 27616 26292 27668
rect 27436 27616 27488 27668
rect 18512 27548 18564 27600
rect 15936 27480 15988 27532
rect 14372 27412 14424 27464
rect 14924 27412 14976 27464
rect 15200 27412 15252 27464
rect 15568 27412 15620 27464
rect 15752 27412 15804 27464
rect 16212 27412 16264 27464
rect 13728 27344 13780 27396
rect 16304 27344 16356 27396
rect 15292 27276 15344 27328
rect 15660 27276 15712 27328
rect 17408 27480 17460 27532
rect 17592 27480 17644 27532
rect 17132 27412 17184 27464
rect 18420 27480 18472 27532
rect 20812 27548 20864 27600
rect 19432 27523 19484 27532
rect 19432 27489 19441 27523
rect 19441 27489 19475 27523
rect 19475 27489 19484 27523
rect 19432 27480 19484 27489
rect 19616 27480 19668 27532
rect 22652 27548 22704 27600
rect 21732 27523 21784 27532
rect 18972 27412 19024 27464
rect 20812 27412 20864 27464
rect 20996 27455 21048 27464
rect 20996 27421 21005 27455
rect 21005 27421 21039 27455
rect 21039 27421 21048 27455
rect 21732 27489 21741 27523
rect 21741 27489 21775 27523
rect 21775 27489 21784 27523
rect 21732 27480 21784 27489
rect 20996 27412 21048 27421
rect 21272 27455 21324 27464
rect 21272 27421 21281 27455
rect 21281 27421 21315 27455
rect 21315 27421 21324 27455
rect 21272 27412 21324 27421
rect 16672 27344 16724 27396
rect 17592 27344 17644 27396
rect 18512 27387 18564 27396
rect 18512 27353 18521 27387
rect 18521 27353 18555 27387
rect 18555 27353 18564 27387
rect 18512 27344 18564 27353
rect 17960 27276 18012 27328
rect 18052 27276 18104 27328
rect 18972 27276 19024 27328
rect 19156 27344 19208 27396
rect 23020 27480 23072 27532
rect 21916 27412 21968 27464
rect 22100 27412 22152 27464
rect 22560 27412 22612 27464
rect 23204 27412 23256 27464
rect 23480 27548 23532 27600
rect 24124 27548 24176 27600
rect 24676 27548 24728 27600
rect 26148 27548 26200 27600
rect 28264 27616 28316 27668
rect 28172 27548 28224 27600
rect 29460 27548 29512 27600
rect 31944 27616 31996 27668
rect 33784 27616 33836 27668
rect 31668 27548 31720 27600
rect 23756 27480 23808 27532
rect 29552 27523 29604 27532
rect 29552 27489 29561 27523
rect 29561 27489 29595 27523
rect 29595 27489 29604 27523
rect 29552 27480 29604 27489
rect 29920 27480 29972 27532
rect 31024 27480 31076 27532
rect 31208 27480 31260 27532
rect 32036 27480 32088 27532
rect 23572 27412 23624 27464
rect 24492 27412 24544 27464
rect 24952 27412 25004 27464
rect 25872 27455 25924 27464
rect 25872 27421 25881 27455
rect 25881 27421 25915 27455
rect 25915 27421 25924 27455
rect 25872 27412 25924 27421
rect 25964 27455 26016 27464
rect 25964 27421 25974 27455
rect 25974 27421 26008 27455
rect 26008 27421 26016 27455
rect 26240 27455 26292 27464
rect 25964 27412 26016 27421
rect 26240 27421 26249 27455
rect 26249 27421 26283 27455
rect 26283 27421 26292 27455
rect 26240 27412 26292 27421
rect 26332 27455 26384 27464
rect 26332 27421 26346 27455
rect 26346 27421 26380 27455
rect 26380 27421 26384 27455
rect 26332 27412 26384 27421
rect 27252 27455 27304 27464
rect 27252 27421 27261 27455
rect 27261 27421 27295 27455
rect 27295 27421 27304 27455
rect 27252 27412 27304 27421
rect 27436 27412 27488 27464
rect 28724 27412 28776 27464
rect 28908 27455 28960 27464
rect 28908 27421 28917 27455
rect 28917 27421 28951 27455
rect 28951 27421 28960 27455
rect 28908 27412 28960 27421
rect 29276 27412 29328 27464
rect 30104 27412 30156 27464
rect 30288 27412 30340 27464
rect 31576 27455 31628 27464
rect 31576 27421 31585 27455
rect 31585 27421 31619 27455
rect 31619 27421 31628 27455
rect 31576 27412 31628 27421
rect 31760 27455 31812 27464
rect 31760 27421 31769 27455
rect 31769 27421 31803 27455
rect 31803 27421 31812 27455
rect 32128 27455 32180 27464
rect 31760 27412 31812 27421
rect 32128 27421 32137 27455
rect 32137 27421 32171 27455
rect 32171 27421 32180 27455
rect 32128 27412 32180 27421
rect 32312 27412 32364 27464
rect 21916 27276 21968 27328
rect 23112 27344 23164 27396
rect 25136 27344 25188 27396
rect 25780 27344 25832 27396
rect 26976 27344 27028 27396
rect 33140 27344 33192 27396
rect 28448 27276 28500 27328
rect 28632 27319 28684 27328
rect 28632 27285 28641 27319
rect 28641 27285 28675 27319
rect 28675 27285 28684 27319
rect 28632 27276 28684 27285
rect 33600 27276 33652 27328
rect 12214 27174 12266 27226
rect 12278 27174 12330 27226
rect 12342 27174 12394 27226
rect 12406 27174 12458 27226
rect 12470 27174 12522 27226
rect 23478 27174 23530 27226
rect 23542 27174 23594 27226
rect 23606 27174 23658 27226
rect 23670 27174 23722 27226
rect 23734 27174 23786 27226
rect 16948 27072 17000 27124
rect 17408 27072 17460 27124
rect 17684 27072 17736 27124
rect 17868 27072 17920 27124
rect 18788 27072 18840 27124
rect 13544 26979 13596 26988
rect 13544 26945 13553 26979
rect 13553 26945 13587 26979
rect 13587 26945 13596 26979
rect 13544 26936 13596 26945
rect 14188 26979 14240 26988
rect 14188 26945 14197 26979
rect 14197 26945 14231 26979
rect 14231 26945 14240 26979
rect 14188 26936 14240 26945
rect 16580 27004 16632 27056
rect 15476 26979 15528 26988
rect 15476 26945 15485 26979
rect 15485 26945 15519 26979
rect 15519 26945 15528 26979
rect 15476 26936 15528 26945
rect 15568 26936 15620 26988
rect 15936 26979 15988 26988
rect 15936 26945 15945 26979
rect 15945 26945 15979 26979
rect 15979 26945 15988 26979
rect 15936 26936 15988 26945
rect 17224 27004 17276 27056
rect 18696 27004 18748 27056
rect 19984 27072 20036 27124
rect 20812 27072 20864 27124
rect 21732 27072 21784 27124
rect 22744 27072 22796 27124
rect 16764 26979 16816 26988
rect 16764 26945 16773 26979
rect 16773 26945 16807 26979
rect 16807 26945 16816 26979
rect 16764 26936 16816 26945
rect 16580 26800 16632 26852
rect 16856 26868 16908 26920
rect 17224 26868 17276 26920
rect 19156 26979 19208 26988
rect 19708 27004 19760 27056
rect 19156 26945 19191 26979
rect 19191 26945 19208 26979
rect 19156 26936 19208 26945
rect 21180 27004 21232 27056
rect 21456 27004 21508 27056
rect 24400 27072 24452 27124
rect 24952 27072 25004 27124
rect 27896 27072 27948 27124
rect 28816 27115 28868 27124
rect 28816 27081 28825 27115
rect 28825 27081 28859 27115
rect 28859 27081 28868 27115
rect 28816 27072 28868 27081
rect 29920 27072 29972 27124
rect 30104 27072 30156 27124
rect 30380 27072 30432 27124
rect 30564 27072 30616 27124
rect 30932 27072 30984 27124
rect 31576 27115 31628 27124
rect 24308 27004 24360 27056
rect 30196 27047 30248 27056
rect 30196 27013 30205 27047
rect 30205 27013 30239 27047
rect 30239 27013 30248 27047
rect 30196 27004 30248 27013
rect 30656 27004 30708 27056
rect 18052 26868 18104 26920
rect 21088 26936 21140 26988
rect 21916 26979 21968 26988
rect 21916 26945 21925 26979
rect 21925 26945 21959 26979
rect 21959 26945 21968 26979
rect 21916 26936 21968 26945
rect 22100 26979 22152 26988
rect 22100 26945 22109 26979
rect 22109 26945 22143 26979
rect 22143 26945 22152 26979
rect 22100 26936 22152 26945
rect 19524 26868 19576 26920
rect 19892 26911 19944 26920
rect 19892 26877 19901 26911
rect 19901 26877 19935 26911
rect 19935 26877 19944 26911
rect 19892 26868 19944 26877
rect 20996 26868 21048 26920
rect 22836 26936 22888 26988
rect 22928 26936 22980 26988
rect 23388 26979 23440 26988
rect 23388 26945 23397 26979
rect 23397 26945 23431 26979
rect 23431 26945 23440 26979
rect 25780 26979 25832 26988
rect 23388 26936 23440 26945
rect 25780 26945 25789 26979
rect 25789 26945 25823 26979
rect 25823 26945 25832 26979
rect 25780 26936 25832 26945
rect 25964 26936 26016 26988
rect 27068 26936 27120 26988
rect 29920 26979 29972 26988
rect 14648 26775 14700 26784
rect 14648 26741 14657 26775
rect 14657 26741 14691 26775
rect 14691 26741 14700 26775
rect 14648 26732 14700 26741
rect 15660 26732 15712 26784
rect 16672 26732 16724 26784
rect 16856 26775 16908 26784
rect 16856 26741 16865 26775
rect 16865 26741 16899 26775
rect 16899 26741 16908 26775
rect 16856 26732 16908 26741
rect 18236 26800 18288 26852
rect 19524 26732 19576 26784
rect 21824 26800 21876 26852
rect 23204 26868 23256 26920
rect 23848 26911 23900 26920
rect 23848 26877 23857 26911
rect 23857 26877 23891 26911
rect 23891 26877 23900 26911
rect 23848 26868 23900 26877
rect 22468 26800 22520 26852
rect 21548 26732 21600 26784
rect 23480 26732 23532 26784
rect 26792 26732 26844 26784
rect 29920 26945 29929 26979
rect 29929 26945 29963 26979
rect 29963 26945 29972 26979
rect 29920 26936 29972 26945
rect 30012 26979 30064 26988
rect 30012 26945 30022 26979
rect 30022 26945 30056 26979
rect 30056 26945 30064 26979
rect 30012 26936 30064 26945
rect 30472 26936 30524 26988
rect 29276 26911 29328 26920
rect 29276 26877 29285 26911
rect 29285 26877 29319 26911
rect 29319 26877 29328 26911
rect 29276 26868 29328 26877
rect 27712 26732 27764 26784
rect 28264 26732 28316 26784
rect 28908 26732 28960 26784
rect 29736 26732 29788 26784
rect 31576 27081 31585 27115
rect 31585 27081 31619 27115
rect 31619 27081 31628 27115
rect 31576 27072 31628 27081
rect 32404 27072 32456 27124
rect 32956 27072 33008 27124
rect 31484 27004 31536 27056
rect 31668 27004 31720 27056
rect 31208 26868 31260 26920
rect 31760 26936 31812 26988
rect 32680 27004 32732 27056
rect 32772 26979 32824 26988
rect 32772 26945 32781 26979
rect 32781 26945 32815 26979
rect 32815 26945 32824 26979
rect 32772 26936 32824 26945
rect 33324 27072 33376 27124
rect 33600 26936 33652 26988
rect 32588 26868 32640 26920
rect 33784 26868 33836 26920
rect 31760 26732 31812 26784
rect 33140 26732 33192 26784
rect 6582 26630 6634 26682
rect 6646 26630 6698 26682
rect 6710 26630 6762 26682
rect 6774 26630 6826 26682
rect 6838 26630 6890 26682
rect 17846 26630 17898 26682
rect 17910 26630 17962 26682
rect 17974 26630 18026 26682
rect 18038 26630 18090 26682
rect 18102 26630 18154 26682
rect 29110 26630 29162 26682
rect 29174 26630 29226 26682
rect 29238 26630 29290 26682
rect 29302 26630 29354 26682
rect 29366 26630 29418 26682
rect 16672 26528 16724 26580
rect 17500 26571 17552 26580
rect 17500 26537 17509 26571
rect 17509 26537 17543 26571
rect 17543 26537 17552 26571
rect 17500 26528 17552 26537
rect 18512 26528 18564 26580
rect 18696 26528 18748 26580
rect 21088 26571 21140 26580
rect 14648 26392 14700 26444
rect 14832 26324 14884 26376
rect 15568 26367 15620 26376
rect 15292 26256 15344 26308
rect 15568 26333 15577 26367
rect 15577 26333 15611 26367
rect 15611 26333 15620 26367
rect 15568 26324 15620 26333
rect 17132 26392 17184 26444
rect 18144 26392 18196 26444
rect 18328 26460 18380 26512
rect 21088 26537 21097 26571
rect 21097 26537 21131 26571
rect 21131 26537 21140 26571
rect 21088 26528 21140 26537
rect 21364 26528 21416 26580
rect 23204 26528 23256 26580
rect 16672 26324 16724 26376
rect 17224 26324 17276 26376
rect 16304 26256 16356 26308
rect 16488 26256 16540 26308
rect 17316 26256 17368 26308
rect 18420 26324 18472 26376
rect 21456 26460 21508 26512
rect 23112 26460 23164 26512
rect 24308 26528 24360 26580
rect 25780 26528 25832 26580
rect 26056 26528 26108 26580
rect 28724 26528 28776 26580
rect 28908 26528 28960 26580
rect 29552 26528 29604 26580
rect 29920 26528 29972 26580
rect 28172 26460 28224 26512
rect 30288 26460 30340 26512
rect 30380 26460 30432 26512
rect 31300 26503 31352 26512
rect 22192 26392 22244 26444
rect 22652 26392 22704 26444
rect 29644 26435 29696 26444
rect 29644 26401 29653 26435
rect 29653 26401 29687 26435
rect 29687 26401 29696 26435
rect 29644 26392 29696 26401
rect 29736 26392 29788 26444
rect 30656 26392 30708 26444
rect 30748 26392 30800 26444
rect 31300 26469 31309 26503
rect 31309 26469 31343 26503
rect 31343 26469 31352 26503
rect 31300 26460 31352 26469
rect 31668 26460 31720 26512
rect 19340 26324 19392 26376
rect 19524 26367 19576 26376
rect 19524 26333 19558 26367
rect 19558 26333 19576 26367
rect 19524 26324 19576 26333
rect 19892 26324 19944 26376
rect 20812 26324 20864 26376
rect 21364 26324 21416 26376
rect 15016 26231 15068 26240
rect 15016 26197 15025 26231
rect 15025 26197 15059 26231
rect 15059 26197 15068 26231
rect 15016 26188 15068 26197
rect 15108 26188 15160 26240
rect 18696 26231 18748 26240
rect 18696 26197 18705 26231
rect 18705 26197 18739 26231
rect 18739 26197 18748 26231
rect 18696 26188 18748 26197
rect 19708 26256 19760 26308
rect 22100 26324 22152 26376
rect 22284 26367 22336 26376
rect 22284 26333 22293 26367
rect 22293 26333 22327 26367
rect 22327 26333 22336 26367
rect 22284 26324 22336 26333
rect 23388 26324 23440 26376
rect 22468 26256 22520 26308
rect 23296 26299 23348 26308
rect 23296 26265 23305 26299
rect 23305 26265 23339 26299
rect 23339 26265 23348 26299
rect 23296 26256 23348 26265
rect 27712 26324 27764 26376
rect 28356 26324 28408 26376
rect 25596 26256 25648 26308
rect 32128 26324 32180 26376
rect 32312 26367 32364 26376
rect 32312 26333 32321 26367
rect 32321 26333 32355 26367
rect 32355 26333 32364 26367
rect 32312 26324 32364 26333
rect 20628 26231 20680 26240
rect 20628 26197 20637 26231
rect 20637 26197 20671 26231
rect 20671 26197 20680 26231
rect 20628 26188 20680 26197
rect 23940 26188 23992 26240
rect 27436 26188 27488 26240
rect 27712 26188 27764 26240
rect 28264 26188 28316 26240
rect 28816 26231 28868 26240
rect 28816 26197 28841 26231
rect 28841 26197 28868 26231
rect 32772 26256 32824 26308
rect 32956 26256 33008 26308
rect 28816 26188 28868 26197
rect 12214 26086 12266 26138
rect 12278 26086 12330 26138
rect 12342 26086 12394 26138
rect 12406 26086 12458 26138
rect 12470 26086 12522 26138
rect 23478 26086 23530 26138
rect 23542 26086 23594 26138
rect 23606 26086 23658 26138
rect 23670 26086 23722 26138
rect 23734 26086 23786 26138
rect 18696 25984 18748 26036
rect 18788 25984 18840 26036
rect 25596 26027 25648 26036
rect 15108 25916 15160 25968
rect 15660 25916 15712 25968
rect 16764 25916 16816 25968
rect 16948 25916 17000 25968
rect 15292 25848 15344 25900
rect 16396 25848 16448 25900
rect 16580 25848 16632 25900
rect 18420 25916 18472 25968
rect 19708 25959 19760 25968
rect 18788 25848 18840 25900
rect 19432 25891 19484 25900
rect 19432 25857 19441 25891
rect 19441 25857 19475 25891
rect 19475 25857 19484 25891
rect 19432 25848 19484 25857
rect 19708 25925 19742 25959
rect 19742 25925 19760 25959
rect 19708 25916 19760 25925
rect 19800 25916 19852 25968
rect 20628 25916 20680 25968
rect 15476 25780 15528 25832
rect 15568 25780 15620 25832
rect 16856 25780 16908 25832
rect 18236 25780 18288 25832
rect 13820 25687 13872 25696
rect 13820 25653 13829 25687
rect 13829 25653 13863 25687
rect 13863 25653 13872 25687
rect 13820 25644 13872 25653
rect 16672 25644 16724 25696
rect 20812 25848 20864 25900
rect 22008 25848 22060 25900
rect 23848 25916 23900 25968
rect 25596 25993 25605 26027
rect 25605 25993 25639 26027
rect 25639 25993 25648 26027
rect 25596 25984 25648 25993
rect 27068 25984 27120 26036
rect 26056 25891 26108 25900
rect 26056 25857 26065 25891
rect 26065 25857 26099 25891
rect 26099 25857 26108 25891
rect 26056 25848 26108 25857
rect 28540 25984 28592 26036
rect 29644 25984 29696 26036
rect 33968 25984 34020 26036
rect 27344 25891 27396 25900
rect 27344 25857 27353 25891
rect 27353 25857 27387 25891
rect 27387 25857 27396 25891
rect 27344 25848 27396 25857
rect 28908 25848 28960 25900
rect 30656 25916 30708 25968
rect 30564 25848 30616 25900
rect 30932 25848 30984 25900
rect 31944 25848 31996 25900
rect 32036 25848 32088 25900
rect 34152 25891 34204 25900
rect 34152 25857 34161 25891
rect 34161 25857 34195 25891
rect 34195 25857 34204 25891
rect 34152 25848 34204 25857
rect 20720 25644 20772 25696
rect 21824 25644 21876 25696
rect 27896 25780 27948 25832
rect 28356 25823 28408 25832
rect 28356 25789 28365 25823
rect 28365 25789 28399 25823
rect 28399 25789 28408 25823
rect 28356 25780 28408 25789
rect 29736 25780 29788 25832
rect 23296 25755 23348 25764
rect 23296 25721 23305 25755
rect 23305 25721 23339 25755
rect 23339 25721 23348 25755
rect 25136 25755 25188 25764
rect 23296 25712 23348 25721
rect 25136 25721 25145 25755
rect 25145 25721 25179 25755
rect 25179 25721 25188 25755
rect 25136 25712 25188 25721
rect 28172 25712 28224 25764
rect 32036 25712 32088 25764
rect 32220 25780 32272 25832
rect 34060 25780 34112 25832
rect 25964 25687 26016 25696
rect 25964 25653 25973 25687
rect 25973 25653 26007 25687
rect 26007 25653 26016 25687
rect 25964 25644 26016 25653
rect 30472 25644 30524 25696
rect 31024 25644 31076 25696
rect 32312 25644 32364 25696
rect 6582 25542 6634 25594
rect 6646 25542 6698 25594
rect 6710 25542 6762 25594
rect 6774 25542 6826 25594
rect 6838 25542 6890 25594
rect 17846 25542 17898 25594
rect 17910 25542 17962 25594
rect 17974 25542 18026 25594
rect 18038 25542 18090 25594
rect 18102 25542 18154 25594
rect 29110 25542 29162 25594
rect 29174 25542 29226 25594
rect 29238 25542 29290 25594
rect 29302 25542 29354 25594
rect 29366 25542 29418 25594
rect 16948 25440 17000 25492
rect 17316 25440 17368 25492
rect 17500 25440 17552 25492
rect 21732 25440 21784 25492
rect 22008 25440 22060 25492
rect 1860 25347 1912 25356
rect 1860 25313 1869 25347
rect 1869 25313 1903 25347
rect 1903 25313 1912 25347
rect 1860 25304 1912 25313
rect 13820 25304 13872 25356
rect 1400 25279 1452 25288
rect 1400 25245 1409 25279
rect 1409 25245 1443 25279
rect 1443 25245 1452 25279
rect 1400 25236 1452 25245
rect 14556 25279 14608 25288
rect 14556 25245 14565 25279
rect 14565 25245 14599 25279
rect 14599 25245 14608 25279
rect 14556 25236 14608 25245
rect 15568 25304 15620 25356
rect 16396 25236 16448 25288
rect 17684 25372 17736 25424
rect 22192 25415 22244 25424
rect 22192 25381 22201 25415
rect 22201 25381 22235 25415
rect 22235 25381 22244 25415
rect 22192 25372 22244 25381
rect 17408 25304 17460 25356
rect 18328 25304 18380 25356
rect 20812 25347 20864 25356
rect 18788 25236 18840 25288
rect 20812 25313 20821 25347
rect 20821 25313 20855 25347
rect 20855 25313 20864 25347
rect 20812 25304 20864 25313
rect 23112 25304 23164 25356
rect 19432 25236 19484 25288
rect 19800 25279 19852 25288
rect 19800 25245 19809 25279
rect 19809 25245 19843 25279
rect 19843 25245 19852 25279
rect 19800 25236 19852 25245
rect 20076 25236 20128 25288
rect 20720 25236 20772 25288
rect 1584 25211 1636 25220
rect 1584 25177 1593 25211
rect 1593 25177 1627 25211
rect 1627 25177 1636 25211
rect 1584 25168 1636 25177
rect 15108 25211 15160 25220
rect 15108 25177 15117 25211
rect 15117 25177 15151 25211
rect 15151 25177 15160 25211
rect 15108 25168 15160 25177
rect 16212 25168 16264 25220
rect 17040 25168 17092 25220
rect 17684 25211 17736 25220
rect 17684 25177 17693 25211
rect 17693 25177 17727 25211
rect 17727 25177 17736 25211
rect 17684 25168 17736 25177
rect 23204 25236 23256 25288
rect 24124 25304 24176 25356
rect 25136 25440 25188 25492
rect 25504 25483 25556 25492
rect 25504 25449 25513 25483
rect 25513 25449 25547 25483
rect 25547 25449 25556 25483
rect 25504 25440 25556 25449
rect 26056 25440 26108 25492
rect 26424 25483 26476 25492
rect 26424 25449 26433 25483
rect 26433 25449 26467 25483
rect 26467 25449 26476 25483
rect 26424 25440 26476 25449
rect 27344 25440 27396 25492
rect 27988 25483 28040 25492
rect 27988 25449 27997 25483
rect 27997 25449 28031 25483
rect 28031 25449 28040 25483
rect 27988 25440 28040 25449
rect 28448 25440 28500 25492
rect 31484 25440 31536 25492
rect 24676 25372 24728 25424
rect 25964 25372 26016 25424
rect 26608 25372 26660 25424
rect 22652 25211 22704 25220
rect 22652 25177 22661 25211
rect 22661 25177 22695 25211
rect 22695 25177 22704 25211
rect 22652 25168 22704 25177
rect 15476 25100 15528 25152
rect 18144 25100 18196 25152
rect 18236 25100 18288 25152
rect 18788 25100 18840 25152
rect 20076 25100 20128 25152
rect 23388 25100 23440 25152
rect 24400 25211 24452 25220
rect 24400 25177 24409 25211
rect 24409 25177 24443 25211
rect 24443 25177 24452 25211
rect 25320 25236 25372 25288
rect 26056 25304 26108 25356
rect 26332 25304 26384 25356
rect 28172 25304 28224 25356
rect 28356 25304 28408 25356
rect 24400 25168 24452 25177
rect 24124 25100 24176 25152
rect 26056 25211 26108 25220
rect 26056 25177 26065 25211
rect 26065 25177 26099 25211
rect 26099 25177 26108 25211
rect 26056 25168 26108 25177
rect 26976 25236 27028 25288
rect 28540 25236 28592 25288
rect 28724 25279 28776 25288
rect 28724 25245 28733 25279
rect 28733 25245 28767 25279
rect 28767 25245 28776 25279
rect 28724 25236 28776 25245
rect 28816 25279 28868 25288
rect 28816 25245 28825 25279
rect 28825 25245 28859 25279
rect 28859 25245 28868 25279
rect 31116 25304 31168 25356
rect 31852 25347 31904 25356
rect 31852 25313 31861 25347
rect 31861 25313 31895 25347
rect 31895 25313 31904 25347
rect 31852 25304 31904 25313
rect 34520 25304 34572 25356
rect 28816 25236 28868 25245
rect 30196 25236 30248 25288
rect 31484 25236 31536 25288
rect 34152 25279 34204 25288
rect 34152 25245 34161 25279
rect 34161 25245 34195 25279
rect 34195 25245 34204 25279
rect 34152 25236 34204 25245
rect 28264 25100 28316 25152
rect 29644 25168 29696 25220
rect 30656 25168 30708 25220
rect 32312 25168 32364 25220
rect 33968 25168 34020 25220
rect 30932 25143 30984 25152
rect 30932 25109 30941 25143
rect 30941 25109 30975 25143
rect 30975 25109 30984 25143
rect 30932 25100 30984 25109
rect 31392 25143 31444 25152
rect 31392 25109 31401 25143
rect 31401 25109 31435 25143
rect 31435 25109 31444 25143
rect 31392 25100 31444 25109
rect 12214 24998 12266 25050
rect 12278 24998 12330 25050
rect 12342 24998 12394 25050
rect 12406 24998 12458 25050
rect 12470 24998 12522 25050
rect 23478 24998 23530 25050
rect 23542 24998 23594 25050
rect 23606 24998 23658 25050
rect 23670 24998 23722 25050
rect 23734 24998 23786 25050
rect 1584 24896 1636 24948
rect 14556 24896 14608 24948
rect 16304 24896 16356 24948
rect 19340 24896 19392 24948
rect 21916 24896 21968 24948
rect 26424 24896 26476 24948
rect 1400 24760 1452 24812
rect 4436 24760 4488 24812
rect 15844 24760 15896 24812
rect 16488 24828 16540 24880
rect 16856 24828 16908 24880
rect 18144 24828 18196 24880
rect 27712 24828 27764 24880
rect 31852 24896 31904 24948
rect 16212 24760 16264 24812
rect 17500 24760 17552 24812
rect 18052 24803 18104 24812
rect 18052 24769 18061 24803
rect 18061 24769 18095 24803
rect 18095 24769 18104 24803
rect 18052 24760 18104 24769
rect 15752 24735 15804 24744
rect 15108 24624 15160 24676
rect 15292 24667 15344 24676
rect 15292 24633 15301 24667
rect 15301 24633 15335 24667
rect 15335 24633 15344 24667
rect 15292 24624 15344 24633
rect 15752 24701 15761 24735
rect 15761 24701 15795 24735
rect 15795 24701 15804 24735
rect 15752 24692 15804 24701
rect 17868 24692 17920 24744
rect 20352 24760 20404 24812
rect 20720 24803 20772 24812
rect 20720 24769 20729 24803
rect 20729 24769 20763 24803
rect 20763 24769 20772 24803
rect 20720 24760 20772 24769
rect 21640 24760 21692 24812
rect 19432 24667 19484 24676
rect 19432 24633 19441 24667
rect 19441 24633 19475 24667
rect 19475 24633 19484 24667
rect 19432 24624 19484 24633
rect 19524 24624 19576 24676
rect 21824 24624 21876 24676
rect 22100 24760 22152 24812
rect 23940 24803 23992 24812
rect 23940 24769 23949 24803
rect 23949 24769 23983 24803
rect 23983 24769 23992 24803
rect 23940 24760 23992 24769
rect 25412 24760 25464 24812
rect 25596 24760 25648 24812
rect 23020 24692 23072 24744
rect 23664 24735 23716 24744
rect 23664 24701 23673 24735
rect 23673 24701 23707 24735
rect 23707 24701 23716 24735
rect 23664 24692 23716 24701
rect 25780 24803 25832 24812
rect 25780 24769 25789 24803
rect 25789 24769 25823 24803
rect 25823 24769 25832 24803
rect 25780 24760 25832 24769
rect 27068 24803 27120 24812
rect 25964 24692 26016 24744
rect 27068 24769 27077 24803
rect 27077 24769 27111 24803
rect 27111 24769 27120 24803
rect 27068 24760 27120 24769
rect 28632 24760 28684 24812
rect 28724 24803 28776 24812
rect 28724 24769 28733 24803
rect 28733 24769 28767 24803
rect 28767 24769 28776 24803
rect 28724 24760 28776 24769
rect 22100 24624 22152 24676
rect 17776 24556 17828 24608
rect 18420 24556 18472 24608
rect 22744 24556 22796 24608
rect 23112 24556 23164 24608
rect 27804 24624 27856 24676
rect 26700 24556 26752 24608
rect 27160 24599 27212 24608
rect 27160 24565 27169 24599
rect 27169 24565 27203 24599
rect 27203 24565 27212 24599
rect 27160 24556 27212 24565
rect 27896 24556 27948 24608
rect 29000 24692 29052 24744
rect 31024 24828 31076 24880
rect 32036 24828 32088 24880
rect 30748 24760 30800 24812
rect 31300 24760 31352 24812
rect 30196 24735 30248 24744
rect 29920 24624 29972 24676
rect 28080 24556 28132 24608
rect 29460 24556 29512 24608
rect 29736 24599 29788 24608
rect 29736 24565 29745 24599
rect 29745 24565 29779 24599
rect 29779 24565 29788 24599
rect 29736 24556 29788 24565
rect 30196 24701 30205 24735
rect 30205 24701 30239 24735
rect 30239 24701 30248 24735
rect 30196 24692 30248 24701
rect 32128 24735 32180 24744
rect 32128 24701 32137 24735
rect 32137 24701 32171 24735
rect 32171 24701 32180 24735
rect 32128 24692 32180 24701
rect 33508 24760 33560 24812
rect 34060 24803 34112 24812
rect 34060 24769 34069 24803
rect 34069 24769 34103 24803
rect 34103 24769 34112 24803
rect 34060 24760 34112 24769
rect 34060 24624 34112 24676
rect 31300 24556 31352 24608
rect 31668 24556 31720 24608
rect 32312 24556 32364 24608
rect 6582 24454 6634 24506
rect 6646 24454 6698 24506
rect 6710 24454 6762 24506
rect 6774 24454 6826 24506
rect 6838 24454 6890 24506
rect 17846 24454 17898 24506
rect 17910 24454 17962 24506
rect 17974 24454 18026 24506
rect 18038 24454 18090 24506
rect 18102 24454 18154 24506
rect 29110 24454 29162 24506
rect 29174 24454 29226 24506
rect 29238 24454 29290 24506
rect 29302 24454 29354 24506
rect 29366 24454 29418 24506
rect 15752 24352 15804 24404
rect 15108 24216 15160 24268
rect 15844 24216 15896 24268
rect 14924 24191 14976 24200
rect 14924 24157 14933 24191
rect 14933 24157 14967 24191
rect 14967 24157 14976 24191
rect 14924 24148 14976 24157
rect 15568 24148 15620 24200
rect 17408 24148 17460 24200
rect 18328 24352 18380 24404
rect 18512 24352 18564 24404
rect 25596 24352 25648 24404
rect 17868 24216 17920 24268
rect 19800 24284 19852 24336
rect 20536 24284 20588 24336
rect 22284 24284 22336 24336
rect 18144 24191 18196 24200
rect 18144 24157 18153 24191
rect 18153 24157 18187 24191
rect 18187 24157 18196 24191
rect 18144 24148 18196 24157
rect 14280 24080 14332 24132
rect 15108 24080 15160 24132
rect 16396 24123 16448 24132
rect 16396 24089 16430 24123
rect 16430 24089 16448 24123
rect 16396 24080 16448 24089
rect 16580 24080 16632 24132
rect 17040 24080 17092 24132
rect 19524 24148 19576 24200
rect 19708 24191 19760 24200
rect 19708 24157 19717 24191
rect 19717 24157 19751 24191
rect 19751 24157 19760 24191
rect 19708 24148 19760 24157
rect 21548 24216 21600 24268
rect 23112 24284 23164 24336
rect 29552 24327 29604 24336
rect 29552 24293 29561 24327
rect 29561 24293 29595 24327
rect 29595 24293 29604 24327
rect 29552 24284 29604 24293
rect 31852 24352 31904 24404
rect 32496 24352 32548 24404
rect 22560 24216 22612 24268
rect 20076 24191 20128 24200
rect 18420 24080 18472 24132
rect 20076 24157 20085 24191
rect 20085 24157 20119 24191
rect 20119 24157 20128 24191
rect 20076 24148 20128 24157
rect 21088 24148 21140 24200
rect 14740 24055 14792 24064
rect 14740 24021 14749 24055
rect 14749 24021 14783 24055
rect 14783 24021 14792 24055
rect 14740 24012 14792 24021
rect 16672 24012 16724 24064
rect 17868 24012 17920 24064
rect 17960 24012 18012 24064
rect 18328 24012 18380 24064
rect 19524 24012 19576 24064
rect 20628 24080 20680 24132
rect 21732 24080 21784 24132
rect 22192 24191 22244 24200
rect 22192 24157 22201 24191
rect 22201 24157 22235 24191
rect 22235 24157 22244 24191
rect 22468 24191 22520 24200
rect 22192 24148 22244 24157
rect 22468 24157 22477 24191
rect 22477 24157 22511 24191
rect 22511 24157 22520 24191
rect 22468 24148 22520 24157
rect 22836 24148 22888 24200
rect 23388 24191 23440 24200
rect 23388 24157 23397 24191
rect 23397 24157 23431 24191
rect 23431 24157 23440 24191
rect 23388 24148 23440 24157
rect 33140 24216 33192 24268
rect 34152 24259 34204 24268
rect 34152 24225 34161 24259
rect 34161 24225 34195 24259
rect 34195 24225 34204 24259
rect 34152 24216 34204 24225
rect 26056 24148 26108 24200
rect 26148 24148 26200 24200
rect 28356 24148 28408 24200
rect 28448 24148 28500 24200
rect 25872 24080 25924 24132
rect 28540 24080 28592 24132
rect 29644 24148 29696 24200
rect 30196 24148 30248 24200
rect 32128 24148 32180 24200
rect 28816 24080 28868 24132
rect 31392 24080 31444 24132
rect 34428 24080 34480 24132
rect 20720 24012 20772 24064
rect 21364 24012 21416 24064
rect 21640 24012 21692 24064
rect 22376 24055 22428 24064
rect 22376 24021 22385 24055
rect 22385 24021 22419 24055
rect 22419 24021 22428 24055
rect 22376 24012 22428 24021
rect 22928 24012 22980 24064
rect 23388 24012 23440 24064
rect 23940 24012 23992 24064
rect 24124 24012 24176 24064
rect 25964 24012 26016 24064
rect 26884 24055 26936 24064
rect 26884 24021 26893 24055
rect 26893 24021 26927 24055
rect 26927 24021 26936 24055
rect 26884 24012 26936 24021
rect 27160 24012 27212 24064
rect 29184 24012 29236 24064
rect 29460 24012 29512 24064
rect 29736 24055 29788 24064
rect 29736 24021 29745 24055
rect 29745 24021 29779 24055
rect 29779 24021 29788 24055
rect 29736 24012 29788 24021
rect 29920 24012 29972 24064
rect 33048 24012 33100 24064
rect 12214 23910 12266 23962
rect 12278 23910 12330 23962
rect 12342 23910 12394 23962
rect 12406 23910 12458 23962
rect 12470 23910 12522 23962
rect 23478 23910 23530 23962
rect 23542 23910 23594 23962
rect 23606 23910 23658 23962
rect 23670 23910 23722 23962
rect 23734 23910 23786 23962
rect 16672 23808 16724 23860
rect 18144 23808 18196 23860
rect 18420 23808 18472 23860
rect 18512 23808 18564 23860
rect 21456 23808 21508 23860
rect 22192 23808 22244 23860
rect 18696 23740 18748 23792
rect 21180 23740 21232 23792
rect 16488 23672 16540 23724
rect 17040 23715 17092 23724
rect 17040 23681 17049 23715
rect 17049 23681 17083 23715
rect 17083 23681 17092 23715
rect 17040 23672 17092 23681
rect 17408 23715 17460 23724
rect 17408 23681 17417 23715
rect 17417 23681 17451 23715
rect 17451 23681 17460 23715
rect 17408 23672 17460 23681
rect 19616 23672 19668 23724
rect 19892 23715 19944 23724
rect 19892 23681 19901 23715
rect 19901 23681 19935 23715
rect 19935 23681 19944 23715
rect 19892 23672 19944 23681
rect 21732 23672 21784 23724
rect 22928 23740 22980 23792
rect 22008 23672 22060 23724
rect 22284 23715 22336 23724
rect 22284 23681 22318 23715
rect 22318 23681 22336 23715
rect 22284 23672 22336 23681
rect 22468 23672 22520 23724
rect 27988 23808 28040 23860
rect 28172 23808 28224 23860
rect 28448 23808 28500 23860
rect 23940 23740 23992 23792
rect 25688 23740 25740 23792
rect 23480 23715 23532 23724
rect 23480 23681 23489 23715
rect 23489 23681 23523 23715
rect 23523 23681 23532 23715
rect 24124 23715 24176 23724
rect 23480 23672 23532 23681
rect 24124 23681 24133 23715
rect 24133 23681 24167 23715
rect 24167 23681 24176 23715
rect 24124 23672 24176 23681
rect 25228 23715 25280 23724
rect 17960 23604 18012 23656
rect 16580 23536 16632 23588
rect 15200 23468 15252 23520
rect 22008 23536 22060 23588
rect 22468 23536 22520 23588
rect 25228 23681 25237 23715
rect 25237 23681 25271 23715
rect 25271 23681 25280 23715
rect 25228 23672 25280 23681
rect 24492 23604 24544 23656
rect 27528 23715 27580 23724
rect 25504 23647 25556 23656
rect 25504 23613 25513 23647
rect 25513 23613 25547 23647
rect 25547 23613 25556 23647
rect 25504 23604 25556 23613
rect 25688 23604 25740 23656
rect 23020 23536 23072 23588
rect 27528 23681 27537 23715
rect 27537 23681 27571 23715
rect 27571 23681 27580 23715
rect 27528 23672 27580 23681
rect 29736 23808 29788 23860
rect 29920 23808 29972 23860
rect 31116 23851 31168 23860
rect 31116 23817 31125 23851
rect 31125 23817 31159 23851
rect 31159 23817 31168 23851
rect 31116 23808 31168 23817
rect 31300 23808 31352 23860
rect 31852 23808 31904 23860
rect 28724 23740 28776 23792
rect 29000 23740 29052 23792
rect 34152 23783 34204 23792
rect 34152 23749 34161 23783
rect 34161 23749 34195 23783
rect 34195 23749 34204 23783
rect 34152 23740 34204 23749
rect 27712 23604 27764 23656
rect 28172 23536 28224 23588
rect 31024 23672 31076 23724
rect 29184 23604 29236 23656
rect 29644 23604 29696 23656
rect 31392 23604 31444 23656
rect 31668 23604 31720 23656
rect 32312 23647 32364 23656
rect 32312 23613 32321 23647
rect 32321 23613 32355 23647
rect 32355 23613 32364 23647
rect 32312 23604 32364 23613
rect 32496 23647 32548 23656
rect 32496 23613 32505 23647
rect 32505 23613 32539 23647
rect 32539 23613 32548 23647
rect 32496 23604 32548 23613
rect 19248 23468 19300 23520
rect 19340 23468 19392 23520
rect 21272 23511 21324 23520
rect 21272 23477 21281 23511
rect 21281 23477 21315 23511
rect 21315 23477 21324 23511
rect 21272 23468 21324 23477
rect 24676 23468 24728 23520
rect 25780 23468 25832 23520
rect 26332 23468 26384 23520
rect 28724 23468 28776 23520
rect 29552 23468 29604 23520
rect 30564 23468 30616 23520
rect 31668 23468 31720 23520
rect 6582 23366 6634 23418
rect 6646 23366 6698 23418
rect 6710 23366 6762 23418
rect 6774 23366 6826 23418
rect 6838 23366 6890 23418
rect 17846 23366 17898 23418
rect 17910 23366 17962 23418
rect 17974 23366 18026 23418
rect 18038 23366 18090 23418
rect 18102 23366 18154 23418
rect 29110 23366 29162 23418
rect 29174 23366 29226 23418
rect 29238 23366 29290 23418
rect 29302 23366 29354 23418
rect 29366 23366 29418 23418
rect 16396 23264 16448 23316
rect 18236 23264 18288 23316
rect 22284 23196 22336 23248
rect 23480 23264 23532 23316
rect 25504 23264 25556 23316
rect 27528 23264 27580 23316
rect 28908 23264 28960 23316
rect 29736 23264 29788 23316
rect 29920 23264 29972 23316
rect 31300 23264 31352 23316
rect 16580 23171 16632 23180
rect 16580 23137 16589 23171
rect 16589 23137 16623 23171
rect 16623 23137 16632 23171
rect 16580 23128 16632 23137
rect 15200 23060 15252 23112
rect 15844 23060 15896 23112
rect 17776 23060 17828 23112
rect 19248 23103 19300 23112
rect 19248 23069 19257 23103
rect 19257 23069 19291 23103
rect 19291 23069 19300 23103
rect 19248 23060 19300 23069
rect 20720 23128 20772 23180
rect 20996 23060 21048 23112
rect 16396 22992 16448 23044
rect 16948 22992 17000 23044
rect 19064 22992 19116 23044
rect 21364 23128 21416 23180
rect 22744 23128 22796 23180
rect 23112 23128 23164 23180
rect 23204 23128 23256 23180
rect 25136 23171 25188 23180
rect 21824 23103 21876 23112
rect 21824 23069 21833 23103
rect 21833 23069 21867 23103
rect 21867 23069 21876 23103
rect 21824 23060 21876 23069
rect 22008 23103 22060 23112
rect 22008 23069 22017 23103
rect 22017 23069 22051 23103
rect 22051 23069 22060 23103
rect 22008 23060 22060 23069
rect 21548 22992 21600 23044
rect 22192 22992 22244 23044
rect 22928 23060 22980 23112
rect 25136 23137 25145 23171
rect 25145 23137 25179 23171
rect 25179 23137 25188 23171
rect 25136 23128 25188 23137
rect 24952 23060 25004 23112
rect 23020 22992 23072 23044
rect 25412 23128 25464 23180
rect 25596 23060 25648 23112
rect 28172 23196 28224 23248
rect 27804 23128 27856 23180
rect 26056 23103 26108 23112
rect 26056 23069 26065 23103
rect 26065 23069 26099 23103
rect 26099 23069 26108 23103
rect 26056 23060 26108 23069
rect 26332 23103 26384 23112
rect 26332 23069 26366 23103
rect 26366 23069 26384 23103
rect 26332 23060 26384 23069
rect 27896 23103 27948 23112
rect 27896 23069 27905 23103
rect 27905 23069 27939 23103
rect 27939 23069 27948 23103
rect 27896 23060 27948 23069
rect 16488 22924 16540 22976
rect 20444 22924 20496 22976
rect 20628 22967 20680 22976
rect 20628 22933 20637 22967
rect 20637 22933 20671 22967
rect 20671 22933 20680 22967
rect 20628 22924 20680 22933
rect 20812 22924 20864 22976
rect 24124 22924 24176 22976
rect 27528 22924 27580 22976
rect 28172 23035 28224 23044
rect 28172 23001 28181 23035
rect 28181 23001 28215 23035
rect 28215 23001 28224 23035
rect 29368 23196 29420 23248
rect 28908 23128 28960 23180
rect 29000 23060 29052 23112
rect 31300 23128 31352 23180
rect 32036 23128 32088 23180
rect 33324 23128 33376 23180
rect 34152 23171 34204 23180
rect 34152 23137 34161 23171
rect 34161 23137 34195 23171
rect 34195 23137 34204 23171
rect 34152 23128 34204 23137
rect 28172 22992 28224 23001
rect 29368 22992 29420 23044
rect 30564 22992 30616 23044
rect 33692 22992 33744 23044
rect 30196 22924 30248 22976
rect 30380 22924 30432 22976
rect 12214 22822 12266 22874
rect 12278 22822 12330 22874
rect 12342 22822 12394 22874
rect 12406 22822 12458 22874
rect 12470 22822 12522 22874
rect 23478 22822 23530 22874
rect 23542 22822 23594 22874
rect 23606 22822 23658 22874
rect 23670 22822 23722 22874
rect 23734 22822 23786 22874
rect 14372 22720 14424 22772
rect 17776 22720 17828 22772
rect 18328 22720 18380 22772
rect 19064 22763 19116 22772
rect 19064 22729 19073 22763
rect 19073 22729 19107 22763
rect 19107 22729 19116 22763
rect 19064 22720 19116 22729
rect 21916 22720 21968 22772
rect 23112 22720 23164 22772
rect 24860 22720 24912 22772
rect 16396 22652 16448 22704
rect 16580 22652 16632 22704
rect 16488 22584 16540 22636
rect 16764 22652 16816 22704
rect 19248 22652 19300 22704
rect 16580 22516 16632 22568
rect 18420 22584 18472 22636
rect 19524 22627 19576 22636
rect 19524 22593 19533 22627
rect 19533 22593 19567 22627
rect 19567 22593 19576 22627
rect 19524 22584 19576 22593
rect 20076 22627 20128 22636
rect 20076 22593 20085 22627
rect 20085 22593 20119 22627
rect 20119 22593 20128 22627
rect 20076 22584 20128 22593
rect 20352 22627 20404 22636
rect 20352 22593 20361 22627
rect 20361 22593 20395 22627
rect 20395 22593 20404 22627
rect 20352 22584 20404 22593
rect 19156 22516 19208 22568
rect 19800 22516 19852 22568
rect 20536 22516 20588 22568
rect 20996 22516 21048 22568
rect 23940 22652 23992 22704
rect 22928 22584 22980 22636
rect 24400 22584 24452 22636
rect 24584 22584 24636 22636
rect 25044 22627 25096 22636
rect 25044 22593 25053 22627
rect 25053 22593 25087 22627
rect 25087 22593 25096 22627
rect 25044 22584 25096 22593
rect 28264 22720 28316 22772
rect 28908 22720 28960 22772
rect 30564 22720 30616 22772
rect 25228 22652 25280 22704
rect 25596 22652 25648 22704
rect 25872 22652 25924 22704
rect 25504 22584 25556 22636
rect 25964 22627 26016 22636
rect 25964 22593 25973 22627
rect 25973 22593 26007 22627
rect 26007 22593 26016 22627
rect 25964 22584 26016 22593
rect 31668 22720 31720 22772
rect 31300 22652 31352 22704
rect 28448 22584 28500 22636
rect 26148 22559 26200 22568
rect 20628 22448 20680 22500
rect 16580 22380 16632 22432
rect 17040 22380 17092 22432
rect 17776 22380 17828 22432
rect 19984 22380 20036 22432
rect 22100 22380 22152 22432
rect 24308 22448 24360 22500
rect 26148 22525 26157 22559
rect 26157 22525 26191 22559
rect 26191 22525 26200 22559
rect 26148 22516 26200 22525
rect 26240 22559 26292 22568
rect 26240 22525 26249 22559
rect 26249 22525 26283 22559
rect 26283 22525 26292 22559
rect 27252 22559 27304 22568
rect 26240 22516 26292 22525
rect 27252 22525 27261 22559
rect 27261 22525 27295 22559
rect 27295 22525 27304 22559
rect 27252 22516 27304 22525
rect 27344 22516 27396 22568
rect 27988 22516 28040 22568
rect 30380 22584 30432 22636
rect 30472 22584 30524 22636
rect 29000 22516 29052 22568
rect 30932 22516 30984 22568
rect 31852 22516 31904 22568
rect 24492 22380 24544 22432
rect 26332 22380 26384 22432
rect 30380 22448 30432 22500
rect 32772 22584 32824 22636
rect 32956 22627 33008 22636
rect 32956 22593 32965 22627
rect 32965 22593 32999 22627
rect 32999 22593 33008 22627
rect 32956 22584 33008 22593
rect 33876 22584 33928 22636
rect 33324 22516 33376 22568
rect 32772 22448 32824 22500
rect 30104 22380 30156 22432
rect 31760 22380 31812 22432
rect 31852 22380 31904 22432
rect 32680 22380 32732 22432
rect 32864 22380 32916 22432
rect 6582 22278 6634 22330
rect 6646 22278 6698 22330
rect 6710 22278 6762 22330
rect 6774 22278 6826 22330
rect 6838 22278 6890 22330
rect 17846 22278 17898 22330
rect 17910 22278 17962 22330
rect 17974 22278 18026 22330
rect 18038 22278 18090 22330
rect 18102 22278 18154 22330
rect 29110 22278 29162 22330
rect 29174 22278 29226 22330
rect 29238 22278 29290 22330
rect 29302 22278 29354 22330
rect 29366 22278 29418 22330
rect 16764 22176 16816 22228
rect 17040 22176 17092 22228
rect 19340 22219 19392 22228
rect 19340 22185 19349 22219
rect 19349 22185 19383 22219
rect 19383 22185 19392 22219
rect 19340 22176 19392 22185
rect 19432 22176 19484 22228
rect 21088 22176 21140 22228
rect 21364 22176 21416 22228
rect 22928 22219 22980 22228
rect 22928 22185 22937 22219
rect 22937 22185 22971 22219
rect 22971 22185 22980 22219
rect 22928 22176 22980 22185
rect 23112 22176 23164 22228
rect 27988 22176 28040 22228
rect 28264 22176 28316 22228
rect 19156 22108 19208 22160
rect 23296 22108 23348 22160
rect 19340 22040 19392 22092
rect 19616 22040 19668 22092
rect 16028 21972 16080 22024
rect 16488 21972 16540 22024
rect 17408 21972 17460 22024
rect 19432 22015 19484 22024
rect 19432 21981 19441 22015
rect 19441 21981 19475 22015
rect 19475 21981 19484 22015
rect 19432 21972 19484 21981
rect 19524 22015 19576 22024
rect 19524 21981 19533 22015
rect 19533 21981 19567 22015
rect 19567 21981 19576 22015
rect 19524 21972 19576 21981
rect 17040 21904 17092 21956
rect 18512 21836 18564 21888
rect 19340 21904 19392 21956
rect 21456 22040 21508 22092
rect 21364 21972 21416 22024
rect 21824 21972 21876 22024
rect 22744 22040 22796 22092
rect 25872 22108 25924 22160
rect 27252 22108 27304 22160
rect 22008 22015 22060 22024
rect 22008 21981 22017 22015
rect 22017 21981 22051 22015
rect 22051 21981 22060 22015
rect 22008 21972 22060 21981
rect 22192 21972 22244 22024
rect 23204 22015 23256 22024
rect 23204 21981 23213 22015
rect 23213 21981 23247 22015
rect 23247 21981 23256 22015
rect 23204 21972 23256 21981
rect 23020 21904 23072 21956
rect 23388 22015 23440 22024
rect 23388 21981 23397 22015
rect 23397 21981 23431 22015
rect 23431 21981 23440 22015
rect 23940 22040 23992 22092
rect 24952 22083 25004 22092
rect 23388 21972 23440 21981
rect 24124 21972 24176 22024
rect 24308 21972 24360 22024
rect 24584 22015 24636 22024
rect 24584 21981 24593 22015
rect 24593 21981 24627 22015
rect 24627 21981 24636 22015
rect 24584 21972 24636 21981
rect 24952 22049 24961 22083
rect 24961 22049 24995 22083
rect 24995 22049 25004 22083
rect 24952 22040 25004 22049
rect 25320 21972 25372 22024
rect 25596 22040 25648 22092
rect 27896 22083 27948 22092
rect 27896 22049 27905 22083
rect 27905 22049 27939 22083
rect 27939 22049 27948 22083
rect 27896 22040 27948 22049
rect 25504 21972 25556 22024
rect 26056 22015 26108 22024
rect 26056 21981 26065 22015
rect 26065 21981 26099 22015
rect 26099 21981 26108 22015
rect 26056 21972 26108 21981
rect 26332 22015 26384 22024
rect 26332 21981 26366 22015
rect 26366 21981 26384 22015
rect 26332 21972 26384 21981
rect 29184 22108 29236 22160
rect 25044 21904 25096 21956
rect 19524 21836 19576 21888
rect 19708 21879 19760 21888
rect 19708 21845 19717 21879
rect 19717 21845 19751 21879
rect 19751 21845 19760 21879
rect 19708 21836 19760 21845
rect 24400 21836 24452 21888
rect 27160 21904 27212 21956
rect 27896 21904 27948 21956
rect 28172 22015 28224 22024
rect 28172 21981 28181 22015
rect 28181 21981 28215 22015
rect 28215 21981 28224 22015
rect 28172 21972 28224 21981
rect 29920 22176 29972 22228
rect 31668 22176 31720 22228
rect 32036 22176 32088 22228
rect 32956 22176 33008 22228
rect 33324 22176 33376 22228
rect 29920 22040 29972 22092
rect 30012 22040 30064 22092
rect 31392 22108 31444 22160
rect 28264 21904 28316 21956
rect 29276 21904 29328 21956
rect 27252 21836 27304 21888
rect 28080 21836 28132 21888
rect 30288 21904 30340 21956
rect 31668 22040 31720 22092
rect 31024 21972 31076 22024
rect 31760 21972 31812 22024
rect 32864 22083 32916 22092
rect 32864 22049 32873 22083
rect 32873 22049 32907 22083
rect 32907 22049 32916 22083
rect 32864 22040 32916 22049
rect 33692 22083 33744 22092
rect 33692 22049 33701 22083
rect 33701 22049 33735 22083
rect 33735 22049 33744 22083
rect 33692 22040 33744 22049
rect 32404 21972 32456 22024
rect 33600 22015 33652 22024
rect 33600 21981 33609 22015
rect 33609 21981 33643 22015
rect 33643 21981 33652 22015
rect 33600 21972 33652 21981
rect 32864 21904 32916 21956
rect 33324 21904 33376 21956
rect 29644 21836 29696 21888
rect 30472 21836 30524 21888
rect 30932 21836 30984 21888
rect 31576 21836 31628 21888
rect 12214 21734 12266 21786
rect 12278 21734 12330 21786
rect 12342 21734 12394 21786
rect 12406 21734 12458 21786
rect 12470 21734 12522 21786
rect 23478 21734 23530 21786
rect 23542 21734 23594 21786
rect 23606 21734 23658 21786
rect 23670 21734 23722 21786
rect 23734 21734 23786 21786
rect 16580 21496 16632 21548
rect 17408 21539 17460 21548
rect 17408 21505 17417 21539
rect 17417 21505 17451 21539
rect 17451 21505 17460 21539
rect 17408 21496 17460 21505
rect 19524 21632 19576 21684
rect 19800 21632 19852 21684
rect 24400 21632 24452 21684
rect 24768 21632 24820 21684
rect 18328 21539 18380 21548
rect 18328 21505 18362 21539
rect 18362 21505 18380 21539
rect 18328 21496 18380 21505
rect 21088 21564 21140 21616
rect 21364 21564 21416 21616
rect 19984 21496 20036 21548
rect 21824 21539 21876 21548
rect 21824 21505 21833 21539
rect 21833 21505 21867 21539
rect 21867 21505 21876 21539
rect 21824 21496 21876 21505
rect 22376 21496 22428 21548
rect 22836 21539 22888 21548
rect 22836 21505 22845 21539
rect 22845 21505 22879 21539
rect 22879 21505 22888 21539
rect 22836 21496 22888 21505
rect 23112 21539 23164 21548
rect 23112 21505 23121 21539
rect 23121 21505 23155 21539
rect 23155 21505 23164 21539
rect 23112 21496 23164 21505
rect 23572 21539 23624 21548
rect 23572 21505 23581 21539
rect 23581 21505 23615 21539
rect 23615 21505 23624 21539
rect 23572 21496 23624 21505
rect 16948 21360 17000 21412
rect 21640 21428 21692 21480
rect 23940 21496 23992 21548
rect 24308 21496 24360 21548
rect 24492 21496 24544 21548
rect 27252 21632 27304 21684
rect 27160 21564 27212 21616
rect 27712 21632 27764 21684
rect 29644 21632 29696 21684
rect 30012 21632 30064 21684
rect 31392 21632 31444 21684
rect 31576 21632 31628 21684
rect 32128 21632 32180 21684
rect 32496 21632 32548 21684
rect 33968 21632 34020 21684
rect 25780 21539 25832 21548
rect 23388 21360 23440 21412
rect 17224 21292 17276 21344
rect 18236 21292 18288 21344
rect 19432 21335 19484 21344
rect 19432 21301 19441 21335
rect 19441 21301 19475 21335
rect 19475 21301 19484 21335
rect 19432 21292 19484 21301
rect 24584 21428 24636 21480
rect 25780 21505 25789 21539
rect 25789 21505 25823 21539
rect 25823 21505 25832 21539
rect 25780 21496 25832 21505
rect 25320 21428 25372 21480
rect 25964 21428 26016 21480
rect 27344 21539 27396 21548
rect 27344 21505 27353 21539
rect 27353 21505 27387 21539
rect 27387 21505 27396 21539
rect 27344 21496 27396 21505
rect 27528 21428 27580 21480
rect 28172 21496 28224 21548
rect 33232 21564 33284 21616
rect 30472 21496 30524 21548
rect 30656 21496 30708 21548
rect 31024 21496 31076 21548
rect 25136 21360 25188 21412
rect 27068 21360 27120 21412
rect 25688 21292 25740 21344
rect 26332 21292 26384 21344
rect 29552 21292 29604 21344
rect 29920 21360 29972 21412
rect 30472 21360 30524 21412
rect 31852 21360 31904 21412
rect 30656 21292 30708 21344
rect 31576 21292 31628 21344
rect 33784 21496 33836 21548
rect 33876 21496 33928 21548
rect 6582 21190 6634 21242
rect 6646 21190 6698 21242
rect 6710 21190 6762 21242
rect 6774 21190 6826 21242
rect 6838 21190 6890 21242
rect 17846 21190 17898 21242
rect 17910 21190 17962 21242
rect 17974 21190 18026 21242
rect 18038 21190 18090 21242
rect 18102 21190 18154 21242
rect 29110 21190 29162 21242
rect 29174 21190 29226 21242
rect 29238 21190 29290 21242
rect 29302 21190 29354 21242
rect 29366 21190 29418 21242
rect 17040 21131 17092 21140
rect 17040 21097 17049 21131
rect 17049 21097 17083 21131
rect 17083 21097 17092 21131
rect 17040 21088 17092 21097
rect 19984 21088 20036 21140
rect 20536 21131 20588 21140
rect 20536 21097 20545 21131
rect 20545 21097 20579 21131
rect 20579 21097 20588 21131
rect 20536 21088 20588 21097
rect 22376 21088 22428 21140
rect 22744 21088 22796 21140
rect 24308 21088 24360 21140
rect 24860 21088 24912 21140
rect 17408 21020 17460 21072
rect 17224 20927 17276 20936
rect 17224 20893 17233 20927
rect 17233 20893 17267 20927
rect 17267 20893 17276 20927
rect 17224 20884 17276 20893
rect 18236 20884 18288 20936
rect 23296 21020 23348 21072
rect 20812 20952 20864 21004
rect 21088 20995 21140 21004
rect 21088 20961 21097 20995
rect 21097 20961 21131 20995
rect 21131 20961 21140 20995
rect 21088 20952 21140 20961
rect 19984 20927 20036 20936
rect 19984 20893 19993 20927
rect 19993 20893 20027 20927
rect 20027 20893 20036 20927
rect 19984 20884 20036 20893
rect 20444 20927 20496 20936
rect 20444 20893 20453 20927
rect 20453 20893 20487 20927
rect 20487 20893 20496 20927
rect 20444 20884 20496 20893
rect 23020 20952 23072 21004
rect 24676 21020 24728 21072
rect 26148 21088 26200 21140
rect 26700 21088 26752 21140
rect 29460 21088 29512 21140
rect 25412 21020 25464 21072
rect 30656 21088 30708 21140
rect 31576 21131 31628 21140
rect 31576 21097 31585 21131
rect 31585 21097 31619 21131
rect 31619 21097 31628 21131
rect 31576 21088 31628 21097
rect 32312 21088 32364 21140
rect 23204 20927 23256 20936
rect 23204 20893 23213 20927
rect 23213 20893 23247 20927
rect 23247 20893 23256 20927
rect 23204 20884 23256 20893
rect 23388 20927 23440 20936
rect 23388 20893 23397 20927
rect 23397 20893 23431 20927
rect 23431 20893 23440 20927
rect 24768 20952 24820 21004
rect 27712 20995 27764 21004
rect 23388 20884 23440 20893
rect 24860 20884 24912 20936
rect 27712 20961 27721 20995
rect 27721 20961 27755 20995
rect 27755 20961 27764 20995
rect 27712 20952 27764 20961
rect 25044 20884 25096 20936
rect 25504 20884 25556 20936
rect 15292 20816 15344 20868
rect 25688 20859 25740 20868
rect 25688 20825 25722 20859
rect 25722 20825 25740 20859
rect 27252 20884 27304 20936
rect 27528 20927 27580 20936
rect 27528 20893 27537 20927
rect 27537 20893 27571 20927
rect 27571 20893 27580 20927
rect 28172 20952 28224 21004
rect 27528 20884 27580 20893
rect 27896 20884 27948 20936
rect 28724 20927 28776 20936
rect 28724 20893 28733 20927
rect 28733 20893 28767 20927
rect 28767 20893 28776 20927
rect 28724 20884 28776 20893
rect 29000 20884 29052 20936
rect 29460 20884 29512 20936
rect 33048 20952 33100 21004
rect 25688 20816 25740 20825
rect 16856 20748 16908 20800
rect 22376 20748 22428 20800
rect 23848 20748 23900 20800
rect 24584 20748 24636 20800
rect 26884 20748 26936 20800
rect 29644 20748 29696 20800
rect 30196 20816 30248 20868
rect 31024 20748 31076 20800
rect 33140 20884 33192 20936
rect 34336 20816 34388 20868
rect 33324 20791 33376 20800
rect 33324 20757 33333 20791
rect 33333 20757 33367 20791
rect 33367 20757 33376 20791
rect 33324 20748 33376 20757
rect 12214 20646 12266 20698
rect 12278 20646 12330 20698
rect 12342 20646 12394 20698
rect 12406 20646 12458 20698
rect 12470 20646 12522 20698
rect 23478 20646 23530 20698
rect 23542 20646 23594 20698
rect 23606 20646 23658 20698
rect 23670 20646 23722 20698
rect 23734 20646 23786 20698
rect 16120 20544 16172 20596
rect 22376 20544 22428 20596
rect 22468 20544 22520 20596
rect 23112 20544 23164 20596
rect 22008 20476 22060 20528
rect 18512 20451 18564 20460
rect 18512 20417 18521 20451
rect 18521 20417 18555 20451
rect 18555 20417 18564 20451
rect 18512 20408 18564 20417
rect 21088 20451 21140 20460
rect 21088 20417 21097 20451
rect 21097 20417 21131 20451
rect 21131 20417 21140 20451
rect 21088 20408 21140 20417
rect 21272 20451 21324 20460
rect 21272 20417 21281 20451
rect 21281 20417 21315 20451
rect 21315 20417 21324 20451
rect 21272 20408 21324 20417
rect 21640 20408 21692 20460
rect 23480 20476 23532 20528
rect 23112 20408 23164 20460
rect 23940 20544 23992 20596
rect 24124 20544 24176 20596
rect 24308 20544 24360 20596
rect 21824 20340 21876 20392
rect 22560 20340 22612 20392
rect 18328 20315 18380 20324
rect 18328 20281 18337 20315
rect 18337 20281 18371 20315
rect 18371 20281 18380 20315
rect 18328 20272 18380 20281
rect 22652 20272 22704 20324
rect 23572 20340 23624 20392
rect 24492 20476 24544 20528
rect 28172 20544 28224 20596
rect 28632 20544 28684 20596
rect 29368 20544 29420 20596
rect 24952 20451 25004 20460
rect 24952 20417 24961 20451
rect 24961 20417 24995 20451
rect 24995 20417 25004 20451
rect 24952 20408 25004 20417
rect 25780 20408 25832 20460
rect 25964 20451 26016 20460
rect 25964 20417 25973 20451
rect 25973 20417 26007 20451
rect 26007 20417 26016 20451
rect 25964 20408 26016 20417
rect 26148 20451 26200 20460
rect 26148 20417 26157 20451
rect 26157 20417 26191 20451
rect 26191 20417 26200 20451
rect 26148 20408 26200 20417
rect 26332 20451 26384 20460
rect 26332 20417 26341 20451
rect 26341 20417 26375 20451
rect 26375 20417 26384 20451
rect 26332 20408 26384 20417
rect 26700 20408 26752 20460
rect 27160 20451 27212 20460
rect 27160 20417 27169 20451
rect 27169 20417 27203 20451
rect 27203 20417 27212 20451
rect 27160 20408 27212 20417
rect 27344 20451 27396 20460
rect 27344 20417 27353 20451
rect 27353 20417 27387 20451
rect 27387 20417 27396 20451
rect 27344 20408 27396 20417
rect 23848 20272 23900 20324
rect 22284 20204 22336 20256
rect 22928 20204 22980 20256
rect 24124 20340 24176 20392
rect 26516 20340 26568 20392
rect 26240 20272 26292 20324
rect 29460 20408 29512 20460
rect 30472 20476 30524 20528
rect 31576 20476 31628 20528
rect 33324 20476 33376 20528
rect 28724 20272 28776 20324
rect 31852 20408 31904 20460
rect 34152 20451 34204 20460
rect 34152 20417 34161 20451
rect 34161 20417 34195 20451
rect 34195 20417 34204 20451
rect 34152 20408 34204 20417
rect 31024 20340 31076 20392
rect 30196 20315 30248 20324
rect 30196 20281 30205 20315
rect 30205 20281 30239 20315
rect 30239 20281 30248 20315
rect 30196 20272 30248 20281
rect 24492 20204 24544 20256
rect 28632 20204 28684 20256
rect 29460 20247 29512 20256
rect 29460 20213 29469 20247
rect 29469 20213 29503 20247
rect 29503 20213 29512 20247
rect 29460 20204 29512 20213
rect 30104 20247 30156 20256
rect 30104 20213 30113 20247
rect 30113 20213 30147 20247
rect 30147 20213 30156 20247
rect 30104 20204 30156 20213
rect 30932 20204 30984 20256
rect 31760 20204 31812 20256
rect 6582 20102 6634 20154
rect 6646 20102 6698 20154
rect 6710 20102 6762 20154
rect 6774 20102 6826 20154
rect 6838 20102 6890 20154
rect 17846 20102 17898 20154
rect 17910 20102 17962 20154
rect 17974 20102 18026 20154
rect 18038 20102 18090 20154
rect 18102 20102 18154 20154
rect 29110 20102 29162 20154
rect 29174 20102 29226 20154
rect 29238 20102 29290 20154
rect 29302 20102 29354 20154
rect 29366 20102 29418 20154
rect 19984 20000 20036 20052
rect 22836 20000 22888 20052
rect 26240 20043 26292 20052
rect 26240 20009 26249 20043
rect 26249 20009 26283 20043
rect 26283 20009 26292 20043
rect 26240 20000 26292 20009
rect 27896 20000 27948 20052
rect 23480 19932 23532 19984
rect 22284 19907 22336 19916
rect 22284 19873 22293 19907
rect 22293 19873 22327 19907
rect 22327 19873 22336 19907
rect 22284 19864 22336 19873
rect 23296 19907 23348 19916
rect 23296 19873 23305 19907
rect 23305 19873 23339 19907
rect 23339 19873 23348 19907
rect 26148 19932 26200 19984
rect 24492 19907 24544 19916
rect 23296 19864 23348 19873
rect 24492 19873 24501 19907
rect 24501 19873 24535 19907
rect 24535 19873 24544 19907
rect 24492 19864 24544 19873
rect 24768 19864 24820 19916
rect 1768 19796 1820 19848
rect 21732 19796 21784 19848
rect 22192 19839 22244 19848
rect 22192 19805 22201 19839
rect 22201 19805 22235 19839
rect 22235 19805 22244 19839
rect 22192 19796 22244 19805
rect 23572 19796 23624 19848
rect 23848 19796 23900 19848
rect 25228 19796 25280 19848
rect 26332 19796 26384 19848
rect 27160 19839 27212 19848
rect 27160 19805 27169 19839
rect 27169 19805 27203 19839
rect 27203 19805 27212 19839
rect 27160 19796 27212 19805
rect 28080 20000 28132 20052
rect 28356 20000 28408 20052
rect 28632 19864 28684 19916
rect 29460 19932 29512 19984
rect 27528 19796 27580 19848
rect 27988 19796 28040 19848
rect 29460 19796 29512 19848
rect 30012 19932 30064 19984
rect 30196 20000 30248 20052
rect 32128 19932 32180 19984
rect 30656 19839 30708 19848
rect 30656 19805 30665 19839
rect 30665 19805 30699 19839
rect 30699 19805 30708 19839
rect 30656 19796 30708 19805
rect 22560 19728 22612 19780
rect 22652 19728 22704 19780
rect 26976 19771 27028 19780
rect 26976 19737 26985 19771
rect 26985 19737 27019 19771
rect 27019 19737 27028 19771
rect 26976 19728 27028 19737
rect 22928 19660 22980 19712
rect 25228 19660 25280 19712
rect 26516 19660 26568 19712
rect 28448 19728 28500 19780
rect 28816 19728 28868 19780
rect 30472 19771 30524 19780
rect 29368 19660 29420 19712
rect 30472 19737 30481 19771
rect 30481 19737 30515 19771
rect 30515 19737 30524 19771
rect 30472 19728 30524 19737
rect 30932 19728 30984 19780
rect 31852 19796 31904 19848
rect 33232 19728 33284 19780
rect 34152 19771 34204 19780
rect 34152 19737 34161 19771
rect 34161 19737 34195 19771
rect 34195 19737 34204 19771
rect 34152 19728 34204 19737
rect 12214 19558 12266 19610
rect 12278 19558 12330 19610
rect 12342 19558 12394 19610
rect 12406 19558 12458 19610
rect 12470 19558 12522 19610
rect 23478 19558 23530 19610
rect 23542 19558 23594 19610
rect 23606 19558 23658 19610
rect 23670 19558 23722 19610
rect 23734 19558 23786 19610
rect 1768 19363 1820 19372
rect 1768 19329 1777 19363
rect 1777 19329 1811 19363
rect 1811 19329 1820 19363
rect 1768 19320 1820 19329
rect 21364 19456 21416 19508
rect 22376 19456 22428 19508
rect 23940 19456 23992 19508
rect 20812 19363 20864 19372
rect 20812 19329 20821 19363
rect 20821 19329 20855 19363
rect 20855 19329 20864 19363
rect 20812 19320 20864 19329
rect 21364 19320 21416 19372
rect 1952 19295 2004 19304
rect 1952 19261 1961 19295
rect 1961 19261 1995 19295
rect 1995 19261 2004 19295
rect 1952 19252 2004 19261
rect 2228 19295 2280 19304
rect 2228 19261 2237 19295
rect 2237 19261 2271 19295
rect 2271 19261 2280 19295
rect 2228 19252 2280 19261
rect 22284 19388 22336 19440
rect 22376 19363 22428 19372
rect 22376 19329 22385 19363
rect 22385 19329 22419 19363
rect 22419 19329 22428 19363
rect 22376 19320 22428 19329
rect 22468 19320 22520 19372
rect 23388 19388 23440 19440
rect 27252 19456 27304 19508
rect 26976 19388 27028 19440
rect 27804 19456 27856 19508
rect 29276 19456 29328 19508
rect 30656 19499 30708 19508
rect 30656 19465 30665 19499
rect 30665 19465 30699 19499
rect 30699 19465 30708 19499
rect 30656 19456 30708 19465
rect 31576 19456 31628 19508
rect 32128 19499 32180 19508
rect 32128 19465 32137 19499
rect 32137 19465 32171 19499
rect 32171 19465 32180 19499
rect 32128 19456 32180 19465
rect 33232 19499 33284 19508
rect 33232 19465 33241 19499
rect 33241 19465 33275 19499
rect 33275 19465 33284 19499
rect 33232 19456 33284 19465
rect 33416 19456 33468 19508
rect 24216 19320 24268 19372
rect 24952 19363 25004 19372
rect 24952 19329 24961 19363
rect 24961 19329 24995 19363
rect 24995 19329 25004 19363
rect 24952 19320 25004 19329
rect 27252 19363 27304 19372
rect 23204 19295 23256 19304
rect 23204 19261 23213 19295
rect 23213 19261 23247 19295
rect 23247 19261 23256 19295
rect 23204 19252 23256 19261
rect 23848 19252 23900 19304
rect 24400 19252 24452 19304
rect 25136 19252 25188 19304
rect 25412 19252 25464 19304
rect 27252 19329 27261 19363
rect 27261 19329 27295 19363
rect 27295 19329 27304 19363
rect 27252 19320 27304 19329
rect 27712 19388 27764 19440
rect 29368 19388 29420 19440
rect 27528 19295 27580 19304
rect 27528 19261 27537 19295
rect 27537 19261 27571 19295
rect 27571 19261 27580 19295
rect 27528 19252 27580 19261
rect 28724 19320 28776 19372
rect 29000 19320 29052 19372
rect 31576 19320 31628 19372
rect 31760 19320 31812 19372
rect 34060 19320 34112 19372
rect 28724 19184 28776 19236
rect 23388 19116 23440 19168
rect 25136 19116 25188 19168
rect 26424 19116 26476 19168
rect 27068 19159 27120 19168
rect 27068 19125 27077 19159
rect 27077 19125 27111 19159
rect 27111 19125 27120 19159
rect 27068 19116 27120 19125
rect 28632 19116 28684 19168
rect 30380 19184 30432 19236
rect 31944 19116 31996 19168
rect 6582 19014 6634 19066
rect 6646 19014 6698 19066
rect 6710 19014 6762 19066
rect 6774 19014 6826 19066
rect 6838 19014 6890 19066
rect 17846 19014 17898 19066
rect 17910 19014 17962 19066
rect 17974 19014 18026 19066
rect 18038 19014 18090 19066
rect 18102 19014 18154 19066
rect 29110 19014 29162 19066
rect 29174 19014 29226 19066
rect 29238 19014 29290 19066
rect 29302 19014 29354 19066
rect 29366 19014 29418 19066
rect 1952 18912 2004 18964
rect 22192 18912 22244 18964
rect 22376 18912 22428 18964
rect 24952 18912 25004 18964
rect 25872 18912 25924 18964
rect 28724 18955 28776 18964
rect 28724 18921 28733 18955
rect 28733 18921 28767 18955
rect 28767 18921 28776 18955
rect 28724 18912 28776 18921
rect 30932 18955 30984 18964
rect 30932 18921 30941 18955
rect 30941 18921 30975 18955
rect 30975 18921 30984 18955
rect 30932 18912 30984 18921
rect 31208 18912 31260 18964
rect 1492 18708 1544 18760
rect 16488 18708 16540 18760
rect 22928 18776 22980 18828
rect 23296 18819 23348 18828
rect 23296 18785 23305 18819
rect 23305 18785 23339 18819
rect 23339 18785 23348 18819
rect 23296 18776 23348 18785
rect 23848 18776 23900 18828
rect 21916 18751 21968 18760
rect 21916 18717 21925 18751
rect 21925 18717 21959 18751
rect 21959 18717 21968 18751
rect 21916 18708 21968 18717
rect 22560 18751 22612 18760
rect 22560 18717 22569 18751
rect 22569 18717 22603 18751
rect 22603 18717 22612 18751
rect 22560 18708 22612 18717
rect 23204 18708 23256 18760
rect 25136 18844 25188 18896
rect 24308 18776 24360 18828
rect 24768 18819 24820 18828
rect 24768 18785 24777 18819
rect 24777 18785 24811 18819
rect 24811 18785 24820 18819
rect 24768 18776 24820 18785
rect 24216 18708 24268 18760
rect 22744 18640 22796 18692
rect 25044 18708 25096 18760
rect 29000 18708 29052 18760
rect 30104 18708 30156 18760
rect 34244 18844 34296 18896
rect 34152 18819 34204 18828
rect 34152 18785 34161 18819
rect 34161 18785 34195 18819
rect 34195 18785 34204 18819
rect 34152 18776 34204 18785
rect 32312 18751 32364 18760
rect 32312 18717 32321 18751
rect 32321 18717 32355 18751
rect 32355 18717 32364 18751
rect 32312 18708 32364 18717
rect 25504 18683 25556 18692
rect 24952 18572 25004 18624
rect 25504 18649 25538 18683
rect 25538 18649 25556 18683
rect 25504 18640 25556 18649
rect 27896 18640 27948 18692
rect 33692 18640 33744 18692
rect 26516 18572 26568 18624
rect 12214 18470 12266 18522
rect 12278 18470 12330 18522
rect 12342 18470 12394 18522
rect 12406 18470 12458 18522
rect 12470 18470 12522 18522
rect 23478 18470 23530 18522
rect 23542 18470 23594 18522
rect 23606 18470 23658 18522
rect 23670 18470 23722 18522
rect 23734 18470 23786 18522
rect 21916 18368 21968 18420
rect 25596 18368 25648 18420
rect 25780 18368 25832 18420
rect 26424 18411 26476 18420
rect 26424 18377 26433 18411
rect 26433 18377 26467 18411
rect 26467 18377 26476 18411
rect 26424 18368 26476 18377
rect 27528 18368 27580 18420
rect 29644 18411 29696 18420
rect 29644 18377 29653 18411
rect 29653 18377 29687 18411
rect 29687 18377 29696 18411
rect 29644 18368 29696 18377
rect 29736 18368 29788 18420
rect 30748 18368 30800 18420
rect 32588 18411 32640 18420
rect 32588 18377 32597 18411
rect 32597 18377 32631 18411
rect 32631 18377 32640 18411
rect 32588 18368 32640 18377
rect 33692 18411 33744 18420
rect 33692 18377 33701 18411
rect 33701 18377 33735 18411
rect 33735 18377 33744 18411
rect 33692 18368 33744 18377
rect 1492 18275 1544 18284
rect 1492 18241 1501 18275
rect 1501 18241 1535 18275
rect 1535 18241 1544 18275
rect 1492 18232 1544 18241
rect 23296 18300 23348 18352
rect 22744 18232 22796 18284
rect 23388 18232 23440 18284
rect 24860 18300 24912 18352
rect 24676 18232 24728 18284
rect 25044 18275 25096 18284
rect 25044 18241 25053 18275
rect 25053 18241 25087 18275
rect 25087 18241 25096 18275
rect 25044 18232 25096 18241
rect 25136 18232 25188 18284
rect 27068 18300 27120 18352
rect 28724 18232 28776 18284
rect 29920 18300 29972 18352
rect 31116 18300 31168 18352
rect 30012 18232 30064 18284
rect 30380 18275 30432 18284
rect 1676 18207 1728 18216
rect 1676 18173 1685 18207
rect 1685 18173 1719 18207
rect 1719 18173 1728 18207
rect 1676 18164 1728 18173
rect 2872 18207 2924 18216
rect 2872 18173 2881 18207
rect 2881 18173 2915 18207
rect 2915 18173 2924 18207
rect 2872 18164 2924 18173
rect 23848 18164 23900 18216
rect 30380 18241 30389 18275
rect 30389 18241 30423 18275
rect 30423 18241 30432 18275
rect 30380 18232 30432 18241
rect 31392 18275 31444 18284
rect 31392 18241 31401 18275
rect 31401 18241 31435 18275
rect 31435 18241 31444 18275
rect 31392 18232 31444 18241
rect 32956 18300 33008 18352
rect 32496 18275 32548 18284
rect 32496 18241 32505 18275
rect 32505 18241 32539 18275
rect 32539 18241 32548 18275
rect 32496 18232 32548 18241
rect 32680 18232 32732 18284
rect 33600 18275 33652 18284
rect 33600 18241 33609 18275
rect 33609 18241 33643 18275
rect 33643 18241 33652 18275
rect 33600 18232 33652 18241
rect 24860 18096 24912 18148
rect 31668 18164 31720 18216
rect 30656 18096 30708 18148
rect 28816 18028 28868 18080
rect 29000 18071 29052 18080
rect 29000 18037 29009 18071
rect 29009 18037 29043 18071
rect 29043 18037 29052 18071
rect 29000 18028 29052 18037
rect 6582 17926 6634 17978
rect 6646 17926 6698 17978
rect 6710 17926 6762 17978
rect 6774 17926 6826 17978
rect 6838 17926 6890 17978
rect 17846 17926 17898 17978
rect 17910 17926 17962 17978
rect 17974 17926 18026 17978
rect 18038 17926 18090 17978
rect 18102 17926 18154 17978
rect 29110 17926 29162 17978
rect 29174 17926 29226 17978
rect 29238 17926 29290 17978
rect 29302 17926 29354 17978
rect 29366 17926 29418 17978
rect 1676 17824 1728 17876
rect 25504 17824 25556 17876
rect 25872 17824 25924 17876
rect 26884 17824 26936 17876
rect 27252 17824 27304 17876
rect 28540 17867 28592 17876
rect 28540 17833 28549 17867
rect 28549 17833 28583 17867
rect 28583 17833 28592 17867
rect 28540 17824 28592 17833
rect 28908 17824 28960 17876
rect 31484 17824 31536 17876
rect 24492 17756 24544 17808
rect 1860 17688 1912 17740
rect 4804 17688 4856 17740
rect 24768 17688 24820 17740
rect 1768 17663 1820 17672
rect 1768 17629 1777 17663
rect 1777 17629 1811 17663
rect 1811 17629 1820 17663
rect 1768 17620 1820 17629
rect 24952 17663 25004 17672
rect 24952 17629 24961 17663
rect 24961 17629 24995 17663
rect 24995 17629 25004 17663
rect 24952 17620 25004 17629
rect 25228 17663 25280 17672
rect 25228 17629 25237 17663
rect 25237 17629 25271 17663
rect 25271 17629 25280 17663
rect 25228 17620 25280 17629
rect 25780 17620 25832 17672
rect 27528 17663 27580 17672
rect 25044 17552 25096 17604
rect 25412 17552 25464 17604
rect 27528 17629 27537 17663
rect 27537 17629 27571 17663
rect 27571 17629 27580 17663
rect 27528 17620 27580 17629
rect 27712 17620 27764 17672
rect 30380 17688 30432 17740
rect 24584 17484 24636 17536
rect 28448 17552 28500 17604
rect 30196 17620 30248 17672
rect 30564 17663 30616 17672
rect 30564 17629 30573 17663
rect 30573 17629 30607 17663
rect 30607 17629 30616 17663
rect 30564 17620 30616 17629
rect 32496 17688 32548 17740
rect 34152 17731 34204 17740
rect 34152 17697 34161 17731
rect 34161 17697 34195 17731
rect 34195 17697 34204 17731
rect 34152 17688 34204 17697
rect 29460 17552 29512 17604
rect 25964 17527 26016 17536
rect 25964 17493 25973 17527
rect 25973 17493 26007 17527
rect 26007 17493 26016 17527
rect 25964 17484 26016 17493
rect 29552 17484 29604 17536
rect 31484 17484 31536 17536
rect 31944 17620 31996 17672
rect 33784 17552 33836 17604
rect 32404 17484 32456 17536
rect 12214 17382 12266 17434
rect 12278 17382 12330 17434
rect 12342 17382 12394 17434
rect 12406 17382 12458 17434
rect 12470 17382 12522 17434
rect 23478 17382 23530 17434
rect 23542 17382 23594 17434
rect 23606 17382 23658 17434
rect 23670 17382 23722 17434
rect 23734 17382 23786 17434
rect 5080 17280 5132 17332
rect 1676 17119 1728 17128
rect 1676 17085 1685 17119
rect 1685 17085 1719 17119
rect 1719 17085 1728 17119
rect 1676 17076 1728 17085
rect 1952 17119 2004 17128
rect 1952 17085 1961 17119
rect 1961 17085 1995 17119
rect 1995 17085 2004 17119
rect 1952 17076 2004 17085
rect 12900 17076 12952 17128
rect 24492 17076 24544 17128
rect 25044 17280 25096 17332
rect 25320 17280 25372 17332
rect 27896 17323 27948 17332
rect 27896 17289 27905 17323
rect 27905 17289 27939 17323
rect 27939 17289 27948 17323
rect 27896 17280 27948 17289
rect 30472 17280 30524 17332
rect 25964 17212 26016 17264
rect 24952 17187 25004 17196
rect 24952 17153 24961 17187
rect 24961 17153 24995 17187
rect 24995 17153 25004 17187
rect 24952 17144 25004 17153
rect 25412 17187 25464 17196
rect 25412 17153 25421 17187
rect 25421 17153 25455 17187
rect 25455 17153 25464 17187
rect 25412 17144 25464 17153
rect 25688 17144 25740 17196
rect 29000 17212 29052 17264
rect 30288 17187 30340 17196
rect 2596 17008 2648 17060
rect 25136 17008 25188 17060
rect 27712 17076 27764 17128
rect 30288 17153 30297 17187
rect 30297 17153 30331 17187
rect 30331 17153 30340 17187
rect 30288 17144 30340 17153
rect 32312 17212 32364 17264
rect 31300 17144 31352 17196
rect 31484 17144 31536 17196
rect 31852 17144 31904 17196
rect 32036 17076 32088 17128
rect 33140 17076 33192 17128
rect 34152 17119 34204 17128
rect 34152 17085 34161 17119
rect 34161 17085 34195 17119
rect 34195 17085 34204 17119
rect 34152 17076 34204 17085
rect 32956 17008 33008 17060
rect 31668 16940 31720 16992
rect 33416 16940 33468 16992
rect 6582 16838 6634 16890
rect 6646 16838 6698 16890
rect 6710 16838 6762 16890
rect 6774 16838 6826 16890
rect 6838 16838 6890 16890
rect 17846 16838 17898 16890
rect 17910 16838 17962 16890
rect 17974 16838 18026 16890
rect 18038 16838 18090 16890
rect 18102 16838 18154 16890
rect 29110 16838 29162 16890
rect 29174 16838 29226 16890
rect 29238 16838 29290 16890
rect 29302 16838 29354 16890
rect 29366 16838 29418 16890
rect 1676 16736 1728 16788
rect 2596 16779 2648 16788
rect 2596 16745 2605 16779
rect 2605 16745 2639 16779
rect 2639 16745 2648 16779
rect 2596 16736 2648 16745
rect 31024 16779 31076 16788
rect 31024 16745 31033 16779
rect 31033 16745 31067 16779
rect 31067 16745 31076 16779
rect 31024 16736 31076 16745
rect 32312 16736 32364 16788
rect 34520 16668 34572 16720
rect 1676 16600 1728 16652
rect 1860 16600 1912 16652
rect 30104 16600 30156 16652
rect 31668 16600 31720 16652
rect 32864 16600 32916 16652
rect 32956 16600 33008 16652
rect 32404 16532 32456 16584
rect 33416 16600 33468 16652
rect 33140 16575 33192 16584
rect 33140 16541 33149 16575
rect 33149 16541 33183 16575
rect 33183 16541 33192 16575
rect 33140 16532 33192 16541
rect 33784 16575 33836 16584
rect 33784 16541 33793 16575
rect 33793 16541 33827 16575
rect 33827 16541 33836 16575
rect 33784 16532 33836 16541
rect 32128 16396 32180 16448
rect 12214 16294 12266 16346
rect 12278 16294 12330 16346
rect 12342 16294 12394 16346
rect 12406 16294 12458 16346
rect 12470 16294 12522 16346
rect 23478 16294 23530 16346
rect 23542 16294 23594 16346
rect 23606 16294 23658 16346
rect 23670 16294 23722 16346
rect 23734 16294 23786 16346
rect 34152 16167 34204 16176
rect 34152 16133 34161 16167
rect 34161 16133 34195 16167
rect 34195 16133 34204 16167
rect 34152 16124 34204 16133
rect 31944 16056 31996 16108
rect 32312 16099 32364 16108
rect 32312 16065 32321 16099
rect 32321 16065 32355 16099
rect 32355 16065 32364 16099
rect 32312 16056 32364 16065
rect 32036 15988 32088 16040
rect 33692 15988 33744 16040
rect 1400 15852 1452 15904
rect 6582 15750 6634 15802
rect 6646 15750 6698 15802
rect 6710 15750 6762 15802
rect 6774 15750 6826 15802
rect 6838 15750 6890 15802
rect 17846 15750 17898 15802
rect 17910 15750 17962 15802
rect 17974 15750 18026 15802
rect 18038 15750 18090 15802
rect 18102 15750 18154 15802
rect 29110 15750 29162 15802
rect 29174 15750 29226 15802
rect 29238 15750 29290 15802
rect 29302 15750 29354 15802
rect 29366 15750 29418 15802
rect 33692 15691 33744 15700
rect 33692 15657 33701 15691
rect 33701 15657 33735 15691
rect 33735 15657 33744 15691
rect 33692 15648 33744 15657
rect 34428 15580 34480 15632
rect 1400 15555 1452 15564
rect 1400 15521 1409 15555
rect 1409 15521 1443 15555
rect 1443 15521 1452 15555
rect 1400 15512 1452 15521
rect 2780 15555 2832 15564
rect 2780 15521 2789 15555
rect 2789 15521 2823 15555
rect 2823 15521 2832 15555
rect 2780 15512 2832 15521
rect 33600 15487 33652 15496
rect 33600 15453 33609 15487
rect 33609 15453 33643 15487
rect 33643 15453 33652 15487
rect 33600 15444 33652 15453
rect 1584 15419 1636 15428
rect 1584 15385 1593 15419
rect 1593 15385 1627 15419
rect 1627 15385 1636 15419
rect 1584 15376 1636 15385
rect 12214 15206 12266 15258
rect 12278 15206 12330 15258
rect 12342 15206 12394 15258
rect 12406 15206 12458 15258
rect 12470 15206 12522 15258
rect 23478 15206 23530 15258
rect 23542 15206 23594 15258
rect 23606 15206 23658 15258
rect 23670 15206 23722 15258
rect 23734 15206 23786 15258
rect 1584 15104 1636 15156
rect 2228 14968 2280 15020
rect 32956 14968 33008 15020
rect 1400 14764 1452 14816
rect 32312 14764 32364 14816
rect 33140 14807 33192 14816
rect 33140 14773 33149 14807
rect 33149 14773 33183 14807
rect 33183 14773 33192 14807
rect 33140 14764 33192 14773
rect 33784 14807 33836 14816
rect 33784 14773 33793 14807
rect 33793 14773 33827 14807
rect 33827 14773 33836 14807
rect 33784 14764 33836 14773
rect 6582 14662 6634 14714
rect 6646 14662 6698 14714
rect 6710 14662 6762 14714
rect 6774 14662 6826 14714
rect 6838 14662 6890 14714
rect 17846 14662 17898 14714
rect 17910 14662 17962 14714
rect 17974 14662 18026 14714
rect 18038 14662 18090 14714
rect 18102 14662 18154 14714
rect 29110 14662 29162 14714
rect 29174 14662 29226 14714
rect 29238 14662 29290 14714
rect 29302 14662 29354 14714
rect 29366 14662 29418 14714
rect 1400 14467 1452 14476
rect 1400 14433 1409 14467
rect 1409 14433 1443 14467
rect 1443 14433 1452 14467
rect 1400 14424 1452 14433
rect 1952 14467 2004 14476
rect 1952 14433 1961 14467
rect 1961 14433 1995 14467
rect 1995 14433 2004 14467
rect 1952 14424 2004 14433
rect 32312 14467 32364 14476
rect 32312 14433 32321 14467
rect 32321 14433 32355 14467
rect 32355 14433 32364 14467
rect 32312 14424 32364 14433
rect 33140 14424 33192 14476
rect 1860 14288 1912 14340
rect 34152 14331 34204 14340
rect 34152 14297 34161 14331
rect 34161 14297 34195 14331
rect 34195 14297 34204 14331
rect 34152 14288 34204 14297
rect 12214 14118 12266 14170
rect 12278 14118 12330 14170
rect 12342 14118 12394 14170
rect 12406 14118 12458 14170
rect 12470 14118 12522 14170
rect 23478 14118 23530 14170
rect 23542 14118 23594 14170
rect 23606 14118 23658 14170
rect 23670 14118 23722 14170
rect 23734 14118 23786 14170
rect 1860 14059 1912 14068
rect 1860 14025 1869 14059
rect 1869 14025 1903 14059
rect 1903 14025 1912 14059
rect 1860 14016 1912 14025
rect 33784 13948 33836 14000
rect 1676 13880 1728 13932
rect 1860 13880 1912 13932
rect 3056 13880 3108 13932
rect 7932 13880 7984 13932
rect 34152 13855 34204 13864
rect 34152 13821 34161 13855
rect 34161 13821 34195 13855
rect 34195 13821 34204 13855
rect 34152 13812 34204 13821
rect 1584 13676 1636 13728
rect 3424 13719 3476 13728
rect 3424 13685 3433 13719
rect 3433 13685 3467 13719
rect 3467 13685 3476 13719
rect 3424 13676 3476 13685
rect 6582 13574 6634 13626
rect 6646 13574 6698 13626
rect 6710 13574 6762 13626
rect 6774 13574 6826 13626
rect 6838 13574 6890 13626
rect 17846 13574 17898 13626
rect 17910 13574 17962 13626
rect 17974 13574 18026 13626
rect 18038 13574 18090 13626
rect 18102 13574 18154 13626
rect 29110 13574 29162 13626
rect 29174 13574 29226 13626
rect 29238 13574 29290 13626
rect 29302 13574 29354 13626
rect 29366 13574 29418 13626
rect 3424 13404 3476 13456
rect 1584 13379 1636 13388
rect 1584 13345 1593 13379
rect 1593 13345 1627 13379
rect 1627 13345 1636 13379
rect 1584 13336 1636 13345
rect 2780 13379 2832 13388
rect 2780 13345 2789 13379
rect 2789 13345 2823 13379
rect 2823 13345 2832 13379
rect 2780 13336 2832 13345
rect 32312 13268 32364 13320
rect 33140 13311 33192 13320
rect 33140 13277 33149 13311
rect 33149 13277 33183 13311
rect 33183 13277 33192 13311
rect 33140 13268 33192 13277
rect 33416 13268 33468 13320
rect 32496 13132 32548 13184
rect 12214 13030 12266 13082
rect 12278 13030 12330 13082
rect 12342 13030 12394 13082
rect 12406 13030 12458 13082
rect 12470 13030 12522 13082
rect 23478 13030 23530 13082
rect 23542 13030 23594 13082
rect 23606 13030 23658 13082
rect 23670 13030 23722 13082
rect 23734 13030 23786 13082
rect 32496 12903 32548 12912
rect 32496 12869 32505 12903
rect 32505 12869 32539 12903
rect 32539 12869 32548 12903
rect 32496 12860 32548 12869
rect 34152 12903 34204 12912
rect 34152 12869 34161 12903
rect 34161 12869 34195 12903
rect 34195 12869 34204 12903
rect 34152 12860 34204 12869
rect 32312 12835 32364 12844
rect 32312 12801 32321 12835
rect 32321 12801 32355 12835
rect 32355 12801 32364 12835
rect 32312 12792 32364 12801
rect 1584 12588 1636 12640
rect 6582 12486 6634 12538
rect 6646 12486 6698 12538
rect 6710 12486 6762 12538
rect 6774 12486 6826 12538
rect 6838 12486 6890 12538
rect 17846 12486 17898 12538
rect 17910 12486 17962 12538
rect 17974 12486 18026 12538
rect 18038 12486 18090 12538
rect 18102 12486 18154 12538
rect 29110 12486 29162 12538
rect 29174 12486 29226 12538
rect 29238 12486 29290 12538
rect 29302 12486 29354 12538
rect 29366 12486 29418 12538
rect 33140 12248 33192 12300
rect 34152 12291 34204 12300
rect 34152 12257 34161 12291
rect 34161 12257 34195 12291
rect 34195 12257 34204 12291
rect 34152 12248 34204 12257
rect 2228 12180 2280 12232
rect 14372 12180 14424 12232
rect 20904 12180 20956 12232
rect 33692 12112 33744 12164
rect 1768 12044 1820 12096
rect 12214 11942 12266 11994
rect 12278 11942 12330 11994
rect 12342 11942 12394 11994
rect 12406 11942 12458 11994
rect 12470 11942 12522 11994
rect 23478 11942 23530 11994
rect 23542 11942 23594 11994
rect 23606 11942 23658 11994
rect 23670 11942 23722 11994
rect 23734 11942 23786 11994
rect 1768 11815 1820 11824
rect 1768 11781 1777 11815
rect 1777 11781 1811 11815
rect 1811 11781 1820 11815
rect 1768 11772 1820 11781
rect 32772 11772 32824 11824
rect 1584 11747 1636 11756
rect 1584 11713 1593 11747
rect 1593 11713 1627 11747
rect 1627 11713 1636 11747
rect 1584 11704 1636 11713
rect 2780 11679 2832 11688
rect 2780 11645 2789 11679
rect 2789 11645 2823 11679
rect 2823 11645 2832 11679
rect 2780 11636 2832 11645
rect 32680 11636 32732 11688
rect 33968 11568 34020 11620
rect 6582 11398 6634 11450
rect 6646 11398 6698 11450
rect 6710 11398 6762 11450
rect 6774 11398 6826 11450
rect 6838 11398 6890 11450
rect 17846 11398 17898 11450
rect 17910 11398 17962 11450
rect 17974 11398 18026 11450
rect 18038 11398 18090 11450
rect 18102 11398 18154 11450
rect 29110 11398 29162 11450
rect 29174 11398 29226 11450
rect 29238 11398 29290 11450
rect 29302 11398 29354 11450
rect 29366 11398 29418 11450
rect 33692 11339 33744 11348
rect 33692 11305 33701 11339
rect 33701 11305 33735 11339
rect 33735 11305 33744 11339
rect 33692 11296 33744 11305
rect 1860 11203 1912 11212
rect 1860 11169 1869 11203
rect 1869 11169 1903 11203
rect 1903 11169 1912 11203
rect 1860 11160 1912 11169
rect 1400 11135 1452 11144
rect 1400 11101 1409 11135
rect 1409 11101 1443 11135
rect 1443 11101 1452 11135
rect 1400 11092 1452 11101
rect 33600 11135 33652 11144
rect 33600 11101 33609 11135
rect 33609 11101 33643 11135
rect 33643 11101 33652 11135
rect 33600 11092 33652 11101
rect 1584 11067 1636 11076
rect 1584 11033 1593 11067
rect 1593 11033 1627 11067
rect 1627 11033 1636 11067
rect 1584 11024 1636 11033
rect 12214 10854 12266 10906
rect 12278 10854 12330 10906
rect 12342 10854 12394 10906
rect 12406 10854 12458 10906
rect 12470 10854 12522 10906
rect 23478 10854 23530 10906
rect 23542 10854 23594 10906
rect 23606 10854 23658 10906
rect 23670 10854 23722 10906
rect 23734 10854 23786 10906
rect 1584 10752 1636 10804
rect 2136 10616 2188 10668
rect 33968 10659 34020 10668
rect 33968 10625 33977 10659
rect 33977 10625 34011 10659
rect 34011 10625 34020 10659
rect 33968 10616 34020 10625
rect 1400 10548 1452 10600
rect 6582 10310 6634 10362
rect 6646 10310 6698 10362
rect 6710 10310 6762 10362
rect 6774 10310 6826 10362
rect 6838 10310 6890 10362
rect 17846 10310 17898 10362
rect 17910 10310 17962 10362
rect 17974 10310 18026 10362
rect 18038 10310 18090 10362
rect 18102 10310 18154 10362
rect 29110 10310 29162 10362
rect 29174 10310 29226 10362
rect 29238 10310 29290 10362
rect 29302 10310 29354 10362
rect 29366 10310 29418 10362
rect 31576 10208 31628 10260
rect 1768 10047 1820 10056
rect 1768 10013 1777 10047
rect 1777 10013 1811 10047
rect 1811 10013 1820 10047
rect 1768 10004 1820 10013
rect 2596 10047 2648 10056
rect 2596 10013 2605 10047
rect 2605 10013 2639 10047
rect 2639 10013 2648 10047
rect 2596 10004 2648 10013
rect 32128 10004 32180 10056
rect 33968 9979 34020 9988
rect 33968 9945 33977 9979
rect 33977 9945 34011 9979
rect 34011 9945 34020 9979
rect 33968 9936 34020 9945
rect 1676 9868 1728 9920
rect 33324 9911 33376 9920
rect 33324 9877 33333 9911
rect 33333 9877 33367 9911
rect 33367 9877 33376 9911
rect 33324 9868 33376 9877
rect 12214 9766 12266 9818
rect 12278 9766 12330 9818
rect 12342 9766 12394 9818
rect 12406 9766 12458 9818
rect 12470 9766 12522 9818
rect 23478 9766 23530 9818
rect 23542 9766 23594 9818
rect 23606 9766 23658 9818
rect 23670 9766 23722 9818
rect 23734 9766 23786 9818
rect 1676 9639 1728 9648
rect 1676 9605 1685 9639
rect 1685 9605 1719 9639
rect 1719 9605 1728 9639
rect 1676 9596 1728 9605
rect 33324 9596 33376 9648
rect 2596 9460 2648 9512
rect 2872 9503 2924 9512
rect 2872 9469 2881 9503
rect 2881 9469 2915 9503
rect 2915 9469 2924 9503
rect 2872 9460 2924 9469
rect 33968 9460 34020 9512
rect 34152 9503 34204 9512
rect 34152 9469 34161 9503
rect 34161 9469 34195 9503
rect 34195 9469 34204 9503
rect 34152 9460 34204 9469
rect 6582 9222 6634 9274
rect 6646 9222 6698 9274
rect 6710 9222 6762 9274
rect 6774 9222 6826 9274
rect 6838 9222 6890 9274
rect 17846 9222 17898 9274
rect 17910 9222 17962 9274
rect 17974 9222 18026 9274
rect 18038 9222 18090 9274
rect 18102 9222 18154 9274
rect 29110 9222 29162 9274
rect 29174 9222 29226 9274
rect 29238 9222 29290 9274
rect 29302 9222 29354 9274
rect 29366 9222 29418 9274
rect 33968 9163 34020 9172
rect 33968 9129 33977 9163
rect 33977 9129 34011 9163
rect 34011 9129 34020 9163
rect 33968 9120 34020 9129
rect 2780 9027 2832 9036
rect 2780 8993 2789 9027
rect 2789 8993 2823 9027
rect 2823 8993 2832 9027
rect 2780 8984 2832 8993
rect 1400 8959 1452 8968
rect 1400 8925 1409 8959
rect 1409 8925 1443 8959
rect 1443 8925 1452 8959
rect 1400 8916 1452 8925
rect 1952 8848 2004 8900
rect 12214 8678 12266 8730
rect 12278 8678 12330 8730
rect 12342 8678 12394 8730
rect 12406 8678 12458 8730
rect 12470 8678 12522 8730
rect 23478 8678 23530 8730
rect 23542 8678 23594 8730
rect 23606 8678 23658 8730
rect 23670 8678 23722 8730
rect 23734 8678 23786 8730
rect 1952 8619 2004 8628
rect 1952 8585 1961 8619
rect 1961 8585 1995 8619
rect 1995 8585 2004 8619
rect 1952 8576 2004 8585
rect 1400 8508 1452 8560
rect 2320 8440 2372 8492
rect 6582 8134 6634 8186
rect 6646 8134 6698 8186
rect 6710 8134 6762 8186
rect 6774 8134 6826 8186
rect 6838 8134 6890 8186
rect 17846 8134 17898 8186
rect 17910 8134 17962 8186
rect 17974 8134 18026 8186
rect 18038 8134 18090 8186
rect 18102 8134 18154 8186
rect 29110 8134 29162 8186
rect 29174 8134 29226 8186
rect 29238 8134 29290 8186
rect 29302 8134 29354 8186
rect 29366 8134 29418 8186
rect 2044 8075 2096 8084
rect 2044 8041 2053 8075
rect 2053 8041 2087 8075
rect 2087 8041 2096 8075
rect 2044 8032 2096 8041
rect 1952 7871 2004 7880
rect 1952 7837 1961 7871
rect 1961 7837 1995 7871
rect 1995 7837 2004 7871
rect 1952 7828 2004 7837
rect 1584 7760 1636 7812
rect 32588 7828 32640 7880
rect 12214 7590 12266 7642
rect 12278 7590 12330 7642
rect 12342 7590 12394 7642
rect 12406 7590 12458 7642
rect 12470 7590 12522 7642
rect 23478 7590 23530 7642
rect 23542 7590 23594 7642
rect 23606 7590 23658 7642
rect 23670 7590 23722 7642
rect 23734 7590 23786 7642
rect 1584 7395 1636 7404
rect 1584 7361 1593 7395
rect 1593 7361 1627 7395
rect 1627 7361 1636 7395
rect 1584 7352 1636 7361
rect 1768 7327 1820 7336
rect 1768 7293 1777 7327
rect 1777 7293 1811 7327
rect 1811 7293 1820 7327
rect 1768 7284 1820 7293
rect 2780 7327 2832 7336
rect 2780 7293 2789 7327
rect 2789 7293 2823 7327
rect 2823 7293 2832 7327
rect 2780 7284 2832 7293
rect 3884 7148 3936 7200
rect 29736 7148 29788 7200
rect 33968 7191 34020 7200
rect 33968 7157 33977 7191
rect 33977 7157 34011 7191
rect 34011 7157 34020 7191
rect 33968 7148 34020 7157
rect 6582 7046 6634 7098
rect 6646 7046 6698 7098
rect 6710 7046 6762 7098
rect 6774 7046 6826 7098
rect 6838 7046 6890 7098
rect 17846 7046 17898 7098
rect 17910 7046 17962 7098
rect 17974 7046 18026 7098
rect 18038 7046 18090 7098
rect 18102 7046 18154 7098
rect 29110 7046 29162 7098
rect 29174 7046 29226 7098
rect 29238 7046 29290 7098
rect 29302 7046 29354 7098
rect 29366 7046 29418 7098
rect 1768 6944 1820 6996
rect 33968 6808 34020 6860
rect 34152 6851 34204 6860
rect 34152 6817 34161 6851
rect 34161 6817 34195 6851
rect 34195 6817 34204 6851
rect 34152 6808 34204 6817
rect 1952 6783 2004 6792
rect 1952 6749 1961 6783
rect 1961 6749 1995 6783
rect 1995 6749 2004 6783
rect 1952 6740 2004 6749
rect 3148 6740 3200 6792
rect 3792 6783 3844 6792
rect 3792 6749 3801 6783
rect 3801 6749 3835 6783
rect 3835 6749 3844 6783
rect 3792 6740 3844 6749
rect 31668 6740 31720 6792
rect 33692 6672 33744 6724
rect 3976 6604 4028 6656
rect 12214 6502 12266 6554
rect 12278 6502 12330 6554
rect 12342 6502 12394 6554
rect 12406 6502 12458 6554
rect 12470 6502 12522 6554
rect 23478 6502 23530 6554
rect 23542 6502 23594 6554
rect 23606 6502 23658 6554
rect 23670 6502 23722 6554
rect 23734 6502 23786 6554
rect 33692 6443 33744 6452
rect 33692 6409 33701 6443
rect 33701 6409 33735 6443
rect 33735 6409 33744 6443
rect 33692 6400 33744 6409
rect 32956 6307 33008 6316
rect 32956 6273 32965 6307
rect 32965 6273 32999 6307
rect 32999 6273 33008 6307
rect 32956 6264 33008 6273
rect 33416 6264 33468 6316
rect 2872 6196 2924 6248
rect 3240 6239 3292 6248
rect 3240 6205 3249 6239
rect 3249 6205 3283 6239
rect 3283 6205 3292 6239
rect 3240 6196 3292 6205
rect 6460 6128 6512 6180
rect 1400 6060 1452 6112
rect 4528 6103 4580 6112
rect 4528 6069 4537 6103
rect 4537 6069 4571 6103
rect 4571 6069 4580 6103
rect 4528 6060 4580 6069
rect 5172 6103 5224 6112
rect 5172 6069 5181 6103
rect 5181 6069 5215 6103
rect 5215 6069 5224 6103
rect 5172 6060 5224 6069
rect 30472 6060 30524 6112
rect 32496 6103 32548 6112
rect 32496 6069 32505 6103
rect 32505 6069 32539 6103
rect 32539 6069 32548 6103
rect 32496 6060 32548 6069
rect 33048 6103 33100 6112
rect 33048 6069 33057 6103
rect 33057 6069 33091 6103
rect 33091 6069 33100 6103
rect 33048 6060 33100 6069
rect 6582 5958 6634 6010
rect 6646 5958 6698 6010
rect 6710 5958 6762 6010
rect 6774 5958 6826 6010
rect 6838 5958 6890 6010
rect 17846 5958 17898 6010
rect 17910 5958 17962 6010
rect 17974 5958 18026 6010
rect 18038 5958 18090 6010
rect 18102 5958 18154 6010
rect 29110 5958 29162 6010
rect 29174 5958 29226 6010
rect 29238 5958 29290 6010
rect 29302 5958 29354 6010
rect 29366 5958 29418 6010
rect 32312 5856 32364 5908
rect 4528 5788 4580 5840
rect 24032 5788 24084 5840
rect 1860 5763 1912 5772
rect 1860 5729 1869 5763
rect 1869 5729 1903 5763
rect 1903 5729 1912 5763
rect 1860 5720 1912 5729
rect 3792 5763 3844 5772
rect 3792 5729 3801 5763
rect 3801 5729 3835 5763
rect 3835 5729 3844 5763
rect 3792 5720 3844 5729
rect 3976 5763 4028 5772
rect 3976 5729 3985 5763
rect 3985 5729 4019 5763
rect 4019 5729 4028 5763
rect 3976 5720 4028 5729
rect 4160 5720 4212 5772
rect 31668 5763 31720 5772
rect 31668 5729 31677 5763
rect 31677 5729 31711 5763
rect 31711 5729 31720 5763
rect 31668 5720 31720 5729
rect 33140 5763 33192 5772
rect 33140 5729 33149 5763
rect 33149 5729 33183 5763
rect 33183 5729 33192 5763
rect 33140 5720 33192 5729
rect 6276 5695 6328 5704
rect 6276 5661 6285 5695
rect 6285 5661 6319 5695
rect 6319 5661 6328 5695
rect 6276 5652 6328 5661
rect 31484 5652 31536 5704
rect 1584 5627 1636 5636
rect 1584 5593 1593 5627
rect 1593 5593 1627 5627
rect 1627 5593 1636 5627
rect 1584 5584 1636 5593
rect 31852 5627 31904 5636
rect 31852 5593 31861 5627
rect 31861 5593 31895 5627
rect 31895 5593 31904 5627
rect 31852 5584 31904 5593
rect 34060 5559 34112 5568
rect 34060 5525 34069 5559
rect 34069 5525 34103 5559
rect 34103 5525 34112 5559
rect 34060 5516 34112 5525
rect 12214 5414 12266 5466
rect 12278 5414 12330 5466
rect 12342 5414 12394 5466
rect 12406 5414 12458 5466
rect 12470 5414 12522 5466
rect 23478 5414 23530 5466
rect 23542 5414 23594 5466
rect 23606 5414 23658 5466
rect 23670 5414 23722 5466
rect 23734 5414 23786 5466
rect 1584 5312 1636 5364
rect 4712 5312 4764 5364
rect 32956 5312 33008 5364
rect 1676 5176 1728 5228
rect 5172 5244 5224 5296
rect 6460 5176 6512 5228
rect 27620 5176 27672 5228
rect 29644 5176 29696 5228
rect 29828 5176 29880 5228
rect 2780 5151 2832 5160
rect 2780 5117 2789 5151
rect 2789 5117 2823 5151
rect 2823 5117 2832 5151
rect 2780 5108 2832 5117
rect 3056 5151 3108 5160
rect 3056 5117 3065 5151
rect 3065 5117 3099 5151
rect 3099 5117 3108 5151
rect 3056 5108 3108 5117
rect 31392 5219 31444 5228
rect 31392 5185 31401 5219
rect 31401 5185 31435 5219
rect 31435 5185 31444 5219
rect 31392 5176 31444 5185
rect 32220 5108 32272 5160
rect 32588 5108 32640 5160
rect 34152 5151 34204 5160
rect 34152 5117 34161 5151
rect 34161 5117 34195 5151
rect 34195 5117 34204 5151
rect 34152 5108 34204 5117
rect 30380 5040 30432 5092
rect 31392 5040 31444 5092
rect 33876 5040 33928 5092
rect 4436 4972 4488 5024
rect 5172 4972 5224 5024
rect 29552 5015 29604 5024
rect 29552 4981 29561 5015
rect 29561 4981 29595 5015
rect 29595 4981 29604 5015
rect 29552 4972 29604 4981
rect 29828 4972 29880 5024
rect 30840 5015 30892 5024
rect 30840 4981 30849 5015
rect 30849 4981 30883 5015
rect 30883 4981 30892 5015
rect 30840 4972 30892 4981
rect 6582 4870 6634 4922
rect 6646 4870 6698 4922
rect 6710 4870 6762 4922
rect 6774 4870 6826 4922
rect 6838 4870 6890 4922
rect 17846 4870 17898 4922
rect 17910 4870 17962 4922
rect 17974 4870 18026 4922
rect 18038 4870 18090 4922
rect 18102 4870 18154 4922
rect 29110 4870 29162 4922
rect 29174 4870 29226 4922
rect 29238 4870 29290 4922
rect 29302 4870 29354 4922
rect 29366 4870 29418 4922
rect 2780 4768 2832 4820
rect 2964 4700 3016 4752
rect 2872 4632 2924 4684
rect 4896 4632 4948 4684
rect 5172 4675 5224 4684
rect 5172 4641 5181 4675
rect 5181 4641 5215 4675
rect 5215 4641 5224 4675
rect 5172 4632 5224 4641
rect 29552 4700 29604 4752
rect 29828 4675 29880 4684
rect 29828 4641 29837 4675
rect 29837 4641 29871 4675
rect 29871 4641 29880 4675
rect 29828 4632 29880 4641
rect 30932 4675 30984 4684
rect 30932 4641 30941 4675
rect 30941 4641 30975 4675
rect 30975 4641 30984 4675
rect 30932 4632 30984 4641
rect 32312 4675 32364 4684
rect 32312 4641 32321 4675
rect 32321 4641 32355 4675
rect 32355 4641 32364 4675
rect 32312 4632 32364 4641
rect 33048 4632 33100 4684
rect 2780 4496 2832 4548
rect 4252 4564 4304 4616
rect 7748 4564 7800 4616
rect 9864 4607 9916 4616
rect 9864 4573 9873 4607
rect 9873 4573 9907 4607
rect 9907 4573 9916 4607
rect 9864 4564 9916 4573
rect 10508 4607 10560 4616
rect 10508 4573 10517 4607
rect 10517 4573 10551 4607
rect 10551 4573 10560 4607
rect 10508 4564 10560 4573
rect 4712 4496 4764 4548
rect 5356 4539 5408 4548
rect 5356 4505 5365 4539
rect 5365 4505 5399 4539
rect 5399 4505 5408 4539
rect 5356 4496 5408 4505
rect 34152 4539 34204 4548
rect 34152 4505 34161 4539
rect 34161 4505 34195 4539
rect 34195 4505 34204 4539
rect 34152 4496 34204 4505
rect 1584 4428 1636 4480
rect 6368 4428 6420 4480
rect 12214 4326 12266 4378
rect 12278 4326 12330 4378
rect 12342 4326 12394 4378
rect 12406 4326 12458 4378
rect 12470 4326 12522 4378
rect 23478 4326 23530 4378
rect 23542 4326 23594 4378
rect 23606 4326 23658 4378
rect 23670 4326 23722 4378
rect 23734 4326 23786 4378
rect 2504 4156 2556 4208
rect 2872 4063 2924 4072
rect 2872 4029 2881 4063
rect 2881 4029 2915 4063
rect 2915 4029 2924 4063
rect 2872 4020 2924 4029
rect 4252 4156 4304 4208
rect 7748 4131 7800 4140
rect 7748 4097 7757 4131
rect 7757 4097 7791 4131
rect 7791 4097 7800 4131
rect 7748 4088 7800 4097
rect 13820 4088 13872 4140
rect 21824 4088 21876 4140
rect 29736 4131 29788 4140
rect 4344 4020 4396 4072
rect 8024 4020 8076 4072
rect 8392 4063 8444 4072
rect 8392 4029 8401 4063
rect 8401 4029 8435 4063
rect 8435 4029 8444 4063
rect 8392 4020 8444 4029
rect 27712 4020 27764 4072
rect 28908 4020 28960 4072
rect 29736 4097 29745 4131
rect 29745 4097 29779 4131
rect 29779 4097 29788 4131
rect 29736 4088 29788 4097
rect 31484 4088 31536 4140
rect 30748 4020 30800 4072
rect 32036 4020 32088 4072
rect 32312 4063 32364 4072
rect 32312 4029 32321 4063
rect 32321 4029 32355 4063
rect 32355 4029 32364 4063
rect 32312 4020 32364 4029
rect 33048 4063 33100 4072
rect 33048 4029 33057 4063
rect 33057 4029 33091 4063
rect 33091 4029 33100 4063
rect 33048 4020 33100 4029
rect 5356 3952 5408 4004
rect 28356 3952 28408 4004
rect 30380 3952 30432 4004
rect 3148 3884 3200 3936
rect 4620 3884 4672 3936
rect 5540 3927 5592 3936
rect 5540 3893 5549 3927
rect 5549 3893 5583 3927
rect 5583 3893 5592 3927
rect 5540 3884 5592 3893
rect 6920 3884 6972 3936
rect 9772 3884 9824 3936
rect 14280 3884 14332 3936
rect 15476 3884 15528 3936
rect 19432 3884 19484 3936
rect 20812 3884 20864 3936
rect 29644 3884 29696 3936
rect 6582 3782 6634 3834
rect 6646 3782 6698 3834
rect 6710 3782 6762 3834
rect 6774 3782 6826 3834
rect 6838 3782 6890 3834
rect 17846 3782 17898 3834
rect 17910 3782 17962 3834
rect 17974 3782 18026 3834
rect 18038 3782 18090 3834
rect 18102 3782 18154 3834
rect 29110 3782 29162 3834
rect 29174 3782 29226 3834
rect 29238 3782 29290 3834
rect 29302 3782 29354 3834
rect 29366 3782 29418 3834
rect 4252 3680 4304 3732
rect 7840 3680 7892 3732
rect 8024 3723 8076 3732
rect 8024 3689 8033 3723
rect 8033 3689 8067 3723
rect 8067 3689 8076 3723
rect 8024 3680 8076 3689
rect 664 3612 716 3664
rect 1400 3587 1452 3596
rect 1400 3553 1409 3587
rect 1409 3553 1443 3587
rect 1443 3553 1452 3587
rect 1400 3544 1452 3553
rect 1584 3587 1636 3596
rect 1584 3553 1593 3587
rect 1593 3553 1627 3587
rect 1627 3553 1636 3587
rect 1584 3544 1636 3553
rect 4436 3587 4488 3596
rect 4436 3553 4445 3587
rect 4445 3553 4479 3587
rect 4479 3553 4488 3587
rect 4436 3544 4488 3553
rect 4620 3587 4672 3596
rect 4620 3553 4629 3587
rect 4629 3553 4663 3587
rect 4663 3553 4672 3587
rect 4620 3544 4672 3553
rect 5172 3587 5224 3596
rect 5172 3553 5181 3587
rect 5181 3553 5215 3587
rect 5215 3553 5224 3587
rect 5172 3544 5224 3553
rect 5264 3544 5316 3596
rect 2780 3476 2832 3528
rect 7932 3519 7984 3528
rect 7932 3485 7941 3519
rect 7941 3485 7975 3519
rect 7975 3485 7984 3519
rect 28356 3680 28408 3732
rect 32312 3680 32364 3732
rect 10508 3612 10560 3664
rect 9772 3587 9824 3596
rect 9772 3553 9781 3587
rect 9781 3553 9815 3587
rect 9815 3553 9824 3587
rect 9772 3544 9824 3553
rect 9956 3544 10008 3596
rect 8944 3519 8996 3528
rect 7932 3476 7984 3485
rect 8944 3485 8953 3519
rect 8953 3485 8987 3519
rect 8987 3485 8996 3519
rect 8944 3476 8996 3485
rect 10968 3476 11020 3528
rect 2504 3340 2556 3392
rect 9312 3340 9364 3392
rect 11980 3408 12032 3460
rect 15476 3587 15528 3596
rect 15476 3553 15485 3587
rect 15485 3553 15519 3587
rect 15519 3553 15528 3587
rect 15476 3544 15528 3553
rect 16120 3587 16172 3596
rect 16120 3553 16129 3587
rect 16129 3553 16163 3587
rect 16163 3553 16172 3587
rect 16120 3544 16172 3553
rect 20812 3587 20864 3596
rect 20812 3553 20821 3587
rect 20821 3553 20855 3587
rect 20855 3553 20864 3587
rect 20812 3544 20864 3553
rect 14372 3476 14424 3528
rect 16856 3476 16908 3528
rect 18420 3476 18472 3528
rect 19248 3476 19300 3528
rect 20352 3519 20404 3528
rect 20352 3485 20361 3519
rect 20361 3485 20395 3519
rect 20395 3485 20404 3519
rect 20352 3476 20404 3485
rect 15660 3451 15712 3460
rect 15660 3417 15669 3451
rect 15669 3417 15703 3451
rect 15703 3417 15712 3451
rect 15660 3408 15712 3417
rect 21916 3408 21968 3460
rect 14464 3340 14516 3392
rect 19616 3340 19668 3392
rect 21272 3340 21324 3392
rect 23848 3476 23900 3528
rect 30196 3612 30248 3664
rect 35440 3544 35492 3596
rect 27896 3476 27948 3528
rect 29460 3476 29512 3528
rect 32220 3476 32272 3528
rect 29000 3408 29052 3460
rect 30656 3451 30708 3460
rect 30656 3417 30665 3451
rect 30665 3417 30699 3451
rect 30699 3417 30708 3451
rect 30656 3408 30708 3417
rect 33784 3451 33836 3460
rect 33784 3417 33793 3451
rect 33793 3417 33827 3451
rect 33827 3417 33836 3451
rect 33784 3408 33836 3417
rect 12214 3238 12266 3290
rect 12278 3238 12330 3290
rect 12342 3238 12394 3290
rect 12406 3238 12458 3290
rect 12470 3238 12522 3290
rect 23478 3238 23530 3290
rect 23542 3238 23594 3290
rect 23606 3238 23658 3290
rect 23670 3238 23722 3290
rect 23734 3238 23786 3290
rect 5540 3136 5592 3188
rect 2504 3111 2556 3120
rect 2504 3077 2513 3111
rect 2513 3077 2547 3111
rect 2547 3077 2556 3111
rect 2504 3068 2556 3077
rect 2596 3068 2648 3120
rect 15752 3136 15804 3188
rect 21916 3179 21968 3188
rect 2596 2932 2648 2984
rect 4252 2932 4304 2984
rect 6276 3000 6328 3052
rect 9864 3068 9916 3120
rect 14464 3111 14516 3120
rect 14464 3077 14473 3111
rect 14473 3077 14507 3111
rect 14507 3077 14516 3111
rect 14464 3068 14516 3077
rect 11980 3043 12032 3052
rect 11980 3009 11989 3043
rect 11989 3009 12023 3043
rect 12023 3009 12032 3043
rect 11980 3000 12032 3009
rect 14280 3043 14332 3052
rect 14280 3009 14289 3043
rect 14289 3009 14323 3043
rect 14323 3009 14332 3043
rect 14280 3000 14332 3009
rect 16856 3043 16908 3052
rect 16856 3009 16865 3043
rect 16865 3009 16899 3043
rect 16899 3009 16908 3043
rect 16856 3000 16908 3009
rect 20352 3068 20404 3120
rect 21916 3145 21925 3179
rect 21925 3145 21959 3179
rect 21959 3145 21968 3179
rect 21916 3136 21968 3145
rect 29000 3136 29052 3188
rect 30656 3136 30708 3188
rect 21824 3043 21876 3052
rect 21824 3009 21833 3043
rect 21833 3009 21867 3043
rect 21867 3009 21876 3043
rect 21824 3000 21876 3009
rect 23848 3043 23900 3052
rect 1584 2796 1636 2848
rect 1952 2796 2004 2848
rect 9680 2975 9732 2984
rect 6460 2864 6512 2916
rect 9680 2941 9689 2975
rect 9689 2941 9723 2975
rect 9723 2941 9732 2975
rect 9680 2932 9732 2941
rect 13176 2932 13228 2984
rect 13544 2975 13596 2984
rect 13544 2941 13553 2975
rect 13553 2941 13587 2975
rect 13587 2941 13596 2975
rect 13544 2932 13596 2941
rect 14832 2975 14884 2984
rect 14832 2941 14841 2975
rect 14841 2941 14875 2975
rect 14875 2941 14884 2975
rect 14832 2932 14884 2941
rect 17040 2975 17092 2984
rect 17040 2941 17049 2975
rect 17049 2941 17083 2975
rect 17083 2941 17092 2975
rect 17040 2932 17092 2941
rect 17408 2975 17460 2984
rect 17408 2941 17417 2975
rect 17417 2941 17451 2975
rect 17451 2941 17460 2975
rect 17408 2932 17460 2941
rect 20628 2975 20680 2984
rect 10876 2864 10928 2916
rect 20628 2941 20637 2975
rect 20637 2941 20671 2975
rect 20671 2941 20680 2975
rect 20628 2932 20680 2941
rect 21916 2864 21968 2916
rect 23848 3009 23857 3043
rect 23857 3009 23891 3043
rect 23891 3009 23900 3043
rect 23848 3000 23900 3009
rect 24492 2975 24544 2984
rect 24492 2941 24501 2975
rect 24501 2941 24535 2975
rect 24535 2941 24544 2975
rect 24492 2932 24544 2941
rect 27712 3043 27764 3052
rect 27712 3009 27721 3043
rect 27721 3009 27755 3043
rect 27755 3009 27764 3043
rect 27712 3000 27764 3009
rect 34060 3068 34112 3120
rect 29644 3043 29696 3052
rect 27896 2932 27948 2984
rect 29644 3009 29653 3043
rect 29653 3009 29687 3043
rect 29687 3009 29696 3043
rect 29644 3000 29696 3009
rect 30288 2975 30340 2984
rect 30288 2941 30297 2975
rect 30297 2941 30331 2975
rect 30331 2941 30340 2975
rect 30288 2932 30340 2941
rect 32496 2932 32548 2984
rect 34796 2932 34848 2984
rect 33232 2864 33284 2916
rect 4712 2839 4764 2848
rect 4712 2805 4721 2839
rect 4721 2805 4755 2839
rect 4755 2805 4764 2839
rect 4712 2796 4764 2805
rect 7840 2796 7892 2848
rect 12440 2796 12492 2848
rect 19248 2796 19300 2848
rect 27712 2796 27764 2848
rect 29920 2796 29972 2848
rect 32220 2796 32272 2848
rect 33140 2796 33192 2848
rect 6582 2694 6634 2746
rect 6646 2694 6698 2746
rect 6710 2694 6762 2746
rect 6774 2694 6826 2746
rect 6838 2694 6890 2746
rect 17846 2694 17898 2746
rect 17910 2694 17962 2746
rect 17974 2694 18026 2746
rect 18038 2694 18090 2746
rect 18102 2694 18154 2746
rect 29110 2694 29162 2746
rect 29174 2694 29226 2746
rect 29238 2694 29290 2746
rect 29302 2694 29354 2746
rect 29366 2694 29418 2746
rect 3424 2592 3476 2644
rect 9680 2592 9732 2644
rect 13176 2592 13228 2644
rect 15660 2592 15712 2644
rect 17040 2592 17092 2644
rect 17500 2592 17552 2644
rect 21916 2635 21968 2644
rect 21916 2601 21925 2635
rect 21925 2601 21959 2635
rect 21959 2601 21968 2635
rect 21916 2592 21968 2601
rect 31852 2592 31904 2644
rect 1584 2499 1636 2508
rect 1584 2465 1593 2499
rect 1593 2465 1627 2499
rect 1627 2465 1636 2499
rect 1584 2456 1636 2465
rect 2780 2499 2832 2508
rect 2780 2465 2789 2499
rect 2789 2465 2823 2499
rect 2823 2465 2832 2499
rect 2780 2456 2832 2465
rect 4344 2524 4396 2576
rect 4528 2524 4580 2576
rect 4712 2456 4764 2508
rect 5264 2320 5316 2372
rect 3240 2252 3292 2304
rect 6920 2456 6972 2508
rect 10968 2524 11020 2576
rect 9312 2499 9364 2508
rect 9312 2465 9321 2499
rect 9321 2465 9355 2499
rect 9355 2465 9364 2499
rect 9312 2456 9364 2465
rect 10324 2499 10376 2508
rect 10324 2465 10333 2499
rect 10333 2465 10367 2499
rect 10367 2465 10376 2499
rect 10324 2456 10376 2465
rect 10876 2456 10928 2508
rect 19432 2499 19484 2508
rect 12440 2388 12492 2440
rect 14096 2431 14148 2440
rect 6368 2320 6420 2372
rect 14096 2397 14105 2431
rect 14105 2397 14139 2431
rect 14139 2397 14148 2431
rect 15752 2431 15804 2440
rect 14096 2388 14148 2397
rect 15752 2397 15761 2431
rect 15761 2397 15795 2431
rect 15795 2397 15804 2431
rect 15752 2388 15804 2397
rect 19432 2465 19441 2499
rect 19441 2465 19475 2499
rect 19475 2465 19484 2499
rect 19432 2456 19484 2465
rect 19616 2499 19668 2508
rect 19616 2465 19625 2499
rect 19625 2465 19659 2499
rect 19659 2465 19668 2499
rect 19616 2456 19668 2465
rect 19984 2499 20036 2508
rect 19984 2465 19993 2499
rect 19993 2465 20027 2499
rect 20027 2465 20036 2499
rect 19984 2456 20036 2465
rect 29552 2456 29604 2508
rect 28816 2431 28868 2440
rect 28816 2397 28825 2431
rect 28825 2397 28859 2431
rect 28859 2397 28868 2431
rect 28816 2388 28868 2397
rect 15384 2320 15436 2372
rect 18052 2320 18104 2372
rect 30472 2524 30524 2576
rect 29920 2499 29972 2508
rect 29920 2465 29929 2499
rect 29929 2465 29963 2499
rect 29963 2465 29972 2499
rect 29920 2456 29972 2465
rect 30196 2456 30248 2508
rect 32864 2456 32916 2508
rect 30840 2320 30892 2372
rect 34428 2320 34480 2372
rect 33600 2252 33652 2304
rect 12214 2150 12266 2202
rect 12278 2150 12330 2202
rect 12342 2150 12394 2202
rect 12406 2150 12458 2202
rect 12470 2150 12522 2202
rect 23478 2150 23530 2202
rect 23542 2150 23594 2202
rect 23606 2150 23658 2202
rect 23670 2150 23722 2202
rect 23734 2150 23786 2202
<< metal2 >>
rect -10 41200 102 42000
rect 634 41200 746 42000
rect 1278 41200 1390 42000
rect 1922 41200 2034 42000
rect 2566 41200 2678 42000
rect 2962 41576 3018 41585
rect 2962 41511 3018 41520
rect 676 38826 704 41200
rect 664 38820 716 38826
rect 664 38762 716 38768
rect 1320 38418 1348 41200
rect 1400 39432 1452 39438
rect 1400 39374 1452 39380
rect 1412 38865 1440 39374
rect 1676 38888 1728 38894
rect 1398 38856 1454 38865
rect 1676 38830 1728 38836
rect 1398 38791 1454 38800
rect 1308 38412 1360 38418
rect 1308 38354 1360 38360
rect 1584 38276 1636 38282
rect 1584 38218 1636 38224
rect 1596 37466 1624 38218
rect 1688 38010 1716 38830
rect 1860 38480 1912 38486
rect 1860 38422 1912 38428
rect 1676 38004 1728 38010
rect 1676 37946 1728 37952
rect 1872 37874 1900 38422
rect 1860 37868 1912 37874
rect 1860 37810 1912 37816
rect 2976 37806 3004 41511
rect 3210 41200 3322 42000
rect 4498 41200 4610 42000
rect 5142 41200 5254 42000
rect 5786 41200 5898 42000
rect 6430 41200 6542 42000
rect 7074 41200 7186 42000
rect 7718 41200 7830 42000
rect 8362 41200 8474 42000
rect 9006 41200 9118 42000
rect 9650 41200 9762 42000
rect 10938 41200 11050 42000
rect 11582 41200 11694 42000
rect 12226 41200 12338 42000
rect 12870 41200 12982 42000
rect 13514 41200 13626 42000
rect 14158 41200 14270 42000
rect 14802 41200 14914 42000
rect 15446 41200 15558 42000
rect 16090 41200 16202 42000
rect 17378 41200 17490 42000
rect 18022 41200 18134 42000
rect 18666 41200 18778 42000
rect 19310 41200 19422 42000
rect 19954 41200 20066 42000
rect 20598 41200 20710 42000
rect 21242 41200 21354 42000
rect 21886 41200 21998 42000
rect 22530 41200 22642 42000
rect 23818 41200 23930 42000
rect 24462 41200 24574 42000
rect 25106 41200 25218 42000
rect 25750 41200 25862 42000
rect 26394 41200 26506 42000
rect 27038 41200 27150 42000
rect 27682 41200 27794 42000
rect 28326 41200 28438 42000
rect 28970 41200 29082 42000
rect 30258 41200 30370 42000
rect 30902 41200 31014 42000
rect 31546 41200 31658 42000
rect 32190 41200 32302 42000
rect 32834 41200 32946 42000
rect 33478 41200 33590 42000
rect 34122 41200 34234 42000
rect 34766 41200 34878 42000
rect 35410 41200 35522 42000
rect 3252 39386 3280 41200
rect 4158 40896 4214 40905
rect 4158 40831 4214 40840
rect 3608 39432 3660 39438
rect 3252 39358 3372 39386
rect 3608 39374 3660 39380
rect 4068 39432 4120 39438
rect 4068 39374 4120 39380
rect 3148 39296 3200 39302
rect 3148 39238 3200 39244
rect 3240 39296 3292 39302
rect 3240 39238 3292 39244
rect 3160 39030 3188 39238
rect 3148 39024 3200 39030
rect 3148 38966 3200 38972
rect 3252 37942 3280 39238
rect 3240 37936 3292 37942
rect 3240 37878 3292 37884
rect 2964 37800 3016 37806
rect 2964 37742 3016 37748
rect 1584 37460 1636 37466
rect 1584 37402 1636 37408
rect 3344 37330 3372 39358
rect 3332 37324 3384 37330
rect 3332 37266 3384 37272
rect 2320 37256 2372 37262
rect 2320 37198 2372 37204
rect 2332 36378 2360 37198
rect 3056 37188 3108 37194
rect 3056 37130 3108 37136
rect 2778 36816 2834 36825
rect 2778 36751 2834 36760
rect 2688 36644 2740 36650
rect 2688 36586 2740 36592
rect 2320 36372 2372 36378
rect 2320 36314 2372 36320
rect 1398 36136 1454 36145
rect 1398 36071 1454 36080
rect 1584 36100 1636 36106
rect 1412 35698 1440 36071
rect 1584 36042 1636 36048
rect 1596 35834 1624 36042
rect 1584 35828 1636 35834
rect 1584 35770 1636 35776
rect 1400 35692 1452 35698
rect 1400 35634 1452 35640
rect 2136 35692 2188 35698
rect 2136 35634 2188 35640
rect 2148 35494 2176 35634
rect 2136 35488 2188 35494
rect 2136 35430 2188 35436
rect 1768 35284 1820 35290
rect 1768 35226 1820 35232
rect 1400 35080 1452 35086
rect 1400 35022 1452 35028
rect 1412 34610 1440 35022
rect 1400 34604 1452 34610
rect 1400 34546 1452 34552
rect 1400 33992 1452 33998
rect 1400 33934 1452 33940
rect 1412 33522 1440 33934
rect 1400 33516 1452 33522
rect 1400 33458 1452 33464
rect 1492 31816 1544 31822
rect 1492 31758 1544 31764
rect 1504 31346 1532 31758
rect 1492 31340 1544 31346
rect 1492 31282 1544 31288
rect 1780 30734 1808 35226
rect 2044 35012 2096 35018
rect 2044 34954 2096 34960
rect 1950 31376 2006 31385
rect 1950 31311 2006 31320
rect 1964 31278 1992 31311
rect 1860 31272 1912 31278
rect 1860 31214 1912 31220
rect 1952 31272 2004 31278
rect 1952 31214 2004 31220
rect 1872 30938 1900 31214
rect 1860 30932 1912 30938
rect 1860 30874 1912 30880
rect 1768 30728 1820 30734
rect 1768 30670 1820 30676
rect 1780 26234 1808 30670
rect 1688 26206 1808 26234
rect 1400 25288 1452 25294
rect 1400 25230 1452 25236
rect 1412 24818 1440 25230
rect 1584 25220 1636 25226
rect 1584 25162 1636 25168
rect 1596 24954 1624 25162
rect 1584 24948 1636 24954
rect 1584 24890 1636 24896
rect 1400 24812 1452 24818
rect 1400 24754 1452 24760
rect 1492 18760 1544 18766
rect 1492 18702 1544 18708
rect 1504 18290 1532 18702
rect 1688 18306 1716 26206
rect 1860 25356 1912 25362
rect 1860 25298 1912 25304
rect 1872 25265 1900 25298
rect 1858 25256 1914 25265
rect 1858 25191 1914 25200
rect 1768 19848 1820 19854
rect 1768 19790 1820 19796
rect 1780 19378 1808 19790
rect 1768 19372 1820 19378
rect 1768 19314 1820 19320
rect 1952 19304 2004 19310
rect 1952 19246 2004 19252
rect 1964 18970 1992 19246
rect 1952 18964 2004 18970
rect 1952 18906 2004 18912
rect 1492 18284 1544 18290
rect 1688 18278 1808 18306
rect 1492 18226 1544 18232
rect 1676 18216 1728 18222
rect 1676 18158 1728 18164
rect 1688 17882 1716 18158
rect 1676 17876 1728 17882
rect 1676 17818 1728 17824
rect 1780 17678 1808 18278
rect 1860 17740 1912 17746
rect 1860 17682 1912 17688
rect 1768 17672 1820 17678
rect 1768 17614 1820 17620
rect 1676 17128 1728 17134
rect 1676 17070 1728 17076
rect 1688 16794 1716 17070
rect 1676 16788 1728 16794
rect 1676 16730 1728 16736
rect 1676 16652 1728 16658
rect 1676 16594 1728 16600
rect 1400 15904 1452 15910
rect 1400 15846 1452 15852
rect 1412 15570 1440 15846
rect 1400 15564 1452 15570
rect 1400 15506 1452 15512
rect 1584 15428 1636 15434
rect 1584 15370 1636 15376
rect 1596 15162 1624 15370
rect 1584 15156 1636 15162
rect 1584 15098 1636 15104
rect 1400 14816 1452 14822
rect 1400 14758 1452 14764
rect 1412 14482 1440 14758
rect 1400 14476 1452 14482
rect 1400 14418 1452 14424
rect 1688 13938 1716 16594
rect 1676 13932 1728 13938
rect 1676 13874 1728 13880
rect 1584 13728 1636 13734
rect 1584 13670 1636 13676
rect 1596 13394 1624 13670
rect 1584 13388 1636 13394
rect 1584 13330 1636 13336
rect 1584 12640 1636 12646
rect 1584 12582 1636 12588
rect 1596 11762 1624 12582
rect 1780 12434 1808 17614
rect 1872 16658 1900 17682
rect 1952 17128 2004 17134
rect 1950 17096 1952 17105
rect 2004 17096 2006 17105
rect 1950 17031 2006 17040
rect 1860 16652 1912 16658
rect 1860 16594 1912 16600
rect 1952 14476 2004 14482
rect 1952 14418 2004 14424
rect 1964 14385 1992 14418
rect 1950 14376 2006 14385
rect 1860 14340 1912 14346
rect 1950 14311 2006 14320
rect 1860 14282 1912 14288
rect 1872 14074 1900 14282
rect 1860 14068 1912 14074
rect 1860 14010 1912 14016
rect 1860 13932 1912 13938
rect 1860 13874 1912 13880
rect 1688 12406 1808 12434
rect 1584 11756 1636 11762
rect 1584 11698 1636 11704
rect 1400 11144 1452 11150
rect 1400 11086 1452 11092
rect 1412 10606 1440 11086
rect 1584 11076 1636 11082
rect 1584 11018 1636 11024
rect 1596 10810 1624 11018
rect 1584 10804 1636 10810
rect 1584 10746 1636 10752
rect 1688 10690 1716 12406
rect 1768 12096 1820 12102
rect 1768 12038 1820 12044
rect 1780 11830 1808 12038
rect 1768 11824 1820 11830
rect 1768 11766 1820 11772
rect 1872 11642 1900 13874
rect 1596 10662 1716 10690
rect 1780 11614 1900 11642
rect 1400 10600 1452 10606
rect 1400 10542 1452 10548
rect 1596 9466 1624 10662
rect 1780 10062 1808 11614
rect 1860 11212 1912 11218
rect 1860 11154 1912 11160
rect 1872 10985 1900 11154
rect 1858 10976 1914 10985
rect 1858 10911 1914 10920
rect 1768 10056 1820 10062
rect 1768 9998 1820 10004
rect 1676 9920 1728 9926
rect 1676 9862 1728 9868
rect 1688 9654 1716 9862
rect 1676 9648 1728 9654
rect 1676 9590 1728 9596
rect 1596 9438 1716 9466
rect 1400 8968 1452 8974
rect 1400 8910 1452 8916
rect 1412 8566 1440 8910
rect 1400 8560 1452 8566
rect 1400 8502 1452 8508
rect 1584 7812 1636 7818
rect 1584 7754 1636 7760
rect 1596 7410 1624 7754
rect 1584 7404 1636 7410
rect 1584 7346 1636 7352
rect 1400 6112 1452 6118
rect 1400 6054 1452 6060
rect 664 3664 716 3670
rect 664 3606 716 3612
rect 676 800 704 3606
rect 1412 3602 1440 6054
rect 1584 5636 1636 5642
rect 1584 5578 1636 5584
rect 1596 5370 1624 5578
rect 1584 5364 1636 5370
rect 1584 5306 1636 5312
rect 1688 5234 1716 9438
rect 1952 8900 2004 8906
rect 1952 8842 2004 8848
rect 1964 8634 1992 8842
rect 1952 8628 2004 8634
rect 1952 8570 2004 8576
rect 2056 8090 2084 34954
rect 2148 10674 2176 35430
rect 2228 19304 2280 19310
rect 2228 19246 2280 19252
rect 2240 19145 2268 19246
rect 2226 19136 2282 19145
rect 2226 19071 2282 19080
rect 2228 15020 2280 15026
rect 2228 14962 2280 14968
rect 2240 12238 2268 14962
rect 2228 12232 2280 12238
rect 2228 12174 2280 12180
rect 2136 10668 2188 10674
rect 2136 10610 2188 10616
rect 2332 8498 2360 36314
rect 2700 36310 2728 36586
rect 2688 36304 2740 36310
rect 2688 36246 2740 36252
rect 2412 36236 2464 36242
rect 2412 36178 2464 36184
rect 2424 34474 2452 36178
rect 2412 34468 2464 34474
rect 2412 34410 2464 34416
rect 2504 34128 2556 34134
rect 2504 34070 2556 34076
rect 2516 33522 2544 34070
rect 2596 33924 2648 33930
rect 2596 33866 2648 33872
rect 2608 33658 2636 33866
rect 2596 33652 2648 33658
rect 2596 33594 2648 33600
rect 2504 33516 2556 33522
rect 2504 33458 2556 33464
rect 2320 8492 2372 8498
rect 2320 8434 2372 8440
rect 2044 8084 2096 8090
rect 2044 8026 2096 8032
rect 1952 7880 2004 7886
rect 1952 7822 2004 7828
rect 1768 7336 1820 7342
rect 1768 7278 1820 7284
rect 1780 7002 1808 7278
rect 1768 6996 1820 7002
rect 1768 6938 1820 6944
rect 1964 6798 1992 7822
rect 1952 6792 2004 6798
rect 1952 6734 2004 6740
rect 1860 5772 1912 5778
rect 1860 5714 1912 5720
rect 1872 5545 1900 5714
rect 1858 5536 1914 5545
rect 1858 5471 1914 5480
rect 1676 5228 1728 5234
rect 1676 5170 1728 5176
rect 1584 4480 1636 4486
rect 1584 4422 1636 4428
rect 1596 3602 1624 4422
rect 1400 3596 1452 3602
rect 1400 3538 1452 3544
rect 1584 3596 1636 3602
rect 1584 3538 1636 3544
rect 1964 2854 1992 6734
rect 2516 4214 2544 33458
rect 2596 17060 2648 17066
rect 2596 17002 2648 17008
rect 2608 16794 2636 17002
rect 2596 16788 2648 16794
rect 2596 16730 2648 16736
rect 2596 10056 2648 10062
rect 2596 9998 2648 10004
rect 2608 9518 2636 9998
rect 2596 9512 2648 9518
rect 2596 9454 2648 9460
rect 2700 6914 2728 36246
rect 2792 36242 2820 36751
rect 2780 36236 2832 36242
rect 2780 36178 2832 36184
rect 2778 35456 2834 35465
rect 2778 35391 2834 35400
rect 2792 35154 2820 35391
rect 2780 35148 2832 35154
rect 2780 35090 2832 35096
rect 2778 34096 2834 34105
rect 2778 34031 2780 34040
rect 2832 34031 2834 34040
rect 2780 34002 2832 34008
rect 2870 18456 2926 18465
rect 2870 18391 2926 18400
rect 2884 18222 2912 18391
rect 2872 18216 2924 18222
rect 2872 18158 2924 18164
rect 2778 15736 2834 15745
rect 2778 15671 2834 15680
rect 2792 15570 2820 15671
rect 2780 15564 2832 15570
rect 2780 15506 2832 15512
rect 3068 13938 3096 37130
rect 3516 36168 3568 36174
rect 3516 36110 3568 36116
rect 3528 35834 3556 36110
rect 3620 35986 3648 39374
rect 4080 39030 4108 39374
rect 4068 39024 4120 39030
rect 4068 38966 4120 38972
rect 4172 38826 4200 40831
rect 4436 40792 4488 40798
rect 4436 40734 4488 40740
rect 4160 38820 4212 38826
rect 4160 38762 4212 38768
rect 3974 37496 4030 37505
rect 3974 37431 4030 37440
rect 3792 37256 3844 37262
rect 3792 37198 3844 37204
rect 3804 36786 3832 37198
rect 3988 36854 4016 37431
rect 3976 36848 4028 36854
rect 3976 36790 4028 36796
rect 3792 36780 3844 36786
rect 3792 36722 3844 36728
rect 3804 36174 3832 36722
rect 3884 36712 3936 36718
rect 3884 36654 3936 36660
rect 3792 36168 3844 36174
rect 3792 36110 3844 36116
rect 3620 35958 3832 35986
rect 3516 35828 3568 35834
rect 3516 35770 3568 35776
rect 3422 32056 3478 32065
rect 3422 31991 3478 32000
rect 3436 24857 3464 31991
rect 3422 24848 3478 24857
rect 3422 24783 3478 24792
rect 3056 13932 3108 13938
rect 3056 13874 3108 13880
rect 3424 13728 3476 13734
rect 2778 13696 2834 13705
rect 3424 13670 3476 13676
rect 2778 13631 2834 13640
rect 2792 13394 2820 13631
rect 3436 13462 3464 13670
rect 3424 13456 3476 13462
rect 3424 13398 3476 13404
rect 2780 13388 2832 13394
rect 2780 13330 2832 13336
rect 2780 11688 2832 11694
rect 2778 11656 2780 11665
rect 2832 11656 2834 11665
rect 2778 11591 2834 11600
rect 2872 9512 2924 9518
rect 2872 9454 2924 9460
rect 2780 9036 2832 9042
rect 2780 8978 2832 8984
rect 2792 8265 2820 8978
rect 2884 8945 2912 9454
rect 2870 8936 2926 8945
rect 2870 8871 2926 8880
rect 2778 8256 2834 8265
rect 2778 8191 2834 8200
rect 2778 7576 2834 7585
rect 2778 7511 2834 7520
rect 2792 7342 2820 7511
rect 2780 7336 2832 7342
rect 2780 7278 2832 7284
rect 2608 6886 2728 6914
rect 2504 4208 2556 4214
rect 2504 4150 2556 4156
rect 2504 3392 2556 3398
rect 2504 3334 2556 3340
rect 2516 3126 2544 3334
rect 2608 3126 2636 6886
rect 3804 6798 3832 35958
rect 3896 35698 3924 36654
rect 4448 36174 4476 40734
rect 4988 39500 5040 39506
rect 4988 39442 5040 39448
rect 4620 39432 4672 39438
rect 4620 39374 4672 39380
rect 4632 39098 4660 39374
rect 4620 39092 4672 39098
rect 4620 39034 4672 39040
rect 4804 37868 4856 37874
rect 4804 37810 4856 37816
rect 4620 37732 4672 37738
rect 4620 37674 4672 37680
rect 4436 36168 4488 36174
rect 4436 36110 4488 36116
rect 3884 35692 3936 35698
rect 3884 35634 3936 35640
rect 4448 24818 4476 36110
rect 4632 35698 4660 37674
rect 4712 37188 4764 37194
rect 4712 37130 4764 37136
rect 4724 36922 4752 37130
rect 4712 36916 4764 36922
rect 4712 36858 4764 36864
rect 4620 35692 4672 35698
rect 4620 35634 4672 35640
rect 4436 24812 4488 24818
rect 4436 24754 4488 24760
rect 3884 7200 3936 7206
rect 3884 7142 3936 7148
rect 3148 6792 3200 6798
rect 3148 6734 3200 6740
rect 3792 6792 3844 6798
rect 3792 6734 3844 6740
rect 2872 6248 2924 6254
rect 2872 6190 2924 6196
rect 2780 5160 2832 5166
rect 2780 5102 2832 5108
rect 2792 4826 2820 5102
rect 2780 4820 2832 4826
rect 2780 4762 2832 4768
rect 2884 4690 2912 6190
rect 3056 5160 3108 5166
rect 3056 5102 3108 5108
rect 3068 4865 3096 5102
rect 3054 4856 3110 4865
rect 3054 4791 3110 4800
rect 2964 4752 3016 4758
rect 2964 4694 3016 4700
rect 2872 4684 2924 4690
rect 2872 4626 2924 4632
rect 2780 4548 2832 4554
rect 2780 4490 2832 4496
rect 2792 3534 2820 4490
rect 2976 4185 3004 4694
rect 2962 4176 3018 4185
rect 2962 4111 3018 4120
rect 2872 4072 2924 4078
rect 2872 4014 2924 4020
rect 2780 3528 2832 3534
rect 2780 3470 2832 3476
rect 2504 3120 2556 3126
rect 2504 3062 2556 3068
rect 2596 3120 2648 3126
rect 2596 3062 2648 3068
rect 2596 2984 2648 2990
rect 2596 2926 2648 2932
rect 1584 2848 1636 2854
rect 1584 2790 1636 2796
rect 1952 2848 2004 2854
rect 1952 2790 2004 2796
rect 1596 2514 1624 2790
rect 1584 2508 1636 2514
rect 1584 2450 1636 2456
rect 2608 800 2636 2926
rect 2778 2816 2834 2825
rect 2778 2751 2834 2760
rect 2792 2514 2820 2751
rect 2780 2508 2832 2514
rect 2780 2450 2832 2456
rect 2884 2145 2912 4014
rect 3160 3942 3188 6734
rect 3896 6338 3924 7142
rect 3976 6656 4028 6662
rect 3976 6598 4028 6604
rect 3804 6310 3924 6338
rect 3240 6248 3292 6254
rect 3240 6190 3292 6196
rect 3148 3936 3200 3942
rect 3148 3878 3200 3884
rect 3252 3505 3280 6190
rect 3804 5778 3832 6310
rect 3988 5778 4016 6598
rect 4528 6112 4580 6118
rect 4528 6054 4580 6060
rect 4540 5846 4568 6054
rect 4528 5840 4580 5846
rect 4528 5782 4580 5788
rect 3792 5772 3844 5778
rect 3792 5714 3844 5720
rect 3976 5772 4028 5778
rect 3976 5714 4028 5720
rect 4160 5772 4212 5778
rect 4160 5714 4212 5720
rect 3238 3496 3294 3505
rect 3238 3431 3294 3440
rect 4172 2802 4200 5714
rect 4724 5370 4752 36858
rect 4816 36650 4844 37810
rect 4804 36644 4856 36650
rect 4804 36586 4856 36592
rect 4816 17746 4844 36586
rect 5000 36378 5028 39442
rect 5264 39432 5316 39438
rect 5264 39374 5316 39380
rect 5356 39432 5408 39438
rect 5356 39374 5408 39380
rect 5276 38214 5304 39374
rect 5368 38894 5396 39374
rect 5356 38888 5408 38894
rect 5356 38830 5408 38836
rect 5828 38418 5856 41200
rect 6582 39740 6890 39760
rect 6582 39738 6588 39740
rect 6644 39738 6668 39740
rect 6724 39738 6748 39740
rect 6804 39738 6828 39740
rect 6884 39738 6890 39740
rect 6644 39686 6646 39738
rect 6826 39686 6828 39738
rect 6582 39684 6588 39686
rect 6644 39684 6668 39686
rect 6724 39684 6748 39686
rect 6804 39684 6828 39686
rect 6884 39684 6890 39686
rect 6582 39664 6890 39684
rect 7012 39364 7064 39370
rect 7012 39306 7064 39312
rect 7024 38894 7052 39306
rect 7012 38888 7064 38894
rect 7012 38830 7064 38836
rect 6460 38752 6512 38758
rect 6460 38694 6512 38700
rect 6472 38418 6500 38694
rect 6582 38652 6890 38672
rect 6582 38650 6588 38652
rect 6644 38650 6668 38652
rect 6724 38650 6748 38652
rect 6804 38650 6828 38652
rect 6884 38650 6890 38652
rect 6644 38598 6646 38650
rect 6826 38598 6828 38650
rect 6582 38596 6588 38598
rect 6644 38596 6668 38598
rect 6724 38596 6748 38598
rect 6804 38596 6828 38598
rect 6884 38596 6890 38598
rect 6582 38576 6890 38596
rect 5632 38412 5684 38418
rect 5632 38354 5684 38360
rect 5816 38412 5868 38418
rect 5816 38354 5868 38360
rect 6460 38412 6512 38418
rect 6460 38354 6512 38360
rect 5356 38276 5408 38282
rect 5356 38218 5408 38224
rect 5264 38208 5316 38214
rect 5264 38150 5316 38156
rect 5368 38010 5396 38218
rect 5356 38004 5408 38010
rect 5356 37946 5408 37952
rect 5540 37868 5592 37874
rect 5540 37810 5592 37816
rect 5172 37324 5224 37330
rect 5172 37266 5224 37272
rect 5080 36848 5132 36854
rect 5080 36790 5132 36796
rect 4988 36372 5040 36378
rect 4988 36314 5040 36320
rect 4804 17740 4856 17746
rect 4804 17682 4856 17688
rect 5092 17338 5120 36790
rect 5184 36174 5212 37266
rect 5552 36854 5580 37810
rect 5540 36848 5592 36854
rect 5540 36790 5592 36796
rect 5644 36786 5672 38354
rect 6736 38276 6788 38282
rect 6736 38218 6788 38224
rect 6748 38010 6776 38218
rect 6736 38004 6788 38010
rect 6736 37946 6788 37952
rect 6582 37564 6890 37584
rect 6582 37562 6588 37564
rect 6644 37562 6668 37564
rect 6724 37562 6748 37564
rect 6804 37562 6828 37564
rect 6884 37562 6890 37564
rect 6644 37510 6646 37562
rect 6826 37510 6828 37562
rect 6582 37508 6588 37510
rect 6644 37508 6668 37510
rect 6724 37508 6748 37510
rect 6804 37508 6828 37510
rect 6884 37508 6890 37510
rect 6582 37488 6890 37508
rect 7024 37194 7052 38830
rect 7116 38418 7144 41200
rect 7196 39432 7248 39438
rect 7196 39374 7248 39380
rect 7104 38412 7156 38418
rect 7104 38354 7156 38360
rect 7208 37874 7236 39374
rect 7196 37868 7248 37874
rect 7196 37810 7248 37816
rect 7760 37806 7788 41200
rect 8300 39568 8352 39574
rect 8300 39510 8352 39516
rect 7932 39364 7984 39370
rect 7932 39306 7984 39312
rect 7944 38962 7972 39306
rect 7932 38956 7984 38962
rect 7932 38898 7984 38904
rect 7380 37800 7432 37806
rect 7380 37742 7432 37748
rect 7748 37800 7800 37806
rect 7748 37742 7800 37748
rect 7392 37466 7420 37742
rect 7380 37460 7432 37466
rect 7380 37402 7432 37408
rect 7012 37188 7064 37194
rect 7012 37130 7064 37136
rect 7944 36922 7972 38898
rect 8312 38826 8340 39510
rect 8300 38820 8352 38826
rect 8300 38762 8352 38768
rect 8404 38486 8432 41200
rect 9048 40066 9076 41200
rect 13636 40928 13688 40934
rect 13636 40870 13688 40876
rect 12072 40860 12124 40866
rect 12072 40802 12124 40808
rect 11704 40656 11756 40662
rect 11058 40624 11114 40633
rect 11704 40598 11756 40604
rect 11058 40559 11114 40568
rect 9770 40216 9826 40225
rect 9770 40151 9826 40160
rect 9048 40038 9352 40066
rect 8576 39432 8628 39438
rect 8576 39374 8628 39380
rect 8588 38962 8616 39374
rect 8576 38956 8628 38962
rect 8576 38898 8628 38904
rect 9324 38894 9352 40038
rect 9588 39568 9640 39574
rect 9586 39536 9588 39545
rect 9640 39536 9642 39545
rect 9586 39471 9642 39480
rect 9220 38888 9272 38894
rect 9220 38830 9272 38836
rect 9312 38888 9364 38894
rect 9312 38830 9364 38836
rect 9232 38758 9260 38830
rect 9128 38752 9180 38758
rect 9128 38694 9180 38700
rect 9220 38752 9272 38758
rect 9220 38694 9272 38700
rect 8392 38480 8444 38486
rect 8392 38422 8444 38428
rect 9140 38418 9168 38694
rect 9128 38412 9180 38418
rect 9128 38354 9180 38360
rect 8116 38344 8168 38350
rect 8116 38286 8168 38292
rect 8128 37466 8156 38286
rect 8116 37460 8168 37466
rect 8116 37402 8168 37408
rect 7932 36916 7984 36922
rect 7932 36858 7984 36864
rect 5632 36780 5684 36786
rect 5632 36722 5684 36728
rect 6582 36476 6890 36496
rect 6582 36474 6588 36476
rect 6644 36474 6668 36476
rect 6724 36474 6748 36476
rect 6804 36474 6828 36476
rect 6884 36474 6890 36476
rect 6644 36422 6646 36474
rect 6826 36422 6828 36474
rect 6582 36420 6588 36422
rect 6644 36420 6668 36422
rect 6724 36420 6748 36422
rect 6804 36420 6828 36422
rect 6884 36420 6890 36422
rect 6582 36400 6890 36420
rect 5172 36168 5224 36174
rect 5172 36110 5224 36116
rect 6582 35388 6890 35408
rect 6582 35386 6588 35388
rect 6644 35386 6668 35388
rect 6724 35386 6748 35388
rect 6804 35386 6828 35388
rect 6884 35386 6890 35388
rect 6644 35334 6646 35386
rect 6826 35334 6828 35386
rect 6582 35332 6588 35334
rect 6644 35332 6668 35334
rect 6724 35332 6748 35334
rect 6804 35332 6828 35334
rect 6884 35332 6890 35334
rect 6582 35312 6890 35332
rect 6582 34300 6890 34320
rect 6582 34298 6588 34300
rect 6644 34298 6668 34300
rect 6724 34298 6748 34300
rect 6804 34298 6828 34300
rect 6884 34298 6890 34300
rect 6644 34246 6646 34298
rect 6826 34246 6828 34298
rect 6582 34244 6588 34246
rect 6644 34244 6668 34246
rect 6724 34244 6748 34246
rect 6804 34244 6828 34246
rect 6884 34244 6890 34246
rect 6582 34224 6890 34244
rect 6582 33212 6890 33232
rect 6582 33210 6588 33212
rect 6644 33210 6668 33212
rect 6724 33210 6748 33212
rect 6804 33210 6828 33212
rect 6884 33210 6890 33212
rect 6644 33158 6646 33210
rect 6826 33158 6828 33210
rect 6582 33156 6588 33158
rect 6644 33156 6668 33158
rect 6724 33156 6748 33158
rect 6804 33156 6828 33158
rect 6884 33156 6890 33158
rect 6582 33136 6890 33156
rect 6582 32124 6890 32144
rect 6582 32122 6588 32124
rect 6644 32122 6668 32124
rect 6724 32122 6748 32124
rect 6804 32122 6828 32124
rect 6884 32122 6890 32124
rect 6644 32070 6646 32122
rect 6826 32070 6828 32122
rect 6582 32068 6588 32070
rect 6644 32068 6668 32070
rect 6724 32068 6748 32070
rect 6804 32068 6828 32070
rect 6884 32068 6890 32070
rect 6582 32048 6890 32068
rect 6582 31036 6890 31056
rect 6582 31034 6588 31036
rect 6644 31034 6668 31036
rect 6724 31034 6748 31036
rect 6804 31034 6828 31036
rect 6884 31034 6890 31036
rect 6644 30982 6646 31034
rect 6826 30982 6828 31034
rect 6582 30980 6588 30982
rect 6644 30980 6668 30982
rect 6724 30980 6748 30982
rect 6804 30980 6828 30982
rect 6884 30980 6890 30982
rect 6582 30960 6890 30980
rect 6582 29948 6890 29968
rect 6582 29946 6588 29948
rect 6644 29946 6668 29948
rect 6724 29946 6748 29948
rect 6804 29946 6828 29948
rect 6884 29946 6890 29948
rect 6644 29894 6646 29946
rect 6826 29894 6828 29946
rect 6582 29892 6588 29894
rect 6644 29892 6668 29894
rect 6724 29892 6748 29894
rect 6804 29892 6828 29894
rect 6884 29892 6890 29894
rect 6582 29872 6890 29892
rect 6582 28860 6890 28880
rect 6582 28858 6588 28860
rect 6644 28858 6668 28860
rect 6724 28858 6748 28860
rect 6804 28858 6828 28860
rect 6884 28858 6890 28860
rect 6644 28806 6646 28858
rect 6826 28806 6828 28858
rect 6582 28804 6588 28806
rect 6644 28804 6668 28806
rect 6724 28804 6748 28806
rect 6804 28804 6828 28806
rect 6884 28804 6890 28806
rect 6582 28784 6890 28804
rect 6582 27772 6890 27792
rect 6582 27770 6588 27772
rect 6644 27770 6668 27772
rect 6724 27770 6748 27772
rect 6804 27770 6828 27772
rect 6884 27770 6890 27772
rect 6644 27718 6646 27770
rect 6826 27718 6828 27770
rect 6582 27716 6588 27718
rect 6644 27716 6668 27718
rect 6724 27716 6748 27718
rect 6804 27716 6828 27718
rect 6884 27716 6890 27718
rect 6582 27696 6890 27716
rect 6582 26684 6890 26704
rect 6582 26682 6588 26684
rect 6644 26682 6668 26684
rect 6724 26682 6748 26684
rect 6804 26682 6828 26684
rect 6884 26682 6890 26684
rect 6644 26630 6646 26682
rect 6826 26630 6828 26682
rect 6582 26628 6588 26630
rect 6644 26628 6668 26630
rect 6724 26628 6748 26630
rect 6804 26628 6828 26630
rect 6884 26628 6890 26630
rect 6582 26608 6890 26628
rect 9232 26234 9260 38694
rect 9678 37768 9734 37777
rect 9678 37703 9680 37712
rect 9732 37703 9734 37712
rect 9680 37674 9732 37680
rect 9784 37466 9812 40151
rect 10322 39944 10378 39953
rect 10322 39879 10378 39888
rect 10336 39642 10364 39879
rect 10324 39636 10376 39642
rect 10324 39578 10376 39584
rect 10968 39432 11020 39438
rect 10966 39400 10968 39409
rect 11020 39400 11022 39409
rect 10966 39335 11022 39344
rect 10322 38992 10378 39001
rect 10322 38927 10378 38936
rect 10336 37874 10364 38927
rect 11072 38654 11100 40559
rect 10980 38626 11100 38654
rect 10874 38312 10930 38321
rect 10874 38247 10930 38256
rect 10416 37936 10468 37942
rect 10416 37878 10468 37884
rect 10782 37904 10838 37913
rect 10324 37868 10376 37874
rect 10324 37810 10376 37816
rect 9772 37460 9824 37466
rect 9772 37402 9824 37408
rect 10230 37360 10286 37369
rect 10230 37295 10232 37304
rect 10284 37295 10286 37304
rect 10232 37266 10284 37272
rect 10428 36786 10456 37878
rect 10782 37839 10838 37848
rect 10796 36786 10824 37839
rect 10888 37466 10916 38247
rect 10980 37874 11008 38626
rect 11336 38412 11388 38418
rect 11336 38354 11388 38360
rect 10968 37868 11020 37874
rect 10968 37810 11020 37816
rect 10876 37460 10928 37466
rect 10876 37402 10928 37408
rect 10876 36916 10928 36922
rect 10876 36858 10928 36864
rect 10416 36780 10468 36786
rect 10416 36722 10468 36728
rect 10784 36780 10836 36786
rect 10784 36722 10836 36728
rect 10888 36378 10916 36858
rect 10876 36372 10928 36378
rect 10876 36314 10928 36320
rect 11348 36174 11376 38354
rect 11612 38208 11664 38214
rect 11612 38150 11664 38156
rect 11624 38010 11652 38150
rect 11612 38004 11664 38010
rect 11612 37946 11664 37952
rect 11716 37754 11744 40598
rect 11796 40044 11848 40050
rect 11796 39986 11848 39992
rect 11808 38962 11836 39986
rect 11796 38956 11848 38962
rect 11796 38898 11848 38904
rect 12084 37874 12112 40802
rect 13174 40760 13230 40769
rect 13174 40695 13230 40704
rect 12992 40656 13044 40662
rect 12992 40598 13044 40604
rect 12624 40588 12676 40594
rect 12624 40530 12676 40536
rect 12256 39976 12308 39982
rect 12256 39918 12308 39924
rect 12268 39574 12296 39918
rect 12256 39568 12308 39574
rect 12256 39510 12308 39516
rect 12214 39196 12522 39216
rect 12214 39194 12220 39196
rect 12276 39194 12300 39196
rect 12356 39194 12380 39196
rect 12436 39194 12460 39196
rect 12516 39194 12522 39196
rect 12276 39142 12278 39194
rect 12458 39142 12460 39194
rect 12214 39140 12220 39142
rect 12276 39140 12300 39142
rect 12356 39140 12380 39142
rect 12436 39140 12460 39142
rect 12516 39140 12522 39142
rect 12214 39120 12522 39140
rect 12636 38962 12664 40530
rect 12716 40112 12768 40118
rect 12716 40054 12768 40060
rect 12728 39370 12756 40054
rect 12900 39840 12952 39846
rect 12900 39782 12952 39788
rect 12716 39364 12768 39370
rect 12716 39306 12768 39312
rect 12912 39098 12940 39782
rect 12900 39092 12952 39098
rect 12900 39034 12952 39040
rect 12624 38956 12676 38962
rect 12624 38898 12676 38904
rect 12254 38584 12310 38593
rect 12254 38519 12310 38528
rect 12268 38486 12296 38519
rect 12256 38480 12308 38486
rect 12256 38422 12308 38428
rect 12900 38344 12952 38350
rect 12900 38286 12952 38292
rect 12624 38208 12676 38214
rect 12912 38185 12940 38286
rect 12624 38150 12676 38156
rect 12898 38176 12954 38185
rect 12214 38108 12522 38128
rect 12214 38106 12220 38108
rect 12276 38106 12300 38108
rect 12356 38106 12380 38108
rect 12436 38106 12460 38108
rect 12516 38106 12522 38108
rect 12276 38054 12278 38106
rect 12458 38054 12460 38106
rect 12214 38052 12220 38054
rect 12276 38052 12300 38054
rect 12356 38052 12380 38054
rect 12436 38052 12460 38054
rect 12516 38052 12522 38054
rect 12214 38032 12522 38052
rect 12072 37868 12124 37874
rect 12072 37810 12124 37816
rect 12440 37868 12492 37874
rect 12440 37810 12492 37816
rect 11624 37726 11744 37754
rect 11426 37496 11482 37505
rect 11426 37431 11482 37440
rect 11440 36310 11468 37431
rect 11624 36394 11652 37726
rect 12346 37632 12402 37641
rect 12346 37567 12402 37576
rect 12360 37466 12388 37567
rect 12452 37466 12480 37810
rect 12348 37460 12400 37466
rect 12348 37402 12400 37408
rect 12440 37460 12492 37466
rect 12440 37402 12492 37408
rect 12636 37398 12664 38150
rect 12898 38111 12954 38120
rect 12716 38004 12768 38010
rect 12716 37946 12768 37952
rect 12728 37738 12756 37946
rect 12716 37732 12768 37738
rect 12716 37674 12768 37680
rect 12624 37392 12676 37398
rect 12624 37334 12676 37340
rect 12900 37324 12952 37330
rect 12900 37266 12952 37272
rect 11978 37224 12034 37233
rect 12452 37194 12756 37210
rect 11978 37159 12034 37168
rect 12440 37188 12756 37194
rect 11992 37126 12020 37159
rect 12492 37182 12756 37188
rect 12440 37130 12492 37136
rect 11980 37120 12032 37126
rect 12624 37120 12676 37126
rect 11980 37062 12032 37068
rect 12622 37088 12624 37097
rect 12676 37088 12678 37097
rect 12214 37020 12522 37040
rect 12622 37023 12678 37032
rect 12214 37018 12220 37020
rect 12276 37018 12300 37020
rect 12356 37018 12380 37020
rect 12436 37018 12460 37020
rect 12516 37018 12522 37020
rect 12276 36966 12278 37018
rect 12458 36966 12460 37018
rect 12214 36964 12220 36966
rect 12276 36964 12300 36966
rect 12356 36964 12380 36966
rect 12436 36964 12460 36966
rect 12516 36964 12522 36966
rect 12214 36944 12522 36964
rect 12440 36780 12492 36786
rect 12440 36722 12492 36728
rect 12070 36680 12126 36689
rect 12070 36615 12072 36624
rect 12124 36615 12126 36624
rect 12072 36586 12124 36592
rect 12164 36576 12216 36582
rect 12164 36518 12216 36524
rect 11624 36366 11744 36394
rect 11428 36304 11480 36310
rect 11612 36304 11664 36310
rect 11428 36246 11480 36252
rect 11610 36272 11612 36281
rect 11664 36272 11666 36281
rect 11610 36207 11666 36216
rect 11336 36168 11388 36174
rect 11336 36110 11388 36116
rect 11716 35834 11744 36366
rect 12176 36145 12204 36518
rect 12346 36408 12402 36417
rect 12346 36343 12402 36352
rect 12360 36242 12388 36343
rect 12452 36242 12480 36722
rect 12728 36582 12756 37182
rect 12806 36952 12862 36961
rect 12806 36887 12862 36896
rect 12716 36576 12768 36582
rect 12716 36518 12768 36524
rect 12348 36236 12400 36242
rect 12348 36178 12400 36184
rect 12440 36236 12492 36242
rect 12440 36178 12492 36184
rect 12820 36174 12848 36887
rect 12912 36854 12940 37266
rect 12900 36848 12952 36854
rect 12900 36790 12952 36796
rect 12900 36304 12952 36310
rect 12900 36246 12952 36252
rect 12912 36174 12940 36246
rect 12808 36168 12860 36174
rect 12162 36136 12218 36145
rect 12808 36110 12860 36116
rect 12900 36168 12952 36174
rect 12900 36110 12952 36116
rect 12162 36071 12218 36080
rect 12716 36032 12768 36038
rect 12714 36000 12716 36009
rect 12768 36000 12770 36009
rect 12214 35932 12522 35952
rect 12714 35935 12770 35944
rect 12214 35930 12220 35932
rect 12276 35930 12300 35932
rect 12356 35930 12380 35932
rect 12436 35930 12460 35932
rect 12516 35930 12522 35932
rect 12276 35878 12278 35930
rect 12458 35878 12460 35930
rect 12214 35876 12220 35878
rect 12276 35876 12300 35878
rect 12356 35876 12380 35878
rect 12436 35876 12460 35878
rect 12516 35876 12522 35878
rect 12214 35856 12522 35876
rect 11704 35828 11756 35834
rect 11704 35770 11756 35776
rect 12530 35592 12586 35601
rect 12530 35527 12532 35536
rect 12584 35527 12586 35536
rect 12532 35498 12584 35504
rect 12808 35080 12860 35086
rect 12808 35022 12860 35028
rect 12214 34844 12522 34864
rect 12214 34842 12220 34844
rect 12276 34842 12300 34844
rect 12356 34842 12380 34844
rect 12436 34842 12460 34844
rect 12516 34842 12522 34844
rect 12276 34790 12278 34842
rect 12458 34790 12460 34842
rect 12214 34788 12220 34790
rect 12276 34788 12300 34790
rect 12356 34788 12380 34790
rect 12436 34788 12460 34790
rect 12516 34788 12522 34790
rect 12214 34768 12522 34788
rect 12714 34776 12770 34785
rect 12714 34711 12716 34720
rect 12768 34711 12770 34720
rect 12716 34682 12768 34688
rect 12820 34626 12848 35022
rect 12636 34598 12848 34626
rect 13004 34610 13032 40598
rect 13082 38448 13138 38457
rect 13082 38383 13084 38392
rect 13136 38383 13138 38392
rect 13084 38354 13136 38360
rect 13084 38208 13136 38214
rect 13084 38150 13136 38156
rect 13096 38049 13124 38150
rect 13082 38040 13138 38049
rect 13082 37975 13138 37984
rect 13188 37346 13216 40695
rect 13544 40180 13596 40186
rect 13544 40122 13596 40128
rect 13556 39506 13584 40122
rect 13544 39500 13596 39506
rect 13544 39442 13596 39448
rect 13452 39432 13504 39438
rect 13648 39386 13676 40870
rect 14740 40724 14792 40730
rect 14740 40666 14792 40672
rect 14464 40384 14516 40390
rect 14278 40352 14334 40361
rect 14464 40326 14516 40332
rect 14278 40287 14334 40296
rect 14002 40080 14058 40089
rect 14002 40015 14058 40024
rect 13912 39908 13964 39914
rect 13912 39850 13964 39856
rect 13452 39374 13504 39380
rect 13464 39273 13492 39374
rect 13556 39358 13676 39386
rect 13820 39432 13872 39438
rect 13820 39374 13872 39380
rect 13450 39264 13506 39273
rect 13450 39199 13506 39208
rect 13266 39128 13322 39137
rect 13266 39063 13322 39072
rect 13452 39092 13504 39098
rect 13280 38282 13308 39063
rect 13452 39034 13504 39040
rect 13464 38729 13492 39034
rect 13450 38720 13506 38729
rect 13556 38706 13584 39358
rect 13728 39092 13780 39098
rect 13728 39034 13780 39040
rect 13740 38758 13768 39034
rect 13832 38962 13860 39374
rect 13820 38956 13872 38962
rect 13820 38898 13872 38904
rect 13728 38752 13780 38758
rect 13556 38678 13676 38706
rect 13728 38694 13780 38700
rect 13820 38752 13872 38758
rect 13820 38694 13872 38700
rect 13450 38655 13506 38664
rect 13358 38584 13414 38593
rect 13358 38519 13414 38528
rect 13268 38276 13320 38282
rect 13268 38218 13320 38224
rect 13096 37318 13216 37346
rect 13096 36689 13124 37318
rect 13176 37256 13228 37262
rect 13176 37198 13228 37204
rect 13268 37256 13320 37262
rect 13268 37198 13320 37204
rect 13082 36680 13138 36689
rect 13082 36615 13138 36624
rect 13096 34626 13124 36615
rect 13188 36553 13216 37198
rect 13174 36544 13230 36553
rect 13174 36479 13230 36488
rect 13280 35766 13308 37198
rect 13372 36038 13400 38519
rect 13452 38480 13504 38486
rect 13452 38422 13504 38428
rect 13464 36922 13492 38422
rect 13452 36916 13504 36922
rect 13452 36858 13504 36864
rect 13450 36680 13506 36689
rect 13450 36615 13506 36624
rect 13360 36032 13412 36038
rect 13360 35974 13412 35980
rect 13268 35760 13320 35766
rect 13268 35702 13320 35708
rect 13176 35692 13228 35698
rect 13176 35634 13228 35640
rect 13188 35562 13216 35634
rect 13176 35556 13228 35562
rect 13176 35498 13228 35504
rect 13280 35329 13308 35702
rect 13464 35494 13492 36615
rect 13648 36530 13676 38678
rect 13728 38208 13780 38214
rect 13728 38150 13780 38156
rect 13740 38049 13768 38150
rect 13726 38040 13782 38049
rect 13726 37975 13782 37984
rect 13832 37874 13860 38694
rect 13924 38010 13952 39850
rect 13912 38004 13964 38010
rect 13912 37946 13964 37952
rect 13820 37868 13872 37874
rect 13820 37810 13872 37816
rect 13912 37800 13964 37806
rect 13740 37748 13912 37754
rect 13740 37742 13964 37748
rect 13740 37738 13952 37742
rect 13728 37732 13952 37738
rect 13780 37726 13952 37732
rect 13728 37674 13780 37680
rect 13818 36816 13874 36825
rect 13818 36751 13874 36760
rect 13912 36780 13964 36786
rect 13556 36502 13676 36530
rect 13556 36258 13584 36502
rect 13832 36394 13860 36751
rect 13912 36722 13964 36728
rect 13648 36378 13860 36394
rect 13924 36378 13952 36722
rect 13636 36372 13860 36378
rect 13688 36366 13860 36372
rect 13912 36372 13964 36378
rect 13636 36314 13688 36320
rect 13912 36314 13964 36320
rect 13556 36230 13676 36258
rect 13544 36168 13596 36174
rect 13544 36110 13596 36116
rect 13556 36038 13584 36110
rect 13544 36032 13596 36038
rect 13544 35974 13596 35980
rect 13452 35488 13504 35494
rect 13452 35430 13504 35436
rect 13266 35320 13322 35329
rect 13266 35255 13322 35264
rect 13176 35216 13228 35222
rect 13176 35158 13228 35164
rect 13188 34921 13216 35158
rect 13556 35086 13584 35974
rect 13544 35080 13596 35086
rect 13544 35022 13596 35028
rect 13174 34912 13230 34921
rect 13648 34898 13676 36230
rect 13728 36100 13780 36106
rect 13728 36042 13780 36048
rect 13174 34847 13230 34856
rect 13556 34870 13676 34898
rect 13358 34776 13414 34785
rect 13358 34711 13360 34720
rect 13412 34711 13414 34720
rect 13360 34682 13412 34688
rect 12992 34604 13044 34610
rect 12254 34504 12310 34513
rect 12254 34439 12256 34448
rect 12308 34439 12310 34448
rect 12256 34410 12308 34416
rect 11888 34400 11940 34406
rect 11888 34342 11940 34348
rect 11796 32360 11848 32366
rect 11794 32328 11796 32337
rect 11848 32328 11850 32337
rect 11794 32263 11850 32272
rect 11796 30252 11848 30258
rect 11796 30194 11848 30200
rect 11808 29782 11836 30194
rect 11796 29776 11848 29782
rect 11796 29718 11848 29724
rect 11900 29646 11928 34342
rect 12214 33756 12522 33776
rect 12214 33754 12220 33756
rect 12276 33754 12300 33756
rect 12356 33754 12380 33756
rect 12436 33754 12460 33756
rect 12516 33754 12522 33756
rect 12276 33702 12278 33754
rect 12458 33702 12460 33754
rect 12214 33700 12220 33702
rect 12276 33700 12300 33702
rect 12356 33700 12380 33702
rect 12436 33700 12460 33702
rect 12516 33700 12522 33702
rect 12214 33680 12522 33700
rect 12636 33561 12664 34598
rect 13096 34598 13492 34626
rect 12992 34546 13044 34552
rect 12898 34368 12954 34377
rect 12898 34303 12954 34312
rect 12714 34232 12770 34241
rect 12912 34202 12940 34303
rect 12714 34167 12770 34176
rect 12900 34196 12952 34202
rect 12622 33552 12678 33561
rect 12728 33522 12756 34167
rect 12900 34138 12952 34144
rect 13084 34196 13136 34202
rect 13084 34138 13136 34144
rect 13096 33522 13124 34138
rect 13464 34134 13492 34598
rect 13452 34128 13504 34134
rect 13266 34096 13322 34105
rect 13452 34070 13504 34076
rect 13266 34031 13268 34040
rect 13320 34031 13322 34040
rect 13268 34002 13320 34008
rect 13450 33960 13506 33969
rect 13268 33924 13320 33930
rect 13450 33895 13506 33904
rect 13268 33866 13320 33872
rect 13176 33652 13228 33658
rect 13176 33594 13228 33600
rect 12622 33487 12678 33496
rect 12716 33516 12768 33522
rect 12164 33448 12216 33454
rect 12164 33390 12216 33396
rect 12176 33114 12204 33390
rect 12164 33108 12216 33114
rect 12164 33050 12216 33056
rect 12214 32668 12522 32688
rect 12214 32666 12220 32668
rect 12276 32666 12300 32668
rect 12356 32666 12380 32668
rect 12436 32666 12460 32668
rect 12516 32666 12522 32668
rect 12276 32614 12278 32666
rect 12458 32614 12460 32666
rect 12214 32612 12220 32614
rect 12276 32612 12300 32614
rect 12356 32612 12380 32614
rect 12436 32612 12460 32614
rect 12516 32612 12522 32614
rect 12214 32592 12522 32612
rect 12636 32434 12664 33487
rect 12716 33458 12768 33464
rect 13084 33516 13136 33522
rect 13084 33458 13136 33464
rect 13188 33318 13216 33594
rect 12808 33312 12860 33318
rect 12806 33280 12808 33289
rect 13176 33312 13228 33318
rect 12860 33280 12862 33289
rect 13176 33254 13228 33260
rect 12806 33215 12862 33224
rect 12900 32904 12952 32910
rect 12900 32846 12952 32852
rect 13176 32904 13228 32910
rect 13176 32846 13228 32852
rect 12808 32836 12860 32842
rect 12808 32778 12860 32784
rect 12820 32570 12848 32778
rect 12912 32570 12940 32846
rect 12990 32736 13046 32745
rect 12990 32671 13046 32680
rect 12808 32564 12860 32570
rect 12808 32506 12860 32512
rect 12900 32564 12952 32570
rect 12900 32506 12952 32512
rect 13004 32502 13032 32671
rect 12992 32496 13044 32502
rect 12806 32464 12862 32473
rect 12624 32428 12676 32434
rect 12992 32438 13044 32444
rect 12806 32399 12862 32408
rect 12900 32428 12952 32434
rect 12624 32370 12676 32376
rect 12348 32292 12400 32298
rect 12348 32234 12400 32240
rect 12360 31822 12388 32234
rect 12348 31816 12400 31822
rect 12348 31758 12400 31764
rect 12214 31580 12522 31600
rect 12214 31578 12220 31580
rect 12276 31578 12300 31580
rect 12356 31578 12380 31580
rect 12436 31578 12460 31580
rect 12516 31578 12522 31580
rect 12276 31526 12278 31578
rect 12458 31526 12460 31578
rect 12214 31524 12220 31526
rect 12276 31524 12300 31526
rect 12356 31524 12380 31526
rect 12436 31524 12460 31526
rect 12516 31524 12522 31526
rect 12214 31504 12522 31524
rect 12256 31340 12308 31346
rect 12256 31282 12308 31288
rect 12070 31104 12126 31113
rect 12070 31039 12126 31048
rect 12084 30938 12112 31039
rect 12072 30932 12124 30938
rect 12072 30874 12124 30880
rect 12268 30870 12296 31282
rect 12256 30864 12308 30870
rect 12256 30806 12308 30812
rect 12636 30734 12664 32370
rect 12820 31822 12848 32399
rect 12900 32370 12952 32376
rect 13084 32428 13136 32434
rect 13084 32370 13136 32376
rect 12808 31816 12860 31822
rect 12912 31793 12940 32370
rect 12992 31816 13044 31822
rect 12808 31758 12860 31764
rect 12898 31784 12954 31793
rect 12992 31758 13044 31764
rect 12898 31719 12954 31728
rect 12716 31680 12768 31686
rect 12716 31622 12768 31628
rect 12728 31521 12756 31622
rect 12714 31512 12770 31521
rect 13004 31482 13032 31758
rect 12714 31447 12770 31456
rect 12992 31476 13044 31482
rect 12992 31418 13044 31424
rect 12900 31340 12952 31346
rect 12952 31300 13032 31328
rect 12900 31282 12952 31288
rect 12806 30832 12862 30841
rect 12806 30767 12808 30776
rect 12860 30767 12862 30776
rect 12808 30738 12860 30744
rect 13004 30734 13032 31300
rect 13096 30938 13124 32370
rect 13188 31090 13216 32846
rect 13280 32201 13308 33866
rect 13464 33522 13492 33895
rect 13360 33516 13412 33522
rect 13360 33458 13412 33464
rect 13452 33516 13504 33522
rect 13452 33458 13504 33464
rect 13372 33017 13400 33458
rect 13556 33046 13584 34870
rect 13636 34672 13688 34678
rect 13636 34614 13688 34620
rect 13648 33658 13676 34614
rect 13636 33652 13688 33658
rect 13636 33594 13688 33600
rect 13740 33538 13768 36042
rect 13910 35864 13966 35873
rect 13910 35799 13966 35808
rect 13924 35630 13952 35799
rect 13912 35624 13964 35630
rect 13912 35566 13964 35572
rect 13820 35488 13872 35494
rect 14016 35442 14044 40015
rect 14094 39672 14150 39681
rect 14094 39607 14150 39616
rect 13820 35430 13872 35436
rect 13832 35018 13860 35430
rect 13924 35414 14044 35442
rect 13924 35086 13952 35414
rect 14108 35290 14136 39607
rect 14188 38888 14240 38894
rect 14188 38830 14240 38836
rect 14200 38554 14228 38830
rect 14188 38548 14240 38554
rect 14188 38490 14240 38496
rect 14292 38162 14320 40287
rect 14476 39438 14504 40326
rect 14464 39432 14516 39438
rect 14464 39374 14516 39380
rect 14372 38888 14424 38894
rect 14372 38830 14424 38836
rect 14384 38554 14412 38830
rect 14372 38548 14424 38554
rect 14372 38490 14424 38496
rect 14648 38548 14700 38554
rect 14648 38490 14700 38496
rect 14384 38406 14596 38434
rect 14660 38418 14688 38490
rect 14384 38350 14412 38406
rect 14372 38344 14424 38350
rect 14372 38286 14424 38292
rect 14464 38344 14516 38350
rect 14464 38286 14516 38292
rect 14200 38134 14320 38162
rect 14200 38010 14228 38134
rect 14278 38040 14334 38049
rect 14188 38004 14240 38010
rect 14278 37975 14334 37984
rect 14188 37946 14240 37952
rect 14096 35284 14148 35290
rect 14096 35226 14148 35232
rect 14002 35184 14058 35193
rect 14002 35119 14058 35128
rect 13912 35080 13964 35086
rect 13912 35022 13964 35028
rect 13820 35012 13872 35018
rect 13820 34954 13872 34960
rect 14016 34474 14044 35119
rect 14200 35034 14228 37946
rect 14292 35154 14320 37975
rect 14476 37942 14504 38286
rect 14464 37936 14516 37942
rect 14464 37878 14516 37884
rect 14372 37868 14424 37874
rect 14372 37810 14424 37816
rect 14384 37262 14412 37810
rect 14372 37256 14424 37262
rect 14372 37198 14424 37204
rect 14384 37126 14412 37198
rect 14372 37120 14424 37126
rect 14372 37062 14424 37068
rect 14384 36786 14412 37062
rect 14372 36780 14424 36786
rect 14372 36722 14424 36728
rect 14384 36174 14412 36722
rect 14568 36718 14596 38406
rect 14648 38412 14700 38418
rect 14648 38354 14700 38360
rect 14556 36712 14608 36718
rect 14556 36654 14608 36660
rect 14372 36168 14424 36174
rect 14372 36110 14424 36116
rect 14464 36168 14516 36174
rect 14464 36110 14516 36116
rect 14372 36032 14424 36038
rect 14372 35974 14424 35980
rect 14384 35698 14412 35974
rect 14372 35692 14424 35698
rect 14372 35634 14424 35640
rect 14476 35578 14504 36110
rect 14384 35550 14504 35578
rect 14280 35148 14332 35154
rect 14280 35090 14332 35096
rect 14200 35006 14320 35034
rect 14188 34604 14240 34610
rect 14188 34546 14240 34552
rect 14004 34468 14056 34474
rect 14004 34410 14056 34416
rect 14200 34406 14228 34546
rect 14188 34400 14240 34406
rect 14188 34342 14240 34348
rect 14004 33992 14056 33998
rect 14004 33934 14056 33940
rect 14188 33992 14240 33998
rect 14188 33934 14240 33940
rect 13740 33510 13860 33538
rect 13634 33144 13690 33153
rect 13634 33079 13690 33088
rect 13544 33040 13596 33046
rect 13358 33008 13414 33017
rect 13544 32982 13596 32988
rect 13358 32943 13414 32952
rect 13648 32910 13676 33079
rect 13832 33028 13860 33510
rect 13912 33448 13964 33454
rect 13910 33416 13912 33425
rect 13964 33416 13966 33425
rect 13910 33351 13966 33360
rect 13832 33000 13952 33028
rect 13636 32904 13688 32910
rect 13688 32864 13860 32892
rect 13636 32846 13688 32852
rect 13636 32224 13688 32230
rect 13266 32192 13322 32201
rect 13636 32166 13688 32172
rect 13266 32127 13322 32136
rect 13648 31929 13676 32166
rect 13634 31920 13690 31929
rect 13634 31855 13690 31864
rect 13728 31680 13780 31686
rect 13728 31622 13780 31628
rect 13634 31376 13690 31385
rect 13740 31346 13768 31622
rect 13832 31346 13860 32864
rect 13634 31311 13690 31320
rect 13728 31340 13780 31346
rect 13544 31136 13596 31142
rect 13188 31062 13400 31090
rect 13544 31078 13596 31084
rect 13266 30968 13322 30977
rect 13084 30932 13136 30938
rect 13266 30903 13322 30912
rect 13084 30874 13136 30880
rect 11980 30728 12032 30734
rect 11980 30670 12032 30676
rect 12624 30728 12676 30734
rect 12624 30670 12676 30676
rect 12992 30728 13044 30734
rect 12992 30670 13044 30676
rect 13174 30696 13230 30705
rect 11888 29640 11940 29646
rect 11888 29582 11940 29588
rect 11992 28801 12020 30670
rect 13174 30631 13176 30640
rect 13228 30631 13230 30640
rect 13176 30602 13228 30608
rect 12214 30492 12522 30512
rect 12214 30490 12220 30492
rect 12276 30490 12300 30492
rect 12356 30490 12380 30492
rect 12436 30490 12460 30492
rect 12516 30490 12522 30492
rect 12276 30438 12278 30490
rect 12458 30438 12460 30490
rect 12214 30436 12220 30438
rect 12276 30436 12300 30438
rect 12356 30436 12380 30438
rect 12436 30436 12460 30438
rect 12516 30436 12522 30438
rect 12214 30416 12522 30436
rect 13280 30258 13308 30903
rect 12440 30252 12492 30258
rect 12624 30252 12676 30258
rect 12492 30212 12624 30240
rect 12440 30194 12492 30200
rect 12624 30194 12676 30200
rect 12808 30252 12860 30258
rect 12808 30194 12860 30200
rect 13268 30252 13320 30258
rect 13268 30194 13320 30200
rect 12714 29880 12770 29889
rect 12714 29815 12770 29824
rect 12728 29646 12756 29815
rect 12716 29640 12768 29646
rect 12716 29582 12768 29588
rect 12214 29404 12522 29424
rect 12214 29402 12220 29404
rect 12276 29402 12300 29404
rect 12356 29402 12380 29404
rect 12436 29402 12460 29404
rect 12516 29402 12522 29404
rect 12276 29350 12278 29402
rect 12458 29350 12460 29402
rect 12214 29348 12220 29350
rect 12276 29348 12300 29350
rect 12356 29348 12380 29350
rect 12436 29348 12460 29350
rect 12516 29348 12522 29350
rect 12214 29328 12522 29348
rect 12164 28960 12216 28966
rect 12164 28902 12216 28908
rect 11978 28792 12034 28801
rect 11978 28727 12034 28736
rect 12176 28626 12204 28902
rect 12164 28620 12216 28626
rect 12164 28562 12216 28568
rect 12214 28316 12522 28336
rect 12214 28314 12220 28316
rect 12276 28314 12300 28316
rect 12356 28314 12380 28316
rect 12436 28314 12460 28316
rect 12516 28314 12522 28316
rect 12276 28262 12278 28314
rect 12458 28262 12460 28314
rect 12214 28260 12220 28262
rect 12276 28260 12300 28262
rect 12356 28260 12380 28262
rect 12436 28260 12460 28262
rect 12516 28260 12522 28262
rect 12214 28240 12522 28260
rect 12214 27228 12522 27248
rect 12214 27226 12220 27228
rect 12276 27226 12300 27228
rect 12356 27226 12380 27228
rect 12436 27226 12460 27228
rect 12516 27226 12522 27228
rect 12276 27174 12278 27226
rect 12458 27174 12460 27226
rect 12214 27172 12220 27174
rect 12276 27172 12300 27174
rect 12356 27172 12380 27174
rect 12436 27172 12460 27174
rect 12516 27172 12522 27174
rect 12214 27152 12522 27172
rect 8956 26206 9260 26234
rect 6582 25596 6890 25616
rect 6582 25594 6588 25596
rect 6644 25594 6668 25596
rect 6724 25594 6748 25596
rect 6804 25594 6828 25596
rect 6884 25594 6890 25596
rect 6644 25542 6646 25594
rect 6826 25542 6828 25594
rect 6582 25540 6588 25542
rect 6644 25540 6668 25542
rect 6724 25540 6748 25542
rect 6804 25540 6828 25542
rect 6884 25540 6890 25542
rect 6582 25520 6890 25540
rect 6582 24508 6890 24528
rect 6582 24506 6588 24508
rect 6644 24506 6668 24508
rect 6724 24506 6748 24508
rect 6804 24506 6828 24508
rect 6884 24506 6890 24508
rect 6644 24454 6646 24506
rect 6826 24454 6828 24506
rect 6582 24452 6588 24454
rect 6644 24452 6668 24454
rect 6724 24452 6748 24454
rect 6804 24452 6828 24454
rect 6884 24452 6890 24454
rect 6582 24432 6890 24452
rect 6582 23420 6890 23440
rect 6582 23418 6588 23420
rect 6644 23418 6668 23420
rect 6724 23418 6748 23420
rect 6804 23418 6828 23420
rect 6884 23418 6890 23420
rect 6644 23366 6646 23418
rect 6826 23366 6828 23418
rect 6582 23364 6588 23366
rect 6644 23364 6668 23366
rect 6724 23364 6748 23366
rect 6804 23364 6828 23366
rect 6884 23364 6890 23366
rect 6582 23344 6890 23364
rect 6582 22332 6890 22352
rect 6582 22330 6588 22332
rect 6644 22330 6668 22332
rect 6724 22330 6748 22332
rect 6804 22330 6828 22332
rect 6884 22330 6890 22332
rect 6644 22278 6646 22330
rect 6826 22278 6828 22330
rect 6582 22276 6588 22278
rect 6644 22276 6668 22278
rect 6724 22276 6748 22278
rect 6804 22276 6828 22278
rect 6884 22276 6890 22278
rect 6582 22256 6890 22276
rect 6582 21244 6890 21264
rect 6582 21242 6588 21244
rect 6644 21242 6668 21244
rect 6724 21242 6748 21244
rect 6804 21242 6828 21244
rect 6884 21242 6890 21244
rect 6644 21190 6646 21242
rect 6826 21190 6828 21242
rect 6582 21188 6588 21190
rect 6644 21188 6668 21190
rect 6724 21188 6748 21190
rect 6804 21188 6828 21190
rect 6884 21188 6890 21190
rect 6582 21168 6890 21188
rect 6582 20156 6890 20176
rect 6582 20154 6588 20156
rect 6644 20154 6668 20156
rect 6724 20154 6748 20156
rect 6804 20154 6828 20156
rect 6884 20154 6890 20156
rect 6644 20102 6646 20154
rect 6826 20102 6828 20154
rect 6582 20100 6588 20102
rect 6644 20100 6668 20102
rect 6724 20100 6748 20102
rect 6804 20100 6828 20102
rect 6884 20100 6890 20102
rect 6582 20080 6890 20100
rect 6582 19068 6890 19088
rect 6582 19066 6588 19068
rect 6644 19066 6668 19068
rect 6724 19066 6748 19068
rect 6804 19066 6828 19068
rect 6884 19066 6890 19068
rect 6644 19014 6646 19066
rect 6826 19014 6828 19066
rect 6582 19012 6588 19014
rect 6644 19012 6668 19014
rect 6724 19012 6748 19014
rect 6804 19012 6828 19014
rect 6884 19012 6890 19014
rect 6582 18992 6890 19012
rect 6582 17980 6890 18000
rect 6582 17978 6588 17980
rect 6644 17978 6668 17980
rect 6724 17978 6748 17980
rect 6804 17978 6828 17980
rect 6884 17978 6890 17980
rect 6644 17926 6646 17978
rect 6826 17926 6828 17978
rect 6582 17924 6588 17926
rect 6644 17924 6668 17926
rect 6724 17924 6748 17926
rect 6804 17924 6828 17926
rect 6884 17924 6890 17926
rect 6582 17904 6890 17924
rect 5080 17332 5132 17338
rect 5080 17274 5132 17280
rect 5092 6914 5120 17274
rect 6582 16892 6890 16912
rect 6582 16890 6588 16892
rect 6644 16890 6668 16892
rect 6724 16890 6748 16892
rect 6804 16890 6828 16892
rect 6884 16890 6890 16892
rect 6644 16838 6646 16890
rect 6826 16838 6828 16890
rect 6582 16836 6588 16838
rect 6644 16836 6668 16838
rect 6724 16836 6748 16838
rect 6804 16836 6828 16838
rect 6884 16836 6890 16838
rect 6582 16816 6890 16836
rect 6582 15804 6890 15824
rect 6582 15802 6588 15804
rect 6644 15802 6668 15804
rect 6724 15802 6748 15804
rect 6804 15802 6828 15804
rect 6884 15802 6890 15804
rect 6644 15750 6646 15802
rect 6826 15750 6828 15802
rect 6582 15748 6588 15750
rect 6644 15748 6668 15750
rect 6724 15748 6748 15750
rect 6804 15748 6828 15750
rect 6884 15748 6890 15750
rect 6582 15728 6890 15748
rect 6582 14716 6890 14736
rect 6582 14714 6588 14716
rect 6644 14714 6668 14716
rect 6724 14714 6748 14716
rect 6804 14714 6828 14716
rect 6884 14714 6890 14716
rect 6644 14662 6646 14714
rect 6826 14662 6828 14714
rect 6582 14660 6588 14662
rect 6644 14660 6668 14662
rect 6724 14660 6748 14662
rect 6804 14660 6828 14662
rect 6884 14660 6890 14662
rect 6582 14640 6890 14660
rect 7932 13932 7984 13938
rect 7932 13874 7984 13880
rect 6582 13628 6890 13648
rect 6582 13626 6588 13628
rect 6644 13626 6668 13628
rect 6724 13626 6748 13628
rect 6804 13626 6828 13628
rect 6884 13626 6890 13628
rect 6644 13574 6646 13626
rect 6826 13574 6828 13626
rect 6582 13572 6588 13574
rect 6644 13572 6668 13574
rect 6724 13572 6748 13574
rect 6804 13572 6828 13574
rect 6884 13572 6890 13574
rect 6582 13552 6890 13572
rect 6582 12540 6890 12560
rect 6582 12538 6588 12540
rect 6644 12538 6668 12540
rect 6724 12538 6748 12540
rect 6804 12538 6828 12540
rect 6884 12538 6890 12540
rect 6644 12486 6646 12538
rect 6826 12486 6828 12538
rect 6582 12484 6588 12486
rect 6644 12484 6668 12486
rect 6724 12484 6748 12486
rect 6804 12484 6828 12486
rect 6884 12484 6890 12486
rect 6582 12464 6890 12484
rect 6582 11452 6890 11472
rect 6582 11450 6588 11452
rect 6644 11450 6668 11452
rect 6724 11450 6748 11452
rect 6804 11450 6828 11452
rect 6884 11450 6890 11452
rect 6644 11398 6646 11450
rect 6826 11398 6828 11450
rect 6582 11396 6588 11398
rect 6644 11396 6668 11398
rect 6724 11396 6748 11398
rect 6804 11396 6828 11398
rect 6884 11396 6890 11398
rect 6582 11376 6890 11396
rect 6582 10364 6890 10384
rect 6582 10362 6588 10364
rect 6644 10362 6668 10364
rect 6724 10362 6748 10364
rect 6804 10362 6828 10364
rect 6884 10362 6890 10364
rect 6644 10310 6646 10362
rect 6826 10310 6828 10362
rect 6582 10308 6588 10310
rect 6644 10308 6668 10310
rect 6724 10308 6748 10310
rect 6804 10308 6828 10310
rect 6884 10308 6890 10310
rect 6582 10288 6890 10308
rect 6582 9276 6890 9296
rect 6582 9274 6588 9276
rect 6644 9274 6668 9276
rect 6724 9274 6748 9276
rect 6804 9274 6828 9276
rect 6884 9274 6890 9276
rect 6644 9222 6646 9274
rect 6826 9222 6828 9274
rect 6582 9220 6588 9222
rect 6644 9220 6668 9222
rect 6724 9220 6748 9222
rect 6804 9220 6828 9222
rect 6884 9220 6890 9222
rect 6582 9200 6890 9220
rect 6582 8188 6890 8208
rect 6582 8186 6588 8188
rect 6644 8186 6668 8188
rect 6724 8186 6748 8188
rect 6804 8186 6828 8188
rect 6884 8186 6890 8188
rect 6644 8134 6646 8186
rect 6826 8134 6828 8186
rect 6582 8132 6588 8134
rect 6644 8132 6668 8134
rect 6724 8132 6748 8134
rect 6804 8132 6828 8134
rect 6884 8132 6890 8134
rect 6582 8112 6890 8132
rect 6582 7100 6890 7120
rect 6582 7098 6588 7100
rect 6644 7098 6668 7100
rect 6724 7098 6748 7100
rect 6804 7098 6828 7100
rect 6884 7098 6890 7100
rect 6644 7046 6646 7098
rect 6826 7046 6828 7098
rect 6582 7044 6588 7046
rect 6644 7044 6668 7046
rect 6724 7044 6748 7046
rect 6804 7044 6828 7046
rect 6884 7044 6890 7046
rect 6582 7024 6890 7044
rect 4908 6886 5120 6914
rect 4712 5364 4764 5370
rect 4712 5306 4764 5312
rect 4436 5024 4488 5030
rect 4436 4966 4488 4972
rect 4252 4616 4304 4622
rect 4252 4558 4304 4564
rect 4264 4214 4292 4558
rect 4252 4208 4304 4214
rect 4252 4150 4304 4156
rect 4264 3738 4292 4150
rect 4344 4072 4396 4078
rect 4344 4014 4396 4020
rect 4252 3732 4304 3738
rect 4252 3674 4304 3680
rect 4264 2990 4292 3674
rect 4252 2984 4304 2990
rect 4252 2926 4304 2932
rect 3896 2774 4200 2802
rect 3424 2644 3476 2650
rect 3424 2586 3476 2592
rect 3240 2304 3292 2310
rect 3240 2246 3292 2252
rect 2870 2136 2926 2145
rect 2870 2071 2926 2080
rect 3252 800 3280 2246
rect 3436 1465 3464 2586
rect 3422 1456 3478 1465
rect 3422 1391 3478 1400
rect 3896 800 3924 2774
rect 4356 2582 4384 4014
rect 4448 3602 4476 4966
rect 4724 4554 4752 5306
rect 4908 4690 4936 6886
rect 6460 6180 6512 6186
rect 6460 6122 6512 6128
rect 5172 6112 5224 6118
rect 5172 6054 5224 6060
rect 5184 5302 5212 6054
rect 6276 5704 6328 5710
rect 6276 5646 6328 5652
rect 5172 5296 5224 5302
rect 5172 5238 5224 5244
rect 5172 5024 5224 5030
rect 5172 4966 5224 4972
rect 5184 4690 5212 4966
rect 4896 4684 4948 4690
rect 4896 4626 4948 4632
rect 5172 4684 5224 4690
rect 5172 4626 5224 4632
rect 4712 4548 4764 4554
rect 4712 4490 4764 4496
rect 5356 4548 5408 4554
rect 5356 4490 5408 4496
rect 5368 4010 5396 4490
rect 5356 4004 5408 4010
rect 5356 3946 5408 3952
rect 4620 3936 4672 3942
rect 4620 3878 4672 3884
rect 5540 3936 5592 3942
rect 5540 3878 5592 3884
rect 4632 3602 4660 3878
rect 4436 3596 4488 3602
rect 4436 3538 4488 3544
rect 4620 3596 4672 3602
rect 4620 3538 4672 3544
rect 5172 3596 5224 3602
rect 5172 3538 5224 3544
rect 5264 3596 5316 3602
rect 5264 3538 5316 3544
rect 4712 2848 4764 2854
rect 4712 2790 4764 2796
rect 4344 2576 4396 2582
rect 4344 2518 4396 2524
rect 4528 2576 4580 2582
rect 4528 2518 4580 2524
rect 4540 800 4568 2518
rect 4724 2514 4752 2790
rect 4712 2508 4764 2514
rect 4712 2450 4764 2456
rect 5184 800 5212 3538
rect 5276 2378 5304 3538
rect 5552 3194 5580 3878
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 6288 3058 6316 5646
rect 6472 5234 6500 6122
rect 6582 6012 6890 6032
rect 6582 6010 6588 6012
rect 6644 6010 6668 6012
rect 6724 6010 6748 6012
rect 6804 6010 6828 6012
rect 6884 6010 6890 6012
rect 6644 5958 6646 6010
rect 6826 5958 6828 6010
rect 6582 5956 6588 5958
rect 6644 5956 6668 5958
rect 6724 5956 6748 5958
rect 6804 5956 6828 5958
rect 6884 5956 6890 5958
rect 6582 5936 6890 5956
rect 6460 5228 6512 5234
rect 6460 5170 6512 5176
rect 6582 4924 6890 4944
rect 6582 4922 6588 4924
rect 6644 4922 6668 4924
rect 6724 4922 6748 4924
rect 6804 4922 6828 4924
rect 6884 4922 6890 4924
rect 6644 4870 6646 4922
rect 6826 4870 6828 4922
rect 6582 4868 6588 4870
rect 6644 4868 6668 4870
rect 6724 4868 6748 4870
rect 6804 4868 6828 4870
rect 6884 4868 6890 4870
rect 6582 4848 6890 4868
rect 7748 4616 7800 4622
rect 7748 4558 7800 4564
rect 6368 4480 6420 4486
rect 6368 4422 6420 4428
rect 6276 3052 6328 3058
rect 6276 2994 6328 3000
rect 6380 2378 6408 4422
rect 7760 4146 7788 4558
rect 7748 4140 7800 4146
rect 7748 4082 7800 4088
rect 6920 3936 6972 3942
rect 6920 3878 6972 3884
rect 6582 3836 6890 3856
rect 6582 3834 6588 3836
rect 6644 3834 6668 3836
rect 6724 3834 6748 3836
rect 6804 3834 6828 3836
rect 6884 3834 6890 3836
rect 6644 3782 6646 3834
rect 6826 3782 6828 3834
rect 6582 3780 6588 3782
rect 6644 3780 6668 3782
rect 6724 3780 6748 3782
rect 6804 3780 6828 3782
rect 6884 3780 6890 3782
rect 6582 3760 6890 3780
rect 6460 2916 6512 2922
rect 6460 2858 6512 2864
rect 5264 2372 5316 2378
rect 5264 2314 5316 2320
rect 6368 2372 6420 2378
rect 6368 2314 6420 2320
rect 6472 800 6500 2858
rect 6582 2748 6890 2768
rect 6582 2746 6588 2748
rect 6644 2746 6668 2748
rect 6724 2746 6748 2748
rect 6804 2746 6828 2748
rect 6884 2746 6890 2748
rect 6644 2694 6646 2746
rect 6826 2694 6828 2746
rect 6582 2692 6588 2694
rect 6644 2692 6668 2694
rect 6724 2692 6748 2694
rect 6804 2692 6828 2694
rect 6884 2692 6890 2694
rect 6582 2672 6890 2692
rect 6932 2514 6960 3878
rect 7840 3732 7892 3738
rect 7840 3674 7892 3680
rect 7852 2854 7880 3674
rect 7944 3534 7972 13874
rect 8024 4072 8076 4078
rect 8024 4014 8076 4020
rect 8392 4072 8444 4078
rect 8392 4014 8444 4020
rect 8036 3738 8064 4014
rect 8024 3732 8076 3738
rect 8024 3674 8076 3680
rect 7932 3528 7984 3534
rect 7932 3470 7984 3476
rect 7840 2848 7892 2854
rect 7840 2790 7892 2796
rect 6920 2508 6972 2514
rect 6920 2450 6972 2456
rect 8404 800 8432 4014
rect 8956 3534 8984 26206
rect 12214 26140 12522 26160
rect 12214 26138 12220 26140
rect 12276 26138 12300 26140
rect 12356 26138 12380 26140
rect 12436 26138 12460 26140
rect 12516 26138 12522 26140
rect 12276 26086 12278 26138
rect 12458 26086 12460 26138
rect 12214 26084 12220 26086
rect 12276 26084 12300 26086
rect 12356 26084 12380 26086
rect 12436 26084 12460 26086
rect 12516 26084 12522 26086
rect 12214 26064 12522 26084
rect 12214 25052 12522 25072
rect 12214 25050 12220 25052
rect 12276 25050 12300 25052
rect 12356 25050 12380 25052
rect 12436 25050 12460 25052
rect 12516 25050 12522 25052
rect 12276 24998 12278 25050
rect 12458 24998 12460 25050
rect 12214 24996 12220 24998
rect 12276 24996 12300 24998
rect 12356 24996 12380 24998
rect 12436 24996 12460 24998
rect 12516 24996 12522 24998
rect 12214 24976 12522 24996
rect 12820 24721 12848 30194
rect 12990 30152 13046 30161
rect 12990 30087 13046 30096
rect 12900 29640 12952 29646
rect 12900 29582 12952 29588
rect 12806 24712 12862 24721
rect 12806 24647 12862 24656
rect 12214 23964 12522 23984
rect 12214 23962 12220 23964
rect 12276 23962 12300 23964
rect 12356 23962 12380 23964
rect 12436 23962 12460 23964
rect 12516 23962 12522 23964
rect 12276 23910 12278 23962
rect 12458 23910 12460 23962
rect 12214 23908 12220 23910
rect 12276 23908 12300 23910
rect 12356 23908 12380 23910
rect 12436 23908 12460 23910
rect 12516 23908 12522 23910
rect 12214 23888 12522 23908
rect 12214 22876 12522 22896
rect 12214 22874 12220 22876
rect 12276 22874 12300 22876
rect 12356 22874 12380 22876
rect 12436 22874 12460 22876
rect 12516 22874 12522 22876
rect 12276 22822 12278 22874
rect 12458 22822 12460 22874
rect 12214 22820 12220 22822
rect 12276 22820 12300 22822
rect 12356 22820 12380 22822
rect 12436 22820 12460 22822
rect 12516 22820 12522 22822
rect 12214 22800 12522 22820
rect 12214 21788 12522 21808
rect 12214 21786 12220 21788
rect 12276 21786 12300 21788
rect 12356 21786 12380 21788
rect 12436 21786 12460 21788
rect 12516 21786 12522 21788
rect 12276 21734 12278 21786
rect 12458 21734 12460 21786
rect 12214 21732 12220 21734
rect 12276 21732 12300 21734
rect 12356 21732 12380 21734
rect 12436 21732 12460 21734
rect 12516 21732 12522 21734
rect 12214 21712 12522 21732
rect 12214 20700 12522 20720
rect 12214 20698 12220 20700
rect 12276 20698 12300 20700
rect 12356 20698 12380 20700
rect 12436 20698 12460 20700
rect 12516 20698 12522 20700
rect 12276 20646 12278 20698
rect 12458 20646 12460 20698
rect 12214 20644 12220 20646
rect 12276 20644 12300 20646
rect 12356 20644 12380 20646
rect 12436 20644 12460 20646
rect 12516 20644 12522 20646
rect 12214 20624 12522 20644
rect 12214 19612 12522 19632
rect 12214 19610 12220 19612
rect 12276 19610 12300 19612
rect 12356 19610 12380 19612
rect 12436 19610 12460 19612
rect 12516 19610 12522 19612
rect 12276 19558 12278 19610
rect 12458 19558 12460 19610
rect 12214 19556 12220 19558
rect 12276 19556 12300 19558
rect 12356 19556 12380 19558
rect 12436 19556 12460 19558
rect 12516 19556 12522 19558
rect 12214 19536 12522 19556
rect 12214 18524 12522 18544
rect 12214 18522 12220 18524
rect 12276 18522 12300 18524
rect 12356 18522 12380 18524
rect 12436 18522 12460 18524
rect 12516 18522 12522 18524
rect 12276 18470 12278 18522
rect 12458 18470 12460 18522
rect 12214 18468 12220 18470
rect 12276 18468 12300 18470
rect 12356 18468 12380 18470
rect 12436 18468 12460 18470
rect 12516 18468 12522 18470
rect 12214 18448 12522 18468
rect 12214 17436 12522 17456
rect 12214 17434 12220 17436
rect 12276 17434 12300 17436
rect 12356 17434 12380 17436
rect 12436 17434 12460 17436
rect 12516 17434 12522 17436
rect 12276 17382 12278 17434
rect 12458 17382 12460 17434
rect 12214 17380 12220 17382
rect 12276 17380 12300 17382
rect 12356 17380 12380 17382
rect 12436 17380 12460 17382
rect 12516 17380 12522 17382
rect 12214 17360 12522 17380
rect 12912 17134 12940 29582
rect 13004 29306 13032 30087
rect 13176 30048 13228 30054
rect 13176 29990 13228 29996
rect 12992 29300 13044 29306
rect 12992 29242 13044 29248
rect 13082 28792 13138 28801
rect 13082 28727 13138 28736
rect 13096 25809 13124 28727
rect 13082 25800 13138 25809
rect 13082 25735 13138 25744
rect 13188 22817 13216 29990
rect 13372 29646 13400 31062
rect 13556 30938 13584 31078
rect 13544 30932 13596 30938
rect 13544 30874 13596 30880
rect 13544 30728 13596 30734
rect 13544 30670 13596 30676
rect 13450 30424 13506 30433
rect 13450 30359 13506 30368
rect 13360 29640 13412 29646
rect 13360 29582 13412 29588
rect 13268 29504 13320 29510
rect 13268 29446 13320 29452
rect 13280 29170 13308 29446
rect 13268 29164 13320 29170
rect 13268 29106 13320 29112
rect 13268 28484 13320 28490
rect 13268 28426 13320 28432
rect 13280 28218 13308 28426
rect 13268 28212 13320 28218
rect 13268 28154 13320 28160
rect 13372 27713 13400 29582
rect 13464 28966 13492 30359
rect 13452 28960 13504 28966
rect 13452 28902 13504 28908
rect 13452 28552 13504 28558
rect 13452 28494 13504 28500
rect 13464 27985 13492 28494
rect 13450 27976 13506 27985
rect 13450 27911 13506 27920
rect 13358 27704 13414 27713
rect 13358 27639 13414 27648
rect 13556 27169 13584 30670
rect 13648 29170 13676 31311
rect 13728 31282 13780 31288
rect 13820 31340 13872 31346
rect 13820 31282 13872 31288
rect 13740 30258 13768 31282
rect 13820 30388 13872 30394
rect 13820 30330 13872 30336
rect 13728 30252 13780 30258
rect 13728 30194 13780 30200
rect 13726 29336 13782 29345
rect 13726 29271 13782 29280
rect 13636 29164 13688 29170
rect 13636 29106 13688 29112
rect 13648 28966 13676 29106
rect 13740 29102 13768 29271
rect 13832 29238 13860 30330
rect 13820 29232 13872 29238
rect 13820 29174 13872 29180
rect 13728 29096 13780 29102
rect 13728 29038 13780 29044
rect 13820 29096 13872 29102
rect 13820 29038 13872 29044
rect 13636 28960 13688 28966
rect 13636 28902 13688 28908
rect 13728 28552 13780 28558
rect 13728 28494 13780 28500
rect 13740 27402 13768 28494
rect 13832 28150 13860 29038
rect 13820 28144 13872 28150
rect 13820 28086 13872 28092
rect 13728 27396 13780 27402
rect 13728 27338 13780 27344
rect 13542 27160 13598 27169
rect 13542 27095 13598 27104
rect 13542 27024 13598 27033
rect 13542 26959 13544 26968
rect 13596 26959 13598 26968
rect 13544 26930 13596 26936
rect 13820 25696 13872 25702
rect 13820 25638 13872 25644
rect 13832 25362 13860 25638
rect 13820 25356 13872 25362
rect 13820 25298 13872 25304
rect 13174 22808 13230 22817
rect 13174 22743 13230 22752
rect 13924 22094 13952 33000
rect 14016 32881 14044 33934
rect 14002 32872 14058 32881
rect 14002 32807 14058 32816
rect 14094 32600 14150 32609
rect 14094 32535 14150 32544
rect 14004 31272 14056 31278
rect 14004 31214 14056 31220
rect 14016 31142 14044 31214
rect 14004 31136 14056 31142
rect 14004 31078 14056 31084
rect 14004 29640 14056 29646
rect 14004 29582 14056 29588
rect 14016 29209 14044 29582
rect 14002 29200 14058 29209
rect 14002 29135 14058 29144
rect 14004 29096 14056 29102
rect 14002 29064 14004 29073
rect 14056 29064 14058 29073
rect 14002 28999 14058 29008
rect 14004 28960 14056 28966
rect 14004 28902 14056 28908
rect 14016 28082 14044 28902
rect 14004 28076 14056 28082
rect 14004 28018 14056 28024
rect 13832 22066 13952 22094
rect 12900 17128 12952 17134
rect 12900 17070 12952 17076
rect 12214 16348 12522 16368
rect 12214 16346 12220 16348
rect 12276 16346 12300 16348
rect 12356 16346 12380 16348
rect 12436 16346 12460 16348
rect 12516 16346 12522 16348
rect 12276 16294 12278 16346
rect 12458 16294 12460 16346
rect 12214 16292 12220 16294
rect 12276 16292 12300 16294
rect 12356 16292 12380 16294
rect 12436 16292 12460 16294
rect 12516 16292 12522 16294
rect 12214 16272 12522 16292
rect 12214 15260 12522 15280
rect 12214 15258 12220 15260
rect 12276 15258 12300 15260
rect 12356 15258 12380 15260
rect 12436 15258 12460 15260
rect 12516 15258 12522 15260
rect 12276 15206 12278 15258
rect 12458 15206 12460 15258
rect 12214 15204 12220 15206
rect 12276 15204 12300 15206
rect 12356 15204 12380 15206
rect 12436 15204 12460 15206
rect 12516 15204 12522 15206
rect 12214 15184 12522 15204
rect 12214 14172 12522 14192
rect 12214 14170 12220 14172
rect 12276 14170 12300 14172
rect 12356 14170 12380 14172
rect 12436 14170 12460 14172
rect 12516 14170 12522 14172
rect 12276 14118 12278 14170
rect 12458 14118 12460 14170
rect 12214 14116 12220 14118
rect 12276 14116 12300 14118
rect 12356 14116 12380 14118
rect 12436 14116 12460 14118
rect 12516 14116 12522 14118
rect 12214 14096 12522 14116
rect 12214 13084 12522 13104
rect 12214 13082 12220 13084
rect 12276 13082 12300 13084
rect 12356 13082 12380 13084
rect 12436 13082 12460 13084
rect 12516 13082 12522 13084
rect 12276 13030 12278 13082
rect 12458 13030 12460 13082
rect 12214 13028 12220 13030
rect 12276 13028 12300 13030
rect 12356 13028 12380 13030
rect 12436 13028 12460 13030
rect 12516 13028 12522 13030
rect 12214 13008 12522 13028
rect 12214 11996 12522 12016
rect 12214 11994 12220 11996
rect 12276 11994 12300 11996
rect 12356 11994 12380 11996
rect 12436 11994 12460 11996
rect 12516 11994 12522 11996
rect 12276 11942 12278 11994
rect 12458 11942 12460 11994
rect 12214 11940 12220 11942
rect 12276 11940 12300 11942
rect 12356 11940 12380 11942
rect 12436 11940 12460 11942
rect 12516 11940 12522 11942
rect 12214 11920 12522 11940
rect 12214 10908 12522 10928
rect 12214 10906 12220 10908
rect 12276 10906 12300 10908
rect 12356 10906 12380 10908
rect 12436 10906 12460 10908
rect 12516 10906 12522 10908
rect 12276 10854 12278 10906
rect 12458 10854 12460 10906
rect 12214 10852 12220 10854
rect 12276 10852 12300 10854
rect 12356 10852 12380 10854
rect 12436 10852 12460 10854
rect 12516 10852 12522 10854
rect 12214 10832 12522 10852
rect 12214 9820 12522 9840
rect 12214 9818 12220 9820
rect 12276 9818 12300 9820
rect 12356 9818 12380 9820
rect 12436 9818 12460 9820
rect 12516 9818 12522 9820
rect 12276 9766 12278 9818
rect 12458 9766 12460 9818
rect 12214 9764 12220 9766
rect 12276 9764 12300 9766
rect 12356 9764 12380 9766
rect 12436 9764 12460 9766
rect 12516 9764 12522 9766
rect 12214 9744 12522 9764
rect 12214 8732 12522 8752
rect 12214 8730 12220 8732
rect 12276 8730 12300 8732
rect 12356 8730 12380 8732
rect 12436 8730 12460 8732
rect 12516 8730 12522 8732
rect 12276 8678 12278 8730
rect 12458 8678 12460 8730
rect 12214 8676 12220 8678
rect 12276 8676 12300 8678
rect 12356 8676 12380 8678
rect 12436 8676 12460 8678
rect 12516 8676 12522 8678
rect 12214 8656 12522 8676
rect 12214 7644 12522 7664
rect 12214 7642 12220 7644
rect 12276 7642 12300 7644
rect 12356 7642 12380 7644
rect 12436 7642 12460 7644
rect 12516 7642 12522 7644
rect 12276 7590 12278 7642
rect 12458 7590 12460 7642
rect 12214 7588 12220 7590
rect 12276 7588 12300 7590
rect 12356 7588 12380 7590
rect 12436 7588 12460 7590
rect 12516 7588 12522 7590
rect 12214 7568 12522 7588
rect 12214 6556 12522 6576
rect 12214 6554 12220 6556
rect 12276 6554 12300 6556
rect 12356 6554 12380 6556
rect 12436 6554 12460 6556
rect 12516 6554 12522 6556
rect 12276 6502 12278 6554
rect 12458 6502 12460 6554
rect 12214 6500 12220 6502
rect 12276 6500 12300 6502
rect 12356 6500 12380 6502
rect 12436 6500 12460 6502
rect 12516 6500 12522 6502
rect 12214 6480 12522 6500
rect 12214 5468 12522 5488
rect 12214 5466 12220 5468
rect 12276 5466 12300 5468
rect 12356 5466 12380 5468
rect 12436 5466 12460 5468
rect 12516 5466 12522 5468
rect 12276 5414 12278 5466
rect 12458 5414 12460 5466
rect 12214 5412 12220 5414
rect 12276 5412 12300 5414
rect 12356 5412 12380 5414
rect 12436 5412 12460 5414
rect 12516 5412 12522 5414
rect 12214 5392 12522 5412
rect 9864 4616 9916 4622
rect 9864 4558 9916 4564
rect 10508 4616 10560 4622
rect 10508 4558 10560 4564
rect 9772 3936 9824 3942
rect 9772 3878 9824 3884
rect 9784 3602 9812 3878
rect 9772 3596 9824 3602
rect 9772 3538 9824 3544
rect 8944 3528 8996 3534
rect 8944 3470 8996 3476
rect 9312 3392 9364 3398
rect 9312 3334 9364 3340
rect 9324 2514 9352 3334
rect 9876 3126 9904 4558
rect 10520 3670 10548 4558
rect 12214 4380 12522 4400
rect 12214 4378 12220 4380
rect 12276 4378 12300 4380
rect 12356 4378 12380 4380
rect 12436 4378 12460 4380
rect 12516 4378 12522 4380
rect 12276 4326 12278 4378
rect 12458 4326 12460 4378
rect 12214 4324 12220 4326
rect 12276 4324 12300 4326
rect 12356 4324 12380 4326
rect 12436 4324 12460 4326
rect 12516 4324 12522 4326
rect 12214 4304 12522 4324
rect 13832 4146 13860 22066
rect 13820 4140 13872 4146
rect 13820 4082 13872 4088
rect 10508 3664 10560 3670
rect 10508 3606 10560 3612
rect 9956 3596 10008 3602
rect 9956 3538 10008 3544
rect 9864 3120 9916 3126
rect 9864 3062 9916 3068
rect 9680 2984 9732 2990
rect 9680 2926 9732 2932
rect 9692 2650 9720 2926
rect 9680 2644 9732 2650
rect 9680 2586 9732 2592
rect 9312 2508 9364 2514
rect 9312 2450 9364 2456
rect 9968 1714 9996 3538
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 10876 2916 10928 2922
rect 10876 2858 10928 2864
rect 10888 2514 10916 2858
rect 10980 2582 11008 3470
rect 11980 3460 12032 3466
rect 11980 3402 12032 3408
rect 11992 3058 12020 3402
rect 12214 3292 12522 3312
rect 12214 3290 12220 3292
rect 12276 3290 12300 3292
rect 12356 3290 12380 3292
rect 12436 3290 12460 3292
rect 12516 3290 12522 3292
rect 12276 3238 12278 3290
rect 12458 3238 12460 3290
rect 12214 3236 12220 3238
rect 12276 3236 12300 3238
rect 12356 3236 12380 3238
rect 12436 3236 12460 3238
rect 12516 3236 12522 3238
rect 12214 3216 12522 3236
rect 11980 3052 12032 3058
rect 11980 2994 12032 3000
rect 13176 2984 13228 2990
rect 13176 2926 13228 2932
rect 13544 2984 13596 2990
rect 13544 2926 13596 2932
rect 12440 2848 12492 2854
rect 12440 2790 12492 2796
rect 10968 2576 11020 2582
rect 10968 2518 11020 2524
rect 10324 2508 10376 2514
rect 10324 2450 10376 2456
rect 10876 2508 10928 2514
rect 10876 2450 10928 2456
rect 9692 1686 9996 1714
rect 9692 800 9720 1686
rect 10336 800 10364 2450
rect 12452 2446 12480 2790
rect 13188 2650 13216 2926
rect 13176 2644 13228 2650
rect 13176 2586 13228 2592
rect 12440 2440 12492 2446
rect 12440 2382 12492 2388
rect 12214 2204 12522 2224
rect 12214 2202 12220 2204
rect 12276 2202 12300 2204
rect 12356 2202 12380 2204
rect 12436 2202 12460 2204
rect 12516 2202 12522 2204
rect 12276 2150 12278 2202
rect 12458 2150 12460 2202
rect 12214 2148 12220 2150
rect 12276 2148 12300 2150
rect 12356 2148 12380 2150
rect 12436 2148 12460 2150
rect 12516 2148 12522 2150
rect 12214 2128 12522 2148
rect 13556 800 13584 2926
rect 14108 2446 14136 32535
rect 14200 31657 14228 33934
rect 14292 32609 14320 35006
rect 14384 34950 14412 35550
rect 14464 35488 14516 35494
rect 14462 35456 14464 35465
rect 14516 35456 14518 35465
rect 14462 35391 14518 35400
rect 14568 35057 14596 36654
rect 14648 35080 14700 35086
rect 14554 35048 14610 35057
rect 14648 35022 14700 35028
rect 14554 34983 14610 34992
rect 14372 34944 14424 34950
rect 14372 34886 14424 34892
rect 14556 34944 14608 34950
rect 14556 34886 14608 34892
rect 14462 34640 14518 34649
rect 14568 34610 14596 34886
rect 14462 34575 14518 34584
rect 14556 34604 14608 34610
rect 14476 34542 14504 34575
rect 14556 34546 14608 34552
rect 14464 34536 14516 34542
rect 14464 34478 14516 34484
rect 14660 34184 14688 35022
rect 14752 34610 14780 40666
rect 14844 38894 14872 41200
rect 16028 40520 16080 40526
rect 15290 40488 15346 40497
rect 16028 40462 16080 40468
rect 15290 40423 15346 40432
rect 15384 40452 15436 40458
rect 14924 39432 14976 39438
rect 15200 39432 15252 39438
rect 14924 39374 14976 39380
rect 15120 39392 15200 39420
rect 14936 39098 14964 39374
rect 14924 39092 14976 39098
rect 14924 39034 14976 39040
rect 14832 38888 14884 38894
rect 14832 38830 14884 38836
rect 14936 38740 14964 39034
rect 15120 38894 15148 39392
rect 15200 39374 15252 39380
rect 15200 39296 15252 39302
rect 15200 39238 15252 39244
rect 15212 39098 15240 39238
rect 15200 39092 15252 39098
rect 15200 39034 15252 39040
rect 15108 38888 15160 38894
rect 15108 38830 15160 38836
rect 14844 38712 14964 38740
rect 14740 34604 14792 34610
rect 14740 34546 14792 34552
rect 14660 34156 14780 34184
rect 14554 34096 14610 34105
rect 14554 34031 14556 34040
rect 14608 34031 14610 34040
rect 14556 34002 14608 34008
rect 14648 33992 14700 33998
rect 14648 33934 14700 33940
rect 14464 33856 14516 33862
rect 14464 33798 14516 33804
rect 14554 33824 14610 33833
rect 14476 33697 14504 33798
rect 14554 33759 14610 33768
rect 14462 33688 14518 33697
rect 14462 33623 14518 33632
rect 14464 33584 14516 33590
rect 14464 33526 14516 33532
rect 14476 33425 14504 33526
rect 14568 33522 14596 33759
rect 14556 33516 14608 33522
rect 14556 33458 14608 33464
rect 14660 33425 14688 33934
rect 14462 33416 14518 33425
rect 14372 33380 14424 33386
rect 14646 33416 14702 33425
rect 14462 33351 14518 33360
rect 14556 33380 14608 33386
rect 14372 33322 14424 33328
rect 14646 33351 14702 33360
rect 14556 33322 14608 33328
rect 14278 32600 14334 32609
rect 14278 32535 14334 32544
rect 14384 31822 14412 33322
rect 14568 32910 14596 33322
rect 14752 32978 14780 34156
rect 14740 32972 14792 32978
rect 14740 32914 14792 32920
rect 14464 32904 14516 32910
rect 14464 32846 14516 32852
rect 14556 32904 14608 32910
rect 14556 32846 14608 32852
rect 14476 32434 14504 32846
rect 14554 32600 14610 32609
rect 14554 32535 14610 32544
rect 14568 32502 14596 32535
rect 14556 32496 14608 32502
rect 14556 32438 14608 32444
rect 14648 32496 14700 32502
rect 14648 32438 14700 32444
rect 14464 32428 14516 32434
rect 14464 32370 14516 32376
rect 14660 32348 14688 32438
rect 14568 32320 14688 32348
rect 14568 32230 14596 32320
rect 14844 32280 14872 38712
rect 15016 38208 15068 38214
rect 15016 38150 15068 38156
rect 15108 38208 15160 38214
rect 15108 38150 15160 38156
rect 15028 37942 15056 38150
rect 15016 37936 15068 37942
rect 15016 37878 15068 37884
rect 14924 37800 14976 37806
rect 14924 37742 14976 37748
rect 14936 36174 14964 37742
rect 15016 37188 15068 37194
rect 15016 37130 15068 37136
rect 15028 36417 15056 37130
rect 15014 36408 15070 36417
rect 15014 36343 15070 36352
rect 14924 36168 14976 36174
rect 14924 36110 14976 36116
rect 15016 36032 15068 36038
rect 15016 35974 15068 35980
rect 14924 35624 14976 35630
rect 14924 35566 14976 35572
rect 14936 35494 14964 35566
rect 14924 35488 14976 35494
rect 14924 35430 14976 35436
rect 15028 35290 15056 35974
rect 15016 35284 15068 35290
rect 15016 35226 15068 35232
rect 14924 35216 14976 35222
rect 14924 35158 14976 35164
rect 14936 34474 14964 35158
rect 15014 35048 15070 35057
rect 15014 34983 15070 34992
rect 15028 34746 15056 34983
rect 15016 34740 15068 34746
rect 15016 34682 15068 34688
rect 15016 34604 15068 34610
rect 15016 34546 15068 34552
rect 14924 34468 14976 34474
rect 14924 34410 14976 34416
rect 14922 34096 14978 34105
rect 14922 34031 14978 34040
rect 14936 32910 14964 34031
rect 14924 32904 14976 32910
rect 14924 32846 14976 32852
rect 14924 32496 14976 32502
rect 14924 32438 14976 32444
rect 14844 32252 14880 32280
rect 14556 32224 14608 32230
rect 14852 32178 14880 32252
rect 14936 32201 14964 32438
rect 15028 32348 15056 34546
rect 14997 32320 15056 32348
rect 15120 32348 15148 38150
rect 15200 36780 15252 36786
rect 15200 36722 15252 36728
rect 15212 36689 15240 36722
rect 15198 36680 15254 36689
rect 15198 36615 15254 36624
rect 15304 36360 15332 40423
rect 15384 40394 15436 40400
rect 15212 36332 15332 36360
rect 15212 36106 15240 36332
rect 15292 36168 15344 36174
rect 15292 36110 15344 36116
rect 15200 36100 15252 36106
rect 15200 36042 15252 36048
rect 15304 35698 15332 36110
rect 15292 35692 15344 35698
rect 15292 35634 15344 35640
rect 15200 35216 15252 35222
rect 15200 35158 15252 35164
rect 15212 34678 15240 35158
rect 15292 35080 15344 35086
rect 15292 35022 15344 35028
rect 15200 34672 15252 34678
rect 15200 34614 15252 34620
rect 15304 34474 15332 35022
rect 15200 34468 15252 34474
rect 15200 34410 15252 34416
rect 15292 34468 15344 34474
rect 15292 34410 15344 34416
rect 15212 32842 15240 34410
rect 15304 34105 15332 34410
rect 15290 34096 15346 34105
rect 15290 34031 15346 34040
rect 15396 33946 15424 40394
rect 15844 40248 15896 40254
rect 15844 40190 15896 40196
rect 15660 39364 15712 39370
rect 15660 39306 15712 39312
rect 15568 39296 15620 39302
rect 15568 39238 15620 39244
rect 15580 38654 15608 39238
rect 15488 38626 15608 38654
rect 15488 36174 15516 38626
rect 15672 38418 15700 39306
rect 15752 38888 15804 38894
rect 15752 38830 15804 38836
rect 15660 38412 15712 38418
rect 15660 38354 15712 38360
rect 15568 37664 15620 37670
rect 15764 37618 15792 38830
rect 15568 37606 15620 37612
rect 15580 36224 15608 37606
rect 15672 37590 15792 37618
rect 15672 37398 15700 37590
rect 15750 37496 15806 37505
rect 15750 37431 15806 37440
rect 15856 37448 15884 40190
rect 15936 40112 15988 40118
rect 15936 40054 15988 40060
rect 15948 37874 15976 40054
rect 16040 37874 16068 40462
rect 16132 39794 16160 41200
rect 16670 40216 16726 40225
rect 16670 40151 16726 40160
rect 16132 39766 16252 39794
rect 16120 39364 16172 39370
rect 16120 39306 16172 39312
rect 16132 39030 16160 39306
rect 16120 39024 16172 39030
rect 16120 38966 16172 38972
rect 16224 38654 16252 39766
rect 16396 39636 16448 39642
rect 16396 39578 16448 39584
rect 16304 39568 16356 39574
rect 16304 39510 16356 39516
rect 16132 38626 16252 38654
rect 16132 38418 16160 38626
rect 16316 38536 16344 39510
rect 16408 39302 16436 39578
rect 16684 39506 16712 40151
rect 17038 39944 17094 39953
rect 17038 39879 17094 39888
rect 17052 39545 17080 39879
rect 17316 39636 17368 39642
rect 17316 39578 17368 39584
rect 16854 39536 16910 39545
rect 16672 39500 16724 39506
rect 16854 39471 16910 39480
rect 17038 39536 17094 39545
rect 17038 39471 17094 39480
rect 16672 39442 16724 39448
rect 16580 39364 16632 39370
rect 16580 39306 16632 39312
rect 16396 39296 16448 39302
rect 16396 39238 16448 39244
rect 16488 39296 16540 39302
rect 16488 39238 16540 39244
rect 16500 38894 16528 39238
rect 16488 38888 16540 38894
rect 16488 38830 16540 38836
rect 16592 38729 16620 39306
rect 16868 39273 16896 39471
rect 17328 39370 17356 39578
rect 17420 39506 17448 41200
rect 17682 40216 17738 40225
rect 17682 40151 17738 40160
rect 17498 39672 17554 39681
rect 17498 39607 17554 39616
rect 17512 39506 17540 39607
rect 17408 39500 17460 39506
rect 17408 39442 17460 39448
rect 17500 39500 17552 39506
rect 17500 39442 17552 39448
rect 17316 39364 17368 39370
rect 17316 39306 17368 39312
rect 16670 39264 16726 39273
rect 16854 39264 16910 39273
rect 16726 39222 16804 39250
rect 16670 39199 16726 39208
rect 16776 39080 16804 39222
rect 16854 39199 16910 39208
rect 16776 39052 17264 39080
rect 17132 38956 17184 38962
rect 17132 38898 17184 38904
rect 16948 38888 17000 38894
rect 16948 38830 17000 38836
rect 17038 38856 17094 38865
rect 16578 38720 16634 38729
rect 16578 38655 16634 38664
rect 16960 38654 16988 38830
rect 17038 38791 17094 38800
rect 16224 38508 16344 38536
rect 16684 38626 16988 38654
rect 16116 38412 16168 38418
rect 16116 38354 16168 38360
rect 15936 37868 15988 37874
rect 15936 37810 15988 37816
rect 16028 37868 16080 37874
rect 16028 37810 16080 37816
rect 16224 37618 16252 38508
rect 16684 38196 16712 38626
rect 16856 38344 16908 38350
rect 16408 38168 16712 38196
rect 16776 38304 16856 38332
rect 16302 38040 16358 38049
rect 16302 37975 16358 37984
rect 16040 37590 16252 37618
rect 15764 37398 15792 37431
rect 15856 37420 15976 37448
rect 15660 37392 15712 37398
rect 15660 37334 15712 37340
rect 15752 37392 15804 37398
rect 15752 37334 15804 37340
rect 15844 37256 15896 37262
rect 15844 37198 15896 37204
rect 15856 36961 15884 37198
rect 15842 36952 15898 36961
rect 15842 36887 15898 36896
rect 15948 36786 15976 37420
rect 16040 36786 16068 37590
rect 16316 37505 16344 37975
rect 16302 37496 16358 37505
rect 16302 37431 16358 37440
rect 16212 37392 16264 37398
rect 16408 37380 16436 38168
rect 16486 38040 16542 38049
rect 16486 37975 16542 37984
rect 16500 37466 16528 37975
rect 16776 37874 16804 38304
rect 16856 38286 16908 38292
rect 16948 38276 17000 38282
rect 16948 38218 17000 38224
rect 16960 37874 16988 38218
rect 16764 37868 16816 37874
rect 16764 37810 16816 37816
rect 16948 37868 17000 37874
rect 16948 37810 17000 37816
rect 16580 37800 16632 37806
rect 16580 37742 16632 37748
rect 16488 37460 16540 37466
rect 16488 37402 16540 37408
rect 16264 37352 16436 37380
rect 16212 37334 16264 37340
rect 16224 37194 16252 37334
rect 16212 37188 16264 37194
rect 16212 37130 16264 37136
rect 16396 37188 16448 37194
rect 16396 37130 16448 37136
rect 16118 36952 16174 36961
rect 16118 36887 16174 36896
rect 15936 36780 15988 36786
rect 15936 36722 15988 36728
rect 16028 36780 16080 36786
rect 16028 36722 16080 36728
rect 15658 36680 15714 36689
rect 15658 36615 15714 36624
rect 15672 36417 15700 36615
rect 15658 36408 15714 36417
rect 15934 36408 15990 36417
rect 15658 36343 15714 36352
rect 15844 36372 15896 36378
rect 15896 36352 15934 36360
rect 16132 36378 16160 36887
rect 16408 36854 16436 37130
rect 16396 36848 16448 36854
rect 16396 36790 16448 36796
rect 16304 36780 16356 36786
rect 16304 36722 16356 36728
rect 16316 36689 16344 36722
rect 16396 36712 16448 36718
rect 16302 36680 16358 36689
rect 16592 36700 16620 37742
rect 17052 37618 17080 38791
rect 17144 38350 17172 38898
rect 17236 38826 17264 39052
rect 17224 38820 17276 38826
rect 17224 38762 17276 38768
rect 17316 38752 17368 38758
rect 17696 38729 17724 40151
rect 18064 40066 18092 41200
rect 18604 40792 18656 40798
rect 18604 40734 18656 40740
rect 18510 40624 18566 40633
rect 18510 40559 18566 40568
rect 18064 40038 18276 40066
rect 17776 39840 17828 39846
rect 17776 39782 17828 39788
rect 17788 38944 17816 39782
rect 17846 39740 18154 39760
rect 17846 39738 17852 39740
rect 17908 39738 17932 39740
rect 17988 39738 18012 39740
rect 18068 39738 18092 39740
rect 18148 39738 18154 39740
rect 17908 39686 17910 39738
rect 18090 39686 18092 39738
rect 17846 39684 17852 39686
rect 17908 39684 17932 39686
rect 17988 39684 18012 39686
rect 18068 39684 18092 39686
rect 18148 39684 18154 39686
rect 17846 39664 18154 39684
rect 18052 39432 18104 39438
rect 18052 39374 18104 39380
rect 18064 39030 18092 39374
rect 18052 39024 18104 39030
rect 18052 38966 18104 38972
rect 17788 38916 18000 38944
rect 17972 38740 18000 38916
rect 18248 38894 18276 40038
rect 18326 39808 18382 39817
rect 18326 39743 18382 39752
rect 18340 39137 18368 39743
rect 18326 39128 18382 39137
rect 18326 39063 18382 39072
rect 18236 38888 18288 38894
rect 18328 38888 18380 38894
rect 18236 38830 18288 38836
rect 18326 38856 18328 38865
rect 18524 38865 18552 40559
rect 18380 38856 18382 38865
rect 18326 38791 18382 38800
rect 18510 38856 18566 38865
rect 18510 38791 18566 38800
rect 17316 38694 17368 38700
rect 17406 38720 17462 38729
rect 17132 38344 17184 38350
rect 17132 38286 17184 38292
rect 16868 37590 17080 37618
rect 16868 37505 16896 37590
rect 16854 37496 16910 37505
rect 16854 37431 16856 37440
rect 16908 37431 16910 37440
rect 17038 37496 17094 37505
rect 17038 37431 17094 37440
rect 16856 37402 16908 37408
rect 16868 37371 16896 37402
rect 17052 37262 17080 37431
rect 17040 37256 17092 37262
rect 17040 37198 17092 37204
rect 16672 37120 16724 37126
rect 16672 37062 16724 37068
rect 16684 36922 16712 37062
rect 16672 36916 16724 36922
rect 16672 36858 16724 36864
rect 17040 36848 17092 36854
rect 16960 36808 17040 36836
rect 16672 36712 16724 36718
rect 16396 36654 16448 36660
rect 16486 36680 16542 36689
rect 16302 36615 16358 36624
rect 16408 36417 16436 36654
rect 16592 36672 16672 36700
rect 16960 36700 16988 36808
rect 17040 36790 17092 36796
rect 17144 36700 17172 38286
rect 17224 37868 17276 37874
rect 17224 37810 17276 37816
rect 17236 37398 17264 37810
rect 17328 37505 17356 38694
rect 17682 38720 17738 38729
rect 17462 38678 17632 38706
rect 17406 38655 17462 38664
rect 17408 38412 17460 38418
rect 17408 38354 17460 38360
rect 17314 37496 17370 37505
rect 17314 37431 17370 37440
rect 17224 37392 17276 37398
rect 17224 37334 17276 37340
rect 17420 37274 17448 38354
rect 17604 38332 17632 38678
rect 17972 38712 18368 38740
rect 18340 38706 18368 38712
rect 18340 38678 18460 38706
rect 17682 38655 17738 38664
rect 17846 38652 18154 38672
rect 17846 38650 17852 38652
rect 17908 38650 17932 38652
rect 17988 38650 18012 38652
rect 18068 38650 18092 38652
rect 18148 38650 18154 38652
rect 17908 38598 17910 38650
rect 18090 38598 18092 38650
rect 17846 38596 17852 38598
rect 17908 38596 17932 38598
rect 17988 38596 18012 38598
rect 18068 38596 18092 38598
rect 18148 38596 18154 38598
rect 17846 38576 18154 38596
rect 18432 38554 18460 38678
rect 18420 38548 18472 38554
rect 18420 38490 18472 38496
rect 17684 38480 17736 38486
rect 17736 38440 17908 38468
rect 17684 38422 17736 38428
rect 17880 38350 17908 38440
rect 18144 38412 18196 38418
rect 18144 38354 18196 38360
rect 17868 38344 17920 38350
rect 17604 38304 17724 38332
rect 17696 37806 17724 38304
rect 17868 38286 17920 38292
rect 18156 37942 18184 38354
rect 18144 37936 18196 37942
rect 18144 37878 18196 37884
rect 18236 37936 18288 37942
rect 18236 37878 18288 37884
rect 18248 37806 18276 37878
rect 18328 37868 18380 37874
rect 18328 37810 18380 37816
rect 17684 37800 17736 37806
rect 17684 37742 17736 37748
rect 18236 37800 18288 37806
rect 18236 37742 18288 37748
rect 17776 37664 17828 37670
rect 17682 37632 17738 37641
rect 18340 37641 18368 37810
rect 18512 37800 18564 37806
rect 18512 37742 18564 37748
rect 17776 37606 17828 37612
rect 18326 37632 18382 37641
rect 17682 37567 17738 37576
rect 17590 37496 17646 37505
rect 17500 37460 17552 37466
rect 17590 37431 17646 37440
rect 17500 37402 17552 37408
rect 17328 37246 17448 37274
rect 17512 37262 17540 37402
rect 17500 37256 17552 37262
rect 17328 37194 17356 37246
rect 17500 37198 17552 37204
rect 17316 37188 17368 37194
rect 17316 37130 17368 37136
rect 17604 37126 17632 37431
rect 17696 37398 17724 37567
rect 17684 37392 17736 37398
rect 17684 37334 17736 37340
rect 17592 37120 17644 37126
rect 17592 37062 17644 37068
rect 17224 36848 17276 36854
rect 17224 36790 17276 36796
rect 16724 36672 16988 36700
rect 17052 36672 17172 36700
rect 16672 36654 16724 36660
rect 16486 36615 16488 36624
rect 16540 36615 16542 36624
rect 16488 36586 16540 36592
rect 16210 36408 16266 36417
rect 15896 36343 15990 36352
rect 16120 36372 16172 36378
rect 15896 36332 15976 36343
rect 15844 36314 15896 36320
rect 16210 36343 16212 36352
rect 16120 36314 16172 36320
rect 16264 36343 16266 36352
rect 16394 36408 16450 36417
rect 16394 36343 16450 36352
rect 16948 36372 17000 36378
rect 16212 36314 16264 36320
rect 16948 36314 17000 36320
rect 16396 36304 16448 36310
rect 16396 36246 16448 36252
rect 15580 36196 16068 36224
rect 15476 36168 15528 36174
rect 15476 36110 15528 36116
rect 15568 36100 15620 36106
rect 15568 36042 15620 36048
rect 15476 35148 15528 35154
rect 15476 35090 15528 35096
rect 15488 35057 15516 35090
rect 15474 35048 15530 35057
rect 15474 34983 15530 34992
rect 15474 34776 15530 34785
rect 15474 34711 15476 34720
rect 15528 34711 15530 34720
rect 15476 34682 15528 34688
rect 15476 34128 15528 34134
rect 15476 34070 15528 34076
rect 15488 33998 15516 34070
rect 15304 33918 15424 33946
rect 15476 33992 15528 33998
rect 15476 33934 15528 33940
rect 15304 33436 15332 33918
rect 15580 33674 15608 36042
rect 15936 35692 15988 35698
rect 15936 35634 15988 35640
rect 15752 35624 15804 35630
rect 15752 35566 15804 35572
rect 15764 35290 15792 35566
rect 15948 35465 15976 35634
rect 15934 35456 15990 35465
rect 15934 35391 15990 35400
rect 15752 35284 15804 35290
rect 15752 35226 15804 35232
rect 15936 35012 15988 35018
rect 15764 34972 15936 35000
rect 15764 34610 15792 34972
rect 15936 34954 15988 34960
rect 15752 34604 15804 34610
rect 15752 34546 15804 34552
rect 15752 34196 15804 34202
rect 15752 34138 15804 34144
rect 15936 34196 15988 34202
rect 15936 34138 15988 34144
rect 15764 34105 15792 34138
rect 15750 34096 15806 34105
rect 15750 34031 15806 34040
rect 15948 33998 15976 34138
rect 15936 33992 15988 33998
rect 15936 33934 15988 33940
rect 16040 33946 16068 36196
rect 16302 35728 16358 35737
rect 16212 35692 16264 35698
rect 16264 35672 16302 35680
rect 16408 35698 16436 36246
rect 16500 36230 16896 36258
rect 16960 36242 16988 36314
rect 16264 35663 16358 35672
rect 16396 35692 16448 35698
rect 16264 35652 16344 35663
rect 16212 35634 16264 35640
rect 16396 35634 16448 35640
rect 16500 35630 16528 36230
rect 16764 36168 16816 36174
rect 16764 36110 16816 36116
rect 16776 35834 16804 36110
rect 16868 36088 16896 36230
rect 16948 36236 17000 36242
rect 16948 36178 17000 36184
rect 16948 36100 17000 36106
rect 16868 36060 16948 36088
rect 16948 36042 17000 36048
rect 16764 35828 16816 35834
rect 16764 35770 16816 35776
rect 16488 35624 16540 35630
rect 16488 35566 16540 35572
rect 16672 35624 16724 35630
rect 16672 35566 16724 35572
rect 16580 35216 16632 35222
rect 16580 35158 16632 35164
rect 16592 35018 16620 35158
rect 16684 35154 16712 35566
rect 16776 35465 16804 35770
rect 17052 35544 17080 36672
rect 17236 36106 17264 36790
rect 17788 36768 17816 37606
rect 17846 37564 18154 37584
rect 18326 37567 18382 37576
rect 17846 37562 17852 37564
rect 17908 37562 17932 37564
rect 17988 37562 18012 37564
rect 18068 37562 18092 37564
rect 18148 37562 18154 37564
rect 17908 37510 17910 37562
rect 18090 37510 18092 37562
rect 17846 37508 17852 37510
rect 17908 37508 17932 37510
rect 17988 37508 18012 37510
rect 18068 37508 18092 37510
rect 18148 37508 18154 37510
rect 17846 37488 18154 37508
rect 18234 37496 18290 37505
rect 18234 37431 18236 37440
rect 18288 37431 18290 37440
rect 18328 37460 18380 37466
rect 18236 37402 18288 37408
rect 18328 37402 18380 37408
rect 18340 37330 18368 37402
rect 18328 37324 18380 37330
rect 18328 37266 18380 37272
rect 18328 37120 18380 37126
rect 18328 37062 18380 37068
rect 17328 36740 17816 36768
rect 18236 36780 18288 36786
rect 17328 36310 17356 36740
rect 18236 36722 18288 36728
rect 17776 36644 17828 36650
rect 17776 36586 17828 36592
rect 17682 36544 17738 36553
rect 17788 36530 17816 36586
rect 18248 36553 18276 36722
rect 17738 36502 17816 36530
rect 18234 36544 18290 36553
rect 17682 36479 17738 36488
rect 17846 36476 18154 36496
rect 18234 36479 18290 36488
rect 17846 36474 17852 36476
rect 17908 36474 17932 36476
rect 17988 36474 18012 36476
rect 18068 36474 18092 36476
rect 18148 36474 18154 36476
rect 17908 36422 17910 36474
rect 18090 36422 18092 36474
rect 17846 36420 17852 36422
rect 17908 36420 17932 36422
rect 17988 36420 18012 36422
rect 18068 36420 18092 36422
rect 18148 36420 18154 36422
rect 17682 36408 17738 36417
rect 17846 36400 18154 36420
rect 18340 36417 18368 37062
rect 18524 36786 18552 37742
rect 18616 37618 18644 40734
rect 18708 38457 18736 41200
rect 19892 40724 19944 40730
rect 19892 40666 19944 40672
rect 19154 40352 19210 40361
rect 19154 40287 19210 40296
rect 18880 39908 18932 39914
rect 18880 39850 18932 39856
rect 18972 39908 19024 39914
rect 18972 39850 19024 39856
rect 18788 39364 18840 39370
rect 18788 39306 18840 39312
rect 18800 39098 18828 39306
rect 18788 39092 18840 39098
rect 18788 39034 18840 39040
rect 18786 38992 18842 39001
rect 18892 38962 18920 39850
rect 18984 39302 19012 39850
rect 19064 39636 19116 39642
rect 19064 39578 19116 39584
rect 18972 39296 19024 39302
rect 18972 39238 19024 39244
rect 18786 38927 18842 38936
rect 18880 38956 18932 38962
rect 18800 38729 18828 38927
rect 18880 38898 18932 38904
rect 18786 38720 18842 38729
rect 18786 38655 18842 38664
rect 18788 38548 18840 38554
rect 18788 38490 18840 38496
rect 18694 38448 18750 38457
rect 18694 38383 18750 38392
rect 18800 37874 18828 38490
rect 19076 38350 19104 39578
rect 19168 38350 19196 40287
rect 19904 40254 19932 40666
rect 19800 40248 19852 40254
rect 19800 40190 19852 40196
rect 19892 40248 19944 40254
rect 19892 40190 19944 40196
rect 19616 40112 19668 40118
rect 19616 40054 19668 40060
rect 19248 40044 19300 40050
rect 19248 39986 19300 39992
rect 19260 38434 19288 39986
rect 19338 39672 19394 39681
rect 19338 39607 19394 39616
rect 19352 39438 19380 39607
rect 19340 39432 19392 39438
rect 19340 39374 19392 39380
rect 19432 39364 19484 39370
rect 19432 39306 19484 39312
rect 19340 38820 19392 38826
rect 19340 38762 19392 38768
rect 19352 38554 19380 38762
rect 19340 38548 19392 38554
rect 19340 38490 19392 38496
rect 19260 38406 19380 38434
rect 19352 38350 19380 38406
rect 19064 38344 19116 38350
rect 19064 38286 19116 38292
rect 19156 38344 19208 38350
rect 19156 38286 19208 38292
rect 19340 38344 19392 38350
rect 19340 38286 19392 38292
rect 18788 37868 18840 37874
rect 18788 37810 18840 37816
rect 18616 37590 18920 37618
rect 18696 37460 18748 37466
rect 18696 37402 18748 37408
rect 18604 37256 18656 37262
rect 18604 37198 18656 37204
rect 18512 36780 18564 36786
rect 18512 36722 18564 36728
rect 18420 36576 18472 36582
rect 18420 36518 18472 36524
rect 18326 36408 18382 36417
rect 17738 36366 17816 36394
rect 17682 36343 17738 36352
rect 17316 36304 17368 36310
rect 17368 36264 17448 36292
rect 17316 36246 17368 36252
rect 17132 36100 17184 36106
rect 17132 36042 17184 36048
rect 17224 36100 17276 36106
rect 17224 36042 17276 36048
rect 17144 35766 17172 36042
rect 17132 35760 17184 35766
rect 17132 35702 17184 35708
rect 16960 35516 17080 35544
rect 16762 35456 16818 35465
rect 16960 35442 16988 35516
rect 16762 35391 16818 35400
rect 16868 35414 16988 35442
rect 17038 35456 17094 35465
rect 16672 35148 16724 35154
rect 16672 35090 16724 35096
rect 16580 35012 16632 35018
rect 16580 34954 16632 34960
rect 16488 34672 16540 34678
rect 16488 34614 16540 34620
rect 16580 34672 16632 34678
rect 16580 34614 16632 34620
rect 16396 34604 16448 34610
rect 16396 34546 16448 34552
rect 16304 34468 16356 34474
rect 16304 34410 16356 34416
rect 16316 34202 16344 34410
rect 16212 34196 16264 34202
rect 16212 34138 16264 34144
rect 16304 34196 16356 34202
rect 16304 34138 16356 34144
rect 16224 34066 16252 34138
rect 16212 34060 16264 34066
rect 16212 34002 16264 34008
rect 16304 33992 16356 33998
rect 16302 33960 16304 33969
rect 16356 33960 16358 33969
rect 16040 33930 16252 33946
rect 16040 33924 16264 33930
rect 16040 33918 16212 33924
rect 16302 33895 16358 33904
rect 16212 33866 16264 33872
rect 15752 33856 15804 33862
rect 15804 33816 16160 33844
rect 15752 33798 15804 33804
rect 15580 33646 15792 33674
rect 15660 33584 15712 33590
rect 15566 33552 15622 33561
rect 15660 33526 15712 33532
rect 15566 33487 15622 33496
rect 15304 33408 15424 33436
rect 15200 32836 15252 32842
rect 15200 32778 15252 32784
rect 15120 32320 15240 32348
rect 14997 32280 15025 32320
rect 14997 32252 15148 32280
rect 15120 32212 15148 32252
rect 14556 32166 14608 32172
rect 14844 32150 14880 32178
rect 14922 32192 14978 32201
rect 14738 32056 14794 32065
rect 14738 31991 14740 32000
rect 14792 31991 14794 32000
rect 14740 31962 14792 31968
rect 14556 31952 14608 31958
rect 14844 31906 14872 32150
rect 14922 32127 14978 32136
rect 15028 32184 15148 32212
rect 14924 32020 14976 32026
rect 14924 31962 14976 31968
rect 14556 31894 14608 31900
rect 14372 31816 14424 31822
rect 14372 31758 14424 31764
rect 14464 31748 14516 31754
rect 14464 31690 14516 31696
rect 14186 31648 14242 31657
rect 14186 31583 14242 31592
rect 14476 30598 14504 31690
rect 14568 31346 14596 31894
rect 14752 31878 14872 31906
rect 14646 31512 14702 31521
rect 14646 31447 14702 31456
rect 14660 31414 14688 31447
rect 14648 31408 14700 31414
rect 14648 31350 14700 31356
rect 14556 31340 14608 31346
rect 14556 31282 14608 31288
rect 14554 31240 14610 31249
rect 14554 31175 14610 31184
rect 14568 31142 14596 31175
rect 14556 31136 14608 31142
rect 14556 31078 14608 31084
rect 14464 30592 14516 30598
rect 14464 30534 14516 30540
rect 14568 30258 14596 31078
rect 14648 30660 14700 30666
rect 14648 30602 14700 30608
rect 14280 30252 14332 30258
rect 14280 30194 14332 30200
rect 14556 30252 14608 30258
rect 14556 30194 14608 30200
rect 14188 30048 14240 30054
rect 14188 29990 14240 29996
rect 14200 29753 14228 29990
rect 14186 29744 14242 29753
rect 14186 29679 14242 29688
rect 14188 29640 14240 29646
rect 14188 29582 14240 29588
rect 14200 29306 14228 29582
rect 14188 29300 14240 29306
rect 14188 29242 14240 29248
rect 14186 29200 14242 29209
rect 14186 29135 14242 29144
rect 14200 28014 14228 29135
rect 14292 28529 14320 30194
rect 14660 30138 14688 30602
rect 14568 30110 14688 30138
rect 14372 29640 14424 29646
rect 14372 29582 14424 29588
rect 14462 29608 14518 29617
rect 14278 28520 14334 28529
rect 14278 28455 14334 28464
rect 14278 28384 14334 28393
rect 14278 28319 14334 28328
rect 14188 28008 14240 28014
rect 14188 27950 14240 27956
rect 14188 26988 14240 26994
rect 14188 26930 14240 26936
rect 14200 26625 14228 26930
rect 14186 26616 14242 26625
rect 14186 26551 14242 26560
rect 14292 24138 14320 28319
rect 14384 27554 14412 29582
rect 14462 29543 14518 29552
rect 14476 29345 14504 29543
rect 14462 29336 14518 29345
rect 14462 29271 14518 29280
rect 14568 29170 14596 30110
rect 14648 29504 14700 29510
rect 14648 29446 14700 29452
rect 14660 29345 14688 29446
rect 14646 29336 14702 29345
rect 14646 29271 14702 29280
rect 14648 29232 14700 29238
rect 14646 29200 14648 29209
rect 14700 29200 14702 29209
rect 14556 29164 14608 29170
rect 14646 29135 14702 29144
rect 14556 29106 14608 29112
rect 14646 28656 14702 28665
rect 14646 28591 14702 28600
rect 14660 28558 14688 28591
rect 14648 28552 14700 28558
rect 14648 28494 14700 28500
rect 14648 28144 14700 28150
rect 14648 28086 14700 28092
rect 14464 28076 14516 28082
rect 14464 28018 14516 28024
rect 14556 28076 14608 28082
rect 14556 28018 14608 28024
rect 14476 27674 14504 28018
rect 14568 27946 14596 28018
rect 14556 27940 14608 27946
rect 14556 27882 14608 27888
rect 14660 27826 14688 28086
rect 14568 27798 14688 27826
rect 14464 27668 14516 27674
rect 14464 27610 14516 27616
rect 14384 27526 14504 27554
rect 14372 27464 14424 27470
rect 14372 27406 14424 27412
rect 14280 24132 14332 24138
rect 14280 24074 14332 24080
rect 14384 22778 14412 27406
rect 14476 25945 14504 27526
rect 14568 26330 14596 27798
rect 14648 26784 14700 26790
rect 14752 26761 14780 31878
rect 14936 31822 14964 31962
rect 14924 31816 14976 31822
rect 14924 31758 14976 31764
rect 14830 31512 14886 31521
rect 14830 31447 14886 31456
rect 14844 30666 14872 31447
rect 14832 30660 14884 30666
rect 14832 30602 14884 30608
rect 14830 30560 14886 30569
rect 14830 30495 14886 30504
rect 14844 30326 14872 30495
rect 14832 30320 14884 30326
rect 14832 30262 14884 30268
rect 14924 30048 14976 30054
rect 14830 30016 14886 30025
rect 14924 29990 14976 29996
rect 14830 29951 14886 29960
rect 14844 29646 14872 29951
rect 14832 29640 14884 29646
rect 14832 29582 14884 29588
rect 14844 29102 14872 29582
rect 14832 29096 14884 29102
rect 14832 29038 14884 29044
rect 14936 28801 14964 29990
rect 15028 28966 15056 32184
rect 15108 31748 15160 31754
rect 15108 31690 15160 31696
rect 15120 31414 15148 31690
rect 15108 31408 15160 31414
rect 15108 31350 15160 31356
rect 15212 31090 15240 32320
rect 15292 31680 15344 31686
rect 15292 31622 15344 31628
rect 15120 31062 15240 31090
rect 15120 30734 15148 31062
rect 15304 30938 15332 31622
rect 15200 30932 15252 30938
rect 15200 30874 15252 30880
rect 15292 30932 15344 30938
rect 15292 30874 15344 30880
rect 15108 30728 15160 30734
rect 15108 30670 15160 30676
rect 15120 30258 15148 30670
rect 15212 30297 15240 30874
rect 15292 30660 15344 30666
rect 15292 30602 15344 30608
rect 15198 30288 15254 30297
rect 15108 30252 15160 30258
rect 15198 30223 15254 30232
rect 15108 30194 15160 30200
rect 15304 29850 15332 30602
rect 15292 29844 15344 29850
rect 15292 29786 15344 29792
rect 15290 29744 15346 29753
rect 15290 29679 15346 29688
rect 15108 29164 15160 29170
rect 15108 29106 15160 29112
rect 15016 28960 15068 28966
rect 15016 28902 15068 28908
rect 14922 28792 14978 28801
rect 14922 28727 14978 28736
rect 15120 28558 15148 29106
rect 15304 29034 15332 29679
rect 15396 29646 15424 33408
rect 15580 32774 15608 33487
rect 15672 33425 15700 33526
rect 15658 33416 15714 33425
rect 15658 33351 15714 33360
rect 15660 32904 15712 32910
rect 15660 32846 15712 32852
rect 15476 32768 15528 32774
rect 15476 32710 15528 32716
rect 15568 32768 15620 32774
rect 15568 32710 15620 32716
rect 15488 32230 15516 32710
rect 15568 32428 15620 32434
rect 15672 32416 15700 32846
rect 15620 32388 15700 32416
rect 15568 32370 15620 32376
rect 15476 32224 15528 32230
rect 15476 32166 15528 32172
rect 15660 32020 15712 32026
rect 15660 31962 15712 31968
rect 15672 30870 15700 31962
rect 15660 30864 15712 30870
rect 15660 30806 15712 30812
rect 15476 30660 15528 30666
rect 15476 30602 15528 30608
rect 15488 30326 15516 30602
rect 15476 30320 15528 30326
rect 15476 30262 15528 30268
rect 15476 30048 15528 30054
rect 15476 29990 15528 29996
rect 15488 29646 15516 29990
rect 15658 29880 15714 29889
rect 15658 29815 15714 29824
rect 15384 29640 15436 29646
rect 15384 29582 15436 29588
rect 15476 29640 15528 29646
rect 15476 29582 15528 29588
rect 15292 29028 15344 29034
rect 15292 28970 15344 28976
rect 15198 28928 15254 28937
rect 15198 28863 15254 28872
rect 14832 28552 14884 28558
rect 14832 28494 14884 28500
rect 15108 28552 15160 28558
rect 15108 28494 15160 28500
rect 14648 26726 14700 26732
rect 14738 26752 14794 26761
rect 14660 26450 14688 26726
rect 14738 26687 14794 26696
rect 14844 26466 14872 28494
rect 15212 28393 15240 28863
rect 15292 28552 15344 28558
rect 15292 28494 15344 28500
rect 14922 28384 14978 28393
rect 14922 28319 14978 28328
rect 15198 28384 15254 28393
rect 15198 28319 15254 28328
rect 14936 28082 14964 28319
rect 15014 28248 15070 28257
rect 15014 28183 15070 28192
rect 14924 28076 14976 28082
rect 14924 28018 14976 28024
rect 15028 27606 15056 28183
rect 15108 28144 15160 28150
rect 15304 28121 15332 28494
rect 15108 28086 15160 28092
rect 15290 28112 15346 28121
rect 15016 27600 15068 27606
rect 15016 27542 15068 27548
rect 14924 27464 14976 27470
rect 14924 27406 14976 27412
rect 14648 26444 14700 26450
rect 14648 26386 14700 26392
rect 14752 26438 14872 26466
rect 14568 26302 14688 26330
rect 14462 25936 14518 25945
rect 14462 25871 14518 25880
rect 14556 25288 14608 25294
rect 14556 25230 14608 25236
rect 14568 24954 14596 25230
rect 14556 24948 14608 24954
rect 14556 24890 14608 24896
rect 14660 24177 14688 26302
rect 14752 25265 14780 26438
rect 14832 26376 14884 26382
rect 14832 26318 14884 26324
rect 14844 25537 14872 26318
rect 14830 25528 14886 25537
rect 14830 25463 14886 25472
rect 14738 25256 14794 25265
rect 14738 25191 14794 25200
rect 14936 24993 14964 27406
rect 15120 27305 15148 28086
rect 15200 28076 15252 28082
rect 15290 28047 15346 28056
rect 15200 28018 15252 28024
rect 15212 27849 15240 28018
rect 15198 27840 15254 27849
rect 15198 27775 15254 27784
rect 15200 27464 15252 27470
rect 15200 27406 15252 27412
rect 15290 27432 15346 27441
rect 15106 27296 15162 27305
rect 15106 27231 15162 27240
rect 15014 26480 15070 26489
rect 15014 26415 15070 26424
rect 15028 26246 15056 26415
rect 15212 26353 15240 27406
rect 15290 27367 15346 27376
rect 15304 27334 15332 27367
rect 15292 27328 15344 27334
rect 15292 27270 15344 27276
rect 15198 26344 15254 26353
rect 15198 26279 15254 26288
rect 15292 26308 15344 26314
rect 15292 26250 15344 26256
rect 15016 26240 15068 26246
rect 15016 26182 15068 26188
rect 15108 26240 15160 26246
rect 15108 26182 15160 26188
rect 15120 25974 15148 26182
rect 15304 26081 15332 26250
rect 15290 26072 15346 26081
rect 15290 26007 15346 26016
rect 15108 25968 15160 25974
rect 15108 25910 15160 25916
rect 15292 25900 15344 25906
rect 15292 25842 15344 25848
rect 15108 25220 15160 25226
rect 15108 25162 15160 25168
rect 14922 24984 14978 24993
rect 14922 24919 14978 24928
rect 15120 24682 15148 25162
rect 15304 24682 15332 25842
rect 15108 24676 15160 24682
rect 15108 24618 15160 24624
rect 15292 24676 15344 24682
rect 15292 24618 15344 24624
rect 14922 24304 14978 24313
rect 15120 24274 15148 24618
rect 14922 24239 14978 24248
rect 15108 24268 15160 24274
rect 14936 24206 14964 24239
rect 15108 24210 15160 24216
rect 14924 24200 14976 24206
rect 14646 24168 14702 24177
rect 14924 24142 14976 24148
rect 14646 24103 14702 24112
rect 15108 24132 15160 24138
rect 15108 24074 15160 24080
rect 14740 24064 14792 24070
rect 14740 24006 14792 24012
rect 14752 23769 14780 24006
rect 15120 23905 15148 24074
rect 15106 23896 15162 23905
rect 15106 23831 15162 23840
rect 14738 23760 14794 23769
rect 14738 23695 14794 23704
rect 15200 23520 15252 23526
rect 15200 23462 15252 23468
rect 15212 23118 15240 23462
rect 15200 23112 15252 23118
rect 15200 23054 15252 23060
rect 14372 22772 14424 22778
rect 14372 22714 14424 22720
rect 15304 20874 15332 24618
rect 15292 20868 15344 20874
rect 15292 20810 15344 20816
rect 14372 12232 14424 12238
rect 14372 12174 14424 12180
rect 14280 3936 14332 3942
rect 14280 3878 14332 3884
rect 14292 3058 14320 3878
rect 14384 3534 14412 12174
rect 14372 3528 14424 3534
rect 14372 3470 14424 3476
rect 14464 3392 14516 3398
rect 14464 3334 14516 3340
rect 14476 3126 14504 3334
rect 14464 3120 14516 3126
rect 14464 3062 14516 3068
rect 14280 3052 14332 3058
rect 14280 2994 14332 3000
rect 14832 2984 14884 2990
rect 14832 2926 14884 2932
rect 14096 2440 14148 2446
rect 14096 2382 14148 2388
rect 14844 800 14872 2926
rect 15396 2378 15424 29582
rect 15672 29306 15700 29815
rect 15764 29646 15792 33646
rect 15934 33416 15990 33425
rect 15934 33351 15990 33360
rect 15948 33318 15976 33351
rect 15936 33312 15988 33318
rect 15936 33254 15988 33260
rect 16028 33312 16080 33318
rect 16028 33254 16080 33260
rect 15844 32360 15896 32366
rect 15844 32302 15896 32308
rect 15856 31754 15884 32302
rect 16040 32230 16068 33254
rect 16132 32978 16160 33816
rect 16408 33504 16436 34546
rect 16500 34474 16528 34614
rect 16592 34542 16620 34614
rect 16580 34536 16632 34542
rect 16580 34478 16632 34484
rect 16488 34468 16540 34474
rect 16488 34410 16540 34416
rect 16592 34354 16620 34478
rect 16500 34326 16620 34354
rect 16500 33946 16528 34326
rect 16580 34196 16632 34202
rect 16580 34138 16632 34144
rect 16592 34048 16620 34138
rect 16684 34066 16712 35090
rect 16764 34672 16816 34678
rect 16868 34660 16896 35414
rect 17038 35391 17094 35400
rect 16948 35284 17000 35290
rect 16948 35226 17000 35232
rect 16816 34632 16896 34660
rect 16764 34614 16816 34620
rect 16960 34592 16988 35226
rect 17052 35086 17080 35391
rect 17130 35320 17186 35329
rect 17130 35255 17132 35264
rect 17184 35255 17186 35264
rect 17132 35226 17184 35232
rect 17236 35154 17264 36042
rect 17224 35148 17276 35154
rect 17224 35090 17276 35096
rect 17316 35148 17368 35154
rect 17316 35090 17368 35096
rect 17040 35080 17092 35086
rect 17040 35022 17092 35028
rect 17224 35012 17276 35018
rect 17224 34954 17276 34960
rect 17040 34944 17092 34950
rect 17040 34886 17092 34892
rect 17052 34728 17080 34886
rect 17052 34700 17172 34728
rect 17040 34604 17092 34610
rect 16960 34564 17040 34592
rect 17040 34546 17092 34552
rect 17040 34400 17092 34406
rect 17040 34342 17092 34348
rect 17144 34354 17172 34700
rect 17236 34474 17264 34954
rect 17224 34468 17276 34474
rect 17224 34410 17276 34416
rect 17328 34354 17356 35090
rect 17420 34950 17448 36264
rect 17788 36106 17816 36366
rect 18326 36343 18382 36352
rect 17776 36100 17828 36106
rect 17776 36042 17828 36048
rect 17684 36032 17736 36038
rect 17604 35992 17684 36020
rect 17604 35329 17632 35992
rect 17684 35974 17736 35980
rect 18432 35698 18460 36518
rect 18524 36242 18552 36722
rect 18512 36236 18564 36242
rect 18512 36178 18564 36184
rect 18512 36032 18564 36038
rect 18512 35974 18564 35980
rect 17776 35692 17828 35698
rect 17696 35652 17776 35680
rect 17590 35320 17646 35329
rect 17590 35255 17646 35264
rect 17696 35136 17724 35652
rect 17776 35634 17828 35640
rect 18420 35692 18472 35698
rect 18420 35634 18472 35640
rect 18524 35601 18552 35974
rect 18616 35816 18644 37198
rect 18708 36378 18736 37402
rect 18788 36780 18840 36786
rect 18788 36722 18840 36728
rect 18800 36689 18828 36722
rect 18786 36680 18842 36689
rect 18786 36615 18842 36624
rect 18696 36372 18748 36378
rect 18696 36314 18748 36320
rect 18696 36236 18748 36242
rect 18696 36178 18748 36184
rect 18708 35894 18736 36178
rect 18786 36136 18842 36145
rect 18786 36071 18842 36080
rect 18800 36038 18828 36071
rect 18788 36032 18840 36038
rect 18788 35974 18840 35980
rect 18708 35866 18828 35894
rect 18696 35828 18748 35834
rect 18616 35788 18696 35816
rect 18696 35770 18748 35776
rect 18708 35698 18736 35770
rect 18696 35692 18748 35698
rect 18696 35634 18748 35640
rect 18326 35592 18382 35601
rect 18510 35592 18566 35601
rect 18382 35550 18460 35578
rect 18326 35527 18382 35536
rect 17776 35488 17828 35494
rect 17776 35430 17828 35436
rect 18432 35442 18460 35550
rect 18510 35527 18566 35536
rect 17604 35108 17724 35136
rect 17500 35080 17552 35086
rect 17604 35068 17632 35108
rect 17788 35086 17816 35430
rect 18432 35414 18644 35442
rect 17846 35388 18154 35408
rect 17846 35386 17852 35388
rect 17908 35386 17932 35388
rect 17988 35386 18012 35388
rect 18068 35386 18092 35388
rect 18148 35386 18154 35388
rect 17908 35334 17910 35386
rect 18090 35334 18092 35386
rect 17846 35332 17852 35334
rect 17908 35332 17932 35334
rect 17988 35332 18012 35334
rect 18068 35332 18092 35334
rect 18148 35332 18154 35334
rect 17846 35312 18154 35332
rect 18326 35320 18382 35329
rect 18326 35255 18328 35264
rect 18380 35255 18382 35264
rect 18328 35226 18380 35232
rect 18340 35142 18552 35170
rect 18340 35136 18368 35142
rect 18156 35108 18368 35136
rect 17552 35040 17632 35068
rect 17500 35022 17552 35028
rect 17408 34944 17460 34950
rect 17408 34886 17460 34892
rect 17420 34406 17448 34886
rect 17604 34610 17632 35040
rect 17776 35080 17828 35086
rect 17696 35028 17776 35034
rect 17696 35022 17828 35028
rect 17696 35006 17816 35022
rect 17592 34604 17644 34610
rect 17592 34546 17644 34552
rect 17696 34542 17724 35006
rect 17776 34944 17828 34950
rect 17776 34886 17828 34892
rect 17684 34536 17736 34542
rect 17684 34478 17736 34484
rect 17788 34456 17816 34886
rect 18052 34672 18104 34678
rect 18052 34614 18104 34620
rect 18064 34456 18092 34614
rect 17788 34428 18092 34456
rect 16946 34232 17002 34241
rect 16946 34167 17002 34176
rect 17052 34184 17080 34342
rect 17144 34326 17356 34354
rect 17408 34400 17460 34406
rect 18156 34388 18184 35108
rect 18420 35080 18472 35086
rect 18234 35048 18290 35057
rect 18524 35057 18552 35142
rect 18616 35086 18644 35414
rect 18604 35080 18656 35086
rect 18420 35022 18472 35028
rect 18510 35048 18566 35057
rect 18234 34983 18290 34992
rect 18248 34678 18276 34983
rect 18236 34672 18288 34678
rect 18236 34614 18288 34620
rect 18236 34468 18288 34474
rect 18236 34410 18288 34416
rect 17696 34377 18184 34388
rect 17408 34342 17460 34348
rect 17682 34368 18184 34377
rect 17738 34360 18184 34368
rect 17682 34303 17738 34312
rect 17846 34300 18154 34320
rect 17846 34298 17852 34300
rect 17908 34298 17932 34300
rect 17988 34298 18012 34300
rect 18068 34298 18092 34300
rect 18148 34298 18154 34300
rect 17908 34246 17910 34298
rect 18090 34246 18092 34298
rect 17846 34244 17852 34246
rect 17908 34244 17932 34246
rect 17988 34244 18012 34246
rect 18068 34244 18092 34246
rect 18148 34244 18154 34246
rect 17846 34224 18154 34244
rect 18248 34184 18276 34410
rect 18326 34368 18382 34377
rect 18326 34303 18382 34312
rect 16960 34116 16988 34167
rect 17052 34156 18276 34184
rect 18340 34116 18368 34303
rect 16960 34088 18368 34116
rect 16672 34060 16724 34066
rect 16592 34020 16672 34048
rect 16724 34020 16988 34048
rect 16672 34002 16724 34008
rect 16500 33918 16712 33946
rect 16580 33584 16632 33590
rect 16580 33526 16632 33532
rect 16408 33476 16528 33504
rect 16396 33380 16448 33386
rect 16396 33322 16448 33328
rect 16212 33312 16264 33318
rect 16212 33254 16264 33260
rect 16120 32972 16172 32978
rect 16120 32914 16172 32920
rect 16224 32570 16252 33254
rect 16408 33114 16436 33322
rect 16500 33114 16528 33476
rect 16396 33108 16448 33114
rect 16396 33050 16448 33056
rect 16488 33108 16540 33114
rect 16488 33050 16540 33056
rect 16592 33046 16620 33526
rect 16580 33040 16632 33046
rect 16580 32982 16632 32988
rect 16304 32904 16356 32910
rect 16304 32846 16356 32852
rect 16212 32564 16264 32570
rect 16212 32506 16264 32512
rect 16120 32496 16172 32502
rect 16120 32438 16172 32444
rect 16028 32224 16080 32230
rect 16028 32166 16080 32172
rect 16040 31822 16068 32166
rect 16028 31816 16080 31822
rect 16028 31758 16080 31764
rect 15856 31748 15988 31754
rect 15856 31726 15936 31748
rect 15936 31690 15988 31696
rect 15842 31376 15898 31385
rect 15842 31311 15898 31320
rect 15856 31278 15884 31311
rect 15844 31272 15896 31278
rect 15844 31214 15896 31220
rect 15948 31210 15976 31690
rect 16132 31464 16160 32438
rect 16212 32360 16264 32366
rect 16212 32302 16264 32308
rect 16224 32026 16252 32302
rect 16212 32020 16264 32026
rect 16212 31962 16264 31968
rect 16212 31680 16264 31686
rect 16212 31622 16264 31628
rect 16040 31436 16160 31464
rect 15936 31204 15988 31210
rect 15936 31146 15988 31152
rect 15936 30932 15988 30938
rect 15936 30874 15988 30880
rect 15844 30796 15896 30802
rect 15844 30738 15896 30744
rect 15856 30666 15884 30738
rect 15948 30734 15976 30874
rect 16040 30802 16068 31436
rect 16118 31376 16174 31385
rect 16118 31311 16174 31320
rect 16028 30796 16080 30802
rect 16028 30738 16080 30744
rect 15936 30728 15988 30734
rect 15936 30670 15988 30676
rect 15844 30660 15896 30666
rect 15844 30602 15896 30608
rect 16026 30424 16082 30433
rect 16026 30359 16082 30368
rect 16040 30258 16068 30359
rect 15844 30252 15896 30258
rect 15844 30194 15896 30200
rect 16028 30252 16080 30258
rect 16028 30194 16080 30200
rect 15752 29640 15804 29646
rect 15752 29582 15804 29588
rect 15752 29504 15804 29510
rect 15752 29446 15804 29452
rect 15660 29300 15712 29306
rect 15660 29242 15712 29248
rect 15476 29164 15528 29170
rect 15476 29106 15528 29112
rect 15660 29164 15712 29170
rect 15660 29106 15712 29112
rect 15488 28937 15516 29106
rect 15568 29096 15620 29102
rect 15568 29038 15620 29044
rect 15474 28928 15530 28937
rect 15474 28863 15530 28872
rect 15580 28665 15608 29038
rect 15566 28656 15622 28665
rect 15566 28591 15622 28600
rect 15476 28552 15528 28558
rect 15528 28512 15608 28540
rect 15476 28494 15528 28500
rect 15580 28064 15608 28512
rect 15488 28036 15608 28064
rect 15488 27985 15516 28036
rect 15672 27996 15700 29106
rect 15764 28937 15792 29446
rect 15750 28928 15806 28937
rect 15750 28863 15806 28872
rect 15750 28656 15806 28665
rect 15750 28591 15806 28600
rect 15764 28082 15792 28591
rect 15752 28076 15804 28082
rect 15752 28018 15804 28024
rect 15474 27976 15530 27985
rect 15474 27911 15530 27920
rect 15580 27968 15700 27996
rect 15580 27470 15608 27968
rect 15752 27872 15804 27878
rect 15752 27814 15804 27820
rect 15764 27606 15792 27814
rect 15752 27600 15804 27606
rect 15856 27577 15884 30194
rect 15934 29880 15990 29889
rect 15934 29815 15990 29824
rect 15948 29782 15976 29815
rect 15936 29776 15988 29782
rect 15936 29718 15988 29724
rect 16028 29776 16080 29782
rect 16028 29718 16080 29724
rect 15936 29640 15988 29646
rect 15936 29582 15988 29588
rect 15948 28234 15976 29582
rect 16040 29510 16068 29718
rect 16028 29504 16080 29510
rect 16028 29446 16080 29452
rect 16132 29322 16160 31311
rect 16224 30580 16252 31622
rect 16316 30734 16344 32846
rect 16396 32768 16448 32774
rect 16396 32710 16448 32716
rect 16488 32768 16540 32774
rect 16488 32710 16540 32716
rect 16408 32570 16436 32710
rect 16396 32564 16448 32570
rect 16396 32506 16448 32512
rect 16500 32434 16528 32710
rect 16580 32496 16632 32502
rect 16580 32438 16632 32444
rect 16488 32428 16540 32434
rect 16488 32370 16540 32376
rect 16396 32020 16448 32026
rect 16396 31962 16448 31968
rect 16408 31686 16436 31962
rect 16500 31958 16528 32370
rect 16592 32026 16620 32438
rect 16580 32020 16632 32026
rect 16580 31962 16632 31968
rect 16488 31952 16540 31958
rect 16488 31894 16540 31900
rect 16580 31884 16632 31890
rect 16580 31826 16632 31832
rect 16592 31754 16620 31826
rect 16580 31748 16632 31754
rect 16580 31690 16632 31696
rect 16396 31680 16448 31686
rect 16684 31634 16712 33918
rect 16856 33516 16908 33522
rect 16856 33458 16908 33464
rect 16868 32910 16896 33458
rect 16960 32910 16988 34020
rect 17972 33918 18276 33946
rect 17972 33862 18000 33918
rect 17316 33856 17368 33862
rect 17052 33816 17316 33844
rect 16856 32904 16908 32910
rect 16856 32846 16908 32852
rect 16948 32904 17000 32910
rect 16948 32846 17000 32852
rect 17052 32502 17080 33816
rect 17316 33798 17368 33804
rect 17960 33856 18012 33862
rect 17960 33798 18012 33804
rect 18052 33856 18104 33862
rect 18052 33798 18104 33804
rect 18064 33658 18092 33798
rect 18052 33652 18104 33658
rect 18052 33594 18104 33600
rect 17328 33522 18184 33538
rect 18248 33522 18276 33918
rect 18432 33674 18460 35022
rect 18604 35022 18656 35028
rect 18510 34983 18566 34992
rect 18708 34610 18736 35634
rect 18800 35154 18828 35866
rect 18788 35148 18840 35154
rect 18788 35090 18840 35096
rect 18696 34604 18748 34610
rect 18696 34546 18748 34552
rect 18892 34542 18920 37590
rect 19340 37460 19392 37466
rect 19340 37402 19392 37408
rect 19156 37324 19208 37330
rect 19156 37266 19208 37272
rect 19168 36786 19196 37266
rect 19248 37256 19300 37262
rect 19248 37198 19300 37204
rect 19156 36780 19208 36786
rect 19156 36722 19208 36728
rect 19062 36680 19118 36689
rect 19062 36615 19118 36624
rect 18972 36168 19024 36174
rect 18970 36136 18972 36145
rect 19024 36136 19026 36145
rect 18970 36071 19026 36080
rect 18972 35012 19024 35018
rect 18972 34954 19024 34960
rect 18984 34678 19012 34954
rect 18972 34672 19024 34678
rect 18972 34614 19024 34620
rect 18788 34536 18840 34542
rect 18788 34478 18840 34484
rect 18880 34536 18932 34542
rect 18880 34478 18932 34484
rect 18512 34128 18564 34134
rect 18512 34070 18564 34076
rect 18340 33646 18460 33674
rect 17328 33516 18196 33522
rect 17328 33510 18144 33516
rect 17224 33380 17276 33386
rect 17224 33322 17276 33328
rect 17236 33130 17264 33322
rect 17328 33318 17356 33510
rect 18144 33458 18196 33464
rect 18236 33516 18288 33522
rect 18236 33458 18288 33464
rect 17408 33448 17460 33454
rect 18052 33448 18104 33454
rect 17408 33390 17460 33396
rect 17498 33416 17554 33425
rect 17420 33318 17448 33390
rect 17604 33408 18052 33436
rect 17604 33402 17632 33408
rect 17554 33374 17632 33402
rect 18340 33402 18368 33646
rect 18420 33584 18472 33590
rect 18524 33572 18552 34070
rect 18800 34066 18828 34478
rect 18696 34060 18748 34066
rect 18696 34002 18748 34008
rect 18788 34060 18840 34066
rect 18788 34002 18840 34008
rect 18708 33697 18736 34002
rect 18892 33998 18920 34478
rect 18972 34128 19024 34134
rect 19076 34116 19104 36615
rect 19260 35306 19288 37198
rect 19352 35834 19380 37402
rect 19444 36961 19472 39306
rect 19628 36961 19656 40054
rect 19708 38888 19760 38894
rect 19708 38830 19760 38836
rect 19720 38486 19748 38830
rect 19708 38480 19760 38486
rect 19812 38457 19840 40190
rect 19996 39506 20024 41200
rect 20168 40928 20220 40934
rect 20168 40870 20220 40876
rect 20074 40080 20130 40089
rect 20074 40015 20130 40024
rect 19984 39500 20036 39506
rect 19984 39442 20036 39448
rect 19892 38888 19944 38894
rect 19892 38830 19944 38836
rect 19708 38422 19760 38428
rect 19798 38448 19854 38457
rect 19798 38383 19854 38392
rect 19904 37942 19932 38830
rect 19982 38584 20038 38593
rect 19982 38519 20038 38528
rect 19996 38418 20024 38519
rect 19984 38412 20036 38418
rect 19984 38354 20036 38360
rect 19892 37936 19944 37942
rect 19892 37878 19944 37884
rect 19800 37324 19852 37330
rect 19800 37266 19852 37272
rect 19708 37120 19760 37126
rect 19708 37062 19760 37068
rect 19430 36952 19486 36961
rect 19430 36887 19486 36896
rect 19614 36952 19670 36961
rect 19614 36887 19670 36896
rect 19524 36712 19576 36718
rect 19444 36672 19524 36700
rect 19340 35828 19392 35834
rect 19340 35770 19392 35776
rect 19444 35630 19472 36672
rect 19524 36654 19576 36660
rect 19614 35864 19670 35873
rect 19614 35799 19670 35808
rect 19432 35624 19484 35630
rect 19432 35566 19484 35572
rect 19524 35488 19576 35494
rect 19524 35430 19576 35436
rect 19260 35278 19472 35306
rect 19340 35216 19392 35222
rect 19340 35158 19392 35164
rect 19156 35148 19208 35154
rect 19208 35108 19288 35136
rect 19156 35090 19208 35096
rect 19156 34944 19208 34950
rect 19156 34886 19208 34892
rect 19024 34088 19104 34116
rect 18972 34070 19024 34076
rect 19168 34082 19196 34886
rect 19260 34610 19288 35108
rect 19352 34950 19380 35158
rect 19340 34944 19392 34950
rect 19340 34886 19392 34892
rect 19248 34604 19300 34610
rect 19248 34546 19300 34552
rect 19444 34406 19472 35278
rect 19536 35086 19564 35430
rect 19628 35222 19656 35799
rect 19720 35766 19748 37062
rect 19708 35760 19760 35766
rect 19708 35702 19760 35708
rect 19812 35698 19840 37266
rect 19892 37256 19944 37262
rect 19892 37198 19944 37204
rect 19904 36718 19932 37198
rect 19892 36712 19944 36718
rect 19892 36654 19944 36660
rect 19904 36582 19932 36654
rect 19892 36576 19944 36582
rect 19892 36518 19944 36524
rect 19984 36032 20036 36038
rect 19984 35974 20036 35980
rect 19892 35760 19944 35766
rect 19892 35702 19944 35708
rect 19800 35692 19852 35698
rect 19800 35634 19852 35640
rect 19904 35612 19932 35702
rect 19996 35612 20024 35974
rect 20088 35834 20116 40015
rect 20180 39001 20208 40870
rect 20534 40216 20590 40225
rect 20534 40151 20590 40160
rect 20444 39364 20496 39370
rect 20444 39306 20496 39312
rect 20166 38992 20222 39001
rect 20166 38927 20222 38936
rect 20076 35828 20128 35834
rect 20076 35770 20128 35776
rect 20076 35624 20128 35630
rect 19904 35584 20076 35612
rect 20076 35566 20128 35572
rect 19616 35216 19668 35222
rect 20074 35184 20130 35193
rect 19616 35158 19668 35164
rect 19720 35142 20024 35170
rect 19524 35080 19576 35086
rect 19524 35022 19576 35028
rect 19616 35012 19668 35018
rect 19720 35000 19748 35142
rect 19892 35080 19944 35086
rect 19892 35022 19944 35028
rect 19668 34972 19748 35000
rect 19616 34954 19668 34960
rect 19706 34776 19762 34785
rect 19706 34711 19762 34720
rect 19720 34610 19748 34711
rect 19904 34610 19932 35022
rect 19996 34785 20024 35142
rect 20074 35119 20130 35128
rect 20088 35018 20116 35119
rect 20076 35012 20128 35018
rect 20076 34954 20128 34960
rect 19982 34776 20038 34785
rect 19982 34711 20038 34720
rect 19708 34604 19760 34610
rect 19708 34546 19760 34552
rect 19892 34604 19944 34610
rect 19892 34546 19944 34552
rect 19524 34536 19576 34542
rect 19524 34478 19576 34484
rect 19432 34400 19484 34406
rect 19432 34342 19484 34348
rect 19168 34054 19380 34082
rect 18880 33992 18932 33998
rect 18880 33934 18932 33940
rect 19248 33992 19300 33998
rect 19248 33934 19300 33940
rect 19156 33856 19208 33862
rect 19156 33798 19208 33804
rect 19260 33810 19288 33934
rect 19352 33930 19380 34054
rect 19340 33924 19392 33930
rect 19536 33912 19564 34478
rect 19536 33884 19748 33912
rect 19340 33866 19392 33872
rect 18694 33688 18750 33697
rect 19168 33674 19196 33798
rect 19260 33782 19472 33810
rect 18694 33623 18750 33632
rect 18892 33646 19104 33674
rect 19168 33658 19380 33674
rect 19168 33652 19392 33658
rect 19168 33646 19340 33652
rect 18472 33544 18552 33572
rect 18696 33584 18748 33590
rect 18420 33526 18472 33532
rect 18892 33572 18920 33646
rect 18748 33544 18920 33572
rect 18972 33584 19024 33590
rect 18696 33526 18748 33532
rect 18972 33526 19024 33532
rect 18052 33390 18104 33396
rect 18248 33374 18368 33402
rect 17498 33351 17554 33360
rect 17316 33312 17368 33318
rect 17316 33254 17368 33260
rect 17408 33312 17460 33318
rect 17408 33254 17460 33260
rect 17846 33212 18154 33232
rect 17846 33210 17852 33212
rect 17908 33210 17932 33212
rect 17988 33210 18012 33212
rect 18068 33210 18092 33212
rect 18148 33210 18154 33212
rect 17908 33158 17910 33210
rect 18090 33158 18092 33210
rect 17846 33156 17852 33158
rect 17908 33156 17932 33158
rect 17988 33156 18012 33158
rect 18068 33156 18092 33158
rect 18148 33156 18154 33158
rect 17406 33144 17462 33153
rect 17236 33102 17356 33130
rect 17132 32972 17184 32978
rect 17132 32914 17184 32920
rect 17040 32496 17092 32502
rect 17040 32438 17092 32444
rect 17040 32360 17092 32366
rect 17040 32302 17092 32308
rect 16762 32056 16818 32065
rect 16762 31991 16764 32000
rect 16816 31991 16818 32000
rect 16764 31962 16816 31968
rect 17052 31940 17080 32302
rect 17144 32065 17172 32914
rect 17224 32768 17276 32774
rect 17224 32710 17276 32716
rect 17236 32609 17264 32710
rect 17222 32600 17278 32609
rect 17328 32570 17356 33102
rect 17846 33136 18154 33156
rect 17462 33102 17816 33130
rect 17406 33079 17462 33088
rect 17788 32892 17816 33102
rect 17788 32881 18000 32892
rect 17682 32872 17738 32881
rect 17788 32872 18014 32881
rect 17788 32864 17958 32872
rect 17682 32807 17684 32816
rect 17736 32807 17738 32816
rect 18248 32824 18276 33374
rect 18432 33300 18460 33526
rect 18512 33380 18564 33386
rect 18512 33322 18564 33328
rect 18708 33374 18920 33402
rect 17958 32807 18014 32816
rect 17684 32778 17736 32784
rect 18064 32796 18276 32824
rect 18340 33272 18460 33300
rect 18064 32722 18092 32796
rect 18340 32756 18368 33272
rect 18524 33114 18552 33322
rect 18602 33144 18658 33153
rect 18512 33108 18564 33114
rect 18602 33079 18604 33088
rect 18512 33050 18564 33056
rect 18656 33079 18658 33088
rect 18604 33050 18656 33056
rect 18708 32960 18736 33374
rect 18892 33318 18920 33374
rect 18788 33312 18840 33318
rect 18788 33254 18840 33260
rect 18880 33312 18932 33318
rect 18880 33254 18932 33260
rect 18800 33114 18828 33254
rect 18984 33130 19012 33526
rect 19076 33318 19104 33646
rect 19340 33594 19392 33600
rect 19156 33380 19208 33386
rect 19444 33368 19472 33782
rect 19616 33516 19668 33522
rect 19616 33458 19668 33464
rect 19524 33448 19576 33454
rect 19524 33390 19576 33396
rect 19156 33322 19208 33328
rect 19260 33340 19472 33368
rect 19064 33312 19116 33318
rect 19064 33254 19116 33260
rect 18788 33108 18840 33114
rect 18788 33050 18840 33056
rect 18892 33102 19012 33130
rect 19064 33108 19116 33114
rect 17512 32694 18092 32722
rect 18156 32728 18368 32756
rect 18524 32932 18736 32960
rect 18418 32736 18474 32745
rect 17222 32535 17278 32544
rect 17316 32564 17368 32570
rect 17316 32506 17368 32512
rect 17512 32434 17540 32694
rect 17868 32564 17920 32570
rect 17868 32506 17920 32512
rect 17500 32428 17552 32434
rect 17500 32370 17552 32376
rect 17776 32428 17828 32434
rect 17776 32370 17828 32376
rect 17788 32314 17816 32370
rect 17512 32286 17816 32314
rect 17316 32224 17368 32230
rect 17222 32192 17278 32201
rect 17316 32166 17368 32172
rect 17222 32127 17278 32136
rect 17130 32056 17186 32065
rect 17130 31991 17186 32000
rect 17052 31912 17172 31940
rect 16856 31748 16908 31754
rect 16856 31690 16908 31696
rect 16396 31622 16448 31628
rect 16592 31606 16712 31634
rect 16394 31512 16450 31521
rect 16394 31447 16450 31456
rect 16408 30802 16436 31447
rect 16488 31340 16540 31346
rect 16488 31282 16540 31288
rect 16500 31210 16528 31282
rect 16488 31204 16540 31210
rect 16488 31146 16540 31152
rect 16592 31090 16620 31606
rect 16764 31408 16816 31414
rect 16764 31350 16816 31356
rect 16500 31062 16620 31090
rect 16672 31136 16724 31142
rect 16672 31078 16724 31084
rect 16396 30796 16448 30802
rect 16396 30738 16448 30744
rect 16304 30728 16356 30734
rect 16304 30670 16356 30676
rect 16224 30552 16436 30580
rect 16210 30424 16266 30433
rect 16210 30359 16266 30368
rect 16224 30054 16252 30359
rect 16304 30252 16356 30258
rect 16304 30194 16356 30200
rect 16316 30054 16344 30194
rect 16212 30048 16264 30054
rect 16212 29990 16264 29996
rect 16304 30048 16356 30054
rect 16304 29990 16356 29996
rect 16408 29578 16436 30552
rect 16396 29572 16448 29578
rect 16396 29514 16448 29520
rect 16040 29294 16160 29322
rect 16040 28370 16068 29294
rect 16120 29164 16172 29170
rect 16120 29106 16172 29112
rect 16132 29034 16160 29106
rect 16120 29028 16172 29034
rect 16120 28970 16172 28976
rect 16212 29028 16264 29034
rect 16500 28994 16528 31062
rect 16684 30734 16712 31078
rect 16672 30728 16724 30734
rect 16672 30670 16724 30676
rect 16580 30320 16632 30326
rect 16580 30262 16632 30268
rect 16592 29345 16620 30262
rect 16672 29572 16724 29578
rect 16672 29514 16724 29520
rect 16578 29336 16634 29345
rect 16578 29271 16634 29280
rect 16580 29232 16632 29238
rect 16684 29209 16712 29514
rect 16776 29288 16804 31350
rect 16868 31210 16896 31690
rect 17040 31340 17092 31346
rect 17040 31282 17092 31288
rect 16856 31204 16908 31210
rect 16856 31146 16908 31152
rect 16948 31136 17000 31142
rect 16948 31078 17000 31084
rect 16960 30394 16988 31078
rect 17052 30682 17080 31282
rect 17144 31278 17172 31912
rect 17236 31754 17264 32127
rect 17328 31906 17356 32166
rect 17512 32042 17540 32286
rect 17684 32224 17736 32230
rect 17682 32192 17684 32201
rect 17880 32212 17908 32506
rect 17960 32428 18012 32434
rect 17960 32370 18012 32376
rect 17972 32298 18000 32370
rect 18156 32314 18184 32728
rect 18418 32671 18474 32680
rect 18328 32564 18380 32570
rect 18432 32552 18460 32671
rect 18380 32524 18460 32552
rect 18328 32506 18380 32512
rect 18236 32428 18288 32434
rect 18524 32416 18552 32932
rect 18616 32830 18828 32858
rect 18616 32774 18644 32830
rect 18800 32774 18828 32830
rect 18604 32768 18656 32774
rect 18604 32710 18656 32716
rect 18788 32768 18840 32774
rect 18788 32710 18840 32716
rect 18892 32586 18920 33102
rect 19064 33050 19116 33056
rect 18972 33040 19024 33046
rect 18972 32982 19024 32988
rect 18984 32842 19012 32982
rect 18972 32836 19024 32842
rect 18972 32778 19024 32784
rect 18288 32388 18552 32416
rect 18800 32558 18920 32586
rect 18236 32370 18288 32376
rect 17960 32292 18012 32298
rect 18156 32286 18368 32314
rect 17960 32234 18012 32240
rect 17736 32192 17738 32201
rect 17682 32127 17738 32136
rect 17788 32184 17908 32212
rect 18340 32212 18368 32286
rect 18234 32192 18290 32201
rect 17682 32056 17738 32065
rect 17512 32014 17632 32042
rect 17328 31878 17540 31906
rect 17236 31726 17448 31754
rect 17420 31521 17448 31726
rect 17406 31512 17462 31521
rect 17406 31447 17462 31456
rect 17512 31362 17540 31878
rect 17604 31464 17632 32014
rect 17682 31991 17738 32000
rect 17696 31668 17724 31991
rect 17788 31822 17816 32184
rect 17846 32124 18154 32144
rect 18340 32184 18552 32212
rect 18234 32127 18290 32136
rect 17846 32122 17852 32124
rect 17908 32122 17932 32124
rect 17988 32122 18012 32124
rect 18068 32122 18092 32124
rect 18148 32122 18154 32124
rect 17908 32070 17910 32122
rect 18090 32070 18092 32122
rect 17846 32068 17852 32070
rect 17908 32068 17932 32070
rect 17988 32068 18012 32070
rect 18068 32068 18092 32070
rect 18148 32068 18154 32070
rect 17846 32048 18154 32068
rect 18248 32026 18276 32127
rect 18524 32026 18552 32184
rect 18236 32020 18288 32026
rect 18236 31962 18288 31968
rect 18512 32020 18564 32026
rect 18604 32020 18656 32026
rect 18564 31980 18604 32008
rect 18512 31962 18564 31968
rect 18604 31962 18656 31968
rect 18800 31906 18828 32558
rect 18970 32464 19026 32473
rect 19076 32434 19104 33050
rect 19168 33046 19196 33322
rect 19156 33040 19208 33046
rect 19156 32982 19208 32988
rect 19260 32978 19288 33340
rect 19536 33318 19564 33390
rect 19524 33312 19576 33318
rect 19430 33280 19486 33289
rect 19628 33289 19656 33458
rect 19524 33254 19576 33260
rect 19614 33280 19670 33289
rect 19430 33215 19486 33224
rect 19614 33215 19670 33224
rect 19444 33114 19472 33215
rect 19432 33108 19484 33114
rect 19432 33050 19484 33056
rect 19248 32972 19300 32978
rect 19248 32914 19300 32920
rect 19156 32768 19208 32774
rect 19156 32710 19208 32716
rect 19168 32473 19196 32710
rect 19260 32502 19288 32914
rect 19524 32836 19576 32842
rect 19524 32778 19576 32784
rect 19248 32496 19300 32502
rect 19154 32464 19210 32473
rect 18970 32399 19026 32408
rect 19064 32428 19116 32434
rect 18984 32280 19012 32399
rect 19248 32438 19300 32444
rect 19154 32399 19210 32408
rect 19064 32370 19116 32376
rect 18984 32252 19104 32280
rect 19076 32026 19104 32252
rect 18972 32020 19024 32026
rect 18972 31962 19024 31968
rect 19064 32020 19116 32026
rect 19064 31962 19116 31968
rect 18144 31884 18196 31890
rect 18524 31878 18828 31906
rect 18880 31884 18932 31890
rect 18196 31844 18368 31872
rect 18144 31826 18196 31832
rect 17776 31816 17828 31822
rect 18340 31804 18368 31844
rect 18524 31804 18552 31878
rect 18880 31826 18932 31832
rect 18340 31776 18552 31804
rect 18604 31816 18656 31822
rect 17776 31758 17828 31764
rect 18656 31776 18736 31804
rect 18604 31758 18656 31764
rect 18512 31680 18564 31686
rect 17696 31640 18368 31668
rect 17604 31436 17809 31464
rect 17781 31362 17809 31436
rect 17972 31436 18184 31464
rect 17224 31340 17276 31346
rect 17512 31334 17724 31362
rect 17781 31334 17816 31362
rect 17224 31282 17276 31288
rect 17132 31272 17184 31278
rect 17132 31214 17184 31220
rect 17236 31113 17264 31282
rect 17696 31278 17724 31334
rect 17788 31328 17816 31334
rect 17972 31328 18000 31436
rect 18156 31396 18184 31436
rect 18236 31408 18288 31414
rect 18156 31368 18236 31396
rect 18236 31350 18288 31356
rect 18340 31346 18368 31640
rect 18512 31622 18564 31628
rect 18604 31680 18656 31686
rect 18604 31622 18656 31628
rect 18524 31482 18552 31622
rect 18512 31476 18564 31482
rect 18512 31418 18564 31424
rect 17788 31300 18000 31328
rect 18052 31340 18104 31346
rect 18052 31282 18104 31288
rect 18328 31340 18380 31346
rect 18328 31282 18380 31288
rect 17500 31272 17552 31278
rect 17500 31214 17552 31220
rect 17684 31272 17736 31278
rect 17684 31214 17736 31220
rect 17222 31104 17278 31113
rect 17222 31039 17278 31048
rect 17512 30920 17540 31214
rect 18064 31192 18092 31282
rect 18064 31164 18552 31192
rect 17696 31113 18368 31124
rect 17682 31104 18368 31113
rect 17738 31096 18368 31104
rect 17682 31039 17738 31048
rect 17846 31036 18154 31056
rect 17846 31034 17852 31036
rect 17908 31034 17932 31036
rect 17988 31034 18012 31036
rect 18068 31034 18092 31036
rect 18148 31034 18154 31036
rect 17908 30982 17910 31034
rect 18090 30982 18092 31034
rect 17846 30980 17852 30982
rect 17908 30980 17932 30982
rect 17988 30980 18012 30982
rect 18068 30980 18092 30982
rect 18148 30980 18154 30982
rect 17846 30960 18154 30980
rect 18340 30977 18368 31096
rect 18326 30968 18382 30977
rect 17236 30892 17448 30920
rect 17512 30892 18276 30920
rect 18326 30903 18382 30912
rect 17132 30864 17184 30870
rect 17236 30852 17264 30892
rect 17184 30824 17264 30852
rect 17420 30852 17448 30892
rect 17420 30824 18184 30852
rect 17132 30806 17184 30812
rect 17316 30796 17368 30802
rect 17368 30756 17540 30784
rect 17316 30738 17368 30744
rect 17052 30654 17448 30682
rect 16948 30388 17000 30394
rect 16948 30330 17000 30336
rect 16856 30252 16908 30258
rect 16856 30194 16908 30200
rect 17132 30252 17184 30258
rect 17316 30252 17368 30258
rect 17184 30212 17264 30240
rect 17132 30194 17184 30200
rect 16868 29458 16896 30194
rect 17040 30116 17092 30122
rect 17092 30076 17172 30104
rect 17040 30058 17092 30064
rect 17038 30016 17094 30025
rect 17038 29951 17094 29960
rect 17052 29782 17080 29951
rect 17040 29776 17092 29782
rect 17040 29718 17092 29724
rect 17144 29714 17172 30076
rect 17236 30025 17264 30212
rect 17316 30194 17368 30200
rect 17328 30161 17356 30194
rect 17314 30152 17370 30161
rect 17314 30087 17370 30096
rect 17222 30016 17278 30025
rect 17420 30002 17448 30654
rect 17512 30580 17540 30756
rect 18156 30734 18184 30824
rect 18144 30728 18196 30734
rect 18248 30716 18276 30892
rect 18420 30728 18472 30734
rect 18248 30688 18420 30716
rect 18144 30670 18196 30676
rect 18420 30670 18472 30676
rect 17512 30552 18460 30580
rect 17684 30388 17736 30394
rect 17972 30382 18359 30410
rect 17972 30376 18000 30382
rect 17736 30348 18000 30376
rect 17684 30330 17736 30336
rect 18234 30288 18290 30297
rect 17592 30252 17644 30258
rect 17960 30252 18012 30258
rect 17644 30212 17960 30240
rect 17592 30194 17644 30200
rect 17960 30194 18012 30200
rect 18156 30246 18234 30274
rect 17958 30152 18014 30161
rect 17500 30116 17552 30122
rect 17552 30076 17632 30104
rect 18156 30138 18184 30246
rect 18331 30274 18359 30382
rect 18432 30326 18460 30552
rect 18420 30320 18472 30326
rect 18331 30258 18368 30274
rect 18420 30262 18472 30268
rect 18234 30223 18290 30232
rect 18328 30252 18380 30258
rect 18328 30194 18380 30200
rect 18014 30110 18184 30138
rect 17958 30087 18014 30096
rect 17500 30058 17552 30064
rect 17604 30036 17632 30076
rect 17604 30008 18276 30036
rect 17420 29974 17540 30002
rect 17222 29951 17278 29960
rect 17132 29708 17184 29714
rect 17132 29650 17184 29656
rect 17236 29594 17264 29951
rect 17406 29880 17462 29889
rect 17406 29815 17462 29824
rect 17040 29572 17092 29578
rect 17144 29566 17264 29594
rect 17316 29640 17368 29646
rect 17316 29582 17368 29588
rect 17144 29560 17172 29566
rect 17092 29532 17172 29560
rect 17040 29514 17092 29520
rect 17224 29504 17276 29510
rect 16868 29430 17080 29458
rect 17224 29446 17276 29452
rect 17052 29345 17080 29430
rect 17038 29336 17094 29345
rect 16776 29260 16988 29288
rect 17038 29271 17094 29280
rect 16580 29174 16632 29180
rect 16670 29200 16726 29209
rect 16592 29084 16620 29174
rect 16670 29135 16726 29144
rect 16854 29200 16910 29209
rect 16960 29186 16988 29260
rect 16960 29158 17080 29186
rect 16854 29135 16910 29144
rect 16868 29084 16896 29135
rect 16592 29056 16896 29084
rect 16948 29096 17000 29102
rect 16948 29038 17000 29044
rect 16212 28970 16264 28976
rect 16224 28694 16252 28970
rect 16316 28966 16528 28994
rect 16212 28688 16264 28694
rect 16212 28630 16264 28636
rect 16120 28620 16172 28626
rect 16120 28562 16172 28568
rect 16132 28472 16160 28562
rect 16316 28540 16344 28966
rect 16580 28756 16632 28762
rect 16580 28698 16632 28704
rect 16672 28756 16724 28762
rect 16672 28698 16724 28704
rect 16592 28540 16620 28698
rect 16684 28665 16712 28698
rect 16670 28656 16726 28665
rect 16670 28591 16726 28600
rect 16960 28558 16988 29038
rect 16948 28552 17000 28558
rect 16316 28512 16528 28540
rect 16592 28512 16712 28540
rect 16132 28444 16436 28472
rect 16040 28342 16160 28370
rect 15948 28206 16068 28234
rect 15752 27542 15804 27548
rect 15842 27568 15898 27577
rect 15842 27503 15898 27512
rect 15936 27532 15988 27538
rect 15568 27464 15620 27470
rect 15568 27406 15620 27412
rect 15752 27464 15804 27470
rect 15752 27406 15804 27412
rect 15660 27328 15712 27334
rect 15660 27270 15712 27276
rect 15566 27160 15622 27169
rect 15566 27095 15622 27104
rect 15580 26994 15608 27095
rect 15476 26988 15528 26994
rect 15476 26930 15528 26936
rect 15568 26988 15620 26994
rect 15568 26930 15620 26936
rect 15488 26217 15516 26930
rect 15672 26790 15700 27270
rect 15660 26784 15712 26790
rect 15660 26726 15712 26732
rect 15568 26376 15620 26382
rect 15568 26318 15620 26324
rect 15474 26208 15530 26217
rect 15474 26143 15530 26152
rect 15580 25838 15608 26318
rect 15660 25968 15712 25974
rect 15660 25910 15712 25916
rect 15476 25832 15528 25838
rect 15476 25774 15528 25780
rect 15568 25832 15620 25838
rect 15568 25774 15620 25780
rect 15488 25158 15516 25774
rect 15580 25362 15608 25774
rect 15568 25356 15620 25362
rect 15568 25298 15620 25304
rect 15476 25152 15528 25158
rect 15476 25094 15528 25100
rect 15568 24200 15620 24206
rect 15672 24188 15700 25910
rect 15764 25129 15792 27406
rect 15750 25120 15806 25129
rect 15750 25055 15806 25064
rect 15856 24818 15884 27503
rect 15936 27474 15988 27480
rect 15948 27169 15976 27474
rect 15934 27160 15990 27169
rect 15934 27095 15990 27104
rect 15936 26988 15988 26994
rect 15936 26930 15988 26936
rect 15948 25673 15976 26930
rect 15934 25664 15990 25673
rect 15934 25599 15990 25608
rect 15844 24812 15896 24818
rect 15844 24754 15896 24760
rect 15752 24744 15804 24750
rect 15752 24686 15804 24692
rect 15764 24410 15792 24686
rect 15752 24404 15804 24410
rect 15752 24346 15804 24352
rect 15844 24268 15896 24274
rect 15844 24210 15896 24216
rect 15620 24160 15700 24188
rect 15568 24142 15620 24148
rect 15856 24041 15884 24210
rect 15842 24032 15898 24041
rect 15842 23967 15898 23976
rect 15856 23118 15884 23967
rect 15844 23112 15896 23118
rect 15844 23054 15896 23060
rect 16040 22030 16068 28206
rect 16132 28082 16160 28342
rect 16212 28144 16264 28150
rect 16212 28086 16264 28092
rect 16120 28076 16172 28082
rect 16120 28018 16172 28024
rect 16224 27577 16252 28086
rect 16304 28076 16356 28082
rect 16304 28018 16356 28024
rect 16210 27568 16266 27577
rect 16210 27503 16266 27512
rect 16224 27470 16252 27503
rect 16212 27464 16264 27470
rect 16212 27406 16264 27412
rect 16316 27402 16344 28018
rect 16408 27946 16436 28444
rect 16396 27940 16448 27946
rect 16396 27882 16448 27888
rect 16500 27520 16528 28512
rect 16684 28150 16712 28512
rect 16948 28494 17000 28500
rect 16856 28416 16908 28422
rect 16856 28358 16908 28364
rect 16672 28144 16724 28150
rect 16672 28086 16724 28092
rect 16764 28008 16816 28014
rect 16764 27950 16816 27956
rect 16408 27492 16528 27520
rect 16304 27396 16356 27402
rect 16304 27338 16356 27344
rect 16302 27160 16358 27169
rect 16302 27095 16358 27104
rect 16316 26897 16344 27095
rect 16302 26888 16358 26897
rect 16302 26823 16358 26832
rect 16118 26752 16174 26761
rect 16118 26687 16174 26696
rect 16028 22024 16080 22030
rect 16028 21966 16080 21972
rect 16132 20602 16160 26687
rect 16408 26432 16436 27492
rect 16672 27396 16724 27402
rect 16592 27356 16672 27384
rect 16592 27062 16620 27356
rect 16672 27338 16724 27344
rect 16776 27112 16804 27950
rect 16868 27305 16896 28358
rect 16854 27296 16910 27305
rect 16854 27231 16910 27240
rect 16948 27124 17000 27130
rect 16776 27084 16896 27112
rect 16580 27056 16632 27062
rect 16580 26998 16632 27004
rect 16764 26988 16816 26994
rect 16764 26930 16816 26936
rect 16580 26852 16632 26858
rect 16580 26794 16632 26800
rect 16224 26404 16436 26432
rect 16224 25226 16252 26404
rect 16304 26308 16356 26314
rect 16304 26250 16356 26256
rect 16488 26308 16540 26314
rect 16488 26250 16540 26256
rect 16212 25220 16264 25226
rect 16212 25162 16264 25168
rect 16224 24818 16252 25162
rect 16316 24954 16344 26250
rect 16396 25900 16448 25906
rect 16396 25842 16448 25848
rect 16408 25294 16436 25842
rect 16396 25288 16448 25294
rect 16396 25230 16448 25236
rect 16304 24948 16356 24954
rect 16304 24890 16356 24896
rect 16500 24886 16528 26250
rect 16592 25906 16620 26794
rect 16672 26784 16724 26790
rect 16670 26752 16672 26761
rect 16724 26752 16726 26761
rect 16670 26687 16726 26696
rect 16672 26580 16724 26586
rect 16672 26522 16724 26528
rect 16684 26382 16712 26522
rect 16672 26376 16724 26382
rect 16672 26318 16724 26324
rect 16776 25974 16804 26930
rect 16868 26926 16896 27084
rect 16948 27066 17000 27072
rect 16856 26920 16908 26926
rect 16856 26862 16908 26868
rect 16856 26784 16908 26790
rect 16856 26726 16908 26732
rect 16764 25968 16816 25974
rect 16764 25910 16816 25916
rect 16580 25900 16632 25906
rect 16580 25842 16632 25848
rect 16868 25838 16896 26726
rect 16960 25974 16988 27066
rect 16948 25968 17000 25974
rect 16948 25910 17000 25916
rect 16856 25832 16908 25838
rect 16856 25774 16908 25780
rect 16672 25696 16724 25702
rect 16672 25638 16724 25644
rect 16684 25401 16712 25638
rect 16670 25392 16726 25401
rect 16670 25327 16726 25336
rect 16868 24886 16896 25774
rect 16948 25492 17000 25498
rect 16948 25434 17000 25440
rect 16488 24880 16540 24886
rect 16488 24822 16540 24828
rect 16856 24880 16908 24886
rect 16856 24822 16908 24828
rect 16212 24812 16264 24818
rect 16212 24754 16264 24760
rect 16396 24132 16448 24138
rect 16396 24074 16448 24080
rect 16580 24132 16632 24138
rect 16580 24074 16632 24080
rect 16408 23322 16436 24074
rect 16488 23724 16540 23730
rect 16488 23666 16540 23672
rect 16396 23316 16448 23322
rect 16396 23258 16448 23264
rect 16396 23044 16448 23050
rect 16396 22986 16448 22992
rect 16408 22710 16436 22986
rect 16500 22982 16528 23666
rect 16592 23594 16620 24074
rect 16672 24064 16724 24070
rect 16672 24006 16724 24012
rect 16684 23866 16712 24006
rect 16672 23860 16724 23866
rect 16672 23802 16724 23808
rect 16580 23588 16632 23594
rect 16580 23530 16632 23536
rect 16592 23186 16620 23530
rect 16580 23180 16632 23186
rect 16632 23140 16804 23168
rect 16580 23122 16632 23128
rect 16488 22976 16540 22982
rect 16488 22918 16540 22924
rect 16396 22704 16448 22710
rect 16396 22646 16448 22652
rect 16500 22642 16528 22918
rect 16776 22710 16804 23140
rect 16960 23050 16988 25434
rect 17052 25226 17080 29158
rect 17132 28076 17184 28082
rect 17132 28018 17184 28024
rect 17144 27470 17172 28018
rect 17236 27690 17264 29446
rect 17328 28558 17356 29582
rect 17420 29238 17448 29815
rect 17512 29510 17540 29974
rect 17846 29948 18154 29968
rect 17846 29946 17852 29948
rect 17908 29946 17932 29948
rect 17988 29946 18012 29948
rect 18068 29946 18092 29948
rect 18148 29946 18154 29948
rect 17908 29894 17910 29946
rect 18090 29894 18092 29946
rect 17846 29892 17852 29894
rect 17908 29892 17932 29894
rect 17988 29892 18012 29894
rect 18068 29892 18092 29894
rect 18148 29892 18154 29894
rect 17682 29880 17738 29889
rect 17846 29872 18154 29892
rect 18248 29889 18276 30008
rect 18234 29880 18290 29889
rect 17682 29815 17738 29824
rect 18234 29815 18290 29824
rect 17696 29730 17724 29815
rect 17696 29702 17908 29730
rect 17776 29640 17828 29646
rect 17776 29582 17828 29588
rect 17500 29504 17552 29510
rect 17500 29446 17552 29452
rect 17408 29232 17460 29238
rect 17408 29174 17460 29180
rect 17682 28928 17738 28937
rect 17682 28863 17738 28872
rect 17500 28688 17552 28694
rect 17498 28656 17500 28665
rect 17552 28656 17554 28665
rect 17498 28591 17554 28600
rect 17316 28552 17368 28558
rect 17316 28494 17368 28500
rect 17328 28082 17356 28494
rect 17408 28212 17460 28218
rect 17408 28154 17460 28160
rect 17316 28076 17368 28082
rect 17316 28018 17368 28024
rect 17316 27872 17368 27878
rect 17420 27860 17448 28154
rect 17592 27940 17644 27946
rect 17592 27882 17644 27888
rect 17368 27832 17448 27860
rect 17604 27849 17632 27882
rect 17696 27860 17724 28863
rect 17788 28490 17816 29582
rect 17880 29458 17908 29702
rect 17972 29702 18184 29730
rect 17972 29578 18000 29702
rect 18156 29646 18184 29702
rect 18052 29640 18104 29646
rect 18052 29582 18104 29588
rect 18144 29640 18196 29646
rect 18144 29582 18196 29588
rect 17960 29572 18012 29578
rect 17960 29514 18012 29520
rect 18064 29458 18092 29582
rect 17880 29430 18092 29458
rect 18236 29504 18288 29510
rect 18236 29446 18288 29452
rect 18064 29170 18092 29430
rect 18052 29164 18104 29170
rect 18052 29106 18104 29112
rect 17846 28860 18154 28880
rect 17846 28858 17852 28860
rect 17908 28858 17932 28860
rect 17988 28858 18012 28860
rect 18068 28858 18092 28860
rect 18148 28858 18154 28860
rect 17908 28806 17910 28858
rect 18090 28806 18092 28858
rect 17846 28804 17852 28806
rect 17908 28804 17932 28806
rect 17988 28804 18012 28806
rect 18068 28804 18092 28806
rect 18148 28804 18154 28806
rect 17846 28784 18154 28804
rect 18248 28608 18276 29446
rect 18328 29232 18380 29238
rect 18328 29174 18380 29180
rect 18340 28937 18368 29174
rect 18326 28928 18382 28937
rect 18326 28863 18382 28872
rect 17972 28580 18276 28608
rect 17776 28484 17828 28490
rect 17776 28426 17828 28432
rect 17972 28014 18000 28580
rect 18432 28540 18460 30262
rect 18524 29889 18552 31164
rect 18616 30036 18644 31622
rect 18708 30938 18736 31776
rect 18892 31754 18920 31826
rect 18800 31726 18920 31754
rect 18800 31346 18828 31726
rect 18880 31680 18932 31686
rect 18880 31622 18932 31628
rect 18788 31340 18840 31346
rect 18788 31282 18840 31288
rect 18892 31278 18920 31622
rect 18880 31272 18932 31278
rect 18880 31214 18932 31220
rect 18788 31136 18840 31142
rect 18786 31104 18788 31113
rect 18880 31136 18932 31142
rect 18840 31104 18842 31113
rect 18880 31078 18932 31084
rect 18786 31039 18842 31048
rect 18696 30932 18748 30938
rect 18696 30874 18748 30880
rect 18708 30734 18736 30874
rect 18696 30728 18748 30734
rect 18696 30670 18748 30676
rect 18696 30048 18748 30054
rect 18616 30008 18696 30036
rect 18892 30036 18920 31078
rect 18984 30734 19012 31962
rect 19156 31884 19208 31890
rect 19156 31826 19208 31832
rect 19064 31748 19116 31754
rect 19168 31736 19196 31826
rect 19168 31708 19222 31736
rect 19064 31690 19116 31696
rect 19076 31657 19104 31690
rect 19062 31648 19118 31657
rect 19062 31583 19118 31592
rect 19194 31498 19222 31708
rect 19076 31470 19222 31498
rect 18972 30728 19024 30734
rect 18972 30670 19024 30676
rect 18696 29990 18748 29996
rect 18800 30008 18920 30036
rect 18510 29880 18566 29889
rect 18510 29815 18566 29824
rect 18604 29640 18656 29646
rect 18604 29582 18656 29588
rect 18512 29232 18564 29238
rect 18512 29174 18564 29180
rect 18524 28694 18552 29174
rect 18616 29170 18644 29582
rect 18604 29164 18656 29170
rect 18800 29152 18828 30008
rect 19076 29866 19104 31470
rect 19260 30258 19288 32438
rect 19340 32428 19392 32434
rect 19340 32370 19392 32376
rect 19352 31958 19380 32370
rect 19340 31952 19392 31958
rect 19340 31894 19392 31900
rect 19536 31686 19564 32778
rect 19720 31890 19748 33884
rect 19800 33516 19852 33522
rect 19800 33458 19852 33464
rect 19812 33386 19840 33458
rect 19800 33380 19852 33386
rect 19800 33322 19852 33328
rect 19812 32570 19840 33322
rect 19892 32836 19944 32842
rect 19892 32778 19944 32784
rect 19800 32564 19852 32570
rect 19800 32506 19852 32512
rect 19904 32473 19932 32778
rect 19996 32745 20024 34711
rect 20180 33946 20208 38927
rect 20456 38654 20484 39306
rect 20272 38626 20484 38654
rect 20272 38418 20300 38626
rect 20260 38412 20312 38418
rect 20260 38354 20312 38360
rect 20548 37874 20576 40151
rect 20640 38418 20668 41200
rect 21638 40896 21694 40905
rect 21638 40831 21694 40840
rect 20812 39840 20864 39846
rect 20812 39782 20864 39788
rect 20720 39296 20772 39302
rect 20720 39238 20772 39244
rect 20628 38412 20680 38418
rect 20628 38354 20680 38360
rect 20732 38049 20760 39238
rect 20718 38040 20774 38049
rect 20718 37975 20774 37984
rect 20260 37868 20312 37874
rect 20536 37868 20588 37874
rect 20312 37828 20484 37856
rect 20260 37810 20312 37816
rect 20260 37256 20312 37262
rect 20260 37198 20312 37204
rect 20352 37256 20404 37262
rect 20352 37198 20404 37204
rect 20272 37126 20300 37198
rect 20260 37120 20312 37126
rect 20260 37062 20312 37068
rect 20364 36122 20392 37198
rect 20272 36094 20392 36122
rect 20272 35086 20300 36094
rect 20456 35737 20484 37828
rect 20588 37828 20668 37856
rect 20536 37810 20588 37816
rect 20640 37274 20668 37828
rect 20824 37505 20852 39782
rect 20996 39092 21048 39098
rect 20996 39034 21048 39040
rect 21008 38826 21036 39034
rect 20996 38820 21048 38826
rect 20996 38762 21048 38768
rect 21088 38752 21140 38758
rect 21088 38694 21140 38700
rect 20996 38004 21048 38010
rect 20996 37946 21048 37952
rect 21008 37806 21036 37946
rect 20996 37800 21048 37806
rect 20996 37742 21048 37748
rect 20810 37496 20866 37505
rect 20810 37431 20866 37440
rect 20994 37496 21050 37505
rect 20994 37431 21050 37440
rect 20640 37262 20852 37274
rect 20640 37256 20864 37262
rect 20640 37246 20812 37256
rect 20640 36786 20668 37246
rect 20812 37198 20864 37204
rect 20720 37188 20772 37194
rect 20720 37130 20772 37136
rect 20732 37097 20760 37130
rect 20718 37088 20774 37097
rect 20718 37023 20774 37032
rect 20810 36816 20866 36825
rect 20628 36780 20680 36786
rect 20810 36751 20866 36760
rect 20628 36722 20680 36728
rect 20640 36258 20668 36722
rect 20720 36576 20772 36582
rect 20720 36518 20772 36524
rect 20732 36378 20760 36518
rect 20720 36372 20772 36378
rect 20720 36314 20772 36320
rect 20536 36236 20588 36242
rect 20640 36230 20760 36258
rect 20536 36178 20588 36184
rect 20548 36009 20576 36178
rect 20534 36000 20590 36009
rect 20534 35935 20590 35944
rect 20732 35850 20760 36230
rect 20824 36009 20852 36751
rect 20902 36408 20958 36417
rect 20902 36343 20958 36352
rect 20810 36000 20866 36009
rect 20810 35935 20866 35944
rect 20536 35828 20588 35834
rect 20536 35770 20588 35776
rect 20640 35822 20760 35850
rect 20442 35728 20498 35737
rect 20442 35663 20498 35672
rect 20350 35592 20406 35601
rect 20350 35527 20406 35536
rect 20364 35494 20392 35527
rect 20352 35488 20404 35494
rect 20352 35430 20404 35436
rect 20260 35080 20312 35086
rect 20260 35022 20312 35028
rect 20444 35080 20496 35086
rect 20548 35068 20576 35770
rect 20640 35698 20668 35822
rect 20628 35692 20680 35698
rect 20628 35634 20680 35640
rect 20916 35290 20944 36343
rect 21008 35766 21036 37431
rect 21100 37330 21128 38694
rect 21454 38176 21510 38185
rect 21454 38111 21510 38120
rect 21468 37466 21496 38111
rect 21456 37460 21508 37466
rect 21456 37402 21508 37408
rect 21088 37324 21140 37330
rect 21088 37266 21140 37272
rect 21364 37256 21416 37262
rect 21364 37198 21416 37204
rect 21376 36922 21404 37198
rect 21548 37120 21600 37126
rect 21548 37062 21600 37068
rect 21364 36916 21416 36922
rect 21364 36858 21416 36864
rect 21560 36854 21588 37062
rect 21548 36848 21600 36854
rect 21548 36790 21600 36796
rect 21180 36780 21232 36786
rect 21180 36722 21232 36728
rect 21086 36408 21142 36417
rect 21086 36343 21142 36352
rect 21100 36145 21128 36343
rect 21086 36136 21142 36145
rect 21086 36071 21142 36080
rect 20996 35760 21048 35766
rect 20996 35702 21048 35708
rect 21086 35592 21142 35601
rect 21086 35527 21142 35536
rect 20994 35456 21050 35465
rect 20994 35391 21050 35400
rect 20904 35284 20956 35290
rect 20904 35226 20956 35232
rect 20812 35216 20864 35222
rect 20812 35158 20864 35164
rect 20824 35086 20852 35158
rect 20628 35080 20680 35086
rect 20548 35040 20628 35068
rect 20444 35022 20496 35028
rect 20628 35022 20680 35028
rect 20812 35080 20864 35086
rect 20812 35022 20864 35028
rect 20456 34202 20484 35022
rect 20444 34196 20496 34202
rect 20444 34138 20496 34144
rect 20258 34096 20314 34105
rect 20258 34031 20260 34040
rect 20312 34031 20314 34040
rect 20260 34002 20312 34008
rect 20180 33918 20300 33946
rect 20074 33688 20130 33697
rect 20074 33623 20130 33632
rect 20088 33522 20116 33623
rect 20076 33516 20128 33522
rect 20076 33458 20128 33464
rect 19982 32736 20038 32745
rect 19982 32671 20038 32680
rect 19890 32464 19946 32473
rect 19890 32399 19946 32408
rect 19708 31884 19760 31890
rect 19708 31826 19760 31832
rect 19616 31748 19668 31754
rect 19616 31690 19668 31696
rect 19708 31748 19760 31754
rect 19708 31690 19760 31696
rect 19524 31680 19576 31686
rect 19430 31648 19486 31657
rect 19524 31622 19576 31628
rect 19430 31583 19486 31592
rect 19338 31376 19394 31385
rect 19338 31311 19340 31320
rect 19392 31311 19394 31320
rect 19340 31282 19392 31288
rect 19444 31142 19472 31583
rect 19628 31385 19656 31690
rect 19614 31376 19670 31385
rect 19614 31311 19670 31320
rect 19432 31136 19484 31142
rect 19432 31078 19484 31084
rect 19616 31136 19668 31142
rect 19616 31078 19668 31084
rect 19628 30802 19656 31078
rect 19616 30796 19668 30802
rect 19616 30738 19668 30744
rect 19340 30728 19392 30734
rect 19340 30670 19392 30676
rect 19248 30252 19300 30258
rect 19248 30194 19300 30200
rect 18892 29838 19104 29866
rect 18800 29124 18844 29152
rect 18604 29106 18656 29112
rect 18816 29050 18844 29124
rect 18800 29022 18844 29050
rect 18512 28688 18564 28694
rect 18512 28630 18564 28636
rect 18604 28688 18656 28694
rect 18604 28630 18656 28636
rect 18064 28512 18460 28540
rect 18064 28082 18092 28512
rect 18328 28416 18380 28422
rect 18512 28416 18564 28422
rect 18380 28376 18460 28404
rect 18328 28358 18380 28364
rect 18052 28076 18104 28082
rect 18052 28018 18104 28024
rect 17960 28008 18012 28014
rect 17960 27950 18012 27956
rect 17590 27840 17646 27849
rect 17316 27814 17368 27820
rect 17696 27832 18276 27860
rect 17590 27775 17646 27784
rect 17846 27772 18154 27792
rect 17846 27770 17852 27772
rect 17908 27770 17932 27772
rect 17988 27770 18012 27772
rect 18068 27770 18092 27772
rect 18148 27770 18154 27772
rect 17908 27718 17910 27770
rect 18090 27718 18092 27770
rect 17846 27716 17852 27718
rect 17908 27716 17932 27718
rect 17988 27716 18012 27718
rect 18068 27716 18092 27718
rect 18148 27716 18154 27718
rect 17682 27704 17738 27713
rect 17236 27662 17448 27690
rect 17420 27538 17448 27662
rect 17846 27696 18154 27716
rect 18248 27713 18276 27832
rect 18326 27840 18382 27849
rect 18326 27775 18382 27784
rect 18234 27704 18290 27713
rect 17682 27639 17738 27648
rect 18234 27639 18290 27648
rect 17696 27588 17724 27639
rect 18052 27600 18104 27606
rect 17696 27560 17816 27588
rect 17408 27532 17460 27538
rect 17408 27474 17460 27480
rect 17592 27532 17644 27538
rect 17644 27492 17724 27520
rect 17592 27474 17644 27480
rect 17132 27464 17184 27470
rect 17132 27406 17184 27412
rect 17144 26450 17172 27406
rect 17222 27296 17278 27305
rect 17222 27231 17278 27240
rect 17236 27062 17264 27231
rect 17420 27130 17448 27474
rect 17592 27396 17644 27402
rect 17592 27338 17644 27344
rect 17408 27124 17460 27130
rect 17460 27084 17540 27112
rect 17408 27066 17460 27072
rect 17224 27056 17276 27062
rect 17224 26998 17276 27004
rect 17224 26920 17276 26926
rect 17224 26862 17276 26868
rect 17132 26444 17184 26450
rect 17132 26386 17184 26392
rect 17236 26382 17264 26862
rect 17406 26752 17462 26761
rect 17406 26687 17462 26696
rect 17224 26376 17276 26382
rect 17224 26318 17276 26324
rect 17316 26308 17368 26314
rect 17316 26250 17368 26256
rect 17328 25498 17356 26250
rect 17316 25492 17368 25498
rect 17316 25434 17368 25440
rect 17420 25362 17448 26687
rect 17512 26586 17540 27084
rect 17604 26761 17632 27338
rect 17696 27130 17724 27492
rect 17684 27124 17736 27130
rect 17788 27112 17816 27560
rect 18340 27577 18368 27775
rect 18432 27674 18460 28376
rect 18512 28358 18564 28364
rect 18524 28150 18552 28358
rect 18512 28144 18564 28150
rect 18512 28086 18564 28092
rect 18420 27668 18472 27674
rect 18420 27610 18472 27616
rect 18512 27600 18564 27606
rect 18052 27542 18104 27548
rect 18326 27568 18382 27577
rect 18064 27334 18092 27542
rect 18510 27568 18512 27577
rect 18564 27568 18566 27577
rect 18326 27503 18382 27512
rect 18420 27532 18472 27538
rect 18510 27503 18566 27512
rect 18420 27474 18472 27480
rect 17960 27328 18012 27334
rect 17960 27270 18012 27276
rect 18052 27328 18104 27334
rect 18052 27270 18104 27276
rect 17868 27124 17920 27130
rect 17788 27084 17868 27112
rect 17684 27066 17736 27072
rect 17868 27066 17920 27072
rect 17590 26752 17646 26761
rect 17590 26687 17646 26696
rect 17500 26580 17552 26586
rect 17500 26522 17552 26528
rect 17696 26466 17724 27066
rect 17972 26908 18000 27270
rect 18052 26920 18104 26926
rect 17972 26880 18052 26908
rect 18052 26862 18104 26868
rect 18236 26852 18288 26858
rect 18236 26794 18288 26800
rect 17846 26684 18154 26704
rect 17846 26682 17852 26684
rect 17908 26682 17932 26684
rect 17988 26682 18012 26684
rect 18068 26682 18092 26684
rect 18148 26682 18154 26684
rect 17908 26630 17910 26682
rect 18090 26630 18092 26682
rect 17846 26628 17852 26630
rect 17908 26628 17932 26630
rect 17988 26628 18012 26630
rect 18068 26628 18092 26630
rect 18148 26628 18154 26630
rect 17846 26608 18154 26628
rect 17512 26438 17724 26466
rect 18144 26444 18196 26450
rect 17512 25498 17540 26438
rect 18248 26432 18276 26794
rect 18328 26512 18380 26518
rect 18328 26454 18380 26460
rect 18196 26404 18276 26432
rect 18144 26386 18196 26392
rect 18248 25838 18276 26404
rect 18236 25832 18288 25838
rect 18236 25774 18288 25780
rect 17696 25673 18276 25684
rect 17682 25664 18290 25673
rect 17738 25656 18234 25664
rect 17682 25599 17738 25608
rect 17846 25596 18154 25616
rect 18234 25599 18290 25608
rect 17846 25594 17852 25596
rect 17908 25594 17932 25596
rect 17988 25594 18012 25596
rect 18068 25594 18092 25596
rect 18148 25594 18154 25596
rect 17908 25542 17910 25594
rect 18090 25542 18092 25594
rect 17846 25540 17852 25542
rect 17908 25540 17932 25542
rect 17988 25540 18012 25542
rect 18068 25540 18092 25542
rect 18148 25540 18154 25542
rect 17682 25528 17738 25537
rect 17500 25492 17552 25498
rect 17846 25520 18154 25540
rect 18340 25480 18368 26454
rect 18432 26382 18460 27474
rect 18512 27396 18564 27402
rect 18512 27338 18564 27344
rect 18524 26586 18552 27338
rect 18512 26580 18564 26586
rect 18512 26522 18564 26528
rect 18420 26376 18472 26382
rect 18420 26318 18472 26324
rect 18420 25968 18472 25974
rect 18420 25910 18472 25916
rect 17682 25463 17738 25472
rect 17500 25434 17552 25440
rect 17696 25430 17724 25463
rect 18064 25452 18368 25480
rect 17684 25424 17736 25430
rect 17684 25366 17736 25372
rect 17408 25356 17460 25362
rect 17408 25298 17460 25304
rect 17040 25220 17092 25226
rect 17040 25162 17092 25168
rect 17684 25220 17736 25226
rect 17684 25162 17736 25168
rect 17500 24812 17552 24818
rect 17500 24754 17552 24760
rect 17408 24200 17460 24206
rect 17408 24142 17460 24148
rect 17040 24132 17092 24138
rect 17040 24074 17092 24080
rect 17052 23730 17080 24074
rect 17420 23730 17448 24142
rect 17040 23724 17092 23730
rect 17040 23666 17092 23672
rect 17408 23724 17460 23730
rect 17408 23666 17460 23672
rect 16948 23044 17000 23050
rect 16948 22986 17000 22992
rect 16580 22704 16632 22710
rect 16764 22704 16816 22710
rect 16632 22652 16712 22658
rect 16580 22646 16712 22652
rect 16764 22646 16816 22652
rect 16488 22636 16540 22642
rect 16592 22630 16712 22646
rect 16488 22578 16540 22584
rect 16500 22216 16528 22578
rect 16580 22568 16632 22574
rect 16580 22510 16632 22516
rect 16592 22438 16620 22510
rect 16580 22432 16632 22438
rect 16580 22374 16632 22380
rect 16500 22188 16620 22216
rect 16488 22024 16540 22030
rect 16488 21966 16540 21972
rect 16120 20596 16172 20602
rect 16120 20538 16172 20544
rect 16500 18766 16528 21966
rect 16592 21554 16620 22188
rect 16684 22094 16712 22630
rect 16776 22234 16804 22646
rect 17052 22438 17080 23666
rect 17040 22432 17092 22438
rect 17040 22374 17092 22380
rect 17052 22234 17080 22374
rect 16764 22228 16816 22234
rect 17040 22228 17092 22234
rect 16816 22188 16988 22216
rect 16764 22170 16816 22176
rect 16684 22066 16896 22094
rect 16580 21548 16632 21554
rect 16580 21490 16632 21496
rect 16868 20806 16896 22066
rect 16960 21418 16988 22188
rect 17040 22170 17092 22176
rect 17408 22024 17460 22030
rect 17408 21966 17460 21972
rect 17040 21956 17092 21962
rect 17040 21898 17092 21904
rect 16948 21412 17000 21418
rect 16948 21354 17000 21360
rect 17052 21146 17080 21898
rect 17420 21554 17448 21966
rect 17408 21548 17460 21554
rect 17408 21490 17460 21496
rect 17224 21344 17276 21350
rect 17224 21286 17276 21292
rect 17040 21140 17092 21146
rect 17040 21082 17092 21088
rect 17236 20942 17264 21286
rect 17420 21078 17448 21490
rect 17408 21072 17460 21078
rect 17408 21014 17460 21020
rect 17224 20936 17276 20942
rect 17224 20878 17276 20884
rect 16856 20800 16908 20806
rect 16856 20742 16908 20748
rect 16488 18760 16540 18766
rect 16488 18702 16540 18708
rect 15476 3936 15528 3942
rect 15476 3878 15528 3884
rect 15488 3602 15516 3878
rect 15476 3596 15528 3602
rect 15476 3538 15528 3544
rect 16120 3596 16172 3602
rect 16120 3538 16172 3544
rect 15660 3460 15712 3466
rect 15660 3402 15712 3408
rect 15672 2650 15700 3402
rect 15752 3188 15804 3194
rect 15752 3130 15804 3136
rect 15660 2644 15712 2650
rect 15660 2586 15712 2592
rect 15764 2446 15792 3130
rect 15752 2440 15804 2446
rect 15752 2382 15804 2388
rect 15384 2372 15436 2378
rect 15384 2314 15436 2320
rect 16132 800 16160 3538
rect 16856 3528 16908 3534
rect 16856 3470 16908 3476
rect 16868 3058 16896 3470
rect 16856 3052 16908 3058
rect 16856 2994 16908 3000
rect 17040 2984 17092 2990
rect 17040 2926 17092 2932
rect 17408 2984 17460 2990
rect 17408 2926 17460 2932
rect 17052 2650 17080 2926
rect 17040 2644 17092 2650
rect 17040 2586 17092 2592
rect 17420 800 17448 2926
rect 17512 2650 17540 24754
rect 17696 24256 17724 25162
rect 18064 24818 18092 25452
rect 18328 25356 18380 25362
rect 18432 25344 18460 25910
rect 18380 25316 18460 25344
rect 18328 25298 18380 25304
rect 18144 25152 18196 25158
rect 18144 25094 18196 25100
rect 18236 25152 18288 25158
rect 18236 25094 18288 25100
rect 18510 25120 18566 25129
rect 18156 24886 18184 25094
rect 18144 24880 18196 24886
rect 18144 24822 18196 24828
rect 18052 24812 18104 24818
rect 18052 24754 18104 24760
rect 17868 24744 17920 24750
rect 17868 24686 17920 24692
rect 17776 24608 17828 24614
rect 17880 24596 17908 24686
rect 17828 24568 17908 24596
rect 17776 24550 17828 24556
rect 17846 24508 18154 24528
rect 17846 24506 17852 24508
rect 17908 24506 17932 24508
rect 17988 24506 18012 24508
rect 18068 24506 18092 24508
rect 18148 24506 18154 24508
rect 17908 24454 17910 24506
rect 18090 24454 18092 24506
rect 17846 24452 17852 24454
rect 17908 24452 17932 24454
rect 17988 24452 18012 24454
rect 18068 24452 18092 24454
rect 18148 24452 18154 24454
rect 17846 24432 18154 24452
rect 18248 24290 18276 25094
rect 18510 25055 18566 25064
rect 18420 24608 18472 24614
rect 18420 24550 18472 24556
rect 18328 24404 18380 24410
rect 18328 24346 18380 24352
rect 17868 24268 17920 24274
rect 17696 24228 17868 24256
rect 17788 23118 17816 24228
rect 17868 24210 17920 24216
rect 17972 24262 18276 24290
rect 17972 24154 18000 24262
rect 17880 24126 18000 24154
rect 18144 24200 18196 24206
rect 18196 24160 18276 24188
rect 18144 24142 18196 24148
rect 17880 24070 17908 24126
rect 17868 24064 17920 24070
rect 17868 24006 17920 24012
rect 17960 24064 18012 24070
rect 17960 24006 18012 24012
rect 17972 23662 18000 24006
rect 18144 23860 18196 23866
rect 18248 23848 18276 24160
rect 18340 24070 18368 24346
rect 18432 24313 18460 24550
rect 18524 24410 18552 25055
rect 18512 24404 18564 24410
rect 18512 24346 18564 24352
rect 18418 24304 18474 24313
rect 18418 24239 18474 24248
rect 18420 24132 18472 24138
rect 18420 24074 18472 24080
rect 18328 24064 18380 24070
rect 18432 24041 18460 24074
rect 18328 24006 18380 24012
rect 18418 24032 18474 24041
rect 18196 23820 18276 23848
rect 18144 23802 18196 23808
rect 17960 23656 18012 23662
rect 17960 23598 18012 23604
rect 17846 23420 18154 23440
rect 17846 23418 17852 23420
rect 17908 23418 17932 23420
rect 17988 23418 18012 23420
rect 18068 23418 18092 23420
rect 18148 23418 18154 23420
rect 17908 23366 17910 23418
rect 18090 23366 18092 23418
rect 17846 23364 17852 23366
rect 17908 23364 17932 23366
rect 17988 23364 18012 23366
rect 18068 23364 18092 23366
rect 18148 23364 18154 23366
rect 17846 23344 18154 23364
rect 18248 23322 18276 23820
rect 18236 23316 18288 23322
rect 18236 23258 18288 23264
rect 17776 23112 17828 23118
rect 17776 23054 17828 23060
rect 18340 22778 18368 24006
rect 18418 23967 18474 23976
rect 18510 23896 18566 23905
rect 18420 23860 18472 23866
rect 18510 23831 18512 23840
rect 18420 23802 18472 23808
rect 18564 23831 18566 23840
rect 18512 23802 18564 23808
rect 17776 22772 17828 22778
rect 17776 22714 17828 22720
rect 18328 22772 18380 22778
rect 18328 22714 18380 22720
rect 17788 22438 17816 22714
rect 18432 22642 18460 23802
rect 18420 22636 18472 22642
rect 18420 22578 18472 22584
rect 17776 22432 17828 22438
rect 17776 22374 17828 22380
rect 17846 22332 18154 22352
rect 17846 22330 17852 22332
rect 17908 22330 17932 22332
rect 17988 22330 18012 22332
rect 18068 22330 18092 22332
rect 18148 22330 18154 22332
rect 17908 22278 17910 22330
rect 18090 22278 18092 22330
rect 17846 22276 17852 22278
rect 17908 22276 17932 22278
rect 17988 22276 18012 22278
rect 18068 22276 18092 22278
rect 18148 22276 18154 22278
rect 17846 22256 18154 22276
rect 18616 22094 18644 28630
rect 18696 28416 18748 28422
rect 18696 28358 18748 28364
rect 18708 27062 18736 28358
rect 18800 27282 18828 29022
rect 18892 28694 18920 29838
rect 18972 29640 19024 29646
rect 19352 29628 19380 30670
rect 19720 30666 19748 31690
rect 19890 31240 19946 31249
rect 19890 31175 19946 31184
rect 19800 30728 19852 30734
rect 19800 30670 19852 30676
rect 19708 30660 19760 30666
rect 19708 30602 19760 30608
rect 19430 30560 19486 30569
rect 19430 30495 19486 30504
rect 19444 29782 19472 30495
rect 19706 30424 19762 30433
rect 19812 30410 19840 30670
rect 19904 30433 19932 31175
rect 19762 30382 19840 30410
rect 19890 30424 19946 30433
rect 19706 30359 19762 30368
rect 19890 30359 19946 30368
rect 19524 30252 19576 30258
rect 19524 30194 19576 30200
rect 19432 29776 19484 29782
rect 19432 29718 19484 29724
rect 19536 29714 19564 30194
rect 19524 29708 19576 29714
rect 19524 29650 19576 29656
rect 19024 29600 19380 29628
rect 18972 29582 19024 29588
rect 18984 29170 19012 29582
rect 18972 29164 19024 29170
rect 18972 29106 19024 29112
rect 18972 29028 19024 29034
rect 18972 28970 19024 28976
rect 19248 29028 19300 29034
rect 19248 28970 19300 28976
rect 18880 28688 18932 28694
rect 18880 28630 18932 28636
rect 18984 28626 19012 28970
rect 19064 28756 19116 28762
rect 19064 28698 19116 28704
rect 19076 28665 19104 28698
rect 19062 28656 19118 28665
rect 18972 28620 19024 28626
rect 19062 28591 19118 28600
rect 18972 28562 19024 28568
rect 18880 28416 18932 28422
rect 18880 28358 18932 28364
rect 18892 28150 18920 28358
rect 18880 28144 18932 28150
rect 18880 28086 18932 28092
rect 18984 27470 19012 28562
rect 19156 28416 19208 28422
rect 19156 28358 19208 28364
rect 19064 28144 19116 28150
rect 19064 28086 19116 28092
rect 18972 27464 19024 27470
rect 18972 27406 19024 27412
rect 18972 27328 19024 27334
rect 18800 27254 18920 27282
rect 18972 27270 19024 27276
rect 18788 27124 18840 27130
rect 18788 27066 18840 27072
rect 18696 27056 18748 27062
rect 18696 26998 18748 27004
rect 18800 26625 18828 27066
rect 18786 26616 18842 26625
rect 18696 26580 18748 26586
rect 18786 26551 18842 26560
rect 18696 26522 18748 26528
rect 18708 26489 18736 26522
rect 18694 26480 18750 26489
rect 18694 26415 18750 26424
rect 18696 26240 18748 26246
rect 18696 26182 18748 26188
rect 18708 26042 18736 26182
rect 18696 26036 18748 26042
rect 18696 25978 18748 25984
rect 18788 26036 18840 26042
rect 18788 25978 18840 25984
rect 18800 25906 18828 25978
rect 18788 25900 18840 25906
rect 18788 25842 18840 25848
rect 18892 25809 18920 27254
rect 18984 26976 19012 27270
rect 19076 27112 19104 28086
rect 19168 27402 19196 28358
rect 19260 27441 19288 28970
rect 19536 28762 19564 29650
rect 19616 29504 19668 29510
rect 19668 29464 19932 29492
rect 19616 29446 19668 29452
rect 19616 29096 19668 29102
rect 19616 29038 19668 29044
rect 19628 28762 19656 29038
rect 19524 28756 19576 28762
rect 19524 28698 19576 28704
rect 19616 28756 19668 28762
rect 19616 28698 19668 28704
rect 19340 28484 19392 28490
rect 19340 28426 19392 28432
rect 19352 27946 19380 28426
rect 19536 28082 19564 28698
rect 19628 28422 19656 28698
rect 19708 28484 19760 28490
rect 19708 28426 19760 28432
rect 19616 28416 19668 28422
rect 19616 28358 19668 28364
rect 19720 28257 19748 28426
rect 19800 28416 19852 28422
rect 19800 28358 19852 28364
rect 19706 28248 19762 28257
rect 19706 28183 19762 28192
rect 19524 28076 19576 28082
rect 19524 28018 19576 28024
rect 19812 28014 19840 28358
rect 19904 28257 19932 29464
rect 19890 28248 19946 28257
rect 19890 28183 19946 28192
rect 19800 28008 19852 28014
rect 19800 27950 19852 27956
rect 19340 27940 19392 27946
rect 19340 27882 19392 27888
rect 19352 27520 19380 27882
rect 19892 27668 19944 27674
rect 19892 27610 19944 27616
rect 19904 27577 19932 27610
rect 19890 27568 19946 27577
rect 19432 27532 19484 27538
rect 19352 27492 19432 27520
rect 19432 27474 19484 27480
rect 19616 27532 19668 27538
rect 19890 27503 19946 27512
rect 19616 27474 19668 27480
rect 19246 27432 19302 27441
rect 19156 27396 19208 27402
rect 19246 27367 19302 27376
rect 19156 27338 19208 27344
rect 19076 27084 19288 27112
rect 19156 26988 19208 26994
rect 18984 26948 19156 26976
rect 19156 26930 19208 26936
rect 18970 26752 19026 26761
rect 18970 26687 19026 26696
rect 18878 25800 18934 25809
rect 18878 25735 18934 25744
rect 18786 25392 18842 25401
rect 18786 25327 18842 25336
rect 18800 25294 18828 25327
rect 18788 25288 18840 25294
rect 18788 25230 18840 25236
rect 18800 25158 18828 25230
rect 18788 25152 18840 25158
rect 18788 25094 18840 25100
rect 18984 24721 19012 26687
rect 18970 24712 19026 24721
rect 18970 24647 19026 24656
rect 19260 24177 19288 27084
rect 19524 26920 19576 26926
rect 19444 26880 19524 26908
rect 19340 26376 19392 26382
rect 19444 26364 19472 26880
rect 19524 26862 19576 26868
rect 19524 26784 19576 26790
rect 19524 26726 19576 26732
rect 19536 26382 19564 26726
rect 19392 26336 19472 26364
rect 19340 26318 19392 26324
rect 19444 25906 19472 26336
rect 19524 26376 19576 26382
rect 19524 26318 19576 26324
rect 19628 26081 19656 27474
rect 19996 27130 20024 32671
rect 20074 32464 20130 32473
rect 20074 32399 20130 32408
rect 20088 31793 20116 32399
rect 20168 32224 20220 32230
rect 20168 32166 20220 32172
rect 20180 32065 20208 32166
rect 20166 32056 20222 32065
rect 20166 31991 20222 32000
rect 20074 31784 20130 31793
rect 20074 31719 20130 31728
rect 20076 31680 20128 31686
rect 20076 31622 20128 31628
rect 19984 27124 20036 27130
rect 19984 27066 20036 27072
rect 19708 27056 19760 27062
rect 19708 26998 19760 27004
rect 19720 26314 19748 26998
rect 19892 26920 19944 26926
rect 19892 26862 19944 26868
rect 19904 26382 19932 26862
rect 19892 26376 19944 26382
rect 19892 26318 19944 26324
rect 19708 26308 19760 26314
rect 19708 26250 19760 26256
rect 19614 26072 19670 26081
rect 19614 26007 19670 26016
rect 19720 25974 19748 26250
rect 19708 25968 19760 25974
rect 19708 25910 19760 25916
rect 19800 25968 19852 25974
rect 19800 25910 19852 25916
rect 19432 25900 19484 25906
rect 19432 25842 19484 25848
rect 19812 25294 19840 25910
rect 19432 25288 19484 25294
rect 19432 25230 19484 25236
rect 19800 25288 19852 25294
rect 19800 25230 19852 25236
rect 19340 24948 19392 24954
rect 19340 24890 19392 24896
rect 19352 24449 19380 24890
rect 19444 24682 19472 25230
rect 19432 24676 19484 24682
rect 19432 24618 19484 24624
rect 19524 24676 19576 24682
rect 19524 24618 19576 24624
rect 19338 24440 19394 24449
rect 19338 24375 19394 24384
rect 19246 24168 19302 24177
rect 19246 24103 19302 24112
rect 18696 23792 18748 23798
rect 18694 23760 18696 23769
rect 18748 23760 18750 23769
rect 18694 23695 18750 23704
rect 19248 23520 19300 23526
rect 19248 23462 19300 23468
rect 19340 23520 19392 23526
rect 19340 23462 19392 23468
rect 19260 23118 19288 23462
rect 19248 23112 19300 23118
rect 19248 23054 19300 23060
rect 19064 23044 19116 23050
rect 19064 22986 19116 22992
rect 19076 22778 19104 22986
rect 19064 22772 19116 22778
rect 19064 22714 19116 22720
rect 19260 22710 19288 23054
rect 19248 22704 19300 22710
rect 19248 22646 19300 22652
rect 19156 22568 19208 22574
rect 19156 22510 19208 22516
rect 19168 22166 19196 22510
rect 19352 22234 19380 23462
rect 19444 22522 19472 24618
rect 19536 24206 19564 24618
rect 19812 24342 19840 25230
rect 19800 24336 19852 24342
rect 19800 24278 19852 24284
rect 19524 24200 19576 24206
rect 19524 24142 19576 24148
rect 19708 24200 19760 24206
rect 19708 24142 19760 24148
rect 19524 24064 19576 24070
rect 19524 24006 19576 24012
rect 19536 22642 19564 24006
rect 19616 23724 19668 23730
rect 19616 23666 19668 23672
rect 19524 22636 19576 22642
rect 19524 22578 19576 22584
rect 19444 22494 19564 22522
rect 19340 22228 19392 22234
rect 19340 22170 19392 22176
rect 19432 22228 19484 22234
rect 19432 22170 19484 22176
rect 19156 22160 19208 22166
rect 19156 22102 19208 22108
rect 19352 22098 19380 22170
rect 18432 22066 18644 22094
rect 19340 22092 19392 22098
rect 18328 21548 18380 21554
rect 18328 21490 18380 21496
rect 18236 21344 18288 21350
rect 18236 21286 18288 21292
rect 17846 21244 18154 21264
rect 17846 21242 17852 21244
rect 17908 21242 17932 21244
rect 17988 21242 18012 21244
rect 18068 21242 18092 21244
rect 18148 21242 18154 21244
rect 17908 21190 17910 21242
rect 18090 21190 18092 21242
rect 17846 21188 17852 21190
rect 17908 21188 17932 21190
rect 17988 21188 18012 21190
rect 18068 21188 18092 21190
rect 18148 21188 18154 21190
rect 17846 21168 18154 21188
rect 18248 20942 18276 21286
rect 18236 20936 18288 20942
rect 18236 20878 18288 20884
rect 18340 20330 18368 21490
rect 18328 20324 18380 20330
rect 18328 20266 18380 20272
rect 17846 20156 18154 20176
rect 17846 20154 17852 20156
rect 17908 20154 17932 20156
rect 17988 20154 18012 20156
rect 18068 20154 18092 20156
rect 18148 20154 18154 20156
rect 17908 20102 17910 20154
rect 18090 20102 18092 20154
rect 17846 20100 17852 20102
rect 17908 20100 17932 20102
rect 17988 20100 18012 20102
rect 18068 20100 18092 20102
rect 18148 20100 18154 20102
rect 17846 20080 18154 20100
rect 17846 19068 18154 19088
rect 17846 19066 17852 19068
rect 17908 19066 17932 19068
rect 17988 19066 18012 19068
rect 18068 19066 18092 19068
rect 18148 19066 18154 19068
rect 17908 19014 17910 19066
rect 18090 19014 18092 19066
rect 17846 19012 17852 19014
rect 17908 19012 17932 19014
rect 17988 19012 18012 19014
rect 18068 19012 18092 19014
rect 18148 19012 18154 19014
rect 17846 18992 18154 19012
rect 17846 17980 18154 18000
rect 17846 17978 17852 17980
rect 17908 17978 17932 17980
rect 17988 17978 18012 17980
rect 18068 17978 18092 17980
rect 18148 17978 18154 17980
rect 17908 17926 17910 17978
rect 18090 17926 18092 17978
rect 17846 17924 17852 17926
rect 17908 17924 17932 17926
rect 17988 17924 18012 17926
rect 18068 17924 18092 17926
rect 18148 17924 18154 17926
rect 17846 17904 18154 17924
rect 17846 16892 18154 16912
rect 17846 16890 17852 16892
rect 17908 16890 17932 16892
rect 17988 16890 18012 16892
rect 18068 16890 18092 16892
rect 18148 16890 18154 16892
rect 17908 16838 17910 16890
rect 18090 16838 18092 16890
rect 17846 16836 17852 16838
rect 17908 16836 17932 16838
rect 17988 16836 18012 16838
rect 18068 16836 18092 16838
rect 18148 16836 18154 16838
rect 17846 16816 18154 16836
rect 17846 15804 18154 15824
rect 17846 15802 17852 15804
rect 17908 15802 17932 15804
rect 17988 15802 18012 15804
rect 18068 15802 18092 15804
rect 18148 15802 18154 15804
rect 17908 15750 17910 15802
rect 18090 15750 18092 15802
rect 17846 15748 17852 15750
rect 17908 15748 17932 15750
rect 17988 15748 18012 15750
rect 18068 15748 18092 15750
rect 18148 15748 18154 15750
rect 17846 15728 18154 15748
rect 17846 14716 18154 14736
rect 17846 14714 17852 14716
rect 17908 14714 17932 14716
rect 17988 14714 18012 14716
rect 18068 14714 18092 14716
rect 18148 14714 18154 14716
rect 17908 14662 17910 14714
rect 18090 14662 18092 14714
rect 17846 14660 17852 14662
rect 17908 14660 17932 14662
rect 17988 14660 18012 14662
rect 18068 14660 18092 14662
rect 18148 14660 18154 14662
rect 17846 14640 18154 14660
rect 17846 13628 18154 13648
rect 17846 13626 17852 13628
rect 17908 13626 17932 13628
rect 17988 13626 18012 13628
rect 18068 13626 18092 13628
rect 18148 13626 18154 13628
rect 17908 13574 17910 13626
rect 18090 13574 18092 13626
rect 17846 13572 17852 13574
rect 17908 13572 17932 13574
rect 17988 13572 18012 13574
rect 18068 13572 18092 13574
rect 18148 13572 18154 13574
rect 17846 13552 18154 13572
rect 17846 12540 18154 12560
rect 17846 12538 17852 12540
rect 17908 12538 17932 12540
rect 17988 12538 18012 12540
rect 18068 12538 18092 12540
rect 18148 12538 18154 12540
rect 17908 12486 17910 12538
rect 18090 12486 18092 12538
rect 17846 12484 17852 12486
rect 17908 12484 17932 12486
rect 17988 12484 18012 12486
rect 18068 12484 18092 12486
rect 18148 12484 18154 12486
rect 17846 12464 18154 12484
rect 17846 11452 18154 11472
rect 17846 11450 17852 11452
rect 17908 11450 17932 11452
rect 17988 11450 18012 11452
rect 18068 11450 18092 11452
rect 18148 11450 18154 11452
rect 17908 11398 17910 11450
rect 18090 11398 18092 11450
rect 17846 11396 17852 11398
rect 17908 11396 17932 11398
rect 17988 11396 18012 11398
rect 18068 11396 18092 11398
rect 18148 11396 18154 11398
rect 17846 11376 18154 11396
rect 17846 10364 18154 10384
rect 17846 10362 17852 10364
rect 17908 10362 17932 10364
rect 17988 10362 18012 10364
rect 18068 10362 18092 10364
rect 18148 10362 18154 10364
rect 17908 10310 17910 10362
rect 18090 10310 18092 10362
rect 17846 10308 17852 10310
rect 17908 10308 17932 10310
rect 17988 10308 18012 10310
rect 18068 10308 18092 10310
rect 18148 10308 18154 10310
rect 17846 10288 18154 10308
rect 17846 9276 18154 9296
rect 17846 9274 17852 9276
rect 17908 9274 17932 9276
rect 17988 9274 18012 9276
rect 18068 9274 18092 9276
rect 18148 9274 18154 9276
rect 17908 9222 17910 9274
rect 18090 9222 18092 9274
rect 17846 9220 17852 9222
rect 17908 9220 17932 9222
rect 17988 9220 18012 9222
rect 18068 9220 18092 9222
rect 18148 9220 18154 9222
rect 17846 9200 18154 9220
rect 17846 8188 18154 8208
rect 17846 8186 17852 8188
rect 17908 8186 17932 8188
rect 17988 8186 18012 8188
rect 18068 8186 18092 8188
rect 18148 8186 18154 8188
rect 17908 8134 17910 8186
rect 18090 8134 18092 8186
rect 17846 8132 17852 8134
rect 17908 8132 17932 8134
rect 17988 8132 18012 8134
rect 18068 8132 18092 8134
rect 18148 8132 18154 8134
rect 17846 8112 18154 8132
rect 17846 7100 18154 7120
rect 17846 7098 17852 7100
rect 17908 7098 17932 7100
rect 17988 7098 18012 7100
rect 18068 7098 18092 7100
rect 18148 7098 18154 7100
rect 17908 7046 17910 7098
rect 18090 7046 18092 7098
rect 17846 7044 17852 7046
rect 17908 7044 17932 7046
rect 17988 7044 18012 7046
rect 18068 7044 18092 7046
rect 18148 7044 18154 7046
rect 17846 7024 18154 7044
rect 17846 6012 18154 6032
rect 17846 6010 17852 6012
rect 17908 6010 17932 6012
rect 17988 6010 18012 6012
rect 18068 6010 18092 6012
rect 18148 6010 18154 6012
rect 17908 5958 17910 6010
rect 18090 5958 18092 6010
rect 17846 5956 17852 5958
rect 17908 5956 17932 5958
rect 17988 5956 18012 5958
rect 18068 5956 18092 5958
rect 18148 5956 18154 5958
rect 17846 5936 18154 5956
rect 17846 4924 18154 4944
rect 17846 4922 17852 4924
rect 17908 4922 17932 4924
rect 17988 4922 18012 4924
rect 18068 4922 18092 4924
rect 18148 4922 18154 4924
rect 17908 4870 17910 4922
rect 18090 4870 18092 4922
rect 17846 4868 17852 4870
rect 17908 4868 17932 4870
rect 17988 4868 18012 4870
rect 18068 4868 18092 4870
rect 18148 4868 18154 4870
rect 17846 4848 18154 4868
rect 17846 3836 18154 3856
rect 17846 3834 17852 3836
rect 17908 3834 17932 3836
rect 17988 3834 18012 3836
rect 18068 3834 18092 3836
rect 18148 3834 18154 3836
rect 17908 3782 17910 3834
rect 18090 3782 18092 3834
rect 17846 3780 17852 3782
rect 17908 3780 17932 3782
rect 17988 3780 18012 3782
rect 18068 3780 18092 3782
rect 18148 3780 18154 3782
rect 17846 3760 18154 3780
rect 18432 3534 18460 22066
rect 19340 22034 19392 22040
rect 19352 21962 19380 22034
rect 19444 22030 19472 22170
rect 19536 22030 19564 22494
rect 19628 22098 19656 23666
rect 19616 22092 19668 22098
rect 19616 22034 19668 22040
rect 19432 22024 19484 22030
rect 19432 21966 19484 21972
rect 19524 22024 19576 22030
rect 19524 21966 19576 21972
rect 19340 21956 19392 21962
rect 19340 21898 19392 21904
rect 18512 21888 18564 21894
rect 18512 21830 18564 21836
rect 18524 20466 18552 21830
rect 19444 21350 19472 21966
rect 19720 21894 19748 24142
rect 19904 23730 19932 26318
rect 20088 25294 20116 31622
rect 20168 31340 20220 31346
rect 20168 31282 20220 31288
rect 20180 30666 20208 31282
rect 20272 31249 20300 33918
rect 20456 33590 20484 34138
rect 20534 34096 20590 34105
rect 20534 34031 20590 34040
rect 20548 33862 20576 34031
rect 20640 33930 20668 35022
rect 21008 34746 21036 35391
rect 21100 35154 21128 35527
rect 21088 35148 21140 35154
rect 21088 35090 21140 35096
rect 20996 34740 21048 34746
rect 20996 34682 21048 34688
rect 21088 34672 21140 34678
rect 21086 34640 21088 34649
rect 21140 34640 21142 34649
rect 21086 34575 21142 34584
rect 20996 34468 21048 34474
rect 20996 34410 21048 34416
rect 20720 34196 20772 34202
rect 20720 34138 20772 34144
rect 20628 33924 20680 33930
rect 20628 33866 20680 33872
rect 20536 33856 20588 33862
rect 20536 33798 20588 33804
rect 20444 33584 20496 33590
rect 20444 33526 20496 33532
rect 20350 33144 20406 33153
rect 20350 33079 20406 33088
rect 20364 31793 20392 33079
rect 20456 32502 20484 33526
rect 20444 32496 20496 32502
rect 20444 32438 20496 32444
rect 20456 31958 20484 32438
rect 20536 32428 20588 32434
rect 20536 32370 20588 32376
rect 20444 31952 20496 31958
rect 20444 31894 20496 31900
rect 20548 31890 20576 32370
rect 20536 31884 20588 31890
rect 20536 31826 20588 31832
rect 20350 31784 20406 31793
rect 20350 31719 20406 31728
rect 20640 31686 20668 33866
rect 20732 33833 20760 34138
rect 20718 33824 20774 33833
rect 20718 33759 20774 33768
rect 20902 33688 20958 33697
rect 20902 33623 20958 33632
rect 20720 33040 20772 33046
rect 20916 33017 20944 33623
rect 20720 32982 20772 32988
rect 20902 33008 20958 33017
rect 20732 32298 20760 32982
rect 20902 32943 20958 32952
rect 20904 32768 20956 32774
rect 20904 32710 20956 32716
rect 20916 32570 20944 32710
rect 21008 32570 21036 34410
rect 21192 33833 21220 36722
rect 21548 36644 21600 36650
rect 21548 36586 21600 36592
rect 21362 36544 21418 36553
rect 21362 36479 21418 36488
rect 21272 36168 21324 36174
rect 21272 36110 21324 36116
rect 21284 35630 21312 36110
rect 21376 35834 21404 36479
rect 21560 36378 21588 36586
rect 21548 36372 21600 36378
rect 21548 36314 21600 36320
rect 21364 35828 21416 35834
rect 21364 35770 21416 35776
rect 21272 35624 21324 35630
rect 21272 35566 21324 35572
rect 21284 35154 21312 35566
rect 21652 35193 21680 40831
rect 22006 40216 22062 40225
rect 22006 40151 22062 40160
rect 22020 39438 22048 40151
rect 22192 39976 22244 39982
rect 22192 39918 22244 39924
rect 21916 39432 21968 39438
rect 21916 39374 21968 39380
rect 22008 39432 22060 39438
rect 22008 39374 22060 39380
rect 21928 38758 21956 39374
rect 22100 39092 22152 39098
rect 22100 39034 22152 39040
rect 22112 38826 22140 39034
rect 22204 38962 22232 39918
rect 22192 38956 22244 38962
rect 22192 38898 22244 38904
rect 22572 38894 22600 41200
rect 22926 40760 22982 40769
rect 22926 40695 22982 40704
rect 22652 40044 22704 40050
rect 22652 39986 22704 39992
rect 22664 39438 22692 39986
rect 22652 39432 22704 39438
rect 22652 39374 22704 39380
rect 22664 39137 22692 39374
rect 22836 39364 22888 39370
rect 22836 39306 22888 39312
rect 22650 39128 22706 39137
rect 22650 39063 22706 39072
rect 22848 39001 22876 39306
rect 22834 38992 22890 39001
rect 22834 38927 22890 38936
rect 22468 38888 22520 38894
rect 22468 38830 22520 38836
rect 22560 38888 22612 38894
rect 22560 38830 22612 38836
rect 22100 38820 22152 38826
rect 22100 38762 22152 38768
rect 21916 38752 21968 38758
rect 21916 38694 21968 38700
rect 22098 38584 22154 38593
rect 22282 38584 22338 38593
rect 22154 38542 22232 38570
rect 22098 38519 22154 38528
rect 21916 38480 21968 38486
rect 21730 38448 21786 38457
rect 21730 38383 21732 38392
rect 21784 38383 21786 38392
rect 21914 38448 21916 38457
rect 21968 38448 21970 38457
rect 21914 38383 21970 38392
rect 21732 38354 21784 38360
rect 22204 38214 22232 38542
rect 22282 38519 22338 38528
rect 22296 38418 22324 38519
rect 22284 38412 22336 38418
rect 22284 38354 22336 38360
rect 22376 38344 22428 38350
rect 22376 38286 22428 38292
rect 22192 38208 22244 38214
rect 22192 38150 22244 38156
rect 22192 37936 22244 37942
rect 22192 37878 22244 37884
rect 22008 37664 22060 37670
rect 22204 37641 22232 37878
rect 22388 37874 22416 38286
rect 22376 37868 22428 37874
rect 22376 37810 22428 37816
rect 22008 37606 22060 37612
rect 22190 37632 22246 37641
rect 21732 37324 21784 37330
rect 21732 37266 21784 37272
rect 21744 36854 21772 37266
rect 22020 36922 22048 37606
rect 22190 37567 22246 37576
rect 22388 37330 22416 37810
rect 22376 37324 22428 37330
rect 22376 37266 22428 37272
rect 22008 36916 22060 36922
rect 22008 36858 22060 36864
rect 21732 36848 21784 36854
rect 21732 36790 21784 36796
rect 21824 36780 21876 36786
rect 21824 36722 21876 36728
rect 21836 36689 21864 36722
rect 21822 36680 21878 36689
rect 21822 36615 21878 36624
rect 22388 36174 22416 37266
rect 22376 36168 22428 36174
rect 22376 36110 22428 36116
rect 22376 36032 22428 36038
rect 22098 36000 22154 36009
rect 22376 35974 22428 35980
rect 22098 35935 22154 35944
rect 22112 35766 22140 35935
rect 22100 35760 22152 35766
rect 22100 35702 22152 35708
rect 22388 35698 22416 35974
rect 22480 35834 22508 38830
rect 22560 38752 22612 38758
rect 22560 38694 22612 38700
rect 22572 36786 22600 38694
rect 22744 38276 22796 38282
rect 22744 38218 22796 38224
rect 22756 36825 22784 38218
rect 22836 37732 22888 37738
rect 22836 37674 22888 37680
rect 22848 36854 22876 37674
rect 22940 36922 22968 40695
rect 23756 39976 23808 39982
rect 23756 39918 23808 39924
rect 23662 39672 23718 39681
rect 23768 39642 23796 39918
rect 23662 39607 23718 39616
rect 23756 39636 23808 39642
rect 23676 39438 23704 39607
rect 23756 39578 23808 39584
rect 23664 39432 23716 39438
rect 23664 39374 23716 39380
rect 24584 39432 24636 39438
rect 24584 39374 24636 39380
rect 23848 39296 23900 39302
rect 23848 39238 23900 39244
rect 23478 39196 23786 39216
rect 23478 39194 23484 39196
rect 23540 39194 23564 39196
rect 23620 39194 23644 39196
rect 23700 39194 23724 39196
rect 23780 39194 23786 39196
rect 23540 39142 23542 39194
rect 23722 39142 23724 39194
rect 23478 39140 23484 39142
rect 23540 39140 23564 39142
rect 23620 39140 23644 39142
rect 23700 39140 23724 39142
rect 23780 39140 23786 39142
rect 23478 39120 23786 39140
rect 23756 38752 23808 38758
rect 23756 38694 23808 38700
rect 23768 38486 23796 38694
rect 23756 38480 23808 38486
rect 23756 38422 23808 38428
rect 23478 38108 23786 38128
rect 23478 38106 23484 38108
rect 23540 38106 23564 38108
rect 23620 38106 23644 38108
rect 23700 38106 23724 38108
rect 23780 38106 23786 38108
rect 23540 38054 23542 38106
rect 23722 38054 23724 38106
rect 23478 38052 23484 38054
rect 23540 38052 23564 38054
rect 23620 38052 23644 38054
rect 23700 38052 23724 38054
rect 23780 38052 23786 38054
rect 23478 38032 23786 38052
rect 23020 38004 23072 38010
rect 23020 37946 23072 37952
rect 23388 38004 23440 38010
rect 23388 37946 23440 37952
rect 23032 37874 23060 37946
rect 23020 37868 23072 37874
rect 23020 37810 23072 37816
rect 22928 36916 22980 36922
rect 22928 36858 22980 36864
rect 22836 36848 22888 36854
rect 22742 36816 22798 36825
rect 22560 36780 22612 36786
rect 22836 36790 22888 36796
rect 22742 36751 22798 36760
rect 22560 36722 22612 36728
rect 23032 36700 23060 37810
rect 23296 37120 23348 37126
rect 23296 37062 23348 37068
rect 23204 36848 23256 36854
rect 23204 36790 23256 36796
rect 22756 36672 23060 36700
rect 22756 36582 22784 36672
rect 22744 36576 22796 36582
rect 22744 36518 22796 36524
rect 22928 36576 22980 36582
rect 22928 36518 22980 36524
rect 23112 36576 23164 36582
rect 23112 36518 23164 36524
rect 22744 36168 22796 36174
rect 22744 36110 22796 36116
rect 22468 35828 22520 35834
rect 22468 35770 22520 35776
rect 22376 35692 22428 35698
rect 22376 35634 22428 35640
rect 22560 35692 22612 35698
rect 22560 35634 22612 35640
rect 21638 35184 21694 35193
rect 21272 35148 21324 35154
rect 21638 35119 21694 35128
rect 21272 35090 21324 35096
rect 21284 34610 21312 35090
rect 22572 34785 22600 35634
rect 22558 34776 22614 34785
rect 22558 34711 22614 34720
rect 21272 34604 21324 34610
rect 22652 34604 22704 34610
rect 21272 34546 21324 34552
rect 22572 34564 22652 34592
rect 22100 34468 22152 34474
rect 22100 34410 22152 34416
rect 21364 34400 21416 34406
rect 21364 34342 21416 34348
rect 21376 34241 21404 34342
rect 21362 34232 21418 34241
rect 21362 34167 21418 34176
rect 21546 34232 21602 34241
rect 21546 34167 21602 34176
rect 21456 33856 21508 33862
rect 21178 33824 21234 33833
rect 21456 33798 21508 33804
rect 21178 33759 21234 33768
rect 21086 33008 21142 33017
rect 21086 32943 21142 32952
rect 21100 32842 21128 32943
rect 21364 32904 21416 32910
rect 21362 32872 21364 32881
rect 21416 32872 21418 32881
rect 21088 32836 21140 32842
rect 21362 32807 21418 32816
rect 21088 32778 21140 32784
rect 20904 32564 20956 32570
rect 20904 32506 20956 32512
rect 20996 32564 21048 32570
rect 20996 32506 21048 32512
rect 21008 32298 21036 32506
rect 20720 32292 20772 32298
rect 20720 32234 20772 32240
rect 20996 32292 21048 32298
rect 20996 32234 21048 32240
rect 20718 32056 20774 32065
rect 20718 31991 20720 32000
rect 20772 31991 20774 32000
rect 20720 31962 20772 31968
rect 21468 31890 21496 33798
rect 21560 33697 21588 34167
rect 21640 33992 21692 33998
rect 21640 33934 21692 33940
rect 21916 33992 21968 33998
rect 21916 33934 21968 33940
rect 21546 33688 21602 33697
rect 21546 33623 21602 33632
rect 21652 33522 21680 33934
rect 21822 33824 21878 33833
rect 21822 33759 21878 33768
rect 21730 33688 21786 33697
rect 21836 33658 21864 33759
rect 21730 33623 21786 33632
rect 21824 33652 21876 33658
rect 21640 33516 21692 33522
rect 21560 33476 21640 33504
rect 21560 32910 21588 33476
rect 21640 33458 21692 33464
rect 21548 32904 21600 32910
rect 21548 32846 21600 32852
rect 21640 32904 21692 32910
rect 21640 32846 21692 32852
rect 21560 32502 21588 32846
rect 21548 32496 21600 32502
rect 21548 32438 21600 32444
rect 21652 32026 21680 32846
rect 21744 32230 21772 33623
rect 21824 33594 21876 33600
rect 21928 33046 21956 33934
rect 22008 33856 22060 33862
rect 22008 33798 22060 33804
rect 21916 33040 21968 33046
rect 21916 32982 21968 32988
rect 21824 32836 21876 32842
rect 21824 32778 21876 32784
rect 21836 32434 21864 32778
rect 21914 32600 21970 32609
rect 21914 32535 21970 32544
rect 21824 32428 21876 32434
rect 21824 32370 21876 32376
rect 21732 32224 21784 32230
rect 21732 32166 21784 32172
rect 21640 32020 21692 32026
rect 21640 31962 21692 31968
rect 21928 31890 21956 32535
rect 20904 31884 20956 31890
rect 20904 31826 20956 31832
rect 21456 31884 21508 31890
rect 21456 31826 21508 31832
rect 21824 31884 21876 31890
rect 21824 31826 21876 31832
rect 21916 31884 21968 31890
rect 21916 31826 21968 31832
rect 20628 31680 20680 31686
rect 20628 31622 20680 31628
rect 20720 31680 20772 31686
rect 20720 31622 20772 31628
rect 20732 31362 20760 31622
rect 20640 31334 20760 31362
rect 20258 31240 20314 31249
rect 20640 31210 20668 31334
rect 20258 31175 20314 31184
rect 20628 31204 20680 31210
rect 20628 31146 20680 31152
rect 20720 31204 20772 31210
rect 20720 31146 20772 31152
rect 20260 30864 20312 30870
rect 20260 30806 20312 30812
rect 20168 30660 20220 30666
rect 20168 30602 20220 30608
rect 20272 30258 20300 30806
rect 20260 30252 20312 30258
rect 20260 30194 20312 30200
rect 20536 30252 20588 30258
rect 20536 30194 20588 30200
rect 20548 30054 20576 30194
rect 20536 30048 20588 30054
rect 20536 29990 20588 29996
rect 20444 29844 20496 29850
rect 20444 29786 20496 29792
rect 20456 29238 20484 29786
rect 20444 29232 20496 29238
rect 20444 29174 20496 29180
rect 20258 29064 20314 29073
rect 20168 29028 20220 29034
rect 20258 28999 20314 29008
rect 20168 28970 20220 28976
rect 20180 27577 20208 28970
rect 20272 28694 20300 28999
rect 20260 28688 20312 28694
rect 20260 28630 20312 28636
rect 20444 28688 20496 28694
rect 20444 28630 20496 28636
rect 20260 28552 20312 28558
rect 20260 28494 20312 28500
rect 20272 28218 20300 28494
rect 20260 28212 20312 28218
rect 20260 28154 20312 28160
rect 20166 27568 20222 27577
rect 20166 27503 20222 27512
rect 20456 25945 20484 28630
rect 20548 28121 20576 29990
rect 20628 29776 20680 29782
rect 20628 29718 20680 29724
rect 20640 29646 20668 29718
rect 20628 29640 20680 29646
rect 20628 29582 20680 29588
rect 20640 28529 20668 29582
rect 20626 28520 20682 28529
rect 20626 28455 20682 28464
rect 20732 28404 20760 31146
rect 20812 30728 20864 30734
rect 20916 30716 20944 31826
rect 21640 31748 21692 31754
rect 21640 31690 21692 31696
rect 21456 31476 21508 31482
rect 21100 31436 21456 31464
rect 21100 31278 21128 31436
rect 21456 31418 21508 31424
rect 21548 31340 21600 31346
rect 21548 31282 21600 31288
rect 21088 31272 21140 31278
rect 21088 31214 21140 31220
rect 21456 31272 21508 31278
rect 21456 31214 21508 31220
rect 21364 31204 21416 31210
rect 21364 31146 21416 31152
rect 21088 31136 21140 31142
rect 21088 31078 21140 31084
rect 21272 31136 21324 31142
rect 21272 31078 21324 31084
rect 20996 30796 21048 30802
rect 20996 30738 21048 30744
rect 20864 30688 20944 30716
rect 20812 30670 20864 30676
rect 21008 30394 21036 30738
rect 20996 30388 21048 30394
rect 20996 30330 21048 30336
rect 20996 30184 21048 30190
rect 20996 30126 21048 30132
rect 20810 30016 20866 30025
rect 20810 29951 20866 29960
rect 20824 28529 20852 29951
rect 21008 29510 21036 30126
rect 21100 29510 21128 31078
rect 21180 30728 21232 30734
rect 21180 30670 21232 30676
rect 20996 29504 21048 29510
rect 20996 29446 21048 29452
rect 21088 29504 21140 29510
rect 21088 29446 21140 29452
rect 20996 29164 21048 29170
rect 20996 29106 21048 29112
rect 20902 29064 20958 29073
rect 20902 28999 20958 29008
rect 20810 28520 20866 28529
rect 20810 28455 20866 28464
rect 20732 28376 20852 28404
rect 20534 28112 20590 28121
rect 20534 28047 20590 28056
rect 20718 28112 20774 28121
rect 20718 28047 20774 28056
rect 20732 27033 20760 28047
rect 20824 27606 20852 28376
rect 20812 27600 20864 27606
rect 20812 27542 20864 27548
rect 20812 27464 20864 27470
rect 20812 27406 20864 27412
rect 20824 27130 20852 27406
rect 20812 27124 20864 27130
rect 20812 27066 20864 27072
rect 20718 27024 20774 27033
rect 20718 26959 20774 26968
rect 20812 26376 20864 26382
rect 20812 26318 20864 26324
rect 20628 26240 20680 26246
rect 20628 26182 20680 26188
rect 20640 25974 20668 26182
rect 20628 25968 20680 25974
rect 20442 25936 20498 25945
rect 20628 25910 20680 25916
rect 20824 25906 20852 26318
rect 20442 25871 20498 25880
rect 20812 25900 20864 25906
rect 20812 25842 20864 25848
rect 20720 25696 20772 25702
rect 20720 25638 20772 25644
rect 20350 25528 20406 25537
rect 20350 25463 20406 25472
rect 20076 25288 20128 25294
rect 20076 25230 20128 25236
rect 20088 25158 20116 25230
rect 20076 25152 20128 25158
rect 20076 25094 20128 25100
rect 20364 24818 20392 25463
rect 20732 25294 20760 25638
rect 20824 25362 20852 25842
rect 20812 25356 20864 25362
rect 20812 25298 20864 25304
rect 20720 25288 20772 25294
rect 20720 25230 20772 25236
rect 20352 24812 20404 24818
rect 20352 24754 20404 24760
rect 20720 24812 20772 24818
rect 20720 24754 20772 24760
rect 20732 24721 20760 24754
rect 20718 24712 20774 24721
rect 20718 24647 20774 24656
rect 20536 24336 20588 24342
rect 20074 24304 20130 24313
rect 20536 24278 20588 24284
rect 20074 24239 20130 24248
rect 20088 24206 20116 24239
rect 20076 24200 20128 24206
rect 20076 24142 20128 24148
rect 19892 23724 19944 23730
rect 19892 23666 19944 23672
rect 20442 23352 20498 23361
rect 20442 23287 20498 23296
rect 20350 23216 20406 23225
rect 20350 23151 20406 23160
rect 20364 22642 20392 23151
rect 20456 22982 20484 23287
rect 20444 22976 20496 22982
rect 20444 22918 20496 22924
rect 20076 22636 20128 22642
rect 20076 22578 20128 22584
rect 20352 22636 20404 22642
rect 20352 22578 20404 22584
rect 19800 22568 19852 22574
rect 19800 22510 19852 22516
rect 19524 21888 19576 21894
rect 19524 21830 19576 21836
rect 19708 21888 19760 21894
rect 19708 21830 19760 21836
rect 19536 21690 19564 21830
rect 19812 21690 19840 22510
rect 19984 22432 20036 22438
rect 20088 22409 20116 22578
rect 20548 22574 20576 24278
rect 20628 24132 20680 24138
rect 20628 24074 20680 24080
rect 20640 22982 20668 24074
rect 20732 24070 20760 24647
rect 20720 24064 20772 24070
rect 20720 24006 20772 24012
rect 20732 23186 20760 24006
rect 20720 23180 20772 23186
rect 20720 23122 20772 23128
rect 20628 22976 20680 22982
rect 20628 22918 20680 22924
rect 20812 22976 20864 22982
rect 20812 22918 20864 22924
rect 20536 22568 20588 22574
rect 20536 22510 20588 22516
rect 20640 22506 20668 22918
rect 20628 22500 20680 22506
rect 20628 22442 20680 22448
rect 19984 22374 20036 22380
rect 20074 22400 20130 22409
rect 19996 22137 20024 22374
rect 20074 22335 20130 22344
rect 19982 22128 20038 22137
rect 19982 22063 20038 22072
rect 19524 21684 19576 21690
rect 19524 21626 19576 21632
rect 19800 21684 19852 21690
rect 19800 21626 19852 21632
rect 19984 21548 20036 21554
rect 19984 21490 20036 21496
rect 19432 21344 19484 21350
rect 19432 21286 19484 21292
rect 19996 21146 20024 21490
rect 20534 21448 20590 21457
rect 20534 21383 20590 21392
rect 20442 21312 20498 21321
rect 20442 21247 20498 21256
rect 19984 21140 20036 21146
rect 19984 21082 20036 21088
rect 20456 20942 20484 21247
rect 20548 21146 20576 21383
rect 20536 21140 20588 21146
rect 20536 21082 20588 21088
rect 20824 21010 20852 22918
rect 20812 21004 20864 21010
rect 20812 20946 20864 20952
rect 19984 20936 20036 20942
rect 19984 20878 20036 20884
rect 20444 20936 20496 20942
rect 20444 20878 20496 20884
rect 18512 20460 18564 20466
rect 18512 20402 18564 20408
rect 19996 20058 20024 20878
rect 19984 20052 20036 20058
rect 19984 19994 20036 20000
rect 20810 19408 20866 19417
rect 20810 19343 20812 19352
rect 20864 19343 20866 19352
rect 20812 19314 20864 19320
rect 20916 12238 20944 28999
rect 21008 27554 21036 29106
rect 21088 28688 21140 28694
rect 21088 28630 21140 28636
rect 21100 28150 21128 28630
rect 21088 28144 21140 28150
rect 21088 28086 21140 28092
rect 21192 28014 21220 30670
rect 21284 28540 21312 31078
rect 21376 30705 21404 31146
rect 21468 30870 21496 31214
rect 21456 30864 21508 30870
rect 21456 30806 21508 30812
rect 21362 30696 21418 30705
rect 21362 30631 21418 30640
rect 21456 29504 21508 29510
rect 21456 29446 21508 29452
rect 21364 29164 21416 29170
rect 21468 29152 21496 29446
rect 21560 29220 21588 31282
rect 21652 31210 21680 31690
rect 21640 31204 21692 31210
rect 21640 31146 21692 31152
rect 21732 30796 21784 30802
rect 21732 30738 21784 30744
rect 21744 30394 21772 30738
rect 21836 30546 21864 31826
rect 22020 31822 22048 33798
rect 22112 33658 22140 34410
rect 22284 33992 22336 33998
rect 22284 33934 22336 33940
rect 22296 33833 22324 33934
rect 22282 33824 22338 33833
rect 22282 33759 22338 33768
rect 22100 33652 22152 33658
rect 22100 33594 22152 33600
rect 22100 33516 22152 33522
rect 22376 33516 22428 33522
rect 22100 33458 22152 33464
rect 22296 33476 22376 33504
rect 22112 33386 22140 33458
rect 22100 33380 22152 33386
rect 22100 33322 22152 33328
rect 22112 32910 22140 33322
rect 22192 33108 22244 33114
rect 22192 33050 22244 33056
rect 22100 32904 22152 32910
rect 22100 32846 22152 32852
rect 22112 32416 22140 32846
rect 22204 32609 22232 33050
rect 22296 32881 22324 33476
rect 22376 33458 22428 33464
rect 22376 33108 22428 33114
rect 22376 33050 22428 33056
rect 22282 32872 22338 32881
rect 22282 32807 22338 32816
rect 22190 32600 22246 32609
rect 22190 32535 22246 32544
rect 22192 32428 22244 32434
rect 22112 32388 22192 32416
rect 22192 32370 22244 32376
rect 22100 32224 22152 32230
rect 22100 32166 22152 32172
rect 22192 32224 22244 32230
rect 22296 32212 22324 32807
rect 22388 32745 22416 33050
rect 22572 33046 22600 34564
rect 22652 34546 22704 34552
rect 22756 33862 22784 36110
rect 22940 36038 22968 36518
rect 22928 36032 22980 36038
rect 22928 35974 22980 35980
rect 22928 35488 22980 35494
rect 22928 35430 22980 35436
rect 22940 34898 22968 35430
rect 23020 34944 23072 34950
rect 22940 34892 23020 34898
rect 22940 34886 23072 34892
rect 22940 34870 23060 34886
rect 22940 33998 22968 34870
rect 23018 34776 23074 34785
rect 23124 34762 23152 36518
rect 23216 35018 23244 36790
rect 23308 36310 23336 37062
rect 23400 36786 23428 37946
rect 23478 37020 23786 37040
rect 23478 37018 23484 37020
rect 23540 37018 23564 37020
rect 23620 37018 23644 37020
rect 23700 37018 23724 37020
rect 23780 37018 23786 37020
rect 23540 36966 23542 37018
rect 23722 36966 23724 37018
rect 23478 36964 23484 36966
rect 23540 36964 23564 36966
rect 23620 36964 23644 36966
rect 23700 36964 23724 36966
rect 23780 36964 23786 36966
rect 23478 36944 23786 36964
rect 23388 36780 23440 36786
rect 23388 36722 23440 36728
rect 23480 36780 23532 36786
rect 23480 36722 23532 36728
rect 23492 36582 23520 36722
rect 23572 36644 23624 36650
rect 23572 36586 23624 36592
rect 23664 36644 23716 36650
rect 23664 36586 23716 36592
rect 23480 36576 23532 36582
rect 23480 36518 23532 36524
rect 23296 36304 23348 36310
rect 23348 36264 23428 36292
rect 23296 36246 23348 36252
rect 23296 35488 23348 35494
rect 23296 35430 23348 35436
rect 23308 35086 23336 35430
rect 23400 35290 23428 36264
rect 23492 36174 23520 36518
rect 23584 36310 23612 36586
rect 23676 36417 23704 36586
rect 23756 36576 23808 36582
rect 23756 36518 23808 36524
rect 23662 36408 23718 36417
rect 23768 36378 23796 36518
rect 23662 36343 23718 36352
rect 23756 36372 23808 36378
rect 23756 36314 23808 36320
rect 23572 36304 23624 36310
rect 23572 36246 23624 36252
rect 23480 36168 23532 36174
rect 23480 36110 23532 36116
rect 23478 35932 23786 35952
rect 23478 35930 23484 35932
rect 23540 35930 23564 35932
rect 23620 35930 23644 35932
rect 23700 35930 23724 35932
rect 23780 35930 23786 35932
rect 23540 35878 23542 35930
rect 23722 35878 23724 35930
rect 23478 35876 23484 35878
rect 23540 35876 23564 35878
rect 23620 35876 23644 35878
rect 23700 35876 23724 35878
rect 23780 35876 23786 35878
rect 23478 35856 23786 35876
rect 23572 35692 23624 35698
rect 23860 35680 23888 39238
rect 24490 38992 24546 39001
rect 24490 38927 24492 38936
rect 24544 38927 24546 38936
rect 24492 38898 24544 38904
rect 24032 38480 24084 38486
rect 24032 38422 24084 38428
rect 24044 38010 24072 38422
rect 24032 38004 24084 38010
rect 24032 37946 24084 37952
rect 24400 37868 24452 37874
rect 24400 37810 24452 37816
rect 24124 37324 24176 37330
rect 24124 37266 24176 37272
rect 23938 36816 23994 36825
rect 23938 36751 23994 36760
rect 23624 35652 23888 35680
rect 23572 35634 23624 35640
rect 23388 35284 23440 35290
rect 23388 35226 23440 35232
rect 23572 35284 23624 35290
rect 23572 35226 23624 35232
rect 23296 35080 23348 35086
rect 23480 35080 23532 35086
rect 23296 35022 23348 35028
rect 23400 35028 23480 35034
rect 23584 35057 23612 35226
rect 23400 35022 23532 35028
rect 23570 35048 23626 35057
rect 23204 35012 23256 35018
rect 23204 34954 23256 34960
rect 23400 35006 23520 35022
rect 23074 34734 23152 34762
rect 23018 34711 23074 34720
rect 22928 33992 22980 33998
rect 22928 33934 22980 33940
rect 22744 33856 22796 33862
rect 22744 33798 22796 33804
rect 22652 33516 22704 33522
rect 22652 33458 22704 33464
rect 22664 33386 22692 33458
rect 22744 33448 22796 33454
rect 22744 33390 22796 33396
rect 22652 33380 22704 33386
rect 22652 33322 22704 33328
rect 22560 33040 22612 33046
rect 22560 32982 22612 32988
rect 22652 33040 22704 33046
rect 22652 32982 22704 32988
rect 22468 32768 22520 32774
rect 22374 32736 22430 32745
rect 22468 32710 22520 32716
rect 22374 32671 22430 32680
rect 22480 32434 22508 32710
rect 22468 32428 22520 32434
rect 22468 32370 22520 32376
rect 22376 32224 22428 32230
rect 22296 32184 22376 32212
rect 22192 32166 22244 32172
rect 22376 32166 22428 32172
rect 22112 31906 22140 32166
rect 22204 32026 22232 32166
rect 22192 32020 22244 32026
rect 22192 31962 22244 31968
rect 22284 32020 22336 32026
rect 22284 31962 22336 31968
rect 22296 31906 22324 31962
rect 22112 31878 22324 31906
rect 22008 31816 22060 31822
rect 22008 31758 22060 31764
rect 22020 31142 22048 31758
rect 22112 31414 22140 31878
rect 22572 31736 22600 32982
rect 22664 32910 22692 32982
rect 22652 32904 22704 32910
rect 22652 32846 22704 32852
rect 22756 32892 22784 33390
rect 22940 33386 22968 33934
rect 23032 33522 23060 34711
rect 23112 34400 23164 34406
rect 23112 34342 23164 34348
rect 23124 34066 23152 34342
rect 23112 34060 23164 34066
rect 23112 34002 23164 34008
rect 23216 33844 23244 34954
rect 23400 34746 23428 35006
rect 23570 34983 23626 34992
rect 23676 35000 23704 35652
rect 23756 35012 23808 35018
rect 23676 34972 23756 35000
rect 23756 34954 23808 34960
rect 23848 34944 23900 34950
rect 23848 34886 23900 34892
rect 23478 34844 23786 34864
rect 23478 34842 23484 34844
rect 23540 34842 23564 34844
rect 23620 34842 23644 34844
rect 23700 34842 23724 34844
rect 23780 34842 23786 34844
rect 23540 34790 23542 34842
rect 23722 34790 23724 34842
rect 23478 34788 23484 34790
rect 23540 34788 23564 34790
rect 23620 34788 23644 34790
rect 23700 34788 23724 34790
rect 23780 34788 23786 34790
rect 23478 34768 23786 34788
rect 23860 34746 23888 34886
rect 23388 34740 23440 34746
rect 23848 34740 23900 34746
rect 23440 34700 23520 34728
rect 23388 34682 23440 34688
rect 23388 34196 23440 34202
rect 23388 34138 23440 34144
rect 23296 33856 23348 33862
rect 23216 33816 23296 33844
rect 23400 33844 23428 34138
rect 23492 33998 23520 34700
rect 23848 34682 23900 34688
rect 23756 34536 23808 34542
rect 23756 34478 23808 34484
rect 23572 34468 23624 34474
rect 23572 34410 23624 34416
rect 23584 34066 23612 34410
rect 23572 34060 23624 34066
rect 23572 34002 23624 34008
rect 23768 33998 23796 34478
rect 23480 33992 23532 33998
rect 23480 33934 23532 33940
rect 23756 33992 23808 33998
rect 23756 33934 23808 33940
rect 23848 33856 23900 33862
rect 23400 33816 23848 33844
rect 23296 33798 23348 33804
rect 23848 33798 23900 33804
rect 23478 33756 23786 33776
rect 23478 33754 23484 33756
rect 23540 33754 23564 33756
rect 23620 33754 23644 33756
rect 23700 33754 23724 33756
rect 23780 33754 23786 33756
rect 23540 33702 23542 33754
rect 23722 33702 23724 33754
rect 23478 33700 23484 33702
rect 23540 33700 23564 33702
rect 23620 33700 23644 33702
rect 23700 33700 23724 33702
rect 23780 33700 23786 33702
rect 23294 33688 23350 33697
rect 23478 33680 23786 33700
rect 23350 33646 23428 33674
rect 23294 33623 23350 33632
rect 23020 33516 23072 33522
rect 23020 33458 23072 33464
rect 23400 33425 23428 33646
rect 23848 33516 23900 33522
rect 23848 33458 23900 33464
rect 23664 33448 23716 33454
rect 23386 33416 23442 33425
rect 22928 33380 22980 33386
rect 23664 33390 23716 33396
rect 23386 33351 23442 33360
rect 22928 33322 22980 33328
rect 23112 33312 23164 33318
rect 23110 33280 23112 33289
rect 23164 33280 23166 33289
rect 23110 33215 23166 33224
rect 22926 33144 22982 33153
rect 22926 33079 22982 33088
rect 22836 32904 22888 32910
rect 22756 32864 22836 32892
rect 22650 32600 22706 32609
rect 22756 32570 22784 32864
rect 22836 32846 22888 32852
rect 22650 32535 22706 32544
rect 22744 32564 22796 32570
rect 22664 32298 22692 32535
rect 22744 32506 22796 32512
rect 22836 32564 22888 32570
rect 22836 32506 22888 32512
rect 22652 32292 22704 32298
rect 22652 32234 22704 32240
rect 22848 31822 22876 32506
rect 22940 32434 22968 33079
rect 23112 32972 23164 32978
rect 23112 32914 23164 32920
rect 23204 32972 23256 32978
rect 23676 32960 23704 33390
rect 23756 32972 23808 32978
rect 23676 32932 23756 32960
rect 23204 32914 23256 32920
rect 23756 32914 23808 32920
rect 23020 32904 23072 32910
rect 23020 32846 23072 32852
rect 23032 32502 23060 32846
rect 23124 32774 23152 32914
rect 23112 32768 23164 32774
rect 23112 32710 23164 32716
rect 23216 32609 23244 32914
rect 23308 32842 23612 32858
rect 23308 32836 23624 32842
rect 23308 32830 23572 32836
rect 23202 32600 23258 32609
rect 23202 32535 23258 32544
rect 23020 32496 23072 32502
rect 23020 32438 23072 32444
rect 23204 32496 23256 32502
rect 23204 32438 23256 32444
rect 22928 32428 22980 32434
rect 22928 32370 22980 32376
rect 22836 31816 22888 31822
rect 22836 31758 22888 31764
rect 22204 31708 22600 31736
rect 22652 31748 22704 31754
rect 22100 31408 22152 31414
rect 22100 31350 22152 31356
rect 22204 31260 22232 31708
rect 22652 31690 22704 31696
rect 22664 31634 22692 31690
rect 22112 31232 22232 31260
rect 22296 31606 22692 31634
rect 22744 31680 22796 31686
rect 22744 31622 22796 31628
rect 22008 31136 22060 31142
rect 22008 31078 22060 31084
rect 22112 30802 22140 31232
rect 22296 30852 22324 31606
rect 22756 31498 22784 31622
rect 22664 31470 22784 31498
rect 22376 31204 22428 31210
rect 22376 31146 22428 31152
rect 22204 30824 22324 30852
rect 22100 30796 22152 30802
rect 22100 30738 22152 30744
rect 22008 30660 22060 30666
rect 22060 30620 22140 30648
rect 22008 30602 22060 30608
rect 21836 30518 22048 30546
rect 21732 30388 21784 30394
rect 21732 30330 21784 30336
rect 21730 30016 21786 30025
rect 21730 29951 21786 29960
rect 21744 29220 21772 29951
rect 21914 29880 21970 29889
rect 21914 29815 21970 29824
rect 21824 29776 21876 29782
rect 21824 29718 21876 29724
rect 21836 29646 21864 29718
rect 21928 29714 21956 29815
rect 21916 29708 21968 29714
rect 21916 29650 21968 29656
rect 21824 29640 21876 29646
rect 21824 29582 21876 29588
rect 22020 29238 22048 30518
rect 21824 29232 21876 29238
rect 21560 29192 21680 29220
rect 21744 29200 21824 29220
rect 22008 29232 22060 29238
rect 21876 29200 21878 29209
rect 21744 29192 21822 29200
rect 21468 29124 21588 29152
rect 21364 29106 21416 29112
rect 21376 28994 21404 29106
rect 21560 29016 21588 29124
rect 21652 29084 21680 29192
rect 22008 29174 22060 29180
rect 21822 29135 21878 29144
rect 21652 29056 21772 29084
rect 21376 28966 21496 28994
rect 21560 28988 21680 29016
rect 21364 28552 21416 28558
rect 21284 28512 21364 28540
rect 21284 28218 21312 28512
rect 21364 28494 21416 28500
rect 21272 28212 21324 28218
rect 21272 28154 21324 28160
rect 21180 28008 21232 28014
rect 21180 27950 21232 27956
rect 21284 27849 21312 28154
rect 21270 27840 21326 27849
rect 21270 27775 21326 27784
rect 21468 27614 21496 28966
rect 21468 27586 21588 27614
rect 21008 27526 21404 27554
rect 20996 27464 21048 27470
rect 21272 27464 21324 27470
rect 20996 27406 21048 27412
rect 21192 27424 21272 27452
rect 21008 27305 21036 27406
rect 20994 27296 21050 27305
rect 20994 27231 21050 27240
rect 21008 26926 21036 27231
rect 21192 27062 21220 27424
rect 21272 27406 21324 27412
rect 21180 27056 21232 27062
rect 21180 26998 21232 27004
rect 21088 26988 21140 26994
rect 21088 26930 21140 26936
rect 20996 26920 21048 26926
rect 20996 26862 21048 26868
rect 21100 26586 21128 26930
rect 21376 26586 21404 27526
rect 21560 27441 21588 27586
rect 21546 27432 21602 27441
rect 21546 27367 21602 27376
rect 21456 27056 21508 27062
rect 21456 26998 21508 27004
rect 21088 26580 21140 26586
rect 21088 26522 21140 26528
rect 21364 26580 21416 26586
rect 21364 26522 21416 26528
rect 21468 26518 21496 26998
rect 21548 26784 21600 26790
rect 21548 26726 21600 26732
rect 21456 26512 21508 26518
rect 21456 26454 21508 26460
rect 21364 26376 21416 26382
rect 21560 26364 21588 26726
rect 21416 26336 21588 26364
rect 21364 26318 21416 26324
rect 21652 26217 21680 28988
rect 21744 28801 21772 29056
rect 21824 29028 21876 29034
rect 21824 28970 21876 28976
rect 21730 28792 21786 28801
rect 21730 28727 21786 28736
rect 21836 27946 21864 28970
rect 21914 28928 21970 28937
rect 21914 28863 21970 28872
rect 21928 28218 21956 28863
rect 22020 28762 22048 29174
rect 22112 29102 22140 30620
rect 22204 30598 22232 30824
rect 22388 30784 22416 31146
rect 22296 30756 22416 30784
rect 22192 30592 22244 30598
rect 22192 30534 22244 30540
rect 22204 30304 22232 30534
rect 22185 30258 22232 30304
rect 22173 30252 22232 30258
rect 22225 30200 22232 30252
rect 22173 30194 22232 30200
rect 22204 29578 22232 30194
rect 22296 29782 22324 30756
rect 22376 30660 22428 30666
rect 22376 30602 22428 30608
rect 22388 30394 22416 30602
rect 22468 30592 22520 30598
rect 22468 30534 22520 30540
rect 22376 30388 22428 30394
rect 22376 30330 22428 30336
rect 22284 29776 22336 29782
rect 22284 29718 22336 29724
rect 22388 29646 22416 30330
rect 22480 30025 22508 30534
rect 22560 30320 22612 30326
rect 22560 30262 22612 30268
rect 22466 30016 22522 30025
rect 22466 29951 22522 29960
rect 22468 29776 22520 29782
rect 22572 29764 22600 30262
rect 22664 30258 22692 31470
rect 22744 31408 22796 31414
rect 22744 31350 22796 31356
rect 22756 31113 22784 31350
rect 22940 31346 22968 32370
rect 23020 32292 23072 32298
rect 23020 32234 23072 32240
rect 22928 31340 22980 31346
rect 22928 31282 22980 31288
rect 22742 31104 22798 31113
rect 22742 31039 22798 31048
rect 22836 30796 22888 30802
rect 22756 30756 22836 30784
rect 22756 30326 22784 30756
rect 22836 30738 22888 30744
rect 22928 30728 22980 30734
rect 22834 30696 22890 30705
rect 22928 30670 22980 30676
rect 22834 30631 22890 30640
rect 22848 30598 22876 30631
rect 22836 30592 22888 30598
rect 22836 30534 22888 30540
rect 22744 30320 22796 30326
rect 22744 30262 22796 30268
rect 22652 30252 22704 30258
rect 22652 30194 22704 30200
rect 22664 29889 22692 30194
rect 22836 30184 22888 30190
rect 22836 30126 22888 30132
rect 22650 29880 22706 29889
rect 22848 29850 22876 30126
rect 22650 29815 22706 29824
rect 22836 29844 22888 29850
rect 22836 29786 22888 29792
rect 22520 29736 22600 29764
rect 22468 29718 22520 29724
rect 22376 29640 22428 29646
rect 22376 29582 22428 29588
rect 22744 29640 22796 29646
rect 22744 29582 22796 29588
rect 22192 29572 22244 29578
rect 22192 29514 22244 29520
rect 22560 29572 22612 29578
rect 22560 29514 22612 29520
rect 22204 29209 22232 29514
rect 22374 29472 22430 29481
rect 22374 29407 22430 29416
rect 22190 29200 22246 29209
rect 22190 29135 22246 29144
rect 22100 29096 22152 29102
rect 22100 29038 22152 29044
rect 22100 28960 22152 28966
rect 22100 28902 22152 28908
rect 22112 28762 22140 28902
rect 22008 28756 22060 28762
rect 22008 28698 22060 28704
rect 22100 28756 22152 28762
rect 22100 28698 22152 28704
rect 22204 28694 22232 29135
rect 22284 28960 22336 28966
rect 22284 28902 22336 28908
rect 22192 28688 22244 28694
rect 22192 28630 22244 28636
rect 22296 28422 22324 28902
rect 22388 28422 22416 29407
rect 22572 29306 22600 29514
rect 22756 29510 22784 29582
rect 22744 29504 22796 29510
rect 22744 29446 22796 29452
rect 22560 29300 22612 29306
rect 22560 29242 22612 29248
rect 22744 29232 22796 29238
rect 22744 29174 22796 29180
rect 22834 29200 22890 29209
rect 22468 29164 22520 29170
rect 22468 29106 22520 29112
rect 22480 28626 22508 29106
rect 22560 29028 22612 29034
rect 22560 28970 22612 28976
rect 22652 29028 22704 29034
rect 22652 28970 22704 28976
rect 22572 28937 22600 28970
rect 22558 28928 22614 28937
rect 22558 28863 22614 28872
rect 22468 28620 22520 28626
rect 22468 28562 22520 28568
rect 22560 28552 22612 28558
rect 22560 28494 22612 28500
rect 22284 28416 22336 28422
rect 22284 28358 22336 28364
rect 22376 28416 22428 28422
rect 22376 28358 22428 28364
rect 21916 28212 21968 28218
rect 21916 28154 21968 28160
rect 22376 28212 22428 28218
rect 22376 28154 22428 28160
rect 22100 28076 22152 28082
rect 22100 28018 22152 28024
rect 22284 28076 22336 28082
rect 22284 28018 22336 28024
rect 21916 28008 21968 28014
rect 21914 27976 21916 27985
rect 21968 27976 21970 27985
rect 21824 27940 21876 27946
rect 21914 27911 21970 27920
rect 21824 27882 21876 27888
rect 22006 27568 22062 27577
rect 21732 27532 21784 27538
rect 22006 27503 22062 27512
rect 21732 27474 21784 27480
rect 21744 27130 21772 27474
rect 21916 27464 21968 27470
rect 21836 27424 21916 27452
rect 21732 27124 21784 27130
rect 21732 27066 21784 27072
rect 21836 26858 21864 27424
rect 21916 27406 21968 27412
rect 21916 27328 21968 27334
rect 21916 27270 21968 27276
rect 21928 26994 21956 27270
rect 21916 26988 21968 26994
rect 21916 26930 21968 26936
rect 21824 26852 21876 26858
rect 21824 26794 21876 26800
rect 21638 26208 21694 26217
rect 21638 26143 21694 26152
rect 21652 25786 21680 26143
rect 22020 25906 22048 27503
rect 22112 27470 22140 28018
rect 22192 27668 22244 27674
rect 22192 27610 22244 27616
rect 22204 27577 22232 27610
rect 22190 27568 22246 27577
rect 22190 27503 22246 27512
rect 22100 27464 22152 27470
rect 22100 27406 22152 27412
rect 22112 26994 22140 27406
rect 22100 26988 22152 26994
rect 22100 26930 22152 26936
rect 22112 26382 22140 26930
rect 22192 26444 22244 26450
rect 22192 26386 22244 26392
rect 22100 26376 22152 26382
rect 22100 26318 22152 26324
rect 22008 25900 22060 25906
rect 22008 25842 22060 25848
rect 21652 25758 22048 25786
rect 21824 25696 21876 25702
rect 21824 25638 21876 25644
rect 21836 25514 21864 25638
rect 21732 25492 21784 25498
rect 21836 25486 21956 25514
rect 22020 25498 22048 25758
rect 21732 25434 21784 25440
rect 21744 25401 21772 25434
rect 21730 25392 21786 25401
rect 21730 25327 21786 25336
rect 21928 25242 21956 25486
rect 22008 25492 22060 25498
rect 22008 25434 22060 25440
rect 22204 25430 22232 26386
rect 22296 26382 22324 28018
rect 22388 27674 22416 28154
rect 22572 28150 22600 28494
rect 22664 28393 22692 28970
rect 22756 28558 22784 29174
rect 22834 29135 22836 29144
rect 22888 29135 22890 29144
rect 22836 29106 22888 29112
rect 22744 28552 22796 28558
rect 22744 28494 22796 28500
rect 22650 28384 22706 28393
rect 22650 28319 22706 28328
rect 22468 28144 22520 28150
rect 22468 28086 22520 28092
rect 22560 28144 22612 28150
rect 22560 28086 22612 28092
rect 22376 27668 22428 27674
rect 22376 27610 22428 27616
rect 22480 26858 22508 28086
rect 22744 28076 22796 28082
rect 22744 28018 22796 28024
rect 22836 28076 22888 28082
rect 22940 28064 22968 30670
rect 23032 29170 23060 32234
rect 23216 32026 23244 32438
rect 23308 32230 23336 32830
rect 23572 32778 23624 32784
rect 23478 32668 23786 32688
rect 23478 32666 23484 32668
rect 23540 32666 23564 32668
rect 23620 32666 23644 32668
rect 23700 32666 23724 32668
rect 23780 32666 23786 32668
rect 23540 32614 23542 32666
rect 23722 32614 23724 32666
rect 23478 32612 23484 32614
rect 23540 32612 23564 32614
rect 23620 32612 23644 32614
rect 23700 32612 23724 32614
rect 23780 32612 23786 32614
rect 23478 32592 23786 32612
rect 23860 32552 23888 33458
rect 23492 32524 23888 32552
rect 23492 32434 23520 32524
rect 23480 32428 23532 32434
rect 23480 32370 23532 32376
rect 23388 32360 23440 32366
rect 23388 32302 23440 32308
rect 23400 32230 23428 32302
rect 23296 32224 23348 32230
rect 23296 32166 23348 32172
rect 23388 32224 23440 32230
rect 23388 32166 23440 32172
rect 23204 32020 23256 32026
rect 23204 31962 23256 31968
rect 23296 32020 23348 32026
rect 23296 31962 23348 31968
rect 23308 31890 23336 31962
rect 23296 31884 23348 31890
rect 23296 31826 23348 31832
rect 23400 31822 23428 32166
rect 23388 31816 23440 31822
rect 23388 31758 23440 31764
rect 23478 31580 23786 31600
rect 23478 31578 23484 31580
rect 23540 31578 23564 31580
rect 23620 31578 23644 31580
rect 23700 31578 23724 31580
rect 23780 31578 23786 31580
rect 23540 31526 23542 31578
rect 23722 31526 23724 31578
rect 23478 31524 23484 31526
rect 23540 31524 23564 31526
rect 23620 31524 23644 31526
rect 23700 31524 23724 31526
rect 23780 31524 23786 31526
rect 23110 31512 23166 31521
rect 23478 31504 23786 31524
rect 23166 31470 23428 31498
rect 23110 31447 23166 31456
rect 23400 31464 23428 31470
rect 23400 31436 23796 31464
rect 23110 31376 23166 31385
rect 23768 31346 23796 31436
rect 23110 31311 23112 31320
rect 23164 31311 23166 31320
rect 23480 31340 23532 31346
rect 23112 31282 23164 31288
rect 23480 31282 23532 31288
rect 23756 31340 23808 31346
rect 23756 31282 23808 31288
rect 23388 30864 23440 30870
rect 23388 30806 23440 30812
rect 23204 30728 23256 30734
rect 23204 30670 23256 30676
rect 23110 30152 23166 30161
rect 23110 30087 23166 30096
rect 23216 30104 23244 30670
rect 23296 30116 23348 30122
rect 23020 29164 23072 29170
rect 23124 29152 23152 30087
rect 23216 30076 23296 30104
rect 23216 29628 23244 30076
rect 23296 30058 23348 30064
rect 23400 29850 23428 30806
rect 23492 30784 23520 31282
rect 23572 31272 23624 31278
rect 23848 31272 23900 31278
rect 23624 31220 23848 31226
rect 23572 31214 23900 31220
rect 23584 31198 23888 31214
rect 23848 31136 23900 31142
rect 23848 31078 23900 31084
rect 23572 30796 23624 30802
rect 23492 30756 23572 30784
rect 23572 30738 23624 30744
rect 23478 30492 23786 30512
rect 23478 30490 23484 30492
rect 23540 30490 23564 30492
rect 23620 30490 23644 30492
rect 23700 30490 23724 30492
rect 23780 30490 23786 30492
rect 23540 30438 23542 30490
rect 23722 30438 23724 30490
rect 23478 30436 23484 30438
rect 23540 30436 23564 30438
rect 23620 30436 23644 30438
rect 23700 30436 23724 30438
rect 23780 30436 23786 30438
rect 23478 30416 23786 30436
rect 23570 30288 23626 30297
rect 23480 30252 23532 30258
rect 23570 30223 23626 30232
rect 23480 30194 23532 30200
rect 23492 29889 23520 30194
rect 23478 29880 23534 29889
rect 23388 29844 23440 29850
rect 23478 29815 23534 29824
rect 23388 29786 23440 29792
rect 23216 29600 23336 29628
rect 23308 29510 23336 29600
rect 23480 29572 23532 29578
rect 23584 29560 23612 30223
rect 23860 29850 23888 31078
rect 23952 30258 23980 36751
rect 24032 36372 24084 36378
rect 24032 36314 24084 36320
rect 24044 32842 24072 36314
rect 24136 36242 24164 37266
rect 24308 37256 24360 37262
rect 24308 37198 24360 37204
rect 24320 36650 24348 37198
rect 24412 36786 24440 37810
rect 24596 37754 24624 39374
rect 25148 38894 25176 41200
rect 25688 39636 25740 39642
rect 25688 39578 25740 39584
rect 25228 39568 25280 39574
rect 25228 39510 25280 39516
rect 25136 38888 25188 38894
rect 25136 38830 25188 38836
rect 25136 38344 25188 38350
rect 25134 38312 25136 38321
rect 25188 38312 25190 38321
rect 24768 38276 24820 38282
rect 25044 38276 25096 38282
rect 24820 38236 25044 38264
rect 24768 38218 24820 38224
rect 25134 38247 25190 38256
rect 25044 38218 25096 38224
rect 24676 38208 24728 38214
rect 24676 38150 24728 38156
rect 24504 37726 24624 37754
rect 24400 36780 24452 36786
rect 24400 36722 24452 36728
rect 24308 36644 24360 36650
rect 24308 36586 24360 36592
rect 24124 36236 24176 36242
rect 24124 36178 24176 36184
rect 24136 35698 24164 36178
rect 24214 35864 24270 35873
rect 24214 35799 24270 35808
rect 24228 35766 24256 35799
rect 24216 35760 24268 35766
rect 24216 35702 24268 35708
rect 24124 35692 24176 35698
rect 24124 35634 24176 35640
rect 24136 33998 24164 35634
rect 24124 33992 24176 33998
rect 24124 33934 24176 33940
rect 24136 33833 24164 33934
rect 24122 33824 24178 33833
rect 24122 33759 24178 33768
rect 24136 33522 24164 33759
rect 24124 33516 24176 33522
rect 24124 33458 24176 33464
rect 24032 32836 24084 32842
rect 24032 32778 24084 32784
rect 24228 32722 24256 35702
rect 24400 34944 24452 34950
rect 24400 34886 24452 34892
rect 24412 34678 24440 34886
rect 24400 34672 24452 34678
rect 24400 34614 24452 34620
rect 24504 33046 24532 37726
rect 24584 37664 24636 37670
rect 24584 37606 24636 37612
rect 24596 35086 24624 37606
rect 24688 37330 24716 38150
rect 24768 37664 24820 37670
rect 24768 37606 24820 37612
rect 24780 37505 24808 37606
rect 24766 37496 24822 37505
rect 24766 37431 24822 37440
rect 24676 37324 24728 37330
rect 24676 37266 24728 37272
rect 24858 37224 24914 37233
rect 24858 37159 24860 37168
rect 24912 37159 24914 37168
rect 24860 37130 24912 37136
rect 24676 36712 24728 36718
rect 24676 36654 24728 36660
rect 24688 35193 24716 36654
rect 24674 35184 24730 35193
rect 24674 35119 24730 35128
rect 24860 35148 24912 35154
rect 24860 35090 24912 35096
rect 25136 35148 25188 35154
rect 25136 35090 25188 35096
rect 24584 35080 24636 35086
rect 24584 35022 24636 35028
rect 24676 35012 24728 35018
rect 24676 34954 24728 34960
rect 24768 35012 24820 35018
rect 24768 34954 24820 34960
rect 24688 34202 24716 34954
rect 24780 34921 24808 34954
rect 24766 34912 24822 34921
rect 24766 34847 24822 34856
rect 24766 34368 24822 34377
rect 24766 34303 24822 34312
rect 24780 34202 24808 34303
rect 24676 34196 24728 34202
rect 24676 34138 24728 34144
rect 24768 34196 24820 34202
rect 24768 34138 24820 34144
rect 24872 34105 24900 35090
rect 24858 34096 24914 34105
rect 25148 34066 25176 35090
rect 24858 34031 24914 34040
rect 25136 34060 25188 34066
rect 24872 33998 24900 34031
rect 25136 34002 25188 34008
rect 24584 33992 24636 33998
rect 24584 33934 24636 33940
rect 24860 33992 24912 33998
rect 24860 33934 24912 33940
rect 24596 33658 24624 33934
rect 25148 33833 25176 34002
rect 25134 33824 25190 33833
rect 25134 33759 25190 33768
rect 24584 33652 24636 33658
rect 24584 33594 24636 33600
rect 24492 33040 24544 33046
rect 24492 32982 24544 32988
rect 24044 32694 24256 32722
rect 23940 30252 23992 30258
rect 23940 30194 23992 30200
rect 23940 30048 23992 30054
rect 23938 30016 23940 30025
rect 23992 30016 23994 30025
rect 23938 29951 23994 29960
rect 23848 29844 23900 29850
rect 23848 29786 23900 29792
rect 23532 29532 23612 29560
rect 23480 29514 23532 29520
rect 23296 29504 23348 29510
rect 23296 29446 23348 29452
rect 23938 29472 23994 29481
rect 23308 29345 23336 29446
rect 23478 29404 23786 29424
rect 23938 29407 23994 29416
rect 23478 29402 23484 29404
rect 23540 29402 23564 29404
rect 23620 29402 23644 29404
rect 23700 29402 23724 29404
rect 23780 29402 23786 29404
rect 23540 29350 23542 29402
rect 23722 29350 23724 29402
rect 23478 29348 23484 29350
rect 23540 29348 23564 29350
rect 23620 29348 23644 29350
rect 23700 29348 23724 29350
rect 23780 29348 23786 29350
rect 23294 29336 23350 29345
rect 23478 29328 23786 29348
rect 23294 29271 23350 29280
rect 23250 29164 23302 29170
rect 23124 29124 23250 29152
rect 23020 29106 23072 29112
rect 23250 29106 23302 29112
rect 23480 29164 23532 29170
rect 23480 29106 23532 29112
rect 23032 29050 23060 29106
rect 23032 29022 23244 29050
rect 23018 28520 23074 28529
rect 23018 28455 23020 28464
rect 23072 28455 23074 28464
rect 23020 28426 23072 28432
rect 23216 28422 23244 29022
rect 23492 28914 23520 29106
rect 23952 28966 23980 29407
rect 23400 28886 23520 28914
rect 23940 28960 23992 28966
rect 23940 28902 23992 28908
rect 23112 28416 23164 28422
rect 23112 28358 23164 28364
rect 23204 28416 23256 28422
rect 23400 28370 23428 28886
rect 23572 28756 23624 28762
rect 23572 28698 23624 28704
rect 23584 28490 23612 28698
rect 23848 28688 23900 28694
rect 23848 28630 23900 28636
rect 23572 28484 23624 28490
rect 23572 28426 23624 28432
rect 23204 28358 23256 28364
rect 23020 28212 23072 28218
rect 23020 28154 23072 28160
rect 23032 28082 23060 28154
rect 23124 28082 23152 28358
rect 22888 28036 22968 28064
rect 23020 28076 23072 28082
rect 22836 28018 22888 28024
rect 23020 28018 23072 28024
rect 23112 28076 23164 28082
rect 23112 28018 23164 28024
rect 22652 27600 22704 27606
rect 22652 27542 22704 27548
rect 22560 27464 22612 27470
rect 22560 27406 22612 27412
rect 22468 26852 22520 26858
rect 22468 26794 22520 26800
rect 22284 26376 22336 26382
rect 22284 26318 22336 26324
rect 22480 26314 22508 26794
rect 22468 26308 22520 26314
rect 22468 26250 22520 26256
rect 22572 25673 22600 27406
rect 22664 26450 22692 27542
rect 22756 27130 22784 28018
rect 22848 27849 22876 28018
rect 22834 27840 22890 27849
rect 22834 27775 22890 27784
rect 23018 27840 23074 27849
rect 23018 27775 23074 27784
rect 22744 27124 22796 27130
rect 22744 27066 22796 27072
rect 22848 26994 22876 27775
rect 23032 27538 23060 27775
rect 23020 27532 23072 27538
rect 23020 27474 23072 27480
rect 23124 27402 23152 28018
rect 23216 27470 23244 28358
rect 23308 28342 23428 28370
rect 23204 27464 23256 27470
rect 23204 27406 23256 27412
rect 23112 27396 23164 27402
rect 23112 27338 23164 27344
rect 22926 27024 22982 27033
rect 22836 26988 22888 26994
rect 22926 26959 22928 26968
rect 22836 26930 22888 26936
rect 22980 26959 22982 26968
rect 22928 26930 22980 26936
rect 23204 26920 23256 26926
rect 23204 26862 23256 26868
rect 23216 26586 23244 26862
rect 23204 26580 23256 26586
rect 23204 26522 23256 26528
rect 23112 26512 23164 26518
rect 23112 26454 23164 26460
rect 22652 26444 22704 26450
rect 22652 26386 22704 26392
rect 22558 25664 22614 25673
rect 22558 25599 22614 25608
rect 22192 25424 22244 25430
rect 22192 25366 22244 25372
rect 23124 25362 23152 26454
rect 23308 26432 23336 28342
rect 23478 28316 23786 28336
rect 23478 28314 23484 28316
rect 23540 28314 23564 28316
rect 23620 28314 23644 28316
rect 23700 28314 23724 28316
rect 23780 28314 23786 28316
rect 23540 28262 23542 28314
rect 23722 28262 23724 28314
rect 23478 28260 23484 28262
rect 23540 28260 23564 28262
rect 23620 28260 23644 28262
rect 23700 28260 23724 28262
rect 23780 28260 23786 28262
rect 23478 28240 23786 28260
rect 23860 28082 23888 28630
rect 23940 28212 23992 28218
rect 23940 28154 23992 28160
rect 23480 28076 23532 28082
rect 23480 28018 23532 28024
rect 23848 28076 23900 28082
rect 23848 28018 23900 28024
rect 23388 27872 23440 27878
rect 23388 27814 23440 27820
rect 23400 27452 23428 27814
rect 23492 27606 23520 28018
rect 23952 27985 23980 28154
rect 23938 27976 23994 27985
rect 23938 27911 23994 27920
rect 23754 27840 23810 27849
rect 23754 27775 23810 27784
rect 23480 27600 23532 27606
rect 23480 27542 23532 27548
rect 23768 27538 23796 27775
rect 23756 27532 23808 27538
rect 23756 27474 23808 27480
rect 23572 27464 23624 27470
rect 23400 27424 23572 27452
rect 23572 27406 23624 27412
rect 23478 27228 23786 27248
rect 23478 27226 23484 27228
rect 23540 27226 23564 27228
rect 23620 27226 23644 27228
rect 23700 27226 23724 27228
rect 23780 27226 23786 27228
rect 23540 27174 23542 27226
rect 23722 27174 23724 27226
rect 23478 27172 23484 27174
rect 23540 27172 23564 27174
rect 23620 27172 23644 27174
rect 23700 27172 23724 27174
rect 23780 27172 23786 27174
rect 23478 27152 23786 27172
rect 23388 26988 23440 26994
rect 23388 26930 23440 26936
rect 23216 26404 23336 26432
rect 23112 25356 23164 25362
rect 23112 25298 23164 25304
rect 23216 25294 23244 26404
rect 23400 26382 23428 26930
rect 23848 26920 23900 26926
rect 23848 26862 23900 26868
rect 23938 26888 23994 26897
rect 23480 26784 23532 26790
rect 23480 26726 23532 26732
rect 23492 26489 23520 26726
rect 23478 26480 23534 26489
rect 23478 26415 23534 26424
rect 23388 26376 23440 26382
rect 23388 26318 23440 26324
rect 23296 26308 23348 26314
rect 23296 26250 23348 26256
rect 23308 25770 23336 26250
rect 23478 26140 23786 26160
rect 23478 26138 23484 26140
rect 23540 26138 23564 26140
rect 23620 26138 23644 26140
rect 23700 26138 23724 26140
rect 23780 26138 23786 26140
rect 23540 26086 23542 26138
rect 23722 26086 23724 26138
rect 23478 26084 23484 26086
rect 23540 26084 23564 26086
rect 23620 26084 23644 26086
rect 23700 26084 23724 26086
rect 23780 26084 23786 26086
rect 23478 26064 23786 26084
rect 23860 25974 23888 26862
rect 23938 26823 23994 26832
rect 23952 26246 23980 26823
rect 23940 26240 23992 26246
rect 23940 26182 23992 26188
rect 23848 25968 23900 25974
rect 23848 25910 23900 25916
rect 23296 25764 23348 25770
rect 23296 25706 23348 25712
rect 23204 25288 23256 25294
rect 21928 25214 22048 25242
rect 23204 25230 23256 25236
rect 21730 24984 21786 24993
rect 21730 24919 21786 24928
rect 21916 24948 21968 24954
rect 21744 24834 21772 24919
rect 21916 24890 21968 24896
rect 21928 24834 21956 24890
rect 21640 24812 21692 24818
rect 21744 24806 21956 24834
rect 22020 24834 22048 25214
rect 22652 25220 22704 25226
rect 22652 25162 22704 25168
rect 22020 24818 22140 24834
rect 22020 24812 22152 24818
rect 22020 24806 22100 24812
rect 21640 24754 21692 24760
rect 21548 24268 21600 24274
rect 21548 24210 21600 24216
rect 21088 24200 21140 24206
rect 21088 24142 21140 24148
rect 20996 23112 21048 23118
rect 20996 23054 21048 23060
rect 21008 22574 21036 23054
rect 20996 22568 21048 22574
rect 20996 22510 21048 22516
rect 21100 22234 21128 24142
rect 21364 24064 21416 24070
rect 21364 24006 21416 24012
rect 21180 23792 21232 23798
rect 21180 23734 21232 23740
rect 21088 22228 21140 22234
rect 21088 22170 21140 22176
rect 21088 21616 21140 21622
rect 21088 21558 21140 21564
rect 21100 21010 21128 21558
rect 21088 21004 21140 21010
rect 21088 20946 21140 20952
rect 21088 20460 21140 20466
rect 21192 20448 21220 23734
rect 21272 23520 21324 23526
rect 21272 23462 21324 23468
rect 21284 20466 21312 23462
rect 21376 23186 21404 24006
rect 21456 23860 21508 23866
rect 21456 23802 21508 23808
rect 21468 23633 21496 23802
rect 21454 23624 21510 23633
rect 21454 23559 21510 23568
rect 21364 23180 21416 23186
rect 21560 23168 21588 24210
rect 21652 24154 21680 24754
rect 21824 24676 21876 24682
rect 21824 24618 21876 24624
rect 21836 24585 21864 24618
rect 21822 24576 21878 24585
rect 21822 24511 21878 24520
rect 21652 24138 21772 24154
rect 21652 24132 21784 24138
rect 21652 24126 21732 24132
rect 21732 24074 21784 24080
rect 21640 24064 21692 24070
rect 21640 24006 21692 24012
rect 21364 23122 21416 23128
rect 21468 23140 21588 23168
rect 21376 22234 21404 23122
rect 21364 22228 21416 22234
rect 21364 22170 21416 22176
rect 21468 22098 21496 23140
rect 21546 23080 21602 23089
rect 21546 23015 21548 23024
rect 21600 23015 21602 23024
rect 21548 22986 21600 22992
rect 21456 22092 21508 22098
rect 21456 22034 21508 22040
rect 21364 22024 21416 22030
rect 21364 21966 21416 21972
rect 21376 21622 21404 21966
rect 21364 21616 21416 21622
rect 21364 21558 21416 21564
rect 21652 21486 21680 24006
rect 21744 23730 21772 24074
rect 22020 23730 22048 24806
rect 22100 24754 22152 24760
rect 22100 24676 22152 24682
rect 22100 24618 22152 24624
rect 21732 23724 21784 23730
rect 21732 23666 21784 23672
rect 22008 23724 22060 23730
rect 22008 23666 22060 23672
rect 22008 23588 22060 23594
rect 22008 23530 22060 23536
rect 22020 23118 22048 23530
rect 21824 23112 21876 23118
rect 21824 23054 21876 23060
rect 22008 23112 22060 23118
rect 22008 23054 22060 23060
rect 21836 22953 21864 23054
rect 21822 22944 21878 22953
rect 21744 22902 21822 22930
rect 21640 21480 21692 21486
rect 21640 21422 21692 21428
rect 21652 20466 21680 21422
rect 21140 20420 21220 20448
rect 21272 20460 21324 20466
rect 21088 20402 21140 20408
rect 21272 20402 21324 20408
rect 21640 20460 21692 20466
rect 21640 20402 21692 20408
rect 21744 19854 21772 22902
rect 21822 22879 21878 22888
rect 21916 22772 21968 22778
rect 21916 22714 21968 22720
rect 21928 22681 21956 22714
rect 21914 22672 21970 22681
rect 21914 22607 21970 22616
rect 22020 22030 22048 23054
rect 22112 22817 22140 24618
rect 22284 24336 22336 24342
rect 22284 24278 22336 24284
rect 22192 24200 22244 24206
rect 22192 24142 22244 24148
rect 22204 23866 22232 24142
rect 22192 23860 22244 23866
rect 22192 23802 22244 23808
rect 22296 23730 22324 24278
rect 22560 24268 22612 24274
rect 22560 24210 22612 24216
rect 22468 24200 22520 24206
rect 22468 24142 22520 24148
rect 22376 24064 22428 24070
rect 22376 24006 22428 24012
rect 22284 23724 22336 23730
rect 22284 23666 22336 23672
rect 22388 23610 22416 24006
rect 22480 23730 22508 24142
rect 22468 23724 22520 23730
rect 22468 23666 22520 23672
rect 22204 23582 22416 23610
rect 22480 23594 22508 23666
rect 22468 23588 22520 23594
rect 22204 23050 22232 23582
rect 22468 23530 22520 23536
rect 22572 23474 22600 24210
rect 22480 23446 22600 23474
rect 22480 23338 22508 23446
rect 22296 23310 22508 23338
rect 22296 23254 22324 23310
rect 22284 23248 22336 23254
rect 22284 23190 22336 23196
rect 22192 23044 22244 23050
rect 22192 22986 22244 22992
rect 22098 22808 22154 22817
rect 22098 22743 22154 22752
rect 22100 22432 22152 22438
rect 22204 22420 22232 22986
rect 22152 22392 22232 22420
rect 22100 22374 22152 22380
rect 21824 22024 21876 22030
rect 21824 21966 21876 21972
rect 22008 22024 22060 22030
rect 22112 22012 22140 22374
rect 22192 22024 22244 22030
rect 22112 21984 22192 22012
rect 22008 21966 22060 21972
rect 22192 21966 22244 21972
rect 21836 21554 21864 21966
rect 21824 21548 21876 21554
rect 21824 21490 21876 21496
rect 21836 20398 21864 21490
rect 22020 20534 22048 21966
rect 22376 21548 22428 21554
rect 22376 21490 22428 21496
rect 22388 21146 22416 21490
rect 22376 21140 22428 21146
rect 22376 21082 22428 21088
rect 22664 20890 22692 25162
rect 23020 24744 23072 24750
rect 23020 24686 23072 24692
rect 22744 24608 22796 24614
rect 22744 24550 22796 24556
rect 22756 23186 22784 24550
rect 22836 24200 22888 24206
rect 22836 24142 22888 24148
rect 22744 23180 22796 23186
rect 22744 23122 22796 23128
rect 22756 22098 22784 23122
rect 22744 22092 22796 22098
rect 22744 22034 22796 22040
rect 22848 21554 22876 24142
rect 22928 24064 22980 24070
rect 22928 24006 22980 24012
rect 22940 23798 22968 24006
rect 22928 23792 22980 23798
rect 22928 23734 22980 23740
rect 23032 23594 23060 24686
rect 23112 24608 23164 24614
rect 23112 24550 23164 24556
rect 23124 24342 23152 24550
rect 23112 24336 23164 24342
rect 23112 24278 23164 24284
rect 23020 23588 23072 23594
rect 23216 23576 23244 25230
rect 23388 25152 23440 25158
rect 23388 25094 23440 25100
rect 23400 24206 23428 25094
rect 23478 25052 23786 25072
rect 23478 25050 23484 25052
rect 23540 25050 23564 25052
rect 23620 25050 23644 25052
rect 23700 25050 23724 25052
rect 23780 25050 23786 25052
rect 23540 24998 23542 25050
rect 23722 24998 23724 25050
rect 23478 24996 23484 24998
rect 23540 24996 23564 24998
rect 23620 24996 23644 24998
rect 23700 24996 23724 24998
rect 23780 24996 23786 24998
rect 23478 24976 23786 24996
rect 23940 24812 23992 24818
rect 23940 24754 23992 24760
rect 23664 24744 23716 24750
rect 23662 24712 23664 24721
rect 23716 24712 23718 24721
rect 23662 24647 23718 24656
rect 23952 24585 23980 24754
rect 23938 24576 23994 24585
rect 23938 24511 23994 24520
rect 23388 24200 23440 24206
rect 23388 24142 23440 24148
rect 23388 24064 23440 24070
rect 23388 24006 23440 24012
rect 23940 24064 23992 24070
rect 23940 24006 23992 24012
rect 23216 23548 23336 23576
rect 23020 23530 23072 23536
rect 22926 23216 22982 23225
rect 22926 23151 22982 23160
rect 23112 23180 23164 23186
rect 22940 23118 22968 23151
rect 23112 23122 23164 23128
rect 23204 23180 23256 23186
rect 23204 23122 23256 23128
rect 22928 23112 22980 23118
rect 22928 23054 22980 23060
rect 23020 23044 23072 23050
rect 23020 22986 23072 22992
rect 23032 22681 23060 22986
rect 23124 22778 23152 23122
rect 23216 22953 23244 23122
rect 23202 22944 23258 22953
rect 23202 22879 23258 22888
rect 23112 22772 23164 22778
rect 23112 22714 23164 22720
rect 23018 22672 23074 22681
rect 22928 22636 22980 22642
rect 23018 22607 23074 22616
rect 22928 22578 22980 22584
rect 22940 22234 22968 22578
rect 23018 22264 23074 22273
rect 22928 22228 22980 22234
rect 23018 22199 23074 22208
rect 23112 22228 23164 22234
rect 22928 22170 22980 22176
rect 23032 21962 23060 22199
rect 23112 22170 23164 22176
rect 23124 22137 23152 22170
rect 23110 22128 23166 22137
rect 23110 22063 23166 22072
rect 23216 22030 23244 22879
rect 23308 22681 23336 23548
rect 23294 22672 23350 22681
rect 23294 22607 23350 22616
rect 23308 22166 23336 22607
rect 23296 22160 23348 22166
rect 23296 22102 23348 22108
rect 23204 22024 23256 22030
rect 23204 21966 23256 21972
rect 23020 21956 23072 21962
rect 23020 21898 23072 21904
rect 22836 21548 22888 21554
rect 22836 21490 22888 21496
rect 23112 21548 23164 21554
rect 23112 21490 23164 21496
rect 22744 21140 22796 21146
rect 22744 21082 22796 21088
rect 22388 20862 22692 20890
rect 22388 20806 22416 20862
rect 22376 20800 22428 20806
rect 22376 20742 22428 20748
rect 22376 20596 22428 20602
rect 22376 20538 22428 20544
rect 22468 20596 22520 20602
rect 22468 20538 22520 20544
rect 22008 20528 22060 20534
rect 22008 20470 22060 20476
rect 21824 20392 21876 20398
rect 21822 20360 21824 20369
rect 21876 20360 21878 20369
rect 21822 20295 21878 20304
rect 21836 20269 21864 20295
rect 22284 20256 22336 20262
rect 22284 20198 22336 20204
rect 22296 19922 22324 20198
rect 22284 19916 22336 19922
rect 22284 19858 22336 19864
rect 21732 19848 21784 19854
rect 21732 19790 21784 19796
rect 22192 19848 22244 19854
rect 22192 19790 22244 19796
rect 22204 19553 22232 19790
rect 22190 19544 22246 19553
rect 21364 19508 21416 19514
rect 22190 19479 22246 19488
rect 21364 19450 21416 19456
rect 21376 19378 21404 19450
rect 21364 19372 21416 19378
rect 21364 19314 21416 19320
rect 22204 18970 22232 19479
rect 22296 19446 22324 19858
rect 22388 19825 22416 20538
rect 22374 19816 22430 19825
rect 22374 19751 22430 19760
rect 22374 19544 22430 19553
rect 22374 19479 22376 19488
rect 22428 19479 22430 19488
rect 22376 19450 22428 19456
rect 22284 19440 22336 19446
rect 22284 19382 22336 19388
rect 22480 19378 22508 20538
rect 22560 20392 22612 20398
rect 22560 20334 22612 20340
rect 22572 19786 22600 20334
rect 22652 20324 22704 20330
rect 22652 20266 22704 20272
rect 22664 19786 22692 20266
rect 22560 19780 22612 19786
rect 22560 19722 22612 19728
rect 22652 19780 22704 19786
rect 22652 19722 22704 19728
rect 22376 19372 22428 19378
rect 22376 19314 22428 19320
rect 22468 19372 22520 19378
rect 22468 19314 22520 19320
rect 22388 18970 22416 19314
rect 22192 18964 22244 18970
rect 22192 18906 22244 18912
rect 22376 18964 22428 18970
rect 22376 18906 22428 18912
rect 22572 18766 22600 19722
rect 21916 18760 21968 18766
rect 21916 18702 21968 18708
rect 22560 18760 22612 18766
rect 22560 18702 22612 18708
rect 21928 18426 21956 18702
rect 22756 18698 22784 21082
rect 22848 20913 22876 21490
rect 23020 21004 23072 21010
rect 23020 20946 23072 20952
rect 22834 20904 22890 20913
rect 22834 20839 22890 20848
rect 23032 20346 23060 20946
rect 23124 20602 23152 21490
rect 23308 21078 23336 22102
rect 23400 22030 23428 24006
rect 23478 23964 23786 23984
rect 23478 23962 23484 23964
rect 23540 23962 23564 23964
rect 23620 23962 23644 23964
rect 23700 23962 23724 23964
rect 23780 23962 23786 23964
rect 23540 23910 23542 23962
rect 23722 23910 23724 23962
rect 23478 23908 23484 23910
rect 23540 23908 23564 23910
rect 23620 23908 23644 23910
rect 23700 23908 23724 23910
rect 23780 23908 23786 23910
rect 23478 23888 23786 23908
rect 23952 23798 23980 24006
rect 23940 23792 23992 23798
rect 23940 23734 23992 23740
rect 23480 23724 23532 23730
rect 23480 23666 23532 23672
rect 23492 23322 23520 23666
rect 23480 23316 23532 23322
rect 23480 23258 23532 23264
rect 23478 22876 23786 22896
rect 23478 22874 23484 22876
rect 23540 22874 23564 22876
rect 23620 22874 23644 22876
rect 23700 22874 23724 22876
rect 23780 22874 23786 22876
rect 23540 22822 23542 22874
rect 23722 22822 23724 22874
rect 23478 22820 23484 22822
rect 23540 22820 23564 22822
rect 23620 22820 23644 22822
rect 23700 22820 23724 22822
rect 23780 22820 23786 22822
rect 23478 22800 23786 22820
rect 23952 22710 23980 23734
rect 23940 22704 23992 22710
rect 23860 22652 23940 22658
rect 23860 22646 23992 22652
rect 23860 22630 23980 22646
rect 23388 22024 23440 22030
rect 23388 21966 23440 21972
rect 23478 21788 23786 21808
rect 23478 21786 23484 21788
rect 23540 21786 23564 21788
rect 23620 21786 23644 21788
rect 23700 21786 23724 21788
rect 23780 21786 23786 21788
rect 23540 21734 23542 21786
rect 23722 21734 23724 21786
rect 23478 21732 23484 21734
rect 23540 21732 23564 21734
rect 23620 21732 23644 21734
rect 23700 21732 23724 21734
rect 23780 21732 23786 21734
rect 23478 21712 23786 21732
rect 23570 21584 23626 21593
rect 23570 21519 23572 21528
rect 23624 21519 23626 21528
rect 23572 21490 23624 21496
rect 23388 21412 23440 21418
rect 23388 21354 23440 21360
rect 23296 21072 23348 21078
rect 23296 21014 23348 21020
rect 23400 20942 23428 21354
rect 23204 20936 23256 20942
rect 23202 20904 23204 20913
rect 23388 20936 23440 20942
rect 23256 20904 23258 20913
rect 23388 20878 23440 20884
rect 23202 20839 23258 20848
rect 23860 20806 23888 22630
rect 23952 22581 23980 22630
rect 23940 22092 23992 22098
rect 23940 22034 23992 22040
rect 23952 21554 23980 22034
rect 23940 21548 23992 21554
rect 23940 21490 23992 21496
rect 23848 20800 23900 20806
rect 23848 20742 23900 20748
rect 23478 20700 23786 20720
rect 23478 20698 23484 20700
rect 23540 20698 23564 20700
rect 23620 20698 23644 20700
rect 23700 20698 23724 20700
rect 23780 20698 23786 20700
rect 23540 20646 23542 20698
rect 23722 20646 23724 20698
rect 23478 20644 23484 20646
rect 23540 20644 23564 20646
rect 23620 20644 23644 20646
rect 23700 20644 23724 20646
rect 23780 20644 23786 20646
rect 23478 20624 23786 20644
rect 23112 20596 23164 20602
rect 23112 20538 23164 20544
rect 23940 20596 23992 20602
rect 23940 20538 23992 20544
rect 23480 20528 23532 20534
rect 23110 20496 23166 20505
rect 23480 20470 23532 20476
rect 23110 20431 23112 20440
rect 23164 20431 23166 20440
rect 23112 20402 23164 20408
rect 22848 20318 23060 20346
rect 22848 20058 22876 20318
rect 22928 20256 22980 20262
rect 22928 20198 22980 20204
rect 22836 20052 22888 20058
rect 22836 19994 22888 20000
rect 22940 19718 22968 20198
rect 23492 19990 23520 20470
rect 23572 20392 23624 20398
rect 23572 20334 23624 20340
rect 23480 19984 23532 19990
rect 23400 19944 23480 19972
rect 23296 19916 23348 19922
rect 23296 19858 23348 19864
rect 22928 19712 22980 19718
rect 22928 19654 22980 19660
rect 22940 18834 22968 19654
rect 23308 19334 23336 19858
rect 23400 19446 23428 19944
rect 23480 19926 23532 19932
rect 23584 19854 23612 20334
rect 23848 20324 23900 20330
rect 23848 20266 23900 20272
rect 23860 19854 23888 20266
rect 23572 19848 23624 19854
rect 23572 19790 23624 19796
rect 23848 19848 23900 19854
rect 23848 19790 23900 19796
rect 23478 19612 23786 19632
rect 23478 19610 23484 19612
rect 23540 19610 23564 19612
rect 23620 19610 23644 19612
rect 23700 19610 23724 19612
rect 23780 19610 23786 19612
rect 23540 19558 23542 19610
rect 23722 19558 23724 19610
rect 23478 19556 23484 19558
rect 23540 19556 23564 19558
rect 23620 19556 23644 19558
rect 23700 19556 23724 19558
rect 23780 19556 23786 19558
rect 23478 19536 23786 19556
rect 23388 19440 23440 19446
rect 23388 19382 23440 19388
rect 23216 19310 23336 19334
rect 23860 19310 23888 19790
rect 23952 19514 23980 20538
rect 23940 19508 23992 19514
rect 23940 19450 23992 19456
rect 23952 19417 23980 19450
rect 23938 19408 23994 19417
rect 23938 19343 23994 19352
rect 23204 19306 23336 19310
rect 23204 19304 23256 19306
rect 23204 19246 23256 19252
rect 23848 19304 23900 19310
rect 23848 19246 23900 19252
rect 22928 18828 22980 18834
rect 22928 18770 22980 18776
rect 23216 18766 23244 19246
rect 23388 19168 23440 19174
rect 23388 19110 23440 19116
rect 23296 18828 23348 18834
rect 23296 18770 23348 18776
rect 23204 18760 23256 18766
rect 23204 18702 23256 18708
rect 22744 18692 22796 18698
rect 22744 18634 22796 18640
rect 21916 18420 21968 18426
rect 21916 18362 21968 18368
rect 22756 18290 22784 18634
rect 23308 18358 23336 18770
rect 23296 18352 23348 18358
rect 23296 18294 23348 18300
rect 22744 18284 22796 18290
rect 22744 18226 22796 18232
rect 23308 17241 23336 18294
rect 23400 18290 23428 19110
rect 23848 18828 23900 18834
rect 23848 18770 23900 18776
rect 23478 18524 23786 18544
rect 23478 18522 23484 18524
rect 23540 18522 23564 18524
rect 23620 18522 23644 18524
rect 23700 18522 23724 18524
rect 23780 18522 23786 18524
rect 23540 18470 23542 18522
rect 23722 18470 23724 18522
rect 23478 18468 23484 18470
rect 23540 18468 23564 18470
rect 23620 18468 23644 18470
rect 23700 18468 23724 18470
rect 23780 18468 23786 18470
rect 23478 18448 23786 18468
rect 23388 18284 23440 18290
rect 23388 18226 23440 18232
rect 23860 18222 23888 18770
rect 23848 18216 23900 18222
rect 23848 18158 23900 18164
rect 23478 17436 23786 17456
rect 23478 17434 23484 17436
rect 23540 17434 23564 17436
rect 23620 17434 23644 17436
rect 23700 17434 23724 17436
rect 23780 17434 23786 17436
rect 23540 17382 23542 17434
rect 23722 17382 23724 17434
rect 23478 17380 23484 17382
rect 23540 17380 23564 17382
rect 23620 17380 23644 17382
rect 23700 17380 23724 17382
rect 23780 17380 23786 17382
rect 23478 17360 23786 17380
rect 23294 17232 23350 17241
rect 23294 17167 23350 17176
rect 23478 16348 23786 16368
rect 23478 16346 23484 16348
rect 23540 16346 23564 16348
rect 23620 16346 23644 16348
rect 23700 16346 23724 16348
rect 23780 16346 23786 16348
rect 23540 16294 23542 16346
rect 23722 16294 23724 16346
rect 23478 16292 23484 16294
rect 23540 16292 23564 16294
rect 23620 16292 23644 16294
rect 23700 16292 23724 16294
rect 23780 16292 23786 16294
rect 23478 16272 23786 16292
rect 23478 15260 23786 15280
rect 23478 15258 23484 15260
rect 23540 15258 23564 15260
rect 23620 15258 23644 15260
rect 23700 15258 23724 15260
rect 23780 15258 23786 15260
rect 23540 15206 23542 15258
rect 23722 15206 23724 15258
rect 23478 15204 23484 15206
rect 23540 15204 23564 15206
rect 23620 15204 23644 15206
rect 23700 15204 23724 15206
rect 23780 15204 23786 15206
rect 23478 15184 23786 15204
rect 23478 14172 23786 14192
rect 23478 14170 23484 14172
rect 23540 14170 23564 14172
rect 23620 14170 23644 14172
rect 23700 14170 23724 14172
rect 23780 14170 23786 14172
rect 23540 14118 23542 14170
rect 23722 14118 23724 14170
rect 23478 14116 23484 14118
rect 23540 14116 23564 14118
rect 23620 14116 23644 14118
rect 23700 14116 23724 14118
rect 23780 14116 23786 14118
rect 23478 14096 23786 14116
rect 23478 13084 23786 13104
rect 23478 13082 23484 13084
rect 23540 13082 23564 13084
rect 23620 13082 23644 13084
rect 23700 13082 23724 13084
rect 23780 13082 23786 13084
rect 23540 13030 23542 13082
rect 23722 13030 23724 13082
rect 23478 13028 23484 13030
rect 23540 13028 23564 13030
rect 23620 13028 23644 13030
rect 23700 13028 23724 13030
rect 23780 13028 23786 13030
rect 23478 13008 23786 13028
rect 20904 12232 20956 12238
rect 20904 12174 20956 12180
rect 23478 11996 23786 12016
rect 23478 11994 23484 11996
rect 23540 11994 23564 11996
rect 23620 11994 23644 11996
rect 23700 11994 23724 11996
rect 23780 11994 23786 11996
rect 23540 11942 23542 11994
rect 23722 11942 23724 11994
rect 23478 11940 23484 11942
rect 23540 11940 23564 11942
rect 23620 11940 23644 11942
rect 23700 11940 23724 11942
rect 23780 11940 23786 11942
rect 23478 11920 23786 11940
rect 23478 10908 23786 10928
rect 23478 10906 23484 10908
rect 23540 10906 23564 10908
rect 23620 10906 23644 10908
rect 23700 10906 23724 10908
rect 23780 10906 23786 10908
rect 23540 10854 23542 10906
rect 23722 10854 23724 10906
rect 23478 10852 23484 10854
rect 23540 10852 23564 10854
rect 23620 10852 23644 10854
rect 23700 10852 23724 10854
rect 23780 10852 23786 10854
rect 23478 10832 23786 10852
rect 23478 9820 23786 9840
rect 23478 9818 23484 9820
rect 23540 9818 23564 9820
rect 23620 9818 23644 9820
rect 23700 9818 23724 9820
rect 23780 9818 23786 9820
rect 23540 9766 23542 9818
rect 23722 9766 23724 9818
rect 23478 9764 23484 9766
rect 23540 9764 23564 9766
rect 23620 9764 23644 9766
rect 23700 9764 23724 9766
rect 23780 9764 23786 9766
rect 23478 9744 23786 9764
rect 23478 8732 23786 8752
rect 23478 8730 23484 8732
rect 23540 8730 23564 8732
rect 23620 8730 23644 8732
rect 23700 8730 23724 8732
rect 23780 8730 23786 8732
rect 23540 8678 23542 8730
rect 23722 8678 23724 8730
rect 23478 8676 23484 8678
rect 23540 8676 23564 8678
rect 23620 8676 23644 8678
rect 23700 8676 23724 8678
rect 23780 8676 23786 8678
rect 23478 8656 23786 8676
rect 23478 7644 23786 7664
rect 23478 7642 23484 7644
rect 23540 7642 23564 7644
rect 23620 7642 23644 7644
rect 23700 7642 23724 7644
rect 23780 7642 23786 7644
rect 23540 7590 23542 7642
rect 23722 7590 23724 7642
rect 23478 7588 23484 7590
rect 23540 7588 23564 7590
rect 23620 7588 23644 7590
rect 23700 7588 23724 7590
rect 23780 7588 23786 7590
rect 23478 7568 23786 7588
rect 23478 6556 23786 6576
rect 23478 6554 23484 6556
rect 23540 6554 23564 6556
rect 23620 6554 23644 6556
rect 23700 6554 23724 6556
rect 23780 6554 23786 6556
rect 23540 6502 23542 6554
rect 23722 6502 23724 6554
rect 23478 6500 23484 6502
rect 23540 6500 23564 6502
rect 23620 6500 23644 6502
rect 23700 6500 23724 6502
rect 23780 6500 23786 6502
rect 23478 6480 23786 6500
rect 24044 5846 24072 32694
rect 24504 32298 24532 32982
rect 24768 32972 24820 32978
rect 24768 32914 24820 32920
rect 24492 32292 24544 32298
rect 24492 32234 24544 32240
rect 24584 31816 24636 31822
rect 24584 31758 24636 31764
rect 24216 31680 24268 31686
rect 24122 31648 24178 31657
rect 24216 31622 24268 31628
rect 24122 31583 24178 31592
rect 24136 31482 24164 31583
rect 24228 31482 24256 31622
rect 24124 31476 24176 31482
rect 24124 31418 24176 31424
rect 24216 31476 24268 31482
rect 24216 31418 24268 31424
rect 24400 31340 24452 31346
rect 24452 31300 24532 31328
rect 24400 31282 24452 31288
rect 24124 31136 24176 31142
rect 24124 31078 24176 31084
rect 24216 31136 24268 31142
rect 24216 31078 24268 31084
rect 24136 30258 24164 31078
rect 24124 30252 24176 30258
rect 24124 30194 24176 30200
rect 24136 29889 24164 30194
rect 24122 29880 24178 29889
rect 24122 29815 24178 29824
rect 24136 29578 24164 29815
rect 24124 29572 24176 29578
rect 24124 29514 24176 29520
rect 24228 28694 24256 31078
rect 24308 30728 24360 30734
rect 24308 30670 24360 30676
rect 24320 29306 24348 30670
rect 24400 30592 24452 30598
rect 24398 30560 24400 30569
rect 24452 30560 24454 30569
rect 24398 30495 24454 30504
rect 24308 29300 24360 29306
rect 24308 29242 24360 29248
rect 24400 29164 24452 29170
rect 24400 29106 24452 29112
rect 24216 28688 24268 28694
rect 24216 28630 24268 28636
rect 24216 28416 24268 28422
rect 24216 28358 24268 28364
rect 24124 28144 24176 28150
rect 24124 28086 24176 28092
rect 24136 27878 24164 28086
rect 24124 27872 24176 27878
rect 24124 27814 24176 27820
rect 24124 27600 24176 27606
rect 24124 27542 24176 27548
rect 24136 25362 24164 27542
rect 24228 25537 24256 28358
rect 24412 28150 24440 29106
rect 24504 28150 24532 31300
rect 24596 29850 24624 31758
rect 24676 31748 24728 31754
rect 24676 31690 24728 31696
rect 24688 31414 24716 31690
rect 24676 31408 24728 31414
rect 24676 31350 24728 31356
rect 24676 30932 24728 30938
rect 24676 30874 24728 30880
rect 24584 29844 24636 29850
rect 24584 29786 24636 29792
rect 24688 29578 24716 30874
rect 24676 29572 24728 29578
rect 24676 29514 24728 29520
rect 24676 29164 24728 29170
rect 24596 29124 24676 29152
rect 24400 28144 24452 28150
rect 24400 28086 24452 28092
rect 24492 28144 24544 28150
rect 24492 28086 24544 28092
rect 24308 28008 24360 28014
rect 24308 27950 24360 27956
rect 24320 27849 24348 27950
rect 24306 27840 24362 27849
rect 24306 27775 24362 27784
rect 24320 27441 24348 27775
rect 24504 27470 24532 28086
rect 24596 28082 24624 29124
rect 24676 29106 24728 29112
rect 24780 29050 24808 32914
rect 25240 32881 25268 39510
rect 25700 37874 25728 39578
rect 25792 38418 25820 41200
rect 26424 40656 26476 40662
rect 26424 40598 26476 40604
rect 26436 39642 26464 40598
rect 26882 39944 26938 39953
rect 26700 39908 26752 39914
rect 26882 39879 26938 39888
rect 26700 39850 26752 39856
rect 26514 39672 26570 39681
rect 26240 39636 26292 39642
rect 26240 39578 26292 39584
rect 26424 39636 26476 39642
rect 26514 39607 26516 39616
rect 26424 39578 26476 39584
rect 26568 39607 26570 39616
rect 26516 39578 26568 39584
rect 26252 39438 26280 39578
rect 26148 39432 26200 39438
rect 26148 39374 26200 39380
rect 26240 39432 26292 39438
rect 26240 39374 26292 39380
rect 26056 39364 26108 39370
rect 26056 39306 26108 39312
rect 25780 38412 25832 38418
rect 25780 38354 25832 38360
rect 25688 37868 25740 37874
rect 25688 37810 25740 37816
rect 25412 37800 25464 37806
rect 25412 37742 25464 37748
rect 25872 37800 25924 37806
rect 25872 37742 25924 37748
rect 25320 37120 25372 37126
rect 25320 37062 25372 37068
rect 25332 36582 25360 37062
rect 25424 36582 25452 37742
rect 25780 36848 25832 36854
rect 25780 36790 25832 36796
rect 25320 36576 25372 36582
rect 25320 36518 25372 36524
rect 25412 36576 25464 36582
rect 25412 36518 25464 36524
rect 25688 36576 25740 36582
rect 25688 36518 25740 36524
rect 25424 36106 25452 36518
rect 25700 36310 25728 36518
rect 25504 36304 25556 36310
rect 25504 36246 25556 36252
rect 25688 36304 25740 36310
rect 25688 36246 25740 36252
rect 25412 36100 25464 36106
rect 25412 36042 25464 36048
rect 25318 35728 25374 35737
rect 25318 35663 25374 35672
rect 25332 35630 25360 35663
rect 25320 35624 25372 35630
rect 25320 35566 25372 35572
rect 25320 35216 25372 35222
rect 25320 35158 25372 35164
rect 25332 34610 25360 35158
rect 25320 34604 25372 34610
rect 25320 34546 25372 34552
rect 25320 34400 25372 34406
rect 25320 34342 25372 34348
rect 25332 33658 25360 34342
rect 25424 33658 25452 36042
rect 25516 35306 25544 36246
rect 25792 35834 25820 36790
rect 25884 36786 25912 37742
rect 25872 36780 25924 36786
rect 25872 36722 25924 36728
rect 25964 36780 26016 36786
rect 25964 36722 26016 36728
rect 25884 36378 25912 36722
rect 25872 36372 25924 36378
rect 25872 36314 25924 36320
rect 25976 36242 26004 36722
rect 25964 36236 26016 36242
rect 25964 36178 26016 36184
rect 25964 36032 26016 36038
rect 25964 35974 26016 35980
rect 25780 35828 25832 35834
rect 25780 35770 25832 35776
rect 25780 35488 25832 35494
rect 25780 35430 25832 35436
rect 25516 35278 25728 35306
rect 25596 34468 25648 34474
rect 25596 34410 25648 34416
rect 25502 34232 25558 34241
rect 25502 34167 25558 34176
rect 25320 33652 25372 33658
rect 25320 33594 25372 33600
rect 25412 33652 25464 33658
rect 25412 33594 25464 33600
rect 25332 33454 25360 33594
rect 25320 33448 25372 33454
rect 25320 33390 25372 33396
rect 25226 32872 25282 32881
rect 25226 32807 25282 32816
rect 25318 32600 25374 32609
rect 25318 32535 25374 32544
rect 25332 32298 25360 32535
rect 25412 32428 25464 32434
rect 25412 32370 25464 32376
rect 25320 32292 25372 32298
rect 25320 32234 25372 32240
rect 24860 32224 24912 32230
rect 24860 32166 24912 32172
rect 24950 32192 25006 32201
rect 24872 32026 24900 32166
rect 24950 32127 25006 32136
rect 24860 32020 24912 32026
rect 24860 31962 24912 31968
rect 24872 31346 24900 31962
rect 24860 31340 24912 31346
rect 24860 31282 24912 31288
rect 24964 30734 24992 32127
rect 25228 31952 25280 31958
rect 25228 31894 25280 31900
rect 25044 31272 25096 31278
rect 25044 31214 25096 31220
rect 24952 30728 25004 30734
rect 24952 30670 25004 30676
rect 24952 30184 25004 30190
rect 24952 30126 25004 30132
rect 24964 29578 24992 30126
rect 25056 29714 25084 31214
rect 25240 30938 25268 31894
rect 25424 31521 25452 32370
rect 25516 32230 25544 34167
rect 25504 32224 25556 32230
rect 25504 32166 25556 32172
rect 25608 31822 25636 34410
rect 25700 32910 25728 35278
rect 25792 33046 25820 35430
rect 25976 34610 26004 35974
rect 25964 34604 26016 34610
rect 25964 34546 26016 34552
rect 26068 34105 26096 39306
rect 26160 36242 26188 39374
rect 26516 38344 26568 38350
rect 26516 38286 26568 38292
rect 26240 37664 26292 37670
rect 26240 37606 26292 37612
rect 26252 37194 26280 37606
rect 26528 37466 26556 38286
rect 26608 37800 26660 37806
rect 26608 37742 26660 37748
rect 26516 37460 26568 37466
rect 26516 37402 26568 37408
rect 26332 37392 26384 37398
rect 26332 37334 26384 37340
rect 26344 37194 26372 37334
rect 26240 37188 26292 37194
rect 26240 37130 26292 37136
rect 26332 37188 26384 37194
rect 26332 37130 26384 37136
rect 26528 36718 26556 37402
rect 26620 36854 26648 37742
rect 26712 36854 26740 39850
rect 26792 39568 26844 39574
rect 26792 39510 26844 39516
rect 26804 39098 26832 39510
rect 26792 39092 26844 39098
rect 26792 39034 26844 39040
rect 26896 39001 26924 39879
rect 27080 39522 27108 41200
rect 27252 40248 27304 40254
rect 27252 40190 27304 40196
rect 27080 39506 27200 39522
rect 27080 39500 27212 39506
rect 27080 39494 27160 39500
rect 27160 39442 27212 39448
rect 26976 39432 27028 39438
rect 26976 39374 27028 39380
rect 26882 38992 26938 39001
rect 26882 38927 26938 38936
rect 26988 38729 27016 39374
rect 27264 39030 27292 40190
rect 27896 39840 27948 39846
rect 27896 39782 27948 39788
rect 27908 39030 27936 39782
rect 27252 39024 27304 39030
rect 27252 38966 27304 38972
rect 27896 39024 27948 39030
rect 27896 38966 27948 38972
rect 26974 38720 27030 38729
rect 26974 38655 27030 38664
rect 27160 37256 27212 37262
rect 27160 37198 27212 37204
rect 26608 36848 26660 36854
rect 26608 36790 26660 36796
rect 26700 36848 26752 36854
rect 26700 36790 26752 36796
rect 26516 36712 26568 36718
rect 26516 36654 26568 36660
rect 26148 36236 26200 36242
rect 26148 36178 26200 36184
rect 26528 36038 26556 36654
rect 26620 36106 26648 36790
rect 27172 36718 27200 37198
rect 27160 36712 27212 36718
rect 27160 36654 27212 36660
rect 26608 36100 26660 36106
rect 26608 36042 26660 36048
rect 26516 36032 26568 36038
rect 26516 35974 26568 35980
rect 26238 35728 26294 35737
rect 27172 35698 27200 36654
rect 26238 35663 26240 35672
rect 26292 35663 26294 35672
rect 27068 35692 27120 35698
rect 26240 35634 26292 35640
rect 27068 35634 27120 35640
rect 27160 35692 27212 35698
rect 27160 35634 27212 35640
rect 26252 35329 26280 35634
rect 26700 35556 26752 35562
rect 26700 35498 26752 35504
rect 26238 35320 26294 35329
rect 26238 35255 26294 35264
rect 26712 35154 26740 35498
rect 27080 35222 27108 35634
rect 27068 35216 27120 35222
rect 27068 35158 27120 35164
rect 26700 35148 26752 35154
rect 26700 35090 26752 35096
rect 26424 35080 26476 35086
rect 26424 35022 26476 35028
rect 26148 34944 26200 34950
rect 26148 34886 26200 34892
rect 26160 34746 26188 34886
rect 26148 34740 26200 34746
rect 26148 34682 26200 34688
rect 26054 34096 26110 34105
rect 25976 34054 26054 34082
rect 25976 33289 26004 34054
rect 26054 34031 26110 34040
rect 26056 33856 26108 33862
rect 26056 33798 26108 33804
rect 26068 33522 26096 33798
rect 26056 33516 26108 33522
rect 26056 33458 26108 33464
rect 26068 33386 26096 33458
rect 26056 33380 26108 33386
rect 26056 33322 26108 33328
rect 25962 33280 26018 33289
rect 25962 33215 26018 33224
rect 26146 33280 26202 33289
rect 26146 33215 26202 33224
rect 25780 33040 25832 33046
rect 25780 32982 25832 32988
rect 25688 32904 25740 32910
rect 25688 32846 25740 32852
rect 26160 32774 26188 33215
rect 26148 32768 26200 32774
rect 26148 32710 26200 32716
rect 25780 32428 25832 32434
rect 25780 32370 25832 32376
rect 25504 31816 25556 31822
rect 25504 31758 25556 31764
rect 25596 31816 25648 31822
rect 25596 31758 25648 31764
rect 25410 31512 25466 31521
rect 25410 31447 25466 31456
rect 25412 31340 25464 31346
rect 25412 31282 25464 31288
rect 25228 30932 25280 30938
rect 25228 30874 25280 30880
rect 25424 30870 25452 31282
rect 25136 30864 25188 30870
rect 25136 30806 25188 30812
rect 25412 30864 25464 30870
rect 25412 30806 25464 30812
rect 25148 30326 25176 30806
rect 25320 30660 25372 30666
rect 25320 30602 25372 30608
rect 25412 30660 25464 30666
rect 25412 30602 25464 30608
rect 25136 30320 25188 30326
rect 25136 30262 25188 30268
rect 25044 29708 25096 29714
rect 25044 29650 25096 29656
rect 24952 29572 25004 29578
rect 24952 29514 25004 29520
rect 24688 29022 24808 29050
rect 24688 28422 24716 29022
rect 24950 28792 25006 28801
rect 24950 28727 25006 28736
rect 24768 28484 24820 28490
rect 24768 28426 24820 28432
rect 24676 28416 24728 28422
rect 24676 28358 24728 28364
rect 24584 28076 24636 28082
rect 24584 28018 24636 28024
rect 24676 28076 24728 28082
rect 24676 28018 24728 28024
rect 24688 27606 24716 28018
rect 24676 27600 24728 27606
rect 24676 27542 24728 27548
rect 24492 27464 24544 27470
rect 24306 27432 24362 27441
rect 24492 27406 24544 27412
rect 24306 27367 24362 27376
rect 24400 27124 24452 27130
rect 24400 27066 24452 27072
rect 24308 27056 24360 27062
rect 24308 26998 24360 27004
rect 24320 26586 24348 26998
rect 24308 26580 24360 26586
rect 24308 26522 24360 26528
rect 24214 25528 24270 25537
rect 24214 25463 24270 25472
rect 24124 25356 24176 25362
rect 24124 25298 24176 25304
rect 24412 25226 24440 27066
rect 24676 25424 24728 25430
rect 24676 25366 24728 25372
rect 24400 25220 24452 25226
rect 24400 25162 24452 25168
rect 24124 25152 24176 25158
rect 24124 25094 24176 25100
rect 24136 24070 24164 25094
rect 24688 24449 24716 25366
rect 24674 24440 24730 24449
rect 24674 24375 24730 24384
rect 24124 24064 24176 24070
rect 24124 24006 24176 24012
rect 24124 23724 24176 23730
rect 24124 23666 24176 23672
rect 24136 22982 24164 23666
rect 24492 23656 24544 23662
rect 24492 23598 24544 23604
rect 24214 23080 24270 23089
rect 24214 23015 24270 23024
rect 24124 22976 24176 22982
rect 24124 22918 24176 22924
rect 24124 22024 24176 22030
rect 24124 21966 24176 21972
rect 24136 20602 24164 21966
rect 24124 20596 24176 20602
rect 24124 20538 24176 20544
rect 24124 20392 24176 20398
rect 24122 20360 24124 20369
rect 24176 20360 24178 20369
rect 24122 20295 24178 20304
rect 24228 19496 24256 23015
rect 24400 22636 24452 22642
rect 24400 22578 24452 22584
rect 24308 22500 24360 22506
rect 24308 22442 24360 22448
rect 24320 22030 24348 22442
rect 24308 22024 24360 22030
rect 24308 21966 24360 21972
rect 24412 21894 24440 22578
rect 24504 22438 24532 23598
rect 24676 23520 24728 23526
rect 24676 23462 24728 23468
rect 24584 22636 24636 22642
rect 24584 22578 24636 22584
rect 24596 22545 24624 22578
rect 24582 22536 24638 22545
rect 24582 22471 24638 22480
rect 24492 22432 24544 22438
rect 24492 22374 24544 22380
rect 24596 22030 24624 22471
rect 24584 22024 24636 22030
rect 24584 21966 24636 21972
rect 24400 21888 24452 21894
rect 24400 21830 24452 21836
rect 24400 21684 24452 21690
rect 24400 21626 24452 21632
rect 24306 21584 24362 21593
rect 24306 21519 24308 21528
rect 24360 21519 24362 21528
rect 24308 21490 24360 21496
rect 24308 21140 24360 21146
rect 24308 21082 24360 21088
rect 24320 20602 24348 21082
rect 24308 20596 24360 20602
rect 24308 20538 24360 20544
rect 24228 19468 24348 19496
rect 24216 19372 24268 19378
rect 24216 19314 24268 19320
rect 24228 18766 24256 19314
rect 24320 18834 24348 19468
rect 24412 19310 24440 21626
rect 24492 21548 24544 21554
rect 24492 21490 24544 21496
rect 24504 20534 24532 21490
rect 24596 21486 24624 21966
rect 24584 21480 24636 21486
rect 24584 21422 24636 21428
rect 24596 21049 24624 21422
rect 24688 21078 24716 23462
rect 24780 21865 24808 28426
rect 24964 28082 24992 28727
rect 25332 28082 25360 30602
rect 25424 30122 25452 30602
rect 25516 30258 25544 31758
rect 25608 30802 25636 31758
rect 25688 31680 25740 31686
rect 25688 31622 25740 31628
rect 25700 31113 25728 31622
rect 25686 31104 25742 31113
rect 25686 31039 25742 31048
rect 25596 30796 25648 30802
rect 25596 30738 25648 30744
rect 25608 30258 25636 30738
rect 25504 30252 25556 30258
rect 25504 30194 25556 30200
rect 25596 30252 25648 30258
rect 25596 30194 25648 30200
rect 25412 30116 25464 30122
rect 25412 30058 25464 30064
rect 25412 29640 25464 29646
rect 25412 29582 25464 29588
rect 25504 29640 25556 29646
rect 25504 29582 25556 29588
rect 25424 29306 25452 29582
rect 25412 29300 25464 29306
rect 25412 29242 25464 29248
rect 24952 28076 25004 28082
rect 24952 28018 25004 28024
rect 25320 28076 25372 28082
rect 25320 28018 25372 28024
rect 24964 27470 24992 28018
rect 25136 28008 25188 28014
rect 25136 27950 25188 27956
rect 24952 27464 25004 27470
rect 24952 27406 25004 27412
rect 24964 27130 24992 27406
rect 25148 27402 25176 27950
rect 25332 27713 25360 28018
rect 25412 28008 25464 28014
rect 25412 27950 25464 27956
rect 25318 27704 25374 27713
rect 25318 27639 25374 27648
rect 25136 27396 25188 27402
rect 25136 27338 25188 27344
rect 24952 27124 25004 27130
rect 24952 27066 25004 27072
rect 25136 25764 25188 25770
rect 25136 25706 25188 25712
rect 25148 25498 25176 25706
rect 25136 25492 25188 25498
rect 25136 25434 25188 25440
rect 25318 25392 25374 25401
rect 25318 25327 25374 25336
rect 25332 25294 25360 25327
rect 25320 25288 25372 25294
rect 25320 25230 25372 25236
rect 25424 24818 25452 27950
rect 25516 26625 25544 29582
rect 25700 28966 25728 31039
rect 25792 30870 25820 32370
rect 26436 32298 26464 35022
rect 26516 33992 26568 33998
rect 26516 33934 26568 33940
rect 26424 32292 26476 32298
rect 26424 32234 26476 32240
rect 26330 32056 26386 32065
rect 26330 31991 26386 32000
rect 26344 31958 26372 31991
rect 26332 31952 26384 31958
rect 26332 31894 26384 31900
rect 26148 31884 26200 31890
rect 26148 31826 26200 31832
rect 26056 31748 26108 31754
rect 26056 31690 26108 31696
rect 25780 30864 25832 30870
rect 25780 30806 25832 30812
rect 25964 30864 26016 30870
rect 25964 30806 26016 30812
rect 25780 30728 25832 30734
rect 25780 30670 25832 30676
rect 25792 30326 25820 30670
rect 25780 30320 25832 30326
rect 25780 30262 25832 30268
rect 25778 30152 25834 30161
rect 25778 30087 25834 30096
rect 25872 30116 25924 30122
rect 25688 28960 25740 28966
rect 25688 28902 25740 28908
rect 25792 27520 25820 30087
rect 25872 30058 25924 30064
rect 25884 29578 25912 30058
rect 25976 30036 26004 30806
rect 26068 30705 26096 31690
rect 26054 30696 26110 30705
rect 26054 30631 26110 30640
rect 26068 30190 26096 30631
rect 26056 30184 26108 30190
rect 26056 30126 26108 30132
rect 25976 30008 26096 30036
rect 25872 29572 25924 29578
rect 25872 29514 25924 29520
rect 25964 29504 26016 29510
rect 25964 29446 26016 29452
rect 25976 29170 26004 29446
rect 25964 29164 26016 29170
rect 25964 29106 26016 29112
rect 26068 27962 26096 30008
rect 26160 29170 26188 31826
rect 26238 31512 26294 31521
rect 26238 31447 26294 31456
rect 26252 31142 26280 31447
rect 26240 31136 26292 31142
rect 26240 31078 26292 31084
rect 26344 30802 26372 31894
rect 26332 30796 26384 30802
rect 26332 30738 26384 30744
rect 26528 30734 26556 33934
rect 27264 33862 27292 38966
rect 28368 38894 28396 41200
rect 28908 39296 28960 39302
rect 28908 39238 28960 39244
rect 27712 38888 27764 38894
rect 27710 38856 27712 38865
rect 28356 38888 28408 38894
rect 27764 38856 27766 38865
rect 27528 38820 27580 38826
rect 28356 38830 28408 38836
rect 28448 38888 28500 38894
rect 28448 38830 28500 38836
rect 27710 38791 27766 38800
rect 27528 38762 27580 38768
rect 27540 38350 27568 38762
rect 28262 38584 28318 38593
rect 28262 38519 28318 38528
rect 27710 38448 27766 38457
rect 27710 38383 27766 38392
rect 27528 38344 27580 38350
rect 27528 38286 27580 38292
rect 27540 37874 27568 38286
rect 27528 37868 27580 37874
rect 27528 37810 27580 37816
rect 27620 36032 27672 36038
rect 27620 35974 27672 35980
rect 27632 35086 27660 35974
rect 27620 35080 27672 35086
rect 27620 35022 27672 35028
rect 27436 34944 27488 34950
rect 27488 34892 27568 34898
rect 27436 34886 27568 34892
rect 27448 34870 27568 34886
rect 27344 34672 27396 34678
rect 27344 34614 27396 34620
rect 27356 33930 27384 34614
rect 27436 34536 27488 34542
rect 27436 34478 27488 34484
rect 27344 33924 27396 33930
rect 27344 33866 27396 33872
rect 27252 33856 27304 33862
rect 27252 33798 27304 33804
rect 27252 33584 27304 33590
rect 27356 33561 27384 33866
rect 27252 33526 27304 33532
rect 27342 33552 27398 33561
rect 27264 32978 27292 33526
rect 27342 33487 27398 33496
rect 27448 33454 27476 34478
rect 27540 34474 27568 34870
rect 27620 34604 27672 34610
rect 27620 34546 27672 34552
rect 27528 34468 27580 34474
rect 27528 34410 27580 34416
rect 27540 33590 27568 34410
rect 27528 33584 27580 33590
rect 27528 33526 27580 33532
rect 27436 33448 27488 33454
rect 27436 33390 27488 33396
rect 27448 33046 27476 33390
rect 27436 33040 27488 33046
rect 27436 32982 27488 32988
rect 27252 32972 27304 32978
rect 27252 32914 27304 32920
rect 27632 32586 27660 34546
rect 27264 32558 27660 32586
rect 27264 32366 27292 32558
rect 27252 32360 27304 32366
rect 27252 32302 27304 32308
rect 27620 32360 27672 32366
rect 27620 32302 27672 32308
rect 26884 31816 26936 31822
rect 26804 31776 26884 31804
rect 26608 31680 26660 31686
rect 26608 31622 26660 31628
rect 26620 30734 26648 31622
rect 26516 30728 26568 30734
rect 26516 30670 26568 30676
rect 26608 30728 26660 30734
rect 26608 30670 26660 30676
rect 26528 30190 26556 30670
rect 26516 30184 26568 30190
rect 26516 30126 26568 30132
rect 26330 29744 26386 29753
rect 26330 29679 26386 29688
rect 26344 29646 26372 29679
rect 26332 29640 26384 29646
rect 26332 29582 26384 29588
rect 26148 29164 26200 29170
rect 26148 29106 26200 29112
rect 26608 29164 26660 29170
rect 26608 29106 26660 29112
rect 26160 28218 26188 29106
rect 26620 28529 26648 29106
rect 26330 28520 26386 28529
rect 26330 28455 26386 28464
rect 26606 28520 26662 28529
rect 26606 28455 26662 28464
rect 26344 28218 26372 28455
rect 26148 28212 26200 28218
rect 26148 28154 26200 28160
rect 26332 28212 26384 28218
rect 26332 28154 26384 28160
rect 26332 28076 26384 28082
rect 26332 28018 26384 28024
rect 26240 28008 26292 28014
rect 26068 27934 26188 27962
rect 26240 27950 26292 27956
rect 25872 27872 25924 27878
rect 25872 27814 25924 27820
rect 25700 27492 25820 27520
rect 25502 26616 25558 26625
rect 25502 26551 25558 26560
rect 25596 26308 25648 26314
rect 25596 26250 25648 26256
rect 25608 26042 25636 26250
rect 25596 26036 25648 26042
rect 25596 25978 25648 25984
rect 25502 25528 25558 25537
rect 25502 25463 25504 25472
rect 25556 25463 25558 25472
rect 25504 25434 25556 25440
rect 25412 24812 25464 24818
rect 25412 24754 25464 24760
rect 25596 24812 25648 24818
rect 25596 24754 25648 24760
rect 25608 24410 25636 24754
rect 25596 24404 25648 24410
rect 25596 24346 25648 24352
rect 25700 23798 25728 27492
rect 25884 27470 25912 27814
rect 25962 27704 26018 27713
rect 25962 27639 26018 27648
rect 25976 27470 26004 27639
rect 26160 27606 26188 27934
rect 26252 27674 26280 27950
rect 26240 27668 26292 27674
rect 26240 27610 26292 27616
rect 26148 27600 26200 27606
rect 26148 27542 26200 27548
rect 26252 27470 26280 27610
rect 26344 27470 26372 28018
rect 26620 27849 26648 28455
rect 26606 27840 26662 27849
rect 26606 27775 26662 27784
rect 25872 27464 25924 27470
rect 25872 27406 25924 27412
rect 25964 27464 26016 27470
rect 25964 27406 26016 27412
rect 26240 27464 26292 27470
rect 26240 27406 26292 27412
rect 26332 27464 26384 27470
rect 26332 27406 26384 27412
rect 25780 27396 25832 27402
rect 25780 27338 25832 27344
rect 25792 26994 25820 27338
rect 25780 26988 25832 26994
rect 25780 26930 25832 26936
rect 25964 26988 26016 26994
rect 25964 26930 26016 26936
rect 25792 26586 25820 26930
rect 25780 26580 25832 26586
rect 25780 26522 25832 26528
rect 25976 25702 26004 26930
rect 26056 26580 26108 26586
rect 26056 26522 26108 26528
rect 26068 25906 26096 26522
rect 26056 25900 26108 25906
rect 26056 25842 26108 25848
rect 25964 25696 26016 25702
rect 25964 25638 26016 25644
rect 25976 25430 26004 25638
rect 26068 25498 26096 25842
rect 26056 25492 26108 25498
rect 26056 25434 26108 25440
rect 25964 25424 26016 25430
rect 25964 25366 26016 25372
rect 26344 25362 26372 27406
rect 26424 25492 26476 25498
rect 26424 25434 26476 25440
rect 26056 25356 26108 25362
rect 26056 25298 26108 25304
rect 26332 25356 26384 25362
rect 26332 25298 26384 25304
rect 26068 25226 26096 25298
rect 26056 25220 26108 25226
rect 26056 25162 26108 25168
rect 26436 24954 26464 25434
rect 26620 25430 26648 27775
rect 26804 26874 26832 31776
rect 26884 31758 26936 31764
rect 27068 31816 27120 31822
rect 27068 31758 27120 31764
rect 27080 31482 27108 31758
rect 27158 31648 27214 31657
rect 27158 31583 27214 31592
rect 27068 31476 27120 31482
rect 27068 31418 27120 31424
rect 27172 30734 27200 31583
rect 27436 31476 27488 31482
rect 27436 31418 27488 31424
rect 27252 31136 27304 31142
rect 27252 31078 27304 31084
rect 27160 30728 27212 30734
rect 27160 30670 27212 30676
rect 27160 30184 27212 30190
rect 27160 30126 27212 30132
rect 26882 29744 26938 29753
rect 27066 29744 27122 29753
rect 26938 29702 27016 29730
rect 26882 29679 26938 29688
rect 26882 29608 26938 29617
rect 26882 29543 26884 29552
rect 26936 29543 26938 29552
rect 26884 29514 26936 29520
rect 26988 28506 27016 29702
rect 27066 29679 27122 29688
rect 27080 29646 27108 29679
rect 27068 29640 27120 29646
rect 27068 29582 27120 29588
rect 27068 29232 27120 29238
rect 27172 29220 27200 30126
rect 27120 29192 27200 29220
rect 27068 29174 27120 29180
rect 27264 28994 27292 31078
rect 27344 30592 27396 30598
rect 27344 30534 27396 30540
rect 27356 29646 27384 30534
rect 27448 29782 27476 31418
rect 27528 31272 27580 31278
rect 27528 31214 27580 31220
rect 27436 29776 27488 29782
rect 27436 29718 27488 29724
rect 27344 29640 27396 29646
rect 27344 29582 27396 29588
rect 27172 28966 27292 28994
rect 26988 28490 27108 28506
rect 26988 28484 27120 28490
rect 26988 28478 27068 28484
rect 27068 28426 27120 28432
rect 27172 27452 27200 28966
rect 27540 28694 27568 31214
rect 27632 29850 27660 32302
rect 27620 29844 27672 29850
rect 27620 29786 27672 29792
rect 27528 28688 27580 28694
rect 27528 28630 27580 28636
rect 27252 28552 27304 28558
rect 27252 28494 27304 28500
rect 27436 28552 27488 28558
rect 27436 28494 27488 28500
rect 27264 28218 27292 28494
rect 27252 28212 27304 28218
rect 27252 28154 27304 28160
rect 27344 28212 27396 28218
rect 27344 28154 27396 28160
rect 27356 27577 27384 28154
rect 27448 27674 27476 28494
rect 27528 28484 27580 28490
rect 27528 28426 27580 28432
rect 27540 28082 27568 28426
rect 27724 28098 27752 38383
rect 27804 38208 27856 38214
rect 27804 38150 27856 38156
rect 27816 36582 27844 38150
rect 28172 36712 28224 36718
rect 28170 36680 28172 36689
rect 28224 36680 28226 36689
rect 28170 36615 28226 36624
rect 27804 36576 27856 36582
rect 27804 36518 27856 36524
rect 27896 36304 27948 36310
rect 27896 36246 27948 36252
rect 27804 36168 27856 36174
rect 27908 36145 27936 36246
rect 27804 36110 27856 36116
rect 27894 36136 27950 36145
rect 27816 35086 27844 36110
rect 27894 36071 27950 36080
rect 27896 36032 27948 36038
rect 27896 35974 27948 35980
rect 27908 35698 27936 35974
rect 27896 35692 27948 35698
rect 27896 35634 27948 35640
rect 27804 35080 27856 35086
rect 27804 35022 27856 35028
rect 27908 34610 27936 35634
rect 27988 35488 28040 35494
rect 27988 35430 28040 35436
rect 28000 35086 28028 35430
rect 27988 35080 28040 35086
rect 27988 35022 28040 35028
rect 28172 35080 28224 35086
rect 28172 35022 28224 35028
rect 28184 34678 28212 35022
rect 28172 34672 28224 34678
rect 28172 34614 28224 34620
rect 27896 34604 27948 34610
rect 27896 34546 27948 34552
rect 28276 34524 28304 38519
rect 28460 37126 28488 38830
rect 28630 38584 28686 38593
rect 28630 38519 28686 38528
rect 28538 38448 28594 38457
rect 28644 38418 28672 38519
rect 28538 38383 28594 38392
rect 28632 38412 28684 38418
rect 28552 37806 28580 38383
rect 28632 38354 28684 38360
rect 28816 38344 28868 38350
rect 28920 38332 28948 39238
rect 29012 38418 29040 41200
rect 30380 40860 30432 40866
rect 30380 40802 30432 40808
rect 29920 40520 29972 40526
rect 29920 40462 29972 40468
rect 29644 40044 29696 40050
rect 29644 39986 29696 39992
rect 29110 39740 29418 39760
rect 29110 39738 29116 39740
rect 29172 39738 29196 39740
rect 29252 39738 29276 39740
rect 29332 39738 29356 39740
rect 29412 39738 29418 39740
rect 29172 39686 29174 39738
rect 29354 39686 29356 39738
rect 29110 39684 29116 39686
rect 29172 39684 29196 39686
rect 29252 39684 29276 39686
rect 29332 39684 29356 39686
rect 29412 39684 29418 39686
rect 29110 39664 29418 39684
rect 29460 39364 29512 39370
rect 29460 39306 29512 39312
rect 29110 38652 29418 38672
rect 29110 38650 29116 38652
rect 29172 38650 29196 38652
rect 29252 38650 29276 38652
rect 29332 38650 29356 38652
rect 29412 38650 29418 38652
rect 29172 38598 29174 38650
rect 29354 38598 29356 38650
rect 29110 38596 29116 38598
rect 29172 38596 29196 38598
rect 29252 38596 29276 38598
rect 29332 38596 29356 38598
rect 29412 38596 29418 38598
rect 29110 38576 29418 38596
rect 29000 38412 29052 38418
rect 29000 38354 29052 38360
rect 28868 38304 28948 38332
rect 28816 38286 28868 38292
rect 28920 37874 28948 38304
rect 28908 37868 28960 37874
rect 28908 37810 28960 37816
rect 28540 37800 28592 37806
rect 28540 37742 28592 37748
rect 28920 37262 28948 37810
rect 29110 37564 29418 37584
rect 29110 37562 29116 37564
rect 29172 37562 29196 37564
rect 29252 37562 29276 37564
rect 29332 37562 29356 37564
rect 29412 37562 29418 37564
rect 29172 37510 29174 37562
rect 29354 37510 29356 37562
rect 29110 37508 29116 37510
rect 29172 37508 29196 37510
rect 29252 37508 29276 37510
rect 29332 37508 29356 37510
rect 29412 37508 29418 37510
rect 29110 37488 29418 37508
rect 28908 37256 28960 37262
rect 28908 37198 28960 37204
rect 28448 37120 28500 37126
rect 28448 37062 28500 37068
rect 28724 37120 28776 37126
rect 28724 37062 28776 37068
rect 28356 36576 28408 36582
rect 28356 36518 28408 36524
rect 28368 36378 28396 36518
rect 28460 36378 28488 37062
rect 28356 36372 28408 36378
rect 28356 36314 28408 36320
rect 28448 36372 28500 36378
rect 28448 36314 28500 36320
rect 28368 36038 28396 36314
rect 28460 36242 28488 36314
rect 28448 36236 28500 36242
rect 28448 36178 28500 36184
rect 28540 36100 28592 36106
rect 28540 36042 28592 36048
rect 28356 36032 28408 36038
rect 28356 35974 28408 35980
rect 28552 35698 28580 36042
rect 28540 35692 28592 35698
rect 28540 35634 28592 35640
rect 28356 35012 28408 35018
rect 28356 34954 28408 34960
rect 28632 35012 28684 35018
rect 28632 34954 28684 34960
rect 28184 34496 28304 34524
rect 27804 33856 27856 33862
rect 27804 33798 27856 33804
rect 27816 33658 27844 33798
rect 27804 33652 27856 33658
rect 27804 33594 27856 33600
rect 27802 33552 27858 33561
rect 27802 33487 27858 33496
rect 27816 33046 27844 33487
rect 27988 33448 28040 33454
rect 27988 33390 28040 33396
rect 27804 33040 27856 33046
rect 27804 32982 27856 32988
rect 27816 32774 27844 32982
rect 28000 32842 28028 33390
rect 28080 32904 28132 32910
rect 28080 32846 28132 32852
rect 27988 32836 28040 32842
rect 27988 32778 28040 32784
rect 27804 32768 27856 32774
rect 27804 32710 27856 32716
rect 27894 32736 27950 32745
rect 27894 32671 27950 32680
rect 27908 32434 27936 32671
rect 27896 32428 27948 32434
rect 27896 32370 27948 32376
rect 27804 32360 27856 32366
rect 27804 32302 27856 32308
rect 27816 32008 27844 32302
rect 27988 32292 28040 32298
rect 27988 32234 28040 32240
rect 27816 31980 27936 32008
rect 27908 31890 27936 31980
rect 27804 31884 27856 31890
rect 27804 31826 27856 31832
rect 27896 31884 27948 31890
rect 27896 31826 27948 31832
rect 27816 30666 27844 31826
rect 27896 31748 27948 31754
rect 27896 31690 27948 31696
rect 27908 30938 27936 31690
rect 28000 31482 28028 32234
rect 28092 32201 28120 32846
rect 28078 32192 28134 32201
rect 28078 32127 28134 32136
rect 28080 31816 28132 31822
rect 28078 31784 28080 31793
rect 28132 31784 28134 31793
rect 28078 31719 28134 31728
rect 28080 31680 28132 31686
rect 28080 31622 28132 31628
rect 27988 31476 28040 31482
rect 27988 31418 28040 31424
rect 27988 31272 28040 31278
rect 27988 31214 28040 31220
rect 28000 31113 28028 31214
rect 27986 31104 28042 31113
rect 27986 31039 28042 31048
rect 27896 30932 27948 30938
rect 27896 30874 27948 30880
rect 27804 30660 27856 30666
rect 27804 30602 27856 30608
rect 27896 30660 27948 30666
rect 27896 30602 27948 30608
rect 27908 30122 27936 30602
rect 27988 30592 28040 30598
rect 27988 30534 28040 30540
rect 27896 30116 27948 30122
rect 27896 30058 27948 30064
rect 27802 30016 27858 30025
rect 27802 29951 27858 29960
rect 27816 29510 27844 29951
rect 27896 29844 27948 29850
rect 27896 29786 27948 29792
rect 27804 29504 27856 29510
rect 27804 29446 27856 29452
rect 27908 29322 27936 29786
rect 27528 28076 27580 28082
rect 27528 28018 27580 28024
rect 27632 28070 27752 28098
rect 27816 29294 27936 29322
rect 27526 27976 27582 27985
rect 27526 27911 27582 27920
rect 27436 27668 27488 27674
rect 27436 27610 27488 27616
rect 27342 27568 27398 27577
rect 27342 27503 27398 27512
rect 27252 27464 27304 27470
rect 26974 27432 27030 27441
rect 27172 27424 27252 27452
rect 27252 27406 27304 27412
rect 27436 27464 27488 27470
rect 27540 27452 27568 27911
rect 27488 27424 27568 27452
rect 27436 27406 27488 27412
rect 26974 27367 26976 27376
rect 27028 27367 27030 27376
rect 26976 27338 27028 27344
rect 26712 26846 26832 26874
rect 26608 25424 26660 25430
rect 26608 25366 26660 25372
rect 26424 24948 26476 24954
rect 26424 24890 26476 24896
rect 25780 24812 25832 24818
rect 25780 24754 25832 24760
rect 25688 23792 25740 23798
rect 25688 23734 25740 23740
rect 25228 23724 25280 23730
rect 25228 23666 25280 23672
rect 25240 23361 25268 23666
rect 25504 23656 25556 23662
rect 25504 23598 25556 23604
rect 25688 23656 25740 23662
rect 25792 23644 25820 24754
rect 25964 24744 26016 24750
rect 25964 24686 26016 24692
rect 25872 24132 25924 24138
rect 25872 24074 25924 24080
rect 25740 23616 25820 23644
rect 25688 23598 25740 23604
rect 25226 23352 25282 23361
rect 25516 23322 25544 23598
rect 25226 23287 25282 23296
rect 25504 23316 25556 23322
rect 25504 23258 25556 23264
rect 25136 23180 25188 23186
rect 25136 23122 25188 23128
rect 25412 23180 25464 23186
rect 25412 23122 25464 23128
rect 24952 23112 25004 23118
rect 24952 23054 25004 23060
rect 24860 22772 24912 22778
rect 24860 22714 24912 22720
rect 24766 21856 24822 21865
rect 24766 21791 24822 21800
rect 24768 21684 24820 21690
rect 24768 21626 24820 21632
rect 24676 21072 24728 21078
rect 24582 21040 24638 21049
rect 24676 21014 24728 21020
rect 24582 20975 24638 20984
rect 24584 20800 24636 20806
rect 24584 20742 24636 20748
rect 24492 20528 24544 20534
rect 24492 20470 24544 20476
rect 24492 20256 24544 20262
rect 24492 20198 24544 20204
rect 24504 19922 24532 20198
rect 24492 19916 24544 19922
rect 24492 19858 24544 19864
rect 24400 19304 24452 19310
rect 24400 19246 24452 19252
rect 24308 18828 24360 18834
rect 24308 18770 24360 18776
rect 24216 18760 24268 18766
rect 24216 18702 24268 18708
rect 24492 17808 24544 17814
rect 24492 17750 24544 17756
rect 24504 17134 24532 17750
rect 24596 17542 24624 20742
rect 24688 18290 24716 21014
rect 24780 21010 24808 21626
rect 24872 21146 24900 22714
rect 24964 22409 24992 23054
rect 25044 22636 25096 22642
rect 25044 22578 25096 22584
rect 24950 22400 25006 22409
rect 24950 22335 25006 22344
rect 24952 22092 25004 22098
rect 24952 22034 25004 22040
rect 24860 21140 24912 21146
rect 24860 21082 24912 21088
rect 24768 21004 24820 21010
rect 24768 20946 24820 20952
rect 24860 20936 24912 20942
rect 24766 20904 24822 20913
rect 24822 20884 24860 20890
rect 24822 20878 24912 20884
rect 24822 20862 24900 20878
rect 24766 20839 24822 20848
rect 24780 19922 24808 20839
rect 24964 20788 24992 22034
rect 25056 21962 25084 22578
rect 25148 22001 25176 23122
rect 25228 22704 25280 22710
rect 25228 22646 25280 22652
rect 25134 21992 25190 22001
rect 25044 21956 25096 21962
rect 25134 21927 25190 21936
rect 25044 21898 25096 21904
rect 25056 21400 25084 21898
rect 25136 21412 25188 21418
rect 25056 21372 25136 21400
rect 25136 21354 25188 21360
rect 25044 20936 25096 20942
rect 25044 20878 25096 20884
rect 24872 20760 24992 20788
rect 24768 19916 24820 19922
rect 24768 19858 24820 19864
rect 24768 18828 24820 18834
rect 24768 18770 24820 18776
rect 24676 18284 24728 18290
rect 24676 18226 24728 18232
rect 24780 17746 24808 18770
rect 24872 18358 24900 20760
rect 24952 20460 25004 20466
rect 24952 20402 25004 20408
rect 24964 19378 24992 20402
rect 24952 19372 25004 19378
rect 24952 19314 25004 19320
rect 24964 18970 24992 19314
rect 24952 18964 25004 18970
rect 24952 18906 25004 18912
rect 25056 18766 25084 20878
rect 25148 19310 25176 21354
rect 25240 19854 25268 22646
rect 25424 22137 25452 23122
rect 25596 23112 25648 23118
rect 25596 23054 25648 23060
rect 25608 22710 25636 23054
rect 25596 22704 25648 22710
rect 25502 22672 25558 22681
rect 25596 22646 25648 22652
rect 25502 22607 25504 22616
rect 25556 22607 25558 22616
rect 25504 22578 25556 22584
rect 25410 22128 25466 22137
rect 25410 22063 25466 22072
rect 25596 22092 25648 22098
rect 25596 22034 25648 22040
rect 25320 22024 25372 22030
rect 25504 22024 25556 22030
rect 25320 21966 25372 21972
rect 25410 21992 25466 22001
rect 25332 21486 25360 21966
rect 25608 22001 25636 22034
rect 25504 21966 25556 21972
rect 25594 21992 25650 22001
rect 25410 21927 25466 21936
rect 25320 21480 25372 21486
rect 25320 21422 25372 21428
rect 25318 21176 25374 21185
rect 25318 21111 25374 21120
rect 25228 19848 25280 19854
rect 25228 19790 25280 19796
rect 25228 19712 25280 19718
rect 25228 19654 25280 19660
rect 25136 19304 25188 19310
rect 25136 19246 25188 19252
rect 25136 19168 25188 19174
rect 25136 19110 25188 19116
rect 25148 18902 25176 19110
rect 25136 18896 25188 18902
rect 25136 18838 25188 18844
rect 25044 18760 25096 18766
rect 25044 18702 25096 18708
rect 24952 18624 25004 18630
rect 24952 18566 25004 18572
rect 24860 18352 24912 18358
rect 24860 18294 24912 18300
rect 24860 18148 24912 18154
rect 24860 18090 24912 18096
rect 24768 17740 24820 17746
rect 24768 17682 24820 17688
rect 24584 17536 24636 17542
rect 24584 17478 24636 17484
rect 24872 17184 24900 18090
rect 24964 17678 24992 18566
rect 25056 18290 25084 18702
rect 25044 18284 25096 18290
rect 25044 18226 25096 18232
rect 25136 18284 25188 18290
rect 25136 18226 25188 18232
rect 24952 17672 25004 17678
rect 24952 17614 25004 17620
rect 25044 17604 25096 17610
rect 25044 17546 25096 17552
rect 25056 17338 25084 17546
rect 25044 17332 25096 17338
rect 25044 17274 25096 17280
rect 24952 17196 25004 17202
rect 24872 17156 24952 17184
rect 24952 17138 25004 17144
rect 24492 17128 24544 17134
rect 24492 17070 24544 17076
rect 25148 17066 25176 18226
rect 25240 17678 25268 19654
rect 25228 17672 25280 17678
rect 25228 17614 25280 17620
rect 25332 17338 25360 21111
rect 25424 21078 25452 21927
rect 25412 21072 25464 21078
rect 25412 21014 25464 21020
rect 25424 20788 25452 21014
rect 25516 20942 25544 21966
rect 25594 21927 25650 21936
rect 25700 21434 25728 23598
rect 25780 23520 25832 23526
rect 25780 23462 25832 23468
rect 25792 21593 25820 23462
rect 25884 22710 25912 24074
rect 25976 24070 26004 24686
rect 26712 24614 26740 26846
rect 26792 26784 26844 26790
rect 26792 26726 26844 26732
rect 26700 24608 26752 24614
rect 26700 24550 26752 24556
rect 26056 24200 26108 24206
rect 26056 24142 26108 24148
rect 26148 24200 26200 24206
rect 26148 24142 26200 24148
rect 25964 24064 26016 24070
rect 25964 24006 26016 24012
rect 26068 23118 26096 24142
rect 26056 23112 26108 23118
rect 26056 23054 26108 23060
rect 25872 22704 25924 22710
rect 25872 22646 25924 22652
rect 25884 22166 25912 22646
rect 25964 22636 26016 22642
rect 25964 22578 26016 22584
rect 25976 22409 26004 22578
rect 25962 22400 26018 22409
rect 25962 22335 26018 22344
rect 25872 22160 25924 22166
rect 25872 22102 25924 22108
rect 25778 21584 25834 21593
rect 25778 21519 25780 21528
rect 25832 21519 25834 21528
rect 25780 21490 25832 21496
rect 25976 21486 26004 22335
rect 26068 22030 26096 23054
rect 26160 22574 26188 24142
rect 26804 23769 26832 26726
rect 26988 25294 27016 27338
rect 27264 27033 27292 27406
rect 27250 27024 27306 27033
rect 27068 26988 27120 26994
rect 27250 26959 27306 26968
rect 27068 26930 27120 26936
rect 27080 26042 27108 26930
rect 27068 26036 27120 26042
rect 27068 25978 27120 25984
rect 26976 25288 27028 25294
rect 26976 25230 27028 25236
rect 27068 24812 27120 24818
rect 27068 24754 27120 24760
rect 26884 24064 26936 24070
rect 26884 24006 26936 24012
rect 26790 23760 26846 23769
rect 26790 23695 26846 23704
rect 26332 23520 26384 23526
rect 26332 23462 26384 23468
rect 26344 23118 26372 23462
rect 26332 23112 26384 23118
rect 26332 23054 26384 23060
rect 26148 22568 26200 22574
rect 26148 22510 26200 22516
rect 26240 22568 26292 22574
rect 26240 22510 26292 22516
rect 26056 22024 26108 22030
rect 26056 21966 26108 21972
rect 25964 21480 26016 21486
rect 25700 21406 25820 21434
rect 25964 21422 26016 21428
rect 25688 21344 25740 21350
rect 25688 21286 25740 21292
rect 25504 20936 25556 20942
rect 25504 20878 25556 20884
rect 25700 20874 25728 21286
rect 25688 20868 25740 20874
rect 25688 20810 25740 20816
rect 25424 20760 25636 20788
rect 25412 19304 25464 19310
rect 25412 19246 25464 19252
rect 25424 17610 25452 19246
rect 25504 18692 25556 18698
rect 25504 18634 25556 18640
rect 25516 17882 25544 18634
rect 25608 18426 25636 20760
rect 25686 20768 25742 20777
rect 25686 20703 25742 20712
rect 25596 18420 25648 18426
rect 25596 18362 25648 18368
rect 25504 17876 25556 17882
rect 25504 17818 25556 17824
rect 25412 17604 25464 17610
rect 25412 17546 25464 17552
rect 25320 17332 25372 17338
rect 25320 17274 25372 17280
rect 25410 17232 25466 17241
rect 25700 17202 25728 20703
rect 25792 20466 25820 21406
rect 26160 21146 26188 22510
rect 26252 21729 26280 22510
rect 26332 22432 26384 22438
rect 26332 22374 26384 22380
rect 26344 22030 26372 22374
rect 26332 22024 26384 22030
rect 26332 21966 26384 21972
rect 26238 21720 26294 21729
rect 26238 21655 26294 21664
rect 26332 21344 26384 21350
rect 26332 21286 26384 21292
rect 26148 21140 26200 21146
rect 26148 21082 26200 21088
rect 25962 20496 26018 20505
rect 25780 20460 25832 20466
rect 26344 20466 26372 21286
rect 26700 21140 26752 21146
rect 26700 21082 26752 21088
rect 26712 20466 26740 21082
rect 26896 20806 26924 24006
rect 27080 22273 27108 24754
rect 27160 24608 27212 24614
rect 27160 24550 27212 24556
rect 27172 24070 27200 24550
rect 27160 24064 27212 24070
rect 27160 24006 27212 24012
rect 27264 22681 27292 26959
rect 27448 26246 27476 27406
rect 27436 26240 27488 26246
rect 27436 26182 27488 26188
rect 27344 25900 27396 25906
rect 27344 25842 27396 25848
rect 27356 25498 27384 25842
rect 27344 25492 27396 25498
rect 27344 25434 27396 25440
rect 27528 23724 27580 23730
rect 27528 23666 27580 23672
rect 27540 23322 27568 23666
rect 27528 23316 27580 23322
rect 27528 23258 27580 23264
rect 27528 22976 27580 22982
rect 27528 22918 27580 22924
rect 27250 22672 27306 22681
rect 27250 22607 27306 22616
rect 27252 22568 27304 22574
rect 27344 22568 27396 22574
rect 27252 22510 27304 22516
rect 27342 22536 27344 22545
rect 27396 22536 27398 22545
rect 27066 22264 27122 22273
rect 26988 22222 27066 22250
rect 26884 20800 26936 20806
rect 26988 20777 27016 22222
rect 27066 22199 27122 22208
rect 27264 22166 27292 22510
rect 27342 22471 27398 22480
rect 27252 22160 27304 22166
rect 27252 22102 27304 22108
rect 27066 21992 27122 22001
rect 27066 21927 27122 21936
rect 27160 21956 27212 21962
rect 27080 21418 27108 21927
rect 27160 21898 27212 21904
rect 27172 21622 27200 21898
rect 27252 21888 27304 21894
rect 27252 21830 27304 21836
rect 27264 21690 27292 21830
rect 27252 21684 27304 21690
rect 27252 21626 27304 21632
rect 27160 21616 27212 21622
rect 27160 21558 27212 21564
rect 27068 21412 27120 21418
rect 27068 21354 27120 21360
rect 27264 20942 27292 21626
rect 27356 21554 27384 22471
rect 27344 21548 27396 21554
rect 27344 21490 27396 21496
rect 27540 21486 27568 22918
rect 27528 21480 27580 21486
rect 27528 21422 27580 21428
rect 27540 20942 27568 21422
rect 27252 20936 27304 20942
rect 27252 20878 27304 20884
rect 27528 20936 27580 20942
rect 27528 20878 27580 20884
rect 26884 20742 26936 20748
rect 26974 20768 27030 20777
rect 26974 20703 27030 20712
rect 26988 20618 27016 20703
rect 26896 20590 27016 20618
rect 25962 20431 25964 20440
rect 25780 20402 25832 20408
rect 26016 20431 26018 20440
rect 26148 20460 26200 20466
rect 25964 20402 26016 20408
rect 26148 20402 26200 20408
rect 26332 20460 26384 20466
rect 26332 20402 26384 20408
rect 26700 20460 26752 20466
rect 26700 20402 26752 20408
rect 26160 19990 26188 20402
rect 26240 20324 26292 20330
rect 26240 20266 26292 20272
rect 26252 20058 26280 20266
rect 26240 20052 26292 20058
rect 26240 19994 26292 20000
rect 26148 19984 26200 19990
rect 26148 19926 26200 19932
rect 26344 19854 26372 20402
rect 26516 20392 26568 20398
rect 26516 20334 26568 20340
rect 26332 19848 26384 19854
rect 26332 19790 26384 19796
rect 26528 19718 26556 20334
rect 26516 19712 26568 19718
rect 26422 19680 26478 19689
rect 26516 19654 26568 19660
rect 26422 19615 26478 19624
rect 26436 19174 26464 19615
rect 26424 19168 26476 19174
rect 26424 19110 26476 19116
rect 25872 18964 25924 18970
rect 25872 18906 25924 18912
rect 25780 18420 25832 18426
rect 25780 18362 25832 18368
rect 25792 17678 25820 18362
rect 25884 17882 25912 18906
rect 26436 18426 26464 19110
rect 26528 18630 26556 19654
rect 26516 18624 26568 18630
rect 26516 18566 26568 18572
rect 26424 18420 26476 18426
rect 26424 18362 26476 18368
rect 26896 17882 26924 20590
rect 27160 20460 27212 20466
rect 27344 20460 27396 20466
rect 27160 20402 27212 20408
rect 27264 20420 27344 20448
rect 27172 19854 27200 20402
rect 27160 19848 27212 19854
rect 27160 19790 27212 19796
rect 26976 19780 27028 19786
rect 26976 19722 27028 19728
rect 26988 19446 27016 19722
rect 27264 19514 27292 20420
rect 27344 20402 27396 20408
rect 27528 19848 27580 19854
rect 27528 19790 27580 19796
rect 27252 19508 27304 19514
rect 27252 19450 27304 19456
rect 26976 19440 27028 19446
rect 26976 19382 27028 19388
rect 27252 19372 27304 19378
rect 27252 19314 27304 19320
rect 27068 19168 27120 19174
rect 27068 19110 27120 19116
rect 27080 18358 27108 19110
rect 27068 18352 27120 18358
rect 27068 18294 27120 18300
rect 27264 17882 27292 19314
rect 27540 19310 27568 19790
rect 27528 19304 27580 19310
rect 27528 19246 27580 19252
rect 27540 18426 27568 19246
rect 27528 18420 27580 18426
rect 27528 18362 27580 18368
rect 25872 17876 25924 17882
rect 25872 17818 25924 17824
rect 26884 17876 26936 17882
rect 26884 17818 26936 17824
rect 27252 17876 27304 17882
rect 27252 17818 27304 17824
rect 27540 17678 27568 18362
rect 25780 17672 25832 17678
rect 25780 17614 25832 17620
rect 27528 17672 27580 17678
rect 27528 17614 27580 17620
rect 25964 17536 26016 17542
rect 25964 17478 26016 17484
rect 25976 17270 26004 17478
rect 25964 17264 26016 17270
rect 25964 17206 26016 17212
rect 25410 17167 25412 17176
rect 25464 17167 25466 17176
rect 25688 17196 25740 17202
rect 25412 17138 25464 17144
rect 25688 17138 25740 17144
rect 25136 17060 25188 17066
rect 25136 17002 25188 17008
rect 24032 5840 24084 5846
rect 24032 5782 24084 5788
rect 23478 5468 23786 5488
rect 23478 5466 23484 5468
rect 23540 5466 23564 5468
rect 23620 5466 23644 5468
rect 23700 5466 23724 5468
rect 23780 5466 23786 5468
rect 23540 5414 23542 5466
rect 23722 5414 23724 5466
rect 23478 5412 23484 5414
rect 23540 5412 23564 5414
rect 23620 5412 23644 5414
rect 23700 5412 23724 5414
rect 23780 5412 23786 5414
rect 23478 5392 23786 5412
rect 27632 5234 27660 28070
rect 27712 28008 27764 28014
rect 27816 27985 27844 29294
rect 28000 28558 28028 30534
rect 28092 28762 28120 31622
rect 28080 28756 28132 28762
rect 28080 28698 28132 28704
rect 27988 28552 28040 28558
rect 27908 28512 27988 28540
rect 27712 27950 27764 27956
rect 27802 27976 27858 27985
rect 27724 26790 27752 27950
rect 27908 27946 27936 28512
rect 27988 28494 28040 28500
rect 27988 28416 28040 28422
rect 27988 28358 28040 28364
rect 27802 27911 27858 27920
rect 27896 27940 27948 27946
rect 27896 27882 27948 27888
rect 27804 27872 27856 27878
rect 27804 27814 27856 27820
rect 27712 26784 27764 26790
rect 27712 26726 27764 26732
rect 27724 26382 27752 26726
rect 27712 26376 27764 26382
rect 27712 26318 27764 26324
rect 27712 26240 27764 26246
rect 27712 26182 27764 26188
rect 27724 24886 27752 26182
rect 27712 24880 27764 24886
rect 27712 24822 27764 24828
rect 27724 24313 27752 24822
rect 27816 24682 27844 27814
rect 27908 27130 27936 27882
rect 27896 27124 27948 27130
rect 27896 27066 27948 27072
rect 27908 25838 27936 27066
rect 27896 25832 27948 25838
rect 27896 25774 27948 25780
rect 28000 25498 28028 28358
rect 28080 28144 28132 28150
rect 28080 28086 28132 28092
rect 27988 25492 28040 25498
rect 27988 25434 28040 25440
rect 28092 25265 28120 28086
rect 28184 27606 28212 34496
rect 28368 34456 28396 34954
rect 28540 34944 28592 34950
rect 28540 34886 28592 34892
rect 28276 34428 28396 34456
rect 28276 32314 28304 34428
rect 28552 34406 28580 34886
rect 28540 34400 28592 34406
rect 28540 34342 28592 34348
rect 28552 33998 28580 34342
rect 28644 34202 28672 34954
rect 28632 34196 28684 34202
rect 28632 34138 28684 34144
rect 28540 33992 28592 33998
rect 28540 33934 28592 33940
rect 28448 33924 28500 33930
rect 28448 33866 28500 33872
rect 28460 33590 28488 33866
rect 28448 33584 28500 33590
rect 28448 33526 28500 33532
rect 28736 33504 28764 37062
rect 28920 36786 28948 37198
rect 28908 36780 28960 36786
rect 28908 36722 28960 36728
rect 29110 36476 29418 36496
rect 29110 36474 29116 36476
rect 29172 36474 29196 36476
rect 29252 36474 29276 36476
rect 29332 36474 29356 36476
rect 29412 36474 29418 36476
rect 29172 36422 29174 36474
rect 29354 36422 29356 36474
rect 29110 36420 29116 36422
rect 29172 36420 29196 36422
rect 29252 36420 29276 36422
rect 29332 36420 29356 36422
rect 29412 36420 29418 36422
rect 29110 36400 29418 36420
rect 29000 36236 29052 36242
rect 29000 36178 29052 36184
rect 29012 35834 29040 36178
rect 29000 35828 29052 35834
rect 29000 35770 29052 35776
rect 29184 35760 29236 35766
rect 28920 35708 29184 35714
rect 29472 35737 29500 39306
rect 29552 38344 29604 38350
rect 29552 38286 29604 38292
rect 29564 37777 29592 38286
rect 29550 37768 29606 37777
rect 29550 37703 29606 37712
rect 29656 36378 29684 39986
rect 29828 39024 29880 39030
rect 29828 38966 29880 38972
rect 29736 37800 29788 37806
rect 29736 37742 29788 37748
rect 29748 37369 29776 37742
rect 29734 37360 29790 37369
rect 29734 37295 29790 37304
rect 29736 36644 29788 36650
rect 29736 36586 29788 36592
rect 29644 36372 29696 36378
rect 29644 36314 29696 36320
rect 29644 36168 29696 36174
rect 29644 36110 29696 36116
rect 29552 36032 29604 36038
rect 29552 35974 29604 35980
rect 28920 35702 29236 35708
rect 29458 35728 29514 35737
rect 28920 35686 29224 35702
rect 28920 35465 28948 35686
rect 29458 35663 29514 35672
rect 29460 35488 29512 35494
rect 28906 35456 28962 35465
rect 29460 35430 29512 35436
rect 28906 35391 28962 35400
rect 29110 35388 29418 35408
rect 29110 35386 29116 35388
rect 29172 35386 29196 35388
rect 29252 35386 29276 35388
rect 29332 35386 29356 35388
rect 29412 35386 29418 35388
rect 29172 35334 29174 35386
rect 29354 35334 29356 35386
rect 29110 35332 29116 35334
rect 29172 35332 29196 35334
rect 29252 35332 29276 35334
rect 29332 35332 29356 35334
rect 29412 35332 29418 35334
rect 29110 35312 29418 35332
rect 29368 35148 29420 35154
rect 29368 35090 29420 35096
rect 29380 34785 29408 35090
rect 29366 34776 29422 34785
rect 29366 34711 29422 34720
rect 29472 34678 29500 35430
rect 29368 34672 29420 34678
rect 29368 34614 29420 34620
rect 29460 34672 29512 34678
rect 29460 34614 29512 34620
rect 28816 34604 28868 34610
rect 28816 34546 28868 34552
rect 28908 34604 28960 34610
rect 28908 34546 28960 34552
rect 28828 33658 28856 34546
rect 28816 33652 28868 33658
rect 28816 33594 28868 33600
rect 28644 33476 28764 33504
rect 28356 33448 28408 33454
rect 28356 33390 28408 33396
rect 28368 33318 28396 33390
rect 28356 33312 28408 33318
rect 28356 33254 28408 33260
rect 28368 32910 28396 33254
rect 28644 33153 28672 33476
rect 28722 33280 28778 33289
rect 28722 33215 28778 33224
rect 28630 33144 28686 33153
rect 28630 33079 28686 33088
rect 28644 32960 28672 33079
rect 28736 33046 28764 33215
rect 28724 33040 28776 33046
rect 28724 32982 28776 32988
rect 28552 32932 28672 32960
rect 28356 32904 28408 32910
rect 28408 32864 28488 32892
rect 28356 32846 28408 32852
rect 28356 32768 28408 32774
rect 28356 32710 28408 32716
rect 28368 32434 28396 32710
rect 28460 32434 28488 32864
rect 28356 32428 28408 32434
rect 28356 32370 28408 32376
rect 28448 32428 28500 32434
rect 28448 32370 28500 32376
rect 28276 32286 28396 32314
rect 28264 31476 28316 31482
rect 28264 31418 28316 31424
rect 28276 30938 28304 31418
rect 28264 30932 28316 30938
rect 28264 30874 28316 30880
rect 28368 30569 28396 32286
rect 28552 31482 28580 32932
rect 28828 32858 28856 33594
rect 28920 33522 28948 34546
rect 29000 34468 29052 34474
rect 29000 34410 29052 34416
rect 28908 33516 28960 33522
rect 28908 33458 28960 33464
rect 29012 33454 29040 34410
rect 29380 34388 29408 34614
rect 29380 34360 29500 34388
rect 29110 34300 29418 34320
rect 29110 34298 29116 34300
rect 29172 34298 29196 34300
rect 29252 34298 29276 34300
rect 29332 34298 29356 34300
rect 29412 34298 29418 34300
rect 29172 34246 29174 34298
rect 29354 34246 29356 34298
rect 29110 34244 29116 34246
rect 29172 34244 29196 34246
rect 29252 34244 29276 34246
rect 29332 34244 29356 34246
rect 29412 34244 29418 34246
rect 29110 34224 29418 34244
rect 29274 34096 29330 34105
rect 29274 34031 29330 34040
rect 29288 33454 29316 34031
rect 29368 33584 29420 33590
rect 29472 33561 29500 34360
rect 29368 33526 29420 33532
rect 29458 33552 29514 33561
rect 29000 33448 29052 33454
rect 29000 33390 29052 33396
rect 29276 33448 29328 33454
rect 29276 33390 29328 33396
rect 29012 32978 29040 33390
rect 29380 33368 29408 33526
rect 29458 33487 29460 33496
rect 29512 33487 29514 33496
rect 29460 33458 29512 33464
rect 29460 33380 29512 33386
rect 29380 33340 29460 33368
rect 29460 33322 29512 33328
rect 29110 33212 29418 33232
rect 29110 33210 29116 33212
rect 29172 33210 29196 33212
rect 29252 33210 29276 33212
rect 29332 33210 29356 33212
rect 29412 33210 29418 33212
rect 29172 33158 29174 33210
rect 29354 33158 29356 33210
rect 29110 33156 29116 33158
rect 29172 33156 29196 33158
rect 29252 33156 29276 33158
rect 29332 33156 29356 33158
rect 29412 33156 29418 33158
rect 29110 33136 29418 33156
rect 29092 33040 29144 33046
rect 29276 33040 29328 33046
rect 29144 33000 29276 33028
rect 29092 32982 29144 32988
rect 29276 32982 29328 32988
rect 29000 32972 29052 32978
rect 29000 32914 29052 32920
rect 28828 32830 28994 32858
rect 28816 32768 28868 32774
rect 28736 32728 28816 32756
rect 28632 32292 28684 32298
rect 28632 32234 28684 32240
rect 28644 31958 28672 32234
rect 28632 31952 28684 31958
rect 28632 31894 28684 31900
rect 28736 31822 28764 32728
rect 28816 32710 28868 32716
rect 28966 32484 28994 32830
rect 29472 32774 29500 33322
rect 29564 33046 29592 35974
rect 29656 35222 29684 36110
rect 29644 35216 29696 35222
rect 29644 35158 29696 35164
rect 29656 35086 29684 35158
rect 29644 35080 29696 35086
rect 29644 35022 29696 35028
rect 29656 33998 29684 35022
rect 29644 33992 29696 33998
rect 29644 33934 29696 33940
rect 29644 33856 29696 33862
rect 29644 33798 29696 33804
rect 29552 33040 29604 33046
rect 29552 32982 29604 32988
rect 29552 32904 29604 32910
rect 29552 32846 29604 32852
rect 29460 32768 29512 32774
rect 29460 32710 29512 32716
rect 28920 32456 28994 32484
rect 28816 32428 28868 32434
rect 28816 32370 28868 32376
rect 28828 32201 28856 32370
rect 28920 32298 28948 32456
rect 28908 32292 28960 32298
rect 28908 32234 28960 32240
rect 29000 32224 29052 32230
rect 28814 32192 28870 32201
rect 29000 32166 29052 32172
rect 28814 32127 28870 32136
rect 28724 31816 28776 31822
rect 28724 31758 28776 31764
rect 28632 31680 28684 31686
rect 28632 31622 28684 31628
rect 28540 31476 28592 31482
rect 28540 31418 28592 31424
rect 28446 31240 28502 31249
rect 28446 31175 28502 31184
rect 28354 30560 28410 30569
rect 28354 30495 28410 30504
rect 28264 30252 28316 30258
rect 28264 30194 28316 30200
rect 28276 29850 28304 30194
rect 28264 29844 28316 29850
rect 28264 29786 28316 29792
rect 28264 28620 28316 28626
rect 28264 28562 28316 28568
rect 28276 28529 28304 28562
rect 28262 28520 28318 28529
rect 28262 28455 28318 28464
rect 28264 27668 28316 27674
rect 28264 27610 28316 27616
rect 28172 27600 28224 27606
rect 28172 27542 28224 27548
rect 28276 26790 28304 27610
rect 28368 27316 28396 30495
rect 28460 30240 28488 31175
rect 28538 30832 28594 30841
rect 28538 30767 28540 30776
rect 28592 30767 28594 30776
rect 28540 30738 28592 30744
rect 28644 30716 28672 31622
rect 28736 30977 28764 31758
rect 28722 30968 28778 30977
rect 28722 30903 28778 30912
rect 28724 30728 28776 30734
rect 28644 30688 28724 30716
rect 28724 30670 28776 30676
rect 28540 30252 28592 30258
rect 28460 30212 28540 30240
rect 28540 30194 28592 30200
rect 28736 30036 28764 30670
rect 28828 30104 28856 32127
rect 29012 31822 29040 32166
rect 29110 32124 29418 32144
rect 29110 32122 29116 32124
rect 29172 32122 29196 32124
rect 29252 32122 29276 32124
rect 29332 32122 29356 32124
rect 29412 32122 29418 32124
rect 29172 32070 29174 32122
rect 29354 32070 29356 32122
rect 29110 32068 29116 32070
rect 29172 32068 29196 32070
rect 29252 32068 29276 32070
rect 29332 32068 29356 32070
rect 29412 32068 29418 32070
rect 29110 32048 29418 32068
rect 29564 32065 29592 32846
rect 29550 32056 29606 32065
rect 29550 31991 29606 32000
rect 29276 31952 29328 31958
rect 29276 31894 29328 31900
rect 29366 31920 29422 31929
rect 29000 31816 29052 31822
rect 29000 31758 29052 31764
rect 29000 31680 29052 31686
rect 28920 31640 29000 31668
rect 28920 30666 28948 31640
rect 29288 31657 29316 31894
rect 29422 31864 29500 31872
rect 29366 31855 29500 31864
rect 29380 31844 29500 31855
rect 29000 31622 29052 31628
rect 29274 31648 29330 31657
rect 29274 31583 29330 31592
rect 29000 31136 29052 31142
rect 29000 31078 29052 31084
rect 28908 30660 28960 30666
rect 28908 30602 28960 30608
rect 29012 30326 29040 31078
rect 29110 31036 29418 31056
rect 29110 31034 29116 31036
rect 29172 31034 29196 31036
rect 29252 31034 29276 31036
rect 29332 31034 29356 31036
rect 29412 31034 29418 31036
rect 29172 30982 29174 31034
rect 29354 30982 29356 31034
rect 29110 30980 29116 30982
rect 29172 30980 29196 30982
rect 29252 30980 29276 30982
rect 29332 30980 29356 30982
rect 29412 30980 29418 30982
rect 29110 30960 29418 30980
rect 29000 30320 29052 30326
rect 29000 30262 29052 30268
rect 29000 30116 29052 30122
rect 28828 30076 29000 30104
rect 28446 30016 28502 30025
rect 28736 30008 28856 30036
rect 28920 30025 28948 30076
rect 29000 30058 29052 30064
rect 28446 29951 28502 29960
rect 28460 29646 28488 29951
rect 28538 29880 28594 29889
rect 28538 29815 28594 29824
rect 28724 29844 28776 29850
rect 28448 29640 28500 29646
rect 28448 29582 28500 29588
rect 28460 29481 28488 29582
rect 28446 29472 28502 29481
rect 28446 29407 28502 29416
rect 28446 29200 28502 29209
rect 28446 29135 28502 29144
rect 28460 27441 28488 29135
rect 28446 27432 28502 27441
rect 28446 27367 28502 27376
rect 28448 27328 28500 27334
rect 28368 27296 28448 27316
rect 28500 27296 28502 27305
rect 28368 27288 28446 27296
rect 28446 27231 28502 27240
rect 28264 26784 28316 26790
rect 28264 26726 28316 26732
rect 28172 26512 28224 26518
rect 28172 26454 28224 26460
rect 28184 25770 28212 26454
rect 28356 26376 28408 26382
rect 28356 26318 28408 26324
rect 28264 26240 28316 26246
rect 28264 26182 28316 26188
rect 28172 25764 28224 25770
rect 28172 25706 28224 25712
rect 28276 25650 28304 26182
rect 28368 25838 28396 26318
rect 28552 26042 28580 29815
rect 28724 29786 28776 29792
rect 28736 29646 28764 29786
rect 28724 29640 28776 29646
rect 28644 29600 28724 29628
rect 28644 28694 28672 29600
rect 28724 29582 28776 29588
rect 28724 28960 28776 28966
rect 28828 28937 28856 30008
rect 28906 30016 28962 30025
rect 28906 29951 28962 29960
rect 29110 29948 29418 29968
rect 29110 29946 29116 29948
rect 29172 29946 29196 29948
rect 29252 29946 29276 29948
rect 29332 29946 29356 29948
rect 29412 29946 29418 29948
rect 29172 29894 29174 29946
rect 29354 29894 29356 29946
rect 29110 29892 29116 29894
rect 29172 29892 29196 29894
rect 29252 29892 29276 29894
rect 29332 29892 29356 29894
rect 29412 29892 29418 29894
rect 29110 29872 29418 29892
rect 29368 29640 29420 29646
rect 29366 29608 29368 29617
rect 29420 29608 29422 29617
rect 29276 29572 29328 29578
rect 29366 29543 29422 29552
rect 29276 29514 29328 29520
rect 29288 29345 29316 29514
rect 29368 29504 29420 29510
rect 29368 29446 29420 29452
rect 29274 29336 29330 29345
rect 29274 29271 29330 29280
rect 29380 29170 29408 29446
rect 29092 29164 29144 29170
rect 29012 29124 29092 29152
rect 28724 28902 28776 28908
rect 28814 28928 28870 28937
rect 28632 28688 28684 28694
rect 28632 28630 28684 28636
rect 28736 27470 28764 28902
rect 28814 28863 28870 28872
rect 28828 28540 28856 28863
rect 29012 28762 29040 29124
rect 29092 29106 29144 29112
rect 29368 29164 29420 29170
rect 29368 29106 29420 29112
rect 29110 28860 29418 28880
rect 29110 28858 29116 28860
rect 29172 28858 29196 28860
rect 29252 28858 29276 28860
rect 29332 28858 29356 28860
rect 29412 28858 29418 28860
rect 29172 28806 29174 28858
rect 29354 28806 29356 28858
rect 29110 28804 29116 28806
rect 29172 28804 29196 28806
rect 29252 28804 29276 28806
rect 29332 28804 29356 28806
rect 29412 28804 29418 28806
rect 29110 28784 29418 28804
rect 29000 28756 29052 28762
rect 29000 28698 29052 28704
rect 29472 28608 29500 31844
rect 29656 31482 29684 33798
rect 29748 33114 29776 36586
rect 29840 33590 29868 38966
rect 29932 37942 29960 40462
rect 30104 40452 30156 40458
rect 30104 40394 30156 40400
rect 30012 40316 30064 40322
rect 30012 40258 30064 40264
rect 29920 37936 29972 37942
rect 29920 37878 29972 37884
rect 30024 37754 30052 40258
rect 29932 37726 30052 37754
rect 29932 35698 29960 37726
rect 30012 36372 30064 36378
rect 30012 36314 30064 36320
rect 29920 35692 29972 35698
rect 29920 35634 29972 35640
rect 29918 34912 29974 34921
rect 29918 34847 29974 34856
rect 29828 33584 29880 33590
rect 29828 33526 29880 33532
rect 29840 33318 29868 33526
rect 29828 33312 29880 33318
rect 29828 33254 29880 33260
rect 29736 33108 29788 33114
rect 29736 33050 29788 33056
rect 29736 32972 29788 32978
rect 29736 32914 29788 32920
rect 29748 32881 29776 32914
rect 29840 32910 29868 33254
rect 29932 33046 29960 34847
rect 30024 33538 30052 36314
rect 30116 33998 30144 40394
rect 30288 40384 30340 40390
rect 30288 40326 30340 40332
rect 30196 39568 30248 39574
rect 30196 39510 30248 39516
rect 30208 35018 30236 39510
rect 30300 38654 30328 40326
rect 30392 39098 30420 40802
rect 31852 40588 31904 40594
rect 31852 40530 31904 40536
rect 31390 39944 31446 39953
rect 31390 39879 31446 39888
rect 30472 39500 30524 39506
rect 30472 39442 30524 39448
rect 30380 39092 30432 39098
rect 30380 39034 30432 39040
rect 30300 38626 30420 38654
rect 30288 36780 30340 36786
rect 30288 36722 30340 36728
rect 30300 36174 30328 36722
rect 30288 36168 30340 36174
rect 30288 36110 30340 36116
rect 30392 36106 30420 38626
rect 30380 36100 30432 36106
rect 30380 36042 30432 36048
rect 30196 35012 30248 35018
rect 30196 34954 30248 34960
rect 30104 33992 30156 33998
rect 30104 33934 30156 33940
rect 30024 33510 30144 33538
rect 30012 33448 30064 33454
rect 30012 33390 30064 33396
rect 29920 33040 29972 33046
rect 29920 32982 29972 32988
rect 29828 32904 29880 32910
rect 29734 32872 29790 32881
rect 29828 32846 29880 32852
rect 29918 32872 29974 32881
rect 29734 32807 29790 32816
rect 29918 32807 29974 32816
rect 29828 32768 29880 32774
rect 29828 32710 29880 32716
rect 29840 31872 29868 32710
rect 29768 31844 29868 31872
rect 29768 31804 29796 31844
rect 29748 31776 29796 31804
rect 29644 31476 29696 31482
rect 29644 31418 29696 31424
rect 29748 31362 29776 31776
rect 29828 31748 29880 31754
rect 29828 31690 29880 31696
rect 29564 31334 29776 31362
rect 29564 28937 29592 31334
rect 29736 31272 29788 31278
rect 29736 31214 29788 31220
rect 29748 30977 29776 31214
rect 29734 30968 29790 30977
rect 29734 30903 29790 30912
rect 29736 30796 29788 30802
rect 29736 30738 29788 30744
rect 29644 30660 29696 30666
rect 29644 30602 29696 30608
rect 29656 30326 29684 30602
rect 29644 30320 29696 30326
rect 29644 30262 29696 30268
rect 29644 30116 29696 30122
rect 29644 30058 29696 30064
rect 29656 30025 29684 30058
rect 29642 30016 29698 30025
rect 29642 29951 29698 29960
rect 29644 29776 29696 29782
rect 29644 29718 29696 29724
rect 29550 28928 29606 28937
rect 29550 28863 29606 28872
rect 29656 28801 29684 29718
rect 29748 29481 29776 30738
rect 29734 29472 29790 29481
rect 29734 29407 29790 29416
rect 29642 28792 29698 28801
rect 29642 28727 29698 28736
rect 29472 28580 29592 28608
rect 29000 28552 29052 28558
rect 28828 28512 29000 28540
rect 29000 28494 29052 28500
rect 29460 28484 29512 28490
rect 29460 28426 29512 28432
rect 28908 28416 28960 28422
rect 28908 28358 28960 28364
rect 29000 28416 29052 28422
rect 29000 28358 29052 28364
rect 28816 28076 28868 28082
rect 28816 28018 28868 28024
rect 28724 27464 28776 27470
rect 28724 27406 28776 27412
rect 28632 27328 28684 27334
rect 28632 27270 28684 27276
rect 28644 26761 28672 27270
rect 28828 27130 28856 28018
rect 28920 27470 28948 28358
rect 28908 27464 28960 27470
rect 28908 27406 28960 27412
rect 28816 27124 28868 27130
rect 28816 27066 28868 27072
rect 28908 26784 28960 26790
rect 28630 26752 28686 26761
rect 28908 26726 28960 26732
rect 28630 26687 28686 26696
rect 28920 26586 28948 26726
rect 28724 26580 28776 26586
rect 28724 26522 28776 26528
rect 28908 26580 28960 26586
rect 28908 26522 28960 26528
rect 28540 26036 28592 26042
rect 28540 25978 28592 25984
rect 28356 25832 28408 25838
rect 28356 25774 28408 25780
rect 28184 25622 28304 25650
rect 28184 25362 28212 25622
rect 28368 25362 28396 25774
rect 28448 25492 28500 25498
rect 28448 25434 28500 25440
rect 28172 25356 28224 25362
rect 28172 25298 28224 25304
rect 28356 25356 28408 25362
rect 28356 25298 28408 25304
rect 28078 25256 28134 25265
rect 28078 25191 28134 25200
rect 27804 24676 27856 24682
rect 27804 24618 27856 24624
rect 27896 24608 27948 24614
rect 27896 24550 27948 24556
rect 28080 24608 28132 24614
rect 28080 24550 28132 24556
rect 27710 24304 27766 24313
rect 27710 24239 27766 24248
rect 27712 23656 27764 23662
rect 27712 23598 27764 23604
rect 27724 21690 27752 23598
rect 27804 23180 27856 23186
rect 27804 23122 27856 23128
rect 27816 21944 27844 23122
rect 27908 23118 27936 24550
rect 27988 23860 28040 23866
rect 27988 23802 28040 23808
rect 27896 23112 27948 23118
rect 27896 23054 27948 23060
rect 28000 22930 28028 23802
rect 27908 22902 28028 22930
rect 27908 22098 27936 22902
rect 27988 22568 28040 22574
rect 27988 22510 28040 22516
rect 28000 22234 28028 22510
rect 27988 22228 28040 22234
rect 27988 22170 28040 22176
rect 27896 22092 27948 22098
rect 28092 22094 28120 24550
rect 28184 23866 28212 25298
rect 28264 25152 28316 25158
rect 28264 25094 28316 25100
rect 28172 23860 28224 23866
rect 28172 23802 28224 23808
rect 28172 23588 28224 23594
rect 28172 23530 28224 23536
rect 28184 23254 28212 23530
rect 28172 23248 28224 23254
rect 28172 23190 28224 23196
rect 28172 23044 28224 23050
rect 28172 22986 28224 22992
rect 27896 22034 27948 22040
rect 28000 22066 28120 22094
rect 27896 21956 27948 21962
rect 27816 21916 27896 21944
rect 27896 21898 27948 21904
rect 27712 21684 27764 21690
rect 27712 21626 27764 21632
rect 27908 21457 27936 21898
rect 27894 21448 27950 21457
rect 27894 21383 27950 21392
rect 27712 21004 27764 21010
rect 27712 20946 27764 20952
rect 27724 20074 27752 20946
rect 27896 20936 27948 20942
rect 27896 20878 27948 20884
rect 27724 20046 27844 20074
rect 27908 20058 27936 20878
rect 28000 20074 28028 22066
rect 28184 22030 28212 22986
rect 28276 22778 28304 25094
rect 28368 24206 28396 25298
rect 28460 24206 28488 25434
rect 28736 25294 28764 26522
rect 28816 26240 28868 26246
rect 28816 26182 28868 26188
rect 28828 25294 28856 26182
rect 28908 25900 28960 25906
rect 28908 25842 28960 25848
rect 28540 25288 28592 25294
rect 28540 25230 28592 25236
rect 28724 25288 28776 25294
rect 28724 25230 28776 25236
rect 28816 25288 28868 25294
rect 28816 25230 28868 25236
rect 28552 25140 28580 25230
rect 28552 25112 28764 25140
rect 28736 24818 28764 25112
rect 28632 24812 28684 24818
rect 28632 24754 28684 24760
rect 28724 24812 28776 24818
rect 28724 24754 28776 24760
rect 28356 24200 28408 24206
rect 28356 24142 28408 24148
rect 28448 24200 28500 24206
rect 28448 24142 28500 24148
rect 28540 24132 28592 24138
rect 28540 24074 28592 24080
rect 28354 24032 28410 24041
rect 28354 23967 28410 23976
rect 28264 22772 28316 22778
rect 28264 22714 28316 22720
rect 28262 22672 28318 22681
rect 28262 22607 28318 22616
rect 28276 22234 28304 22607
rect 28264 22228 28316 22234
rect 28264 22170 28316 22176
rect 28172 22024 28224 22030
rect 28172 21966 28224 21972
rect 28264 21956 28316 21962
rect 28264 21898 28316 21904
rect 28080 21888 28132 21894
rect 28276 21865 28304 21898
rect 28080 21830 28132 21836
rect 28262 21856 28318 21865
rect 28092 21321 28120 21830
rect 28262 21791 28318 21800
rect 28172 21548 28224 21554
rect 28172 21490 28224 21496
rect 28078 21312 28134 21321
rect 28078 21247 28134 21256
rect 28184 21010 28212 21490
rect 28172 21004 28224 21010
rect 28172 20946 28224 20952
rect 28172 20596 28224 20602
rect 28172 20538 28224 20544
rect 28000 20058 28120 20074
rect 27816 19514 27844 20046
rect 27896 20052 27948 20058
rect 28000 20052 28132 20058
rect 28000 20046 28080 20052
rect 27896 19994 27948 20000
rect 28080 19994 28132 20000
rect 27988 19848 28040 19854
rect 28184 19836 28212 20538
rect 28368 20058 28396 23967
rect 28448 23860 28500 23866
rect 28448 23802 28500 23808
rect 28460 23225 28488 23802
rect 28446 23216 28502 23225
rect 28446 23151 28502 23160
rect 28448 22636 28500 22642
rect 28448 22578 28500 22584
rect 28460 21457 28488 22578
rect 28446 21448 28502 21457
rect 28446 21383 28502 21392
rect 28356 20052 28408 20058
rect 28356 19994 28408 20000
rect 28040 19808 28212 19836
rect 27988 19790 28040 19796
rect 28000 19689 28028 19790
rect 28448 19780 28500 19786
rect 28448 19722 28500 19728
rect 27986 19680 28042 19689
rect 27986 19615 28042 19624
rect 27804 19508 27856 19514
rect 27804 19450 27856 19456
rect 27712 19440 27764 19446
rect 27712 19382 27764 19388
rect 27724 17678 27752 19382
rect 27896 18692 27948 18698
rect 27896 18634 27948 18640
rect 27712 17672 27764 17678
rect 27712 17614 27764 17620
rect 27724 17134 27752 17614
rect 27908 17338 27936 18634
rect 28460 17610 28488 19722
rect 28552 17882 28580 24074
rect 28644 20602 28672 24754
rect 28736 24041 28764 24754
rect 28816 24132 28868 24138
rect 28816 24074 28868 24080
rect 28722 24032 28778 24041
rect 28722 23967 28778 23976
rect 28724 23792 28776 23798
rect 28724 23734 28776 23740
rect 28736 23633 28764 23734
rect 28722 23624 28778 23633
rect 28722 23559 28778 23568
rect 28724 23520 28776 23526
rect 28724 23462 28776 23468
rect 28736 20942 28764 23462
rect 28724 20936 28776 20942
rect 28724 20878 28776 20884
rect 28632 20596 28684 20602
rect 28632 20538 28684 20544
rect 28724 20324 28776 20330
rect 28724 20266 28776 20272
rect 28632 20256 28684 20262
rect 28632 20198 28684 20204
rect 28644 19922 28672 20198
rect 28632 19916 28684 19922
rect 28632 19858 28684 19864
rect 28630 19816 28686 19825
rect 28630 19751 28686 19760
rect 28644 19174 28672 19751
rect 28736 19378 28764 20266
rect 28828 19786 28856 24074
rect 28920 23322 28948 25842
rect 29012 24750 29040 28358
rect 29110 27772 29418 27792
rect 29110 27770 29116 27772
rect 29172 27770 29196 27772
rect 29252 27770 29276 27772
rect 29332 27770 29356 27772
rect 29412 27770 29418 27772
rect 29172 27718 29174 27770
rect 29354 27718 29356 27770
rect 29110 27716 29116 27718
rect 29172 27716 29196 27718
rect 29252 27716 29276 27718
rect 29332 27716 29356 27718
rect 29412 27716 29418 27718
rect 29110 27696 29418 27716
rect 29472 27606 29500 28426
rect 29564 28257 29592 28580
rect 29550 28248 29606 28257
rect 29550 28183 29606 28192
rect 29644 28144 29696 28150
rect 29644 28086 29696 28092
rect 29552 27940 29604 27946
rect 29552 27882 29604 27888
rect 29460 27600 29512 27606
rect 29460 27542 29512 27548
rect 29564 27538 29592 27882
rect 29552 27532 29604 27538
rect 29552 27474 29604 27480
rect 29276 27464 29328 27470
rect 29276 27406 29328 27412
rect 29288 26926 29316 27406
rect 29276 26920 29328 26926
rect 29276 26862 29328 26868
rect 29550 26888 29606 26897
rect 29550 26823 29606 26832
rect 29110 26684 29418 26704
rect 29110 26682 29116 26684
rect 29172 26682 29196 26684
rect 29252 26682 29276 26684
rect 29332 26682 29356 26684
rect 29412 26682 29418 26684
rect 29172 26630 29174 26682
rect 29354 26630 29356 26682
rect 29110 26628 29116 26630
rect 29172 26628 29196 26630
rect 29252 26628 29276 26630
rect 29332 26628 29356 26630
rect 29412 26628 29418 26630
rect 29110 26608 29418 26628
rect 29564 26586 29592 26823
rect 29552 26580 29604 26586
rect 29552 26522 29604 26528
rect 29656 26450 29684 28086
rect 29736 26784 29788 26790
rect 29736 26726 29788 26732
rect 29748 26450 29776 26726
rect 29644 26444 29696 26450
rect 29644 26386 29696 26392
rect 29736 26444 29788 26450
rect 29736 26386 29788 26392
rect 29656 26042 29684 26386
rect 29644 26036 29696 26042
rect 29644 25978 29696 25984
rect 29736 25832 29788 25838
rect 29736 25774 29788 25780
rect 29110 25596 29418 25616
rect 29110 25594 29116 25596
rect 29172 25594 29196 25596
rect 29252 25594 29276 25596
rect 29332 25594 29356 25596
rect 29412 25594 29418 25596
rect 29172 25542 29174 25594
rect 29354 25542 29356 25594
rect 29110 25540 29116 25542
rect 29172 25540 29196 25542
rect 29252 25540 29276 25542
rect 29332 25540 29356 25542
rect 29412 25540 29418 25542
rect 29110 25520 29418 25540
rect 29644 25220 29696 25226
rect 29748 25208 29776 25774
rect 29696 25180 29776 25208
rect 29644 25162 29696 25168
rect 29000 24744 29052 24750
rect 29000 24686 29052 24692
rect 29458 24712 29514 24721
rect 29458 24647 29514 24656
rect 29472 24614 29500 24647
rect 29748 24614 29776 25180
rect 29460 24608 29512 24614
rect 29736 24608 29788 24614
rect 29460 24550 29512 24556
rect 29734 24576 29736 24585
rect 29788 24576 29790 24585
rect 29110 24508 29418 24528
rect 29734 24511 29790 24520
rect 29110 24506 29116 24508
rect 29172 24506 29196 24508
rect 29252 24506 29276 24508
rect 29332 24506 29356 24508
rect 29412 24506 29418 24508
rect 29172 24454 29174 24506
rect 29354 24454 29356 24506
rect 29110 24452 29116 24454
rect 29172 24452 29196 24454
rect 29252 24452 29276 24454
rect 29332 24452 29356 24454
rect 29412 24452 29418 24454
rect 29110 24432 29418 24452
rect 29552 24336 29604 24342
rect 29552 24278 29604 24284
rect 29184 24064 29236 24070
rect 29184 24006 29236 24012
rect 29460 24064 29512 24070
rect 29460 24006 29512 24012
rect 29000 23792 29052 23798
rect 29000 23734 29052 23740
rect 29012 23633 29040 23734
rect 29196 23662 29224 24006
rect 29184 23656 29236 23662
rect 28998 23624 29054 23633
rect 29184 23598 29236 23604
rect 28998 23559 29054 23568
rect 29110 23420 29418 23440
rect 29110 23418 29116 23420
rect 29172 23418 29196 23420
rect 29252 23418 29276 23420
rect 29332 23418 29356 23420
rect 29412 23418 29418 23420
rect 29172 23366 29174 23418
rect 29354 23366 29356 23418
rect 29110 23364 29116 23366
rect 29172 23364 29196 23366
rect 29252 23364 29276 23366
rect 29332 23364 29356 23366
rect 29412 23364 29418 23366
rect 29110 23344 29418 23364
rect 28908 23316 28960 23322
rect 28908 23258 28960 23264
rect 29368 23248 29420 23254
rect 28906 23216 28962 23225
rect 29368 23190 29420 23196
rect 28906 23151 28908 23160
rect 28960 23151 28962 23160
rect 28908 23122 28960 23128
rect 29000 23112 29052 23118
rect 29000 23054 29052 23060
rect 28908 22772 28960 22778
rect 28908 22714 28960 22720
rect 28816 19780 28868 19786
rect 28816 19722 28868 19728
rect 28724 19372 28776 19378
rect 28776 19332 28856 19360
rect 28724 19314 28776 19320
rect 28724 19236 28776 19242
rect 28724 19178 28776 19184
rect 28632 19168 28684 19174
rect 28632 19110 28684 19116
rect 28736 18970 28764 19178
rect 28724 18964 28776 18970
rect 28724 18906 28776 18912
rect 28736 18290 28764 18906
rect 28724 18284 28776 18290
rect 28724 18226 28776 18232
rect 28828 18086 28856 19332
rect 28816 18080 28868 18086
rect 28816 18022 28868 18028
rect 28920 17882 28948 22714
rect 29012 22574 29040 23054
rect 29380 23050 29408 23190
rect 29368 23044 29420 23050
rect 29368 22986 29420 22992
rect 29000 22568 29052 22574
rect 29000 22510 29052 22516
rect 29012 20942 29040 22510
rect 29110 22332 29418 22352
rect 29110 22330 29116 22332
rect 29172 22330 29196 22332
rect 29252 22330 29276 22332
rect 29332 22330 29356 22332
rect 29412 22330 29418 22332
rect 29172 22278 29174 22330
rect 29354 22278 29356 22330
rect 29110 22276 29116 22278
rect 29172 22276 29196 22278
rect 29252 22276 29276 22278
rect 29332 22276 29356 22278
rect 29412 22276 29418 22278
rect 29110 22256 29418 22276
rect 29184 22160 29236 22166
rect 29184 22102 29236 22108
rect 29196 21865 29224 22102
rect 29276 21956 29328 21962
rect 29276 21898 29328 21904
rect 29182 21856 29238 21865
rect 29182 21791 29238 21800
rect 29288 21593 29316 21898
rect 29274 21584 29330 21593
rect 29274 21519 29330 21528
rect 29110 21244 29418 21264
rect 29110 21242 29116 21244
rect 29172 21242 29196 21244
rect 29252 21242 29276 21244
rect 29332 21242 29356 21244
rect 29412 21242 29418 21244
rect 29172 21190 29174 21242
rect 29354 21190 29356 21242
rect 29110 21188 29116 21190
rect 29172 21188 29196 21190
rect 29252 21188 29276 21190
rect 29332 21188 29356 21190
rect 29412 21188 29418 21190
rect 29110 21168 29418 21188
rect 29472 21146 29500 24006
rect 29564 23526 29592 24278
rect 29644 24200 29696 24206
rect 29644 24142 29696 24148
rect 29656 23662 29684 24142
rect 29736 24064 29788 24070
rect 29736 24006 29788 24012
rect 29748 23866 29776 24006
rect 29736 23860 29788 23866
rect 29736 23802 29788 23808
rect 29644 23656 29696 23662
rect 29644 23598 29696 23604
rect 29552 23520 29604 23526
rect 29552 23462 29604 23468
rect 29656 21894 29684 23598
rect 29736 23316 29788 23322
rect 29736 23258 29788 23264
rect 29644 21888 29696 21894
rect 29644 21830 29696 21836
rect 29656 21690 29684 21830
rect 29644 21684 29696 21690
rect 29644 21626 29696 21632
rect 29552 21344 29604 21350
rect 29552 21286 29604 21292
rect 29460 21140 29512 21146
rect 29460 21082 29512 21088
rect 29564 21026 29592 21286
rect 29380 20998 29592 21026
rect 29000 20936 29052 20942
rect 29000 20878 29052 20884
rect 29012 19378 29040 20878
rect 29380 20602 29408 20998
rect 29460 20936 29512 20942
rect 29460 20878 29512 20884
rect 29368 20596 29420 20602
rect 29368 20538 29420 20544
rect 29472 20466 29500 20878
rect 29460 20460 29512 20466
rect 29460 20402 29512 20408
rect 29460 20256 29512 20262
rect 29460 20198 29512 20204
rect 29110 20156 29418 20176
rect 29110 20154 29116 20156
rect 29172 20154 29196 20156
rect 29252 20154 29276 20156
rect 29332 20154 29356 20156
rect 29412 20154 29418 20156
rect 29172 20102 29174 20154
rect 29354 20102 29356 20154
rect 29110 20100 29116 20102
rect 29172 20100 29196 20102
rect 29252 20100 29276 20102
rect 29332 20100 29356 20102
rect 29412 20100 29418 20102
rect 29110 20080 29418 20100
rect 29472 19990 29500 20198
rect 29460 19984 29512 19990
rect 29460 19926 29512 19932
rect 29460 19848 29512 19854
rect 29564 19836 29592 20998
rect 29644 20800 29696 20806
rect 29644 20742 29696 20748
rect 29512 19825 29592 19836
rect 29512 19816 29606 19825
rect 29512 19808 29550 19816
rect 29460 19790 29512 19796
rect 29550 19751 29606 19760
rect 29368 19712 29420 19718
rect 29368 19654 29420 19660
rect 29458 19680 29514 19689
rect 29274 19544 29330 19553
rect 29274 19479 29276 19488
rect 29328 19479 29330 19488
rect 29276 19450 29328 19456
rect 29380 19446 29408 19654
rect 29458 19615 29514 19624
rect 29368 19440 29420 19446
rect 29368 19382 29420 19388
rect 29000 19372 29052 19378
rect 29000 19314 29052 19320
rect 29012 18766 29040 19314
rect 29110 19068 29418 19088
rect 29110 19066 29116 19068
rect 29172 19066 29196 19068
rect 29252 19066 29276 19068
rect 29332 19066 29356 19068
rect 29412 19066 29418 19068
rect 29172 19014 29174 19066
rect 29354 19014 29356 19066
rect 29110 19012 29116 19014
rect 29172 19012 29196 19014
rect 29252 19012 29276 19014
rect 29332 19012 29356 19014
rect 29412 19012 29418 19014
rect 29110 18992 29418 19012
rect 29000 18760 29052 18766
rect 29000 18702 29052 18708
rect 29000 18080 29052 18086
rect 29000 18022 29052 18028
rect 28540 17876 28592 17882
rect 28540 17818 28592 17824
rect 28908 17876 28960 17882
rect 28908 17818 28960 17824
rect 28448 17604 28500 17610
rect 28448 17546 28500 17552
rect 27896 17332 27948 17338
rect 27896 17274 27948 17280
rect 29012 17270 29040 18022
rect 29110 17980 29418 18000
rect 29110 17978 29116 17980
rect 29172 17978 29196 17980
rect 29252 17978 29276 17980
rect 29332 17978 29356 17980
rect 29412 17978 29418 17980
rect 29172 17926 29174 17978
rect 29354 17926 29356 17978
rect 29110 17924 29116 17926
rect 29172 17924 29196 17926
rect 29252 17924 29276 17926
rect 29332 17924 29356 17926
rect 29412 17924 29418 17926
rect 29110 17904 29418 17924
rect 29472 17610 29500 19615
rect 29550 19408 29606 19417
rect 29550 19343 29606 19352
rect 29460 17604 29512 17610
rect 29460 17546 29512 17552
rect 29564 17542 29592 19343
rect 29656 18426 29684 20742
rect 29748 18426 29776 23258
rect 29644 18420 29696 18426
rect 29644 18362 29696 18368
rect 29736 18420 29788 18426
rect 29736 18362 29788 18368
rect 29552 17536 29604 17542
rect 29552 17478 29604 17484
rect 29000 17264 29052 17270
rect 29000 17206 29052 17212
rect 27712 17128 27764 17134
rect 27712 17070 27764 17076
rect 29110 16892 29418 16912
rect 29110 16890 29116 16892
rect 29172 16890 29196 16892
rect 29252 16890 29276 16892
rect 29332 16890 29356 16892
rect 29412 16890 29418 16892
rect 29172 16838 29174 16890
rect 29354 16838 29356 16890
rect 29110 16836 29116 16838
rect 29172 16836 29196 16838
rect 29252 16836 29276 16838
rect 29332 16836 29356 16838
rect 29412 16836 29418 16838
rect 29110 16816 29418 16836
rect 29110 15804 29418 15824
rect 29110 15802 29116 15804
rect 29172 15802 29196 15804
rect 29252 15802 29276 15804
rect 29332 15802 29356 15804
rect 29412 15802 29418 15804
rect 29172 15750 29174 15802
rect 29354 15750 29356 15802
rect 29110 15748 29116 15750
rect 29172 15748 29196 15750
rect 29252 15748 29276 15750
rect 29332 15748 29356 15750
rect 29412 15748 29418 15750
rect 29110 15728 29418 15748
rect 29110 14716 29418 14736
rect 29110 14714 29116 14716
rect 29172 14714 29196 14716
rect 29252 14714 29276 14716
rect 29332 14714 29356 14716
rect 29412 14714 29418 14716
rect 29172 14662 29174 14714
rect 29354 14662 29356 14714
rect 29110 14660 29116 14662
rect 29172 14660 29196 14662
rect 29252 14660 29276 14662
rect 29332 14660 29356 14662
rect 29412 14660 29418 14662
rect 29110 14640 29418 14660
rect 29110 13628 29418 13648
rect 29110 13626 29116 13628
rect 29172 13626 29196 13628
rect 29252 13626 29276 13628
rect 29332 13626 29356 13628
rect 29412 13626 29418 13628
rect 29172 13574 29174 13626
rect 29354 13574 29356 13626
rect 29110 13572 29116 13574
rect 29172 13572 29196 13574
rect 29252 13572 29276 13574
rect 29332 13572 29356 13574
rect 29412 13572 29418 13574
rect 29110 13552 29418 13572
rect 29110 12540 29418 12560
rect 29110 12538 29116 12540
rect 29172 12538 29196 12540
rect 29252 12538 29276 12540
rect 29332 12538 29356 12540
rect 29412 12538 29418 12540
rect 29172 12486 29174 12538
rect 29354 12486 29356 12538
rect 29110 12484 29116 12486
rect 29172 12484 29196 12486
rect 29252 12484 29276 12486
rect 29332 12484 29356 12486
rect 29412 12484 29418 12486
rect 29110 12464 29418 12484
rect 29110 11452 29418 11472
rect 29110 11450 29116 11452
rect 29172 11450 29196 11452
rect 29252 11450 29276 11452
rect 29332 11450 29356 11452
rect 29412 11450 29418 11452
rect 29172 11398 29174 11450
rect 29354 11398 29356 11450
rect 29110 11396 29116 11398
rect 29172 11396 29196 11398
rect 29252 11396 29276 11398
rect 29332 11396 29356 11398
rect 29412 11396 29418 11398
rect 29110 11376 29418 11396
rect 29110 10364 29418 10384
rect 29110 10362 29116 10364
rect 29172 10362 29196 10364
rect 29252 10362 29276 10364
rect 29332 10362 29356 10364
rect 29412 10362 29418 10364
rect 29172 10310 29174 10362
rect 29354 10310 29356 10362
rect 29110 10308 29116 10310
rect 29172 10308 29196 10310
rect 29252 10308 29276 10310
rect 29332 10308 29356 10310
rect 29412 10308 29418 10310
rect 29110 10288 29418 10308
rect 29110 9276 29418 9296
rect 29110 9274 29116 9276
rect 29172 9274 29196 9276
rect 29252 9274 29276 9276
rect 29332 9274 29356 9276
rect 29412 9274 29418 9276
rect 29172 9222 29174 9274
rect 29354 9222 29356 9274
rect 29110 9220 29116 9222
rect 29172 9220 29196 9222
rect 29252 9220 29276 9222
rect 29332 9220 29356 9222
rect 29412 9220 29418 9222
rect 29110 9200 29418 9220
rect 29110 8188 29418 8208
rect 29110 8186 29116 8188
rect 29172 8186 29196 8188
rect 29252 8186 29276 8188
rect 29332 8186 29356 8188
rect 29412 8186 29418 8188
rect 29172 8134 29174 8186
rect 29354 8134 29356 8186
rect 29110 8132 29116 8134
rect 29172 8132 29196 8134
rect 29252 8132 29276 8134
rect 29332 8132 29356 8134
rect 29412 8132 29418 8134
rect 29110 8112 29418 8132
rect 29736 7200 29788 7206
rect 29736 7142 29788 7148
rect 29110 7100 29418 7120
rect 29110 7098 29116 7100
rect 29172 7098 29196 7100
rect 29252 7098 29276 7100
rect 29332 7098 29356 7100
rect 29412 7098 29418 7100
rect 29172 7046 29174 7098
rect 29354 7046 29356 7098
rect 29110 7044 29116 7046
rect 29172 7044 29196 7046
rect 29252 7044 29276 7046
rect 29332 7044 29356 7046
rect 29412 7044 29418 7046
rect 29110 7024 29418 7044
rect 29110 6012 29418 6032
rect 29110 6010 29116 6012
rect 29172 6010 29196 6012
rect 29252 6010 29276 6012
rect 29332 6010 29356 6012
rect 29412 6010 29418 6012
rect 29172 5958 29174 6010
rect 29354 5958 29356 6010
rect 29110 5956 29116 5958
rect 29172 5956 29196 5958
rect 29252 5956 29276 5958
rect 29332 5956 29356 5958
rect 29412 5956 29418 5958
rect 29110 5936 29418 5956
rect 27620 5228 27672 5234
rect 27620 5170 27672 5176
rect 29644 5228 29696 5234
rect 29644 5170 29696 5176
rect 29552 5024 29604 5030
rect 29552 4966 29604 4972
rect 29110 4924 29418 4944
rect 29110 4922 29116 4924
rect 29172 4922 29196 4924
rect 29252 4922 29276 4924
rect 29332 4922 29356 4924
rect 29412 4922 29418 4924
rect 29172 4870 29174 4922
rect 29354 4870 29356 4922
rect 29110 4868 29116 4870
rect 29172 4868 29196 4870
rect 29252 4868 29276 4870
rect 29332 4868 29356 4870
rect 29412 4868 29418 4870
rect 29110 4848 29418 4868
rect 29564 4758 29592 4966
rect 29552 4752 29604 4758
rect 29552 4694 29604 4700
rect 29656 4570 29684 5170
rect 29564 4542 29684 4570
rect 23478 4380 23786 4400
rect 23478 4378 23484 4380
rect 23540 4378 23564 4380
rect 23620 4378 23644 4380
rect 23700 4378 23724 4380
rect 23780 4378 23786 4380
rect 23540 4326 23542 4378
rect 23722 4326 23724 4378
rect 23478 4324 23484 4326
rect 23540 4324 23564 4326
rect 23620 4324 23644 4326
rect 23700 4324 23724 4326
rect 23780 4324 23786 4326
rect 23478 4304 23786 4324
rect 21824 4140 21876 4146
rect 21824 4082 21876 4088
rect 19432 3936 19484 3942
rect 19432 3878 19484 3884
rect 20812 3936 20864 3942
rect 20812 3878 20864 3884
rect 18420 3528 18472 3534
rect 18420 3470 18472 3476
rect 19248 3528 19300 3534
rect 19248 3470 19300 3476
rect 19260 2854 19288 3470
rect 19248 2848 19300 2854
rect 19248 2790 19300 2796
rect 17846 2748 18154 2768
rect 17846 2746 17852 2748
rect 17908 2746 17932 2748
rect 17988 2746 18012 2748
rect 18068 2746 18092 2748
rect 18148 2746 18154 2748
rect 17908 2694 17910 2746
rect 18090 2694 18092 2746
rect 17846 2692 17852 2694
rect 17908 2692 17932 2694
rect 17988 2692 18012 2694
rect 18068 2692 18092 2694
rect 18148 2692 18154 2694
rect 17846 2672 18154 2692
rect 17500 2644 17552 2650
rect 17500 2586 17552 2592
rect 19444 2514 19472 3878
rect 20824 3602 20852 3878
rect 20812 3596 20864 3602
rect 20812 3538 20864 3544
rect 20352 3528 20404 3534
rect 20352 3470 20404 3476
rect 19616 3392 19668 3398
rect 19616 3334 19668 3340
rect 19628 2514 19656 3334
rect 20364 3126 20392 3470
rect 21272 3392 21324 3398
rect 21272 3334 21324 3340
rect 20352 3120 20404 3126
rect 20352 3062 20404 3068
rect 20628 2984 20680 2990
rect 20628 2926 20680 2932
rect 19432 2508 19484 2514
rect 19432 2450 19484 2456
rect 19616 2508 19668 2514
rect 19616 2450 19668 2456
rect 19984 2508 20036 2514
rect 19984 2450 20036 2456
rect 18052 2372 18104 2378
rect 18052 2314 18104 2320
rect 18064 800 18092 2314
rect 19996 800 20024 2450
rect 20640 800 20668 2926
rect 21284 800 21312 3334
rect 21836 3058 21864 4082
rect 27712 4072 27764 4078
rect 27712 4014 27764 4020
rect 28908 4072 28960 4078
rect 28908 4014 28960 4020
rect 23848 3528 23900 3534
rect 23848 3470 23900 3476
rect 21916 3460 21968 3466
rect 21916 3402 21968 3408
rect 21928 3194 21956 3402
rect 23478 3292 23786 3312
rect 23478 3290 23484 3292
rect 23540 3290 23564 3292
rect 23620 3290 23644 3292
rect 23700 3290 23724 3292
rect 23780 3290 23786 3292
rect 23540 3238 23542 3290
rect 23722 3238 23724 3290
rect 23478 3236 23484 3238
rect 23540 3236 23564 3238
rect 23620 3236 23644 3238
rect 23700 3236 23724 3238
rect 23780 3236 23786 3238
rect 23478 3216 23786 3236
rect 21916 3188 21968 3194
rect 21916 3130 21968 3136
rect 23860 3058 23888 3470
rect 27724 3058 27752 4014
rect 28356 4004 28408 4010
rect 28356 3946 28408 3952
rect 28368 3738 28396 3946
rect 28356 3732 28408 3738
rect 28356 3674 28408 3680
rect 27896 3528 27948 3534
rect 27896 3470 27948 3476
rect 21824 3052 21876 3058
rect 21824 2994 21876 3000
rect 23848 3052 23900 3058
rect 23848 2994 23900 3000
rect 27712 3052 27764 3058
rect 27712 2994 27764 3000
rect 27908 2990 27936 3470
rect 24492 2984 24544 2990
rect 27896 2984 27948 2990
rect 24492 2926 24544 2932
rect 27724 2932 27896 2938
rect 27724 2926 27948 2932
rect 21916 2916 21968 2922
rect 21916 2858 21968 2864
rect 21928 2650 21956 2858
rect 21916 2644 21968 2650
rect 21916 2586 21968 2592
rect 23478 2204 23786 2224
rect 23478 2202 23484 2204
rect 23540 2202 23564 2204
rect 23620 2202 23644 2204
rect 23700 2202 23724 2204
rect 23780 2202 23786 2204
rect 23540 2150 23542 2202
rect 23722 2150 23724 2202
rect 23478 2148 23484 2150
rect 23540 2148 23564 2150
rect 23620 2148 23644 2150
rect 23700 2148 23724 2150
rect 23780 2148 23786 2150
rect 23478 2128 23786 2148
rect 24504 800 24532 2926
rect 27724 2910 27936 2926
rect 27724 2854 27752 2910
rect 27712 2848 27764 2854
rect 27712 2790 27764 2796
rect 28920 2774 28948 4014
rect 29110 3836 29418 3856
rect 29110 3834 29116 3836
rect 29172 3834 29196 3836
rect 29252 3834 29276 3836
rect 29332 3834 29356 3836
rect 29412 3834 29418 3836
rect 29172 3782 29174 3834
rect 29354 3782 29356 3834
rect 29110 3780 29116 3782
rect 29172 3780 29196 3782
rect 29252 3780 29276 3782
rect 29332 3780 29356 3782
rect 29412 3780 29418 3782
rect 29110 3760 29418 3780
rect 29460 3528 29512 3534
rect 29564 3482 29592 4542
rect 29748 4146 29776 7142
rect 29840 5234 29868 31690
rect 29932 28422 29960 32807
rect 30024 32774 30052 33390
rect 30116 33114 30144 33510
rect 30104 33108 30156 33114
rect 30104 33050 30156 33056
rect 30012 32768 30064 32774
rect 30012 32710 30064 32716
rect 30012 32428 30064 32434
rect 30012 32370 30064 32376
rect 30024 30802 30052 32370
rect 30104 32224 30156 32230
rect 30104 32166 30156 32172
rect 30116 31890 30144 32166
rect 30104 31884 30156 31890
rect 30104 31826 30156 31832
rect 30208 31754 30236 34954
rect 30288 34400 30340 34406
rect 30288 34342 30340 34348
rect 30300 33318 30328 34342
rect 30288 33312 30340 33318
rect 30288 33254 30340 33260
rect 30392 32881 30420 36042
rect 30484 35873 30512 39442
rect 30840 39432 30892 39438
rect 30760 39392 30840 39420
rect 30656 38752 30708 38758
rect 30656 38694 30708 38700
rect 30668 37262 30696 38694
rect 30656 37256 30708 37262
rect 30656 37198 30708 37204
rect 30564 37188 30616 37194
rect 30564 37130 30616 37136
rect 30576 36718 30604 37130
rect 30564 36712 30616 36718
rect 30564 36654 30616 36660
rect 30668 36582 30696 37198
rect 30564 36576 30616 36582
rect 30564 36518 30616 36524
rect 30656 36576 30708 36582
rect 30656 36518 30708 36524
rect 30470 35864 30526 35873
rect 30470 35799 30526 35808
rect 30472 35488 30524 35494
rect 30472 35430 30524 35436
rect 30484 35222 30512 35430
rect 30472 35216 30524 35222
rect 30472 35158 30524 35164
rect 30472 35080 30524 35086
rect 30472 35022 30524 35028
rect 30484 34678 30512 35022
rect 30472 34672 30524 34678
rect 30472 34614 30524 34620
rect 30472 33924 30524 33930
rect 30472 33866 30524 33872
rect 30378 32872 30434 32881
rect 30378 32807 30434 32816
rect 30380 32768 30432 32774
rect 30380 32710 30432 32716
rect 30288 32564 30340 32570
rect 30288 32506 30340 32512
rect 30196 31748 30248 31754
rect 30196 31690 30248 31696
rect 30196 31476 30248 31482
rect 30196 31418 30248 31424
rect 30208 30841 30236 31418
rect 30300 31278 30328 32506
rect 30392 32008 30420 32710
rect 30484 32201 30512 33866
rect 30576 32450 30604 36518
rect 30760 34728 30788 39392
rect 30840 39374 30892 39380
rect 30932 39364 30984 39370
rect 30932 39306 30984 39312
rect 30840 39296 30892 39302
rect 30840 39238 30892 39244
rect 30668 34700 30788 34728
rect 30668 32745 30696 34700
rect 30748 34604 30800 34610
rect 30748 34546 30800 34552
rect 30760 34202 30788 34546
rect 30748 34196 30800 34202
rect 30748 34138 30800 34144
rect 30748 34060 30800 34066
rect 30748 34002 30800 34008
rect 30760 33454 30788 34002
rect 30748 33448 30800 33454
rect 30748 33390 30800 33396
rect 30748 33312 30800 33318
rect 30748 33254 30800 33260
rect 30654 32736 30710 32745
rect 30654 32671 30710 32680
rect 30668 32570 30696 32671
rect 30656 32564 30708 32570
rect 30656 32506 30708 32512
rect 30576 32422 30696 32450
rect 30470 32192 30526 32201
rect 30470 32127 30526 32136
rect 30668 32042 30696 32422
rect 30760 32366 30788 33254
rect 30748 32360 30800 32366
rect 30748 32302 30800 32308
rect 30760 32230 30788 32302
rect 30748 32224 30800 32230
rect 30852 32201 30880 39238
rect 30748 32166 30800 32172
rect 30838 32192 30894 32201
rect 30838 32127 30894 32136
rect 30564 32020 30616 32026
rect 30392 31980 30512 32008
rect 30380 31884 30432 31890
rect 30380 31826 30432 31832
rect 30392 31346 30420 31826
rect 30380 31340 30432 31346
rect 30380 31282 30432 31288
rect 30288 31272 30340 31278
rect 30288 31214 30340 31220
rect 30194 30832 30250 30841
rect 30012 30796 30064 30802
rect 30194 30767 30250 30776
rect 30012 30738 30064 30744
rect 30104 30728 30156 30734
rect 30104 30670 30156 30676
rect 30012 30388 30064 30394
rect 30012 30330 30064 30336
rect 30024 30297 30052 30330
rect 30010 30288 30066 30297
rect 30010 30223 30066 30232
rect 30116 29730 30144 30670
rect 30286 30560 30342 30569
rect 30286 30495 30342 30504
rect 30300 30122 30328 30495
rect 30392 30433 30420 31282
rect 30484 31192 30512 31980
rect 30668 32014 30880 32042
rect 30944 32026 30972 39306
rect 31208 37460 31260 37466
rect 31208 37402 31260 37408
rect 31116 36916 31168 36922
rect 31116 36858 31168 36864
rect 31024 36712 31076 36718
rect 31024 36654 31076 36660
rect 31036 34490 31064 36654
rect 31128 36242 31156 36858
rect 31116 36236 31168 36242
rect 31116 36178 31168 36184
rect 31036 34462 31156 34490
rect 31024 34400 31076 34406
rect 31024 34342 31076 34348
rect 31036 33998 31064 34342
rect 31024 33992 31076 33998
rect 31024 33934 31076 33940
rect 30564 31962 30616 31968
rect 30576 31346 30604 31962
rect 30746 31920 30802 31929
rect 30852 31906 30880 32014
rect 30932 32020 30984 32026
rect 30932 31962 30984 31968
rect 30852 31878 30972 31906
rect 30746 31855 30802 31864
rect 30656 31816 30708 31822
rect 30656 31758 30708 31764
rect 30564 31340 30616 31346
rect 30564 31282 30616 31288
rect 30564 31204 30616 31210
rect 30484 31164 30564 31192
rect 30564 31146 30616 31152
rect 30668 30598 30696 31758
rect 30656 30592 30708 30598
rect 30576 30552 30656 30580
rect 30378 30424 30434 30433
rect 30576 30394 30604 30552
rect 30656 30534 30708 30540
rect 30654 30424 30710 30433
rect 30378 30359 30434 30368
rect 30564 30388 30616 30394
rect 30654 30359 30656 30368
rect 30564 30330 30616 30336
rect 30708 30359 30710 30368
rect 30656 30330 30708 30336
rect 30760 30326 30788 31855
rect 30840 31340 30892 31346
rect 30840 31282 30892 31288
rect 30852 30938 30880 31282
rect 30840 30932 30892 30938
rect 30840 30874 30892 30880
rect 30748 30320 30800 30326
rect 30654 30288 30710 30297
rect 30748 30262 30800 30268
rect 30840 30320 30892 30326
rect 30840 30262 30892 30268
rect 30654 30223 30656 30232
rect 30708 30223 30710 30232
rect 30656 30194 30708 30200
rect 30760 30161 30788 30262
rect 30746 30152 30802 30161
rect 30288 30116 30340 30122
rect 30746 30087 30802 30096
rect 30288 30058 30340 30064
rect 30300 29850 30328 30058
rect 30852 30054 30880 30262
rect 30380 30048 30432 30054
rect 30840 30048 30892 30054
rect 30380 29990 30432 29996
rect 30838 30016 30840 30025
rect 30892 30016 30894 30025
rect 30288 29844 30340 29850
rect 30288 29786 30340 29792
rect 30196 29776 30248 29782
rect 30116 29724 30196 29730
rect 30116 29718 30248 29724
rect 30116 29702 30236 29718
rect 30012 29504 30064 29510
rect 30012 29446 30064 29452
rect 29920 28416 29972 28422
rect 29920 28358 29972 28364
rect 29920 28076 29972 28082
rect 29920 28018 29972 28024
rect 29932 27946 29960 28018
rect 29920 27940 29972 27946
rect 29920 27882 29972 27888
rect 29920 27532 29972 27538
rect 29920 27474 29972 27480
rect 29932 27130 29960 27474
rect 29920 27124 29972 27130
rect 29920 27066 29972 27072
rect 30024 26994 30052 29446
rect 30116 29238 30144 29702
rect 30104 29232 30156 29238
rect 30104 29174 30156 29180
rect 30116 28626 30144 29174
rect 30392 29170 30420 29990
rect 30838 29951 30894 29960
rect 30838 29880 30894 29889
rect 30838 29815 30894 29824
rect 30852 29714 30880 29815
rect 30472 29708 30524 29714
rect 30472 29650 30524 29656
rect 30840 29708 30892 29714
rect 30840 29650 30892 29656
rect 30380 29164 30432 29170
rect 30380 29106 30432 29112
rect 30196 28960 30248 28966
rect 30196 28902 30248 28908
rect 30104 28620 30156 28626
rect 30104 28562 30156 28568
rect 30208 28558 30236 28902
rect 30286 28656 30342 28665
rect 30286 28591 30342 28600
rect 30196 28552 30248 28558
rect 30196 28494 30248 28500
rect 30300 28098 30328 28591
rect 30300 28082 30420 28098
rect 30300 28076 30432 28082
rect 30300 28070 30380 28076
rect 30380 28018 30432 28024
rect 30196 27940 30248 27946
rect 30196 27882 30248 27888
rect 30104 27464 30156 27470
rect 30104 27406 30156 27412
rect 30116 27130 30144 27406
rect 30104 27124 30156 27130
rect 30104 27066 30156 27072
rect 30208 27062 30236 27882
rect 30288 27464 30340 27470
rect 30288 27406 30340 27412
rect 30196 27056 30248 27062
rect 30196 26998 30248 27004
rect 29920 26988 29972 26994
rect 29920 26930 29972 26936
rect 30012 26988 30064 26994
rect 30012 26930 30064 26936
rect 29932 26586 29960 26930
rect 29920 26580 29972 26586
rect 29920 26522 29972 26528
rect 30300 26518 30328 27406
rect 30380 27124 30432 27130
rect 30380 27066 30432 27072
rect 30392 26874 30420 27066
rect 30484 26994 30512 29650
rect 30656 29640 30708 29646
rect 30562 29608 30618 29617
rect 30656 29582 30708 29588
rect 30562 29543 30618 29552
rect 30576 27130 30604 29543
rect 30668 29481 30696 29582
rect 30654 29472 30710 29481
rect 30654 29407 30710 29416
rect 30564 27124 30616 27130
rect 30564 27066 30616 27072
rect 30668 27062 30696 29407
rect 30748 28076 30800 28082
rect 30748 28018 30800 28024
rect 30656 27056 30708 27062
rect 30656 26998 30708 27004
rect 30472 26988 30524 26994
rect 30524 26948 30604 26976
rect 30472 26930 30524 26936
rect 30392 26846 30512 26874
rect 30288 26512 30340 26518
rect 30288 26454 30340 26460
rect 30380 26512 30432 26518
rect 30380 26454 30432 26460
rect 30196 25288 30248 25294
rect 30196 25230 30248 25236
rect 30208 24750 30236 25230
rect 30196 24744 30248 24750
rect 30196 24686 30248 24692
rect 29920 24676 29972 24682
rect 29920 24618 29972 24624
rect 29932 24070 29960 24618
rect 30208 24206 30236 24686
rect 30196 24200 30248 24206
rect 30196 24142 30248 24148
rect 29920 24064 29972 24070
rect 29920 24006 29972 24012
rect 29920 23860 29972 23866
rect 29920 23802 29972 23808
rect 29932 23322 29960 23802
rect 29920 23316 29972 23322
rect 29920 23258 29972 23264
rect 29932 22234 29960 23258
rect 30392 23066 30420 26454
rect 30484 25702 30512 26846
rect 30576 25906 30604 26948
rect 30760 26450 30788 28018
rect 30852 27169 30880 29650
rect 30838 27160 30894 27169
rect 30944 27130 30972 31878
rect 31036 31657 31064 33934
rect 31022 31648 31078 31657
rect 31022 31583 31078 31592
rect 31024 30592 31076 30598
rect 31024 30534 31076 30540
rect 31036 28082 31064 30534
rect 31024 28076 31076 28082
rect 31024 28018 31076 28024
rect 31024 27532 31076 27538
rect 31024 27474 31076 27480
rect 31036 27305 31064 27474
rect 31022 27296 31078 27305
rect 31022 27231 31078 27240
rect 30838 27095 30894 27104
rect 30932 27124 30984 27130
rect 30932 27066 30984 27072
rect 31128 27010 31156 34462
rect 31220 34134 31248 37402
rect 31300 37188 31352 37194
rect 31300 37130 31352 37136
rect 31312 35766 31340 37130
rect 31404 36786 31432 39879
rect 31576 39636 31628 39642
rect 31576 39578 31628 39584
rect 31484 38820 31536 38826
rect 31484 38762 31536 38768
rect 31392 36780 31444 36786
rect 31392 36722 31444 36728
rect 31300 35760 31352 35766
rect 31300 35702 31352 35708
rect 31312 35601 31340 35702
rect 31298 35592 31354 35601
rect 31298 35527 31354 35536
rect 31300 34944 31352 34950
rect 31300 34886 31352 34892
rect 31208 34128 31260 34134
rect 31208 34070 31260 34076
rect 31208 33992 31260 33998
rect 31208 33934 31260 33940
rect 31220 33658 31248 33934
rect 31208 33652 31260 33658
rect 31208 33594 31260 33600
rect 31312 33522 31340 34886
rect 31392 34196 31444 34202
rect 31392 34138 31444 34144
rect 31404 33998 31432 34138
rect 31392 33992 31444 33998
rect 31392 33934 31444 33940
rect 31300 33516 31352 33522
rect 31300 33458 31352 33464
rect 31300 33380 31352 33386
rect 31300 33322 31352 33328
rect 31208 33108 31260 33114
rect 31208 33050 31260 33056
rect 31220 30122 31248 33050
rect 31208 30116 31260 30122
rect 31208 30058 31260 30064
rect 31312 30054 31340 33322
rect 31404 31929 31432 33934
rect 31496 33046 31524 38762
rect 31588 35193 31616 39578
rect 31864 38418 31892 40530
rect 31944 40180 31996 40186
rect 31944 40122 31996 40128
rect 31956 38962 31984 40122
rect 32496 39976 32548 39982
rect 32496 39918 32548 39924
rect 32126 39536 32182 39545
rect 32126 39471 32182 39480
rect 32034 39400 32090 39409
rect 32034 39335 32090 39344
rect 31944 38956 31996 38962
rect 31944 38898 31996 38904
rect 31852 38412 31904 38418
rect 31852 38354 31904 38360
rect 31942 37904 31998 37913
rect 32048 37874 32076 39335
rect 31942 37839 31998 37848
rect 32036 37868 32088 37874
rect 31668 37120 31720 37126
rect 31668 37062 31720 37068
rect 31574 35184 31630 35193
rect 31574 35119 31630 35128
rect 31576 34740 31628 34746
rect 31576 34682 31628 34688
rect 31588 34610 31616 34682
rect 31576 34604 31628 34610
rect 31576 34546 31628 34552
rect 31574 33416 31630 33425
rect 31574 33351 31630 33360
rect 31484 33040 31536 33046
rect 31484 32982 31536 32988
rect 31484 32428 31536 32434
rect 31484 32370 31536 32376
rect 31496 31958 31524 32370
rect 31484 31952 31536 31958
rect 31390 31920 31446 31929
rect 31484 31894 31536 31900
rect 31390 31855 31446 31864
rect 31484 31816 31536 31822
rect 31482 31784 31484 31793
rect 31536 31784 31538 31793
rect 31404 31742 31482 31770
rect 31404 30580 31432 31742
rect 31482 31719 31538 31728
rect 31588 31736 31616 33351
rect 31680 32910 31708 37062
rect 31852 36780 31904 36786
rect 31852 36722 31904 36728
rect 31864 34490 31892 36722
rect 31956 36718 31984 37839
rect 32036 37810 32088 37816
rect 32140 37262 32168 39471
rect 32312 39432 32364 39438
rect 32312 39374 32364 39380
rect 32324 39001 32352 39374
rect 32508 39030 32536 39918
rect 32496 39024 32548 39030
rect 32310 38992 32366 39001
rect 32496 38966 32548 38972
rect 32310 38927 32366 38936
rect 32496 38276 32548 38282
rect 32496 38218 32548 38224
rect 32128 37256 32180 37262
rect 32128 37198 32180 37204
rect 32312 37188 32364 37194
rect 32312 37130 32364 37136
rect 32324 36854 32352 37130
rect 32508 36922 32536 38218
rect 32876 37330 32904 41200
rect 32954 39536 33010 39545
rect 32954 39471 33010 39480
rect 32864 37324 32916 37330
rect 32864 37266 32916 37272
rect 32496 36916 32548 36922
rect 32496 36858 32548 36864
rect 32312 36848 32364 36854
rect 32312 36790 32364 36796
rect 31944 36712 31996 36718
rect 31944 36654 31996 36660
rect 32310 36272 32366 36281
rect 32968 36242 32996 39471
rect 33520 38894 33548 41200
rect 34164 41018 34192 41200
rect 34072 40990 34192 41018
rect 33508 38888 33560 38894
rect 33508 38830 33560 38836
rect 33046 38176 33102 38185
rect 33046 38111 33102 38120
rect 33060 37942 33088 38111
rect 34072 37942 34100 40990
rect 34150 40896 34206 40905
rect 34150 40831 34206 40840
rect 34164 39506 34192 40831
rect 34152 39500 34204 39506
rect 34152 39442 34204 39448
rect 34150 38856 34206 38865
rect 34150 38791 34206 38800
rect 34164 38418 34192 38791
rect 34152 38412 34204 38418
rect 34152 38354 34204 38360
rect 33048 37936 33100 37942
rect 33048 37878 33100 37884
rect 34060 37936 34112 37942
rect 34060 37878 34112 37884
rect 33416 37120 33468 37126
rect 33416 37062 33468 37068
rect 32310 36207 32312 36216
rect 32364 36207 32366 36216
rect 32956 36236 33008 36242
rect 32312 36178 32364 36184
rect 32956 36178 33008 36184
rect 33322 36136 33378 36145
rect 33322 36071 33378 36080
rect 32496 35760 32548 35766
rect 32496 35702 32548 35708
rect 32036 35692 32088 35698
rect 32036 35634 32088 35640
rect 32404 35692 32456 35698
rect 32404 35634 32456 35640
rect 31944 35080 31996 35086
rect 31944 35022 31996 35028
rect 31772 34462 31892 34490
rect 31668 32904 31720 32910
rect 31668 32846 31720 32852
rect 31668 32360 31720 32366
rect 31668 32302 31720 32308
rect 31680 32026 31708 32302
rect 31668 32020 31720 32026
rect 31668 31962 31720 31968
rect 31588 31708 31708 31736
rect 31576 31136 31628 31142
rect 31576 31078 31628 31084
rect 31588 30734 31616 31078
rect 31484 30728 31536 30734
rect 31482 30696 31484 30705
rect 31576 30728 31628 30734
rect 31536 30696 31538 30705
rect 31576 30670 31628 30676
rect 31482 30631 31538 30640
rect 31404 30552 31616 30580
rect 31300 30048 31352 30054
rect 31484 30048 31536 30054
rect 31300 29990 31352 29996
rect 31404 29996 31484 30002
rect 31404 29990 31536 29996
rect 31404 29974 31524 29990
rect 31300 29504 31352 29510
rect 31300 29446 31352 29452
rect 31312 29102 31340 29446
rect 31300 29096 31352 29102
rect 31404 29073 31432 29974
rect 31300 29038 31352 29044
rect 31390 29064 31446 29073
rect 31390 28999 31446 29008
rect 31588 28626 31616 30552
rect 31680 30326 31708 31708
rect 31668 30320 31720 30326
rect 31668 30262 31720 30268
rect 31666 29744 31722 29753
rect 31666 29679 31722 29688
rect 31680 29306 31708 29679
rect 31668 29300 31720 29306
rect 31668 29242 31720 29248
rect 31666 29200 31722 29209
rect 31666 29135 31668 29144
rect 31720 29135 31722 29144
rect 31668 29106 31720 29112
rect 31576 28620 31628 28626
rect 31576 28562 31628 28568
rect 31392 28416 31444 28422
rect 31392 28358 31444 28364
rect 31404 28218 31432 28358
rect 31392 28212 31444 28218
rect 31392 28154 31444 28160
rect 31300 27872 31352 27878
rect 31300 27814 31352 27820
rect 31208 27532 31260 27538
rect 31208 27474 31260 27480
rect 30852 26982 31156 27010
rect 30656 26444 30708 26450
rect 30656 26386 30708 26392
rect 30748 26444 30800 26450
rect 30748 26386 30800 26392
rect 30668 25974 30696 26386
rect 30656 25968 30708 25974
rect 30654 25936 30656 25945
rect 30708 25936 30710 25945
rect 30564 25900 30616 25906
rect 30654 25871 30710 25880
rect 30564 25842 30616 25848
rect 30472 25696 30524 25702
rect 30524 25656 30604 25684
rect 30472 25638 30524 25644
rect 30576 23526 30604 25656
rect 30656 25220 30708 25226
rect 30656 25162 30708 25168
rect 30564 23520 30616 23526
rect 30564 23462 30616 23468
rect 30300 23038 30420 23066
rect 30564 23044 30616 23050
rect 30196 22976 30248 22982
rect 30196 22918 30248 22924
rect 30010 22536 30066 22545
rect 30010 22471 30066 22480
rect 29920 22228 29972 22234
rect 29920 22170 29972 22176
rect 30024 22098 30052 22471
rect 30104 22432 30156 22438
rect 30102 22400 30104 22409
rect 30156 22400 30158 22409
rect 30102 22335 30158 22344
rect 30102 22264 30158 22273
rect 30102 22199 30158 22208
rect 29920 22092 29972 22098
rect 29920 22034 29972 22040
rect 30012 22092 30064 22098
rect 30012 22034 30064 22040
rect 29932 21672 29960 22034
rect 30012 21684 30064 21690
rect 29932 21644 30012 21672
rect 30012 21626 30064 21632
rect 29920 21412 29972 21418
rect 29920 21354 29972 21360
rect 29932 18358 29960 21354
rect 30024 20097 30052 21626
rect 30116 20448 30144 22199
rect 30208 20874 30236 22918
rect 30300 22094 30328 23038
rect 30564 22986 30616 22992
rect 30380 22976 30432 22982
rect 30380 22918 30432 22924
rect 30392 22642 30420 22918
rect 30576 22778 30604 22986
rect 30564 22772 30616 22778
rect 30564 22714 30616 22720
rect 30562 22672 30618 22681
rect 30380 22636 30432 22642
rect 30380 22578 30432 22584
rect 30472 22636 30524 22642
rect 30562 22607 30618 22616
rect 30472 22578 30524 22584
rect 30378 22536 30434 22545
rect 30378 22471 30380 22480
rect 30432 22471 30434 22480
rect 30380 22442 30432 22448
rect 30300 22066 30436 22094
rect 30408 22012 30436 22066
rect 30286 21992 30342 22001
rect 30286 21927 30288 21936
rect 30340 21927 30342 21936
rect 30392 21984 30436 22012
rect 30288 21898 30340 21904
rect 30196 20868 30248 20874
rect 30196 20810 30248 20816
rect 30116 20420 30328 20448
rect 30196 20324 30248 20330
rect 30196 20266 30248 20272
rect 30104 20256 30156 20262
rect 30104 20198 30156 20204
rect 30010 20088 30066 20097
rect 30010 20023 30066 20032
rect 30012 19984 30064 19990
rect 30012 19926 30064 19932
rect 30024 19825 30052 19926
rect 30010 19816 30066 19825
rect 30010 19751 30066 19760
rect 29920 18352 29972 18358
rect 29920 18294 29972 18300
rect 30024 18290 30052 19751
rect 30116 18766 30144 20198
rect 30208 20058 30236 20266
rect 30196 20052 30248 20058
rect 30196 19994 30248 20000
rect 30194 19952 30250 19961
rect 30194 19887 30250 19896
rect 30104 18760 30156 18766
rect 30104 18702 30156 18708
rect 30102 18592 30158 18601
rect 30102 18527 30158 18536
rect 30012 18284 30064 18290
rect 30012 18226 30064 18232
rect 30116 16658 30144 18527
rect 30208 17678 30236 19887
rect 30196 17672 30248 17678
rect 30196 17614 30248 17620
rect 30300 17202 30328 20420
rect 30392 19334 30420 21984
rect 30484 21894 30512 22578
rect 30472 21888 30524 21894
rect 30472 21830 30524 21836
rect 30484 21554 30512 21830
rect 30472 21548 30524 21554
rect 30472 21490 30524 21496
rect 30472 21412 30524 21418
rect 30472 21354 30524 21360
rect 30484 21321 30512 21354
rect 30470 21312 30526 21321
rect 30470 21247 30526 21256
rect 30472 20528 30524 20534
rect 30472 20470 30524 20476
rect 30484 19786 30512 20470
rect 30472 19780 30524 19786
rect 30472 19722 30524 19728
rect 30392 19306 30512 19334
rect 30380 19236 30432 19242
rect 30380 19178 30432 19184
rect 30392 18290 30420 19178
rect 30380 18284 30432 18290
rect 30380 18226 30432 18232
rect 30392 17746 30420 18226
rect 30380 17740 30432 17746
rect 30380 17682 30432 17688
rect 30484 17338 30512 19306
rect 30576 17678 30604 22607
rect 30668 21554 30696 25162
rect 30748 24812 30800 24818
rect 30748 24754 30800 24760
rect 30656 21548 30708 21554
rect 30656 21490 30708 21496
rect 30656 21344 30708 21350
rect 30656 21286 30708 21292
rect 30668 21146 30696 21286
rect 30656 21140 30708 21146
rect 30656 21082 30708 21088
rect 30656 19848 30708 19854
rect 30656 19790 30708 19796
rect 30668 19514 30696 19790
rect 30656 19508 30708 19514
rect 30656 19450 30708 19456
rect 30654 19408 30710 19417
rect 30654 19343 30710 19352
rect 30668 18154 30696 19343
rect 30760 18426 30788 24754
rect 30748 18420 30800 18426
rect 30748 18362 30800 18368
rect 30656 18148 30708 18154
rect 30656 18090 30708 18096
rect 30564 17672 30616 17678
rect 30564 17614 30616 17620
rect 30472 17332 30524 17338
rect 30472 17274 30524 17280
rect 30288 17196 30340 17202
rect 30288 17138 30340 17144
rect 30104 16652 30156 16658
rect 30104 16594 30156 16600
rect 30852 12434 30880 26982
rect 31220 26926 31248 27474
rect 31208 26920 31260 26926
rect 31208 26862 31260 26868
rect 30932 25900 30984 25906
rect 30932 25842 30984 25848
rect 30944 25158 30972 25842
rect 31024 25696 31076 25702
rect 31024 25638 31076 25644
rect 30932 25152 30984 25158
rect 30932 25094 30984 25100
rect 30944 22574 30972 25094
rect 31036 24886 31064 25638
rect 31116 25356 31168 25362
rect 31116 25298 31168 25304
rect 31024 24880 31076 24886
rect 31024 24822 31076 24828
rect 31036 23730 31064 24822
rect 31128 23866 31156 25298
rect 31116 23860 31168 23866
rect 31116 23802 31168 23808
rect 31024 23724 31076 23730
rect 31024 23666 31076 23672
rect 30932 22568 30984 22574
rect 30932 22510 30984 22516
rect 30930 22400 30986 22409
rect 30930 22335 30986 22344
rect 30944 21894 30972 22335
rect 31036 22030 31064 23666
rect 31024 22024 31076 22030
rect 31024 21966 31076 21972
rect 30932 21888 30984 21894
rect 30932 21830 30984 21836
rect 31036 21554 31064 21966
rect 31024 21548 31076 21554
rect 31024 21490 31076 21496
rect 30930 21448 30986 21457
rect 30930 21383 30986 21392
rect 30944 20262 30972 21383
rect 31024 20800 31076 20806
rect 31022 20768 31024 20777
rect 31076 20768 31078 20777
rect 31022 20703 31078 20712
rect 31024 20392 31076 20398
rect 31024 20334 31076 20340
rect 30932 20256 30984 20262
rect 30932 20198 30984 20204
rect 30932 19780 30984 19786
rect 30932 19722 30984 19728
rect 30944 18970 30972 19722
rect 30932 18964 30984 18970
rect 30932 18906 30984 18912
rect 31036 16794 31064 20334
rect 31128 18358 31156 23802
rect 31220 18970 31248 26862
rect 31312 26518 31340 27814
rect 31300 26512 31352 26518
rect 31300 26454 31352 26460
rect 31404 26364 31432 28154
rect 31772 27878 31800 34462
rect 31850 33960 31906 33969
rect 31850 33895 31906 33904
rect 31864 33590 31892 33895
rect 31852 33584 31904 33590
rect 31852 33526 31904 33532
rect 31956 33046 31984 35022
rect 32048 33318 32076 35634
rect 32220 35488 32272 35494
rect 32220 35430 32272 35436
rect 32128 35012 32180 35018
rect 32128 34954 32180 34960
rect 32140 34746 32168 34954
rect 32128 34740 32180 34746
rect 32128 34682 32180 34688
rect 32036 33312 32088 33318
rect 32036 33254 32088 33260
rect 31944 33040 31996 33046
rect 31944 32982 31996 32988
rect 32034 33008 32090 33017
rect 32034 32943 32090 32952
rect 32048 32910 32076 32943
rect 32036 32904 32088 32910
rect 32036 32846 32088 32852
rect 31852 32768 31904 32774
rect 31852 32710 31904 32716
rect 31864 30190 31892 32710
rect 32036 31952 32088 31958
rect 32036 31894 32088 31900
rect 31944 31884 31996 31890
rect 31944 31826 31996 31832
rect 31956 30870 31984 31826
rect 31944 30864 31996 30870
rect 31944 30806 31996 30812
rect 32048 30802 32076 31894
rect 32128 31476 32180 31482
rect 32128 31418 32180 31424
rect 32036 30796 32088 30802
rect 32036 30738 32088 30744
rect 31944 30728 31996 30734
rect 31944 30670 31996 30676
rect 31956 30598 31984 30670
rect 31944 30592 31996 30598
rect 31944 30534 31996 30540
rect 31956 30190 31984 30534
rect 31852 30184 31904 30190
rect 31852 30126 31904 30132
rect 31944 30184 31996 30190
rect 31944 30126 31996 30132
rect 32036 29844 32088 29850
rect 32036 29786 32088 29792
rect 31850 29744 31906 29753
rect 31850 29679 31906 29688
rect 31864 29170 31892 29679
rect 32048 29492 32076 29786
rect 32140 29646 32168 31418
rect 32232 30802 32260 35430
rect 32416 35222 32444 35634
rect 32404 35216 32456 35222
rect 32324 35176 32404 35204
rect 32324 34610 32352 35176
rect 32404 35158 32456 35164
rect 32404 34944 32456 34950
rect 32404 34886 32456 34892
rect 32312 34604 32364 34610
rect 32312 34546 32364 34552
rect 32310 34504 32366 34513
rect 32310 34439 32366 34448
rect 32324 33522 32352 34439
rect 32312 33516 32364 33522
rect 32312 33458 32364 33464
rect 32310 32464 32366 32473
rect 32310 32399 32312 32408
rect 32364 32399 32366 32408
rect 32312 32370 32364 32376
rect 32310 32328 32366 32337
rect 32310 32263 32366 32272
rect 32324 31890 32352 32263
rect 32312 31884 32364 31890
rect 32312 31826 32364 31832
rect 32312 31272 32364 31278
rect 32310 31240 32312 31249
rect 32364 31240 32366 31249
rect 32310 31175 32366 31184
rect 32310 30832 32366 30841
rect 32220 30796 32272 30802
rect 32310 30767 32366 30776
rect 32220 30738 32272 30744
rect 32324 30734 32352 30767
rect 32312 30728 32364 30734
rect 32312 30670 32364 30676
rect 32128 29640 32180 29646
rect 32128 29582 32180 29588
rect 32048 29464 32260 29492
rect 31852 29164 31904 29170
rect 31852 29106 31904 29112
rect 31944 28552 31996 28558
rect 31944 28494 31996 28500
rect 32128 28552 32180 28558
rect 32128 28494 32180 28500
rect 31484 27872 31536 27878
rect 31484 27814 31536 27820
rect 31760 27872 31812 27878
rect 31760 27814 31812 27820
rect 31496 27062 31524 27814
rect 31956 27674 31984 28494
rect 32036 28416 32088 28422
rect 32036 28358 32088 28364
rect 31944 27668 31996 27674
rect 31944 27610 31996 27616
rect 31668 27600 31720 27606
rect 31668 27542 31720 27548
rect 31576 27464 31628 27470
rect 31576 27406 31628 27412
rect 31588 27130 31616 27406
rect 31576 27124 31628 27130
rect 31576 27066 31628 27072
rect 31680 27062 31708 27542
rect 32048 27538 32076 28358
rect 32036 27532 32088 27538
rect 32036 27474 32088 27480
rect 31760 27464 31812 27470
rect 31760 27406 31812 27412
rect 31484 27056 31536 27062
rect 31484 26998 31536 27004
rect 31668 27056 31720 27062
rect 31668 26998 31720 27004
rect 31772 26994 31800 27406
rect 31760 26988 31812 26994
rect 31812 26948 31892 26976
rect 31760 26930 31812 26936
rect 31760 26784 31812 26790
rect 31760 26726 31812 26732
rect 31668 26512 31720 26518
rect 31668 26454 31720 26460
rect 31312 26336 31432 26364
rect 31312 24818 31340 26336
rect 31484 25492 31536 25498
rect 31484 25434 31536 25440
rect 31496 25401 31524 25434
rect 31482 25392 31538 25401
rect 31482 25327 31538 25336
rect 31484 25288 31536 25294
rect 31484 25230 31536 25236
rect 31392 25152 31444 25158
rect 31392 25094 31444 25100
rect 31300 24812 31352 24818
rect 31300 24754 31352 24760
rect 31300 24608 31352 24614
rect 31300 24550 31352 24556
rect 31312 23866 31340 24550
rect 31404 24138 31432 25094
rect 31392 24132 31444 24138
rect 31392 24074 31444 24080
rect 31300 23860 31352 23866
rect 31300 23802 31352 23808
rect 31298 23760 31354 23769
rect 31298 23695 31354 23704
rect 31312 23322 31340 23695
rect 31392 23656 31444 23662
rect 31392 23598 31444 23604
rect 31300 23316 31352 23322
rect 31300 23258 31352 23264
rect 31300 23180 31352 23186
rect 31300 23122 31352 23128
rect 31312 23089 31340 23122
rect 31298 23080 31354 23089
rect 31298 23015 31354 23024
rect 31300 22704 31352 22710
rect 31300 22646 31352 22652
rect 31208 18964 31260 18970
rect 31208 18906 31260 18912
rect 31116 18352 31168 18358
rect 31116 18294 31168 18300
rect 31312 17202 31340 22646
rect 31404 22166 31432 23598
rect 31392 22160 31444 22166
rect 31392 22102 31444 22108
rect 31392 21684 31444 21690
rect 31392 21626 31444 21632
rect 31404 18290 31432 21626
rect 31392 18284 31444 18290
rect 31392 18226 31444 18232
rect 31496 17882 31524 25230
rect 31680 24721 31708 26454
rect 31666 24712 31722 24721
rect 31666 24647 31722 24656
rect 31680 24614 31708 24647
rect 31668 24608 31720 24614
rect 31668 24550 31720 24556
rect 31680 23662 31708 24550
rect 31668 23656 31720 23662
rect 31668 23598 31720 23604
rect 31668 23520 31720 23526
rect 31668 23462 31720 23468
rect 31680 22778 31708 23462
rect 31668 22772 31720 22778
rect 31668 22714 31720 22720
rect 31680 22681 31708 22714
rect 31666 22672 31722 22681
rect 31666 22607 31722 22616
rect 31772 22556 31800 26726
rect 31864 25362 31892 26948
rect 32048 25906 32076 27474
rect 32140 27470 32168 28494
rect 32128 27464 32180 27470
rect 32128 27406 32180 27412
rect 32128 26376 32180 26382
rect 32128 26318 32180 26324
rect 31944 25900 31996 25906
rect 31944 25842 31996 25848
rect 32036 25900 32088 25906
rect 32036 25842 32088 25848
rect 31852 25356 31904 25362
rect 31852 25298 31904 25304
rect 31864 24954 31892 25298
rect 31852 24948 31904 24954
rect 31852 24890 31904 24896
rect 31864 24410 31892 24890
rect 31852 24404 31904 24410
rect 31852 24346 31904 24352
rect 31852 23860 31904 23866
rect 31852 23802 31904 23808
rect 31864 22574 31892 23802
rect 31680 22528 31800 22556
rect 31852 22568 31904 22574
rect 31850 22536 31852 22545
rect 31904 22536 31906 22545
rect 31680 22234 31708 22528
rect 31850 22471 31906 22480
rect 31760 22432 31812 22438
rect 31758 22400 31760 22409
rect 31852 22432 31904 22438
rect 31812 22400 31814 22409
rect 31852 22374 31904 22380
rect 31758 22335 31814 22344
rect 31668 22228 31720 22234
rect 31668 22170 31720 22176
rect 31668 22092 31720 22098
rect 31668 22034 31720 22040
rect 31576 21888 31628 21894
rect 31680 21865 31708 22034
rect 31772 22030 31800 22335
rect 31760 22024 31812 22030
rect 31760 21966 31812 21972
rect 31576 21830 31628 21836
rect 31666 21856 31722 21865
rect 31588 21690 31616 21830
rect 31666 21791 31722 21800
rect 31576 21684 31628 21690
rect 31576 21626 31628 21632
rect 31576 21344 31628 21350
rect 31576 21286 31628 21292
rect 31588 21146 31616 21286
rect 31576 21140 31628 21146
rect 31576 21082 31628 21088
rect 31588 20534 31616 21082
rect 31576 20528 31628 20534
rect 31576 20470 31628 20476
rect 31772 20380 31800 21966
rect 31864 21418 31892 22374
rect 31956 22094 31984 25842
rect 32036 25764 32088 25770
rect 32036 25706 32088 25712
rect 32048 24886 32076 25706
rect 32036 24880 32088 24886
rect 32036 24822 32088 24828
rect 32140 24750 32168 26318
rect 32232 26234 32260 29464
rect 32310 28112 32366 28121
rect 32310 28047 32312 28056
rect 32364 28047 32366 28056
rect 32312 28018 32364 28024
rect 32312 27464 32364 27470
rect 32312 27406 32364 27412
rect 32324 26382 32352 27406
rect 32416 27130 32444 34886
rect 32508 34746 32536 35702
rect 33336 35698 33364 36071
rect 33324 35692 33376 35698
rect 33324 35634 33376 35640
rect 33230 34776 33286 34785
rect 32496 34740 32548 34746
rect 33230 34711 33286 34720
rect 32496 34682 32548 34688
rect 33244 34678 33272 34711
rect 32680 34672 32732 34678
rect 32680 34614 32732 34620
rect 33232 34672 33284 34678
rect 33232 34614 33284 34620
rect 32496 34604 32548 34610
rect 32496 34546 32548 34552
rect 32508 34066 32536 34546
rect 32496 34060 32548 34066
rect 32496 34002 32548 34008
rect 32496 33924 32548 33930
rect 32496 33866 32548 33872
rect 32508 29850 32536 33866
rect 32692 33658 32720 34614
rect 33428 34610 33456 37062
rect 34150 36816 34206 36825
rect 34150 36751 34152 36760
rect 34204 36751 34206 36760
rect 34152 36722 34204 36728
rect 34336 36576 34388 36582
rect 34336 36518 34388 36524
rect 33508 35216 33560 35222
rect 33508 35158 33560 35164
rect 32772 34604 32824 34610
rect 32772 34546 32824 34552
rect 33416 34604 33468 34610
rect 33416 34546 33468 34552
rect 32784 34202 32812 34546
rect 32772 34196 32824 34202
rect 32772 34138 32824 34144
rect 33232 33856 33284 33862
rect 33232 33798 33284 33804
rect 32680 33652 32732 33658
rect 32680 33594 32732 33600
rect 32586 33280 32642 33289
rect 32586 33215 32642 33224
rect 32600 31890 32628 33215
rect 33048 32768 33100 32774
rect 33048 32710 33100 32716
rect 32588 31884 32640 31890
rect 32588 31826 32640 31832
rect 33060 30666 33088 32710
rect 33138 32600 33194 32609
rect 33138 32535 33194 32544
rect 33048 30660 33100 30666
rect 33048 30602 33100 30608
rect 33152 30258 33180 32535
rect 33140 30252 33192 30258
rect 33140 30194 33192 30200
rect 33140 30048 33192 30054
rect 33140 29990 33192 29996
rect 32496 29844 32548 29850
rect 32496 29786 32548 29792
rect 33048 29844 33100 29850
rect 33048 29786 33100 29792
rect 32864 29572 32916 29578
rect 32864 29514 32916 29520
rect 32876 29306 32904 29514
rect 32864 29300 32916 29306
rect 32864 29242 32916 29248
rect 33060 29170 33088 29786
rect 33048 29164 33100 29170
rect 33048 29106 33100 29112
rect 32496 29028 32548 29034
rect 32496 28970 32548 28976
rect 32404 27124 32456 27130
rect 32404 27066 32456 27072
rect 32312 26376 32364 26382
rect 32312 26318 32364 26324
rect 32232 26206 32444 26234
rect 32220 25832 32272 25838
rect 32220 25774 32272 25780
rect 32128 24744 32180 24750
rect 32128 24686 32180 24692
rect 32140 24206 32168 24686
rect 32128 24200 32180 24206
rect 32128 24142 32180 24148
rect 32036 23180 32088 23186
rect 32036 23122 32088 23128
rect 32048 22234 32076 23122
rect 32036 22228 32088 22234
rect 32036 22170 32088 22176
rect 31956 22066 32076 22094
rect 31852 21412 31904 21418
rect 31852 21354 31904 21360
rect 31850 20496 31906 20505
rect 31850 20431 31852 20440
rect 31904 20431 31906 20440
rect 31852 20402 31904 20408
rect 31588 20352 31800 20380
rect 31588 19666 31616 20352
rect 31760 20256 31812 20262
rect 31760 20198 31812 20204
rect 31588 19638 31708 19666
rect 31574 19544 31630 19553
rect 31574 19479 31576 19488
rect 31628 19479 31630 19488
rect 31576 19450 31628 19456
rect 31576 19372 31628 19378
rect 31576 19314 31628 19320
rect 31484 17876 31536 17882
rect 31484 17818 31536 17824
rect 31484 17536 31536 17542
rect 31484 17478 31536 17484
rect 31496 17202 31524 17478
rect 31300 17196 31352 17202
rect 31300 17138 31352 17144
rect 31484 17196 31536 17202
rect 31484 17138 31536 17144
rect 31024 16788 31076 16794
rect 31024 16730 31076 16736
rect 30760 12406 30880 12434
rect 30472 6112 30524 6118
rect 30472 6054 30524 6060
rect 29828 5228 29880 5234
rect 29828 5170 29880 5176
rect 30380 5092 30432 5098
rect 30380 5034 30432 5040
rect 29828 5024 29880 5030
rect 29828 4966 29880 4972
rect 29840 4690 29868 4966
rect 29828 4684 29880 4690
rect 29828 4626 29880 4632
rect 29736 4140 29788 4146
rect 29736 4082 29788 4088
rect 30392 4010 30420 5034
rect 30380 4004 30432 4010
rect 30380 3946 30432 3952
rect 29644 3936 29696 3942
rect 29644 3878 29696 3884
rect 29512 3476 29592 3482
rect 29460 3470 29592 3476
rect 29000 3460 29052 3466
rect 29472 3454 29592 3470
rect 29000 3402 29052 3408
rect 29012 3194 29040 3402
rect 29000 3188 29052 3194
rect 29000 3130 29052 3136
rect 28828 2746 28948 2774
rect 29110 2748 29418 2768
rect 29110 2746 29116 2748
rect 29172 2746 29196 2748
rect 29252 2746 29276 2748
rect 29332 2746 29356 2748
rect 29412 2746 29418 2748
rect 28828 2446 28856 2746
rect 29172 2694 29174 2746
rect 29354 2694 29356 2746
rect 29110 2692 29116 2694
rect 29172 2692 29196 2694
rect 29252 2692 29276 2694
rect 29332 2692 29356 2694
rect 29412 2692 29418 2694
rect 29110 2672 29418 2692
rect 29564 2514 29592 3454
rect 29656 3058 29684 3878
rect 30196 3664 30248 3670
rect 30196 3606 30248 3612
rect 29644 3052 29696 3058
rect 29644 2994 29696 3000
rect 29920 2848 29972 2854
rect 29920 2790 29972 2796
rect 29932 2514 29960 2790
rect 30208 2514 30236 3606
rect 30288 2984 30340 2990
rect 30288 2926 30340 2932
rect 29552 2508 29604 2514
rect 29552 2450 29604 2456
rect 29920 2508 29972 2514
rect 29920 2450 29972 2456
rect 30196 2508 30248 2514
rect 30196 2450 30248 2456
rect 28816 2440 28868 2446
rect 28816 2382 28868 2388
rect 30300 800 30328 2926
rect 30484 2582 30512 6054
rect 30760 4078 30788 12406
rect 31588 10266 31616 19314
rect 31680 18222 31708 19638
rect 31772 19378 31800 20198
rect 31864 19938 31892 20402
rect 31864 19910 31984 19938
rect 31852 19848 31904 19854
rect 31852 19790 31904 19796
rect 31760 19372 31812 19378
rect 31760 19314 31812 19320
rect 31668 18216 31720 18222
rect 31668 18158 31720 18164
rect 31864 17202 31892 19790
rect 31956 19174 31984 19910
rect 32048 19258 32076 22066
rect 32140 21690 32168 24142
rect 32232 22273 32260 25774
rect 32312 25696 32364 25702
rect 32312 25638 32364 25644
rect 32324 25226 32352 25638
rect 32312 25220 32364 25226
rect 32312 25162 32364 25168
rect 32324 24614 32352 25162
rect 32312 24608 32364 24614
rect 32312 24550 32364 24556
rect 32416 23905 32444 26206
rect 32508 24410 32536 28970
rect 32956 28620 33008 28626
rect 32956 28562 33008 28568
rect 32588 28552 32640 28558
rect 32588 28494 32640 28500
rect 32600 26926 32628 28494
rect 32772 28416 32824 28422
rect 32772 28358 32824 28364
rect 32680 27056 32732 27062
rect 32680 26998 32732 27004
rect 32588 26920 32640 26926
rect 32588 26862 32640 26868
rect 32496 24404 32548 24410
rect 32496 24346 32548 24352
rect 32402 23896 32458 23905
rect 32402 23831 32458 23840
rect 32508 23746 32536 24346
rect 32416 23718 32536 23746
rect 32312 23656 32364 23662
rect 32312 23598 32364 23604
rect 32218 22264 32274 22273
rect 32218 22199 32274 22208
rect 32218 22128 32274 22137
rect 32218 22063 32274 22072
rect 32128 21684 32180 21690
rect 32128 21626 32180 21632
rect 32128 19984 32180 19990
rect 32128 19926 32180 19932
rect 32140 19514 32168 19926
rect 32128 19508 32180 19514
rect 32128 19450 32180 19456
rect 32048 19230 32168 19258
rect 31944 19168 31996 19174
rect 31944 19110 31996 19116
rect 31944 17672 31996 17678
rect 31944 17614 31996 17620
rect 31852 17196 31904 17202
rect 31852 17138 31904 17144
rect 31668 16992 31720 16998
rect 31668 16934 31720 16940
rect 31680 16658 31708 16934
rect 31668 16652 31720 16658
rect 31668 16594 31720 16600
rect 31956 16114 31984 17614
rect 32036 17128 32088 17134
rect 32036 17070 32088 17076
rect 31944 16108 31996 16114
rect 31944 16050 31996 16056
rect 32048 16046 32076 17070
rect 32140 16454 32168 19230
rect 32128 16448 32180 16454
rect 32128 16390 32180 16396
rect 32036 16040 32088 16046
rect 32036 15982 32088 15988
rect 32232 12434 32260 22063
rect 32324 21146 32352 23598
rect 32416 22953 32444 23718
rect 32496 23656 32548 23662
rect 32496 23598 32548 23604
rect 32402 22944 32458 22953
rect 32402 22879 32458 22888
rect 32402 22808 32458 22817
rect 32402 22743 32458 22752
rect 32416 22030 32444 22743
rect 32404 22024 32456 22030
rect 32404 21966 32456 21972
rect 32402 21856 32458 21865
rect 32402 21791 32458 21800
rect 32312 21140 32364 21146
rect 32312 21082 32364 21088
rect 32312 18760 32364 18766
rect 32312 18702 32364 18708
rect 32324 17270 32352 18702
rect 32416 17542 32444 21791
rect 32508 21690 32536 23598
rect 32496 21684 32548 21690
rect 32496 21626 32548 21632
rect 32600 18426 32628 26862
rect 32692 22545 32720 26998
rect 32784 26994 32812 28358
rect 32864 27872 32916 27878
rect 32864 27814 32916 27820
rect 32772 26988 32824 26994
rect 32772 26930 32824 26936
rect 32772 26308 32824 26314
rect 32772 26250 32824 26256
rect 32784 22642 32812 26250
rect 32772 22636 32824 22642
rect 32772 22578 32824 22584
rect 32678 22536 32734 22545
rect 32678 22471 32734 22480
rect 32772 22500 32824 22506
rect 32772 22442 32824 22448
rect 32680 22432 32732 22438
rect 32680 22374 32732 22380
rect 32588 18420 32640 18426
rect 32588 18362 32640 18368
rect 32692 18290 32720 22374
rect 32496 18284 32548 18290
rect 32496 18226 32548 18232
rect 32680 18284 32732 18290
rect 32680 18226 32732 18232
rect 32508 17746 32536 18226
rect 32496 17740 32548 17746
rect 32496 17682 32548 17688
rect 32404 17536 32456 17542
rect 32404 17478 32456 17484
rect 32312 17264 32364 17270
rect 32312 17206 32364 17212
rect 32312 16788 32364 16794
rect 32312 16730 32364 16736
rect 32324 16114 32352 16730
rect 32416 16590 32444 17478
rect 32404 16584 32456 16590
rect 32404 16526 32456 16532
rect 32312 16108 32364 16114
rect 32312 16050 32364 16056
rect 32312 14816 32364 14822
rect 32312 14758 32364 14764
rect 32324 14482 32352 14758
rect 32312 14476 32364 14482
rect 32312 14418 32364 14424
rect 32312 13320 32364 13326
rect 32312 13262 32364 13268
rect 32324 12850 32352 13262
rect 32496 13184 32548 13190
rect 32496 13126 32548 13132
rect 32508 12918 32536 13126
rect 32496 12912 32548 12918
rect 32496 12854 32548 12860
rect 32312 12844 32364 12850
rect 32312 12786 32364 12792
rect 32140 12406 32260 12434
rect 31576 10260 31628 10266
rect 31576 10202 31628 10208
rect 32140 10062 32168 12406
rect 32784 11830 32812 22442
rect 32876 22438 32904 27814
rect 32968 27130 32996 28562
rect 32956 27124 33008 27130
rect 32956 27066 33008 27072
rect 32968 26314 32996 27066
rect 32956 26308 33008 26314
rect 32956 26250 33008 26256
rect 32954 25392 33010 25401
rect 32954 25327 33010 25336
rect 32968 22642 32996 25327
rect 33060 24154 33088 29106
rect 33152 27402 33180 29990
rect 33244 28694 33272 33798
rect 33324 32904 33376 32910
rect 33324 32846 33376 32852
rect 33336 29306 33364 32846
rect 33428 31958 33456 34546
rect 33416 31952 33468 31958
rect 33416 31894 33468 31900
rect 33520 30802 33548 35158
rect 34152 35012 34204 35018
rect 34152 34954 34204 34960
rect 34164 34785 34192 34954
rect 34150 34776 34206 34785
rect 34150 34711 34206 34720
rect 33692 34604 33744 34610
rect 33692 34546 33744 34552
rect 33704 33454 33732 34546
rect 34150 34096 34206 34105
rect 34150 34031 34152 34040
rect 34204 34031 34206 34040
rect 34152 34002 34204 34008
rect 33692 33448 33744 33454
rect 34152 33448 34204 33454
rect 33692 33390 33744 33396
rect 34150 33416 34152 33425
rect 34204 33416 34206 33425
rect 34150 33351 34206 33360
rect 34150 32736 34206 32745
rect 34150 32671 34206 32680
rect 34164 32502 34192 32671
rect 34152 32496 34204 32502
rect 34152 32438 34204 32444
rect 33784 32292 33836 32298
rect 33784 32234 33836 32240
rect 33508 30796 33560 30802
rect 33508 30738 33560 30744
rect 33796 30258 33824 32234
rect 34150 32056 34206 32065
rect 34150 31991 34206 32000
rect 34164 31890 34192 31991
rect 34152 31884 34204 31890
rect 34152 31826 34204 31832
rect 34150 31376 34206 31385
rect 34150 31311 34152 31320
rect 34204 31311 34206 31320
rect 34152 31282 34204 31288
rect 34060 31272 34112 31278
rect 34060 31214 34112 31220
rect 33874 30968 33930 30977
rect 33874 30903 33930 30912
rect 33888 30734 33916 30903
rect 33876 30728 33928 30734
rect 33876 30670 33928 30676
rect 33968 30728 34020 30734
rect 33968 30670 34020 30676
rect 33876 30320 33928 30326
rect 33876 30262 33928 30268
rect 33784 30252 33836 30258
rect 33784 30194 33836 30200
rect 33506 30152 33562 30161
rect 33506 30087 33562 30096
rect 33416 30048 33468 30054
rect 33416 29990 33468 29996
rect 33324 29300 33376 29306
rect 33324 29242 33376 29248
rect 33232 28688 33284 28694
rect 33232 28630 33284 28636
rect 33324 28552 33376 28558
rect 33324 28494 33376 28500
rect 33140 27396 33192 27402
rect 33140 27338 33192 27344
rect 33336 27130 33364 28494
rect 33324 27124 33376 27130
rect 33324 27066 33376 27072
rect 33428 26897 33456 29990
rect 33520 29170 33548 30087
rect 33692 29504 33744 29510
rect 33692 29446 33744 29452
rect 33600 29232 33652 29238
rect 33600 29174 33652 29180
rect 33508 29164 33560 29170
rect 33508 29106 33560 29112
rect 33508 28416 33560 28422
rect 33508 28358 33560 28364
rect 33414 26888 33470 26897
rect 33414 26823 33470 26832
rect 33140 26784 33192 26790
rect 33520 26738 33548 28358
rect 33612 27334 33640 29174
rect 33704 28490 33732 29446
rect 33796 28558 33824 30194
rect 33888 29170 33916 30262
rect 33876 29164 33928 29170
rect 33876 29106 33928 29112
rect 33784 28552 33836 28558
rect 33784 28494 33836 28500
rect 33692 28484 33744 28490
rect 33692 28426 33744 28432
rect 33600 27328 33652 27334
rect 33600 27270 33652 27276
rect 33600 26988 33652 26994
rect 33704 26976 33732 28426
rect 33796 27674 33824 28494
rect 33784 27668 33836 27674
rect 33784 27610 33836 27616
rect 33652 26948 33732 26976
rect 33600 26930 33652 26936
rect 33140 26726 33192 26732
rect 33152 24274 33180 26726
rect 33336 26710 33548 26738
rect 33140 24268 33192 24274
rect 33140 24210 33192 24216
rect 33060 24126 33180 24154
rect 33048 24064 33100 24070
rect 33048 24006 33100 24012
rect 33060 22681 33088 24006
rect 33046 22672 33102 22681
rect 32956 22636 33008 22642
rect 33046 22607 33102 22616
rect 32956 22578 33008 22584
rect 32864 22432 32916 22438
rect 32864 22374 32916 22380
rect 32968 22234 32996 22578
rect 33152 22488 33180 24126
rect 33336 23644 33364 26710
rect 33612 26602 33640 26930
rect 33796 26926 33824 27610
rect 33784 26920 33836 26926
rect 33784 26862 33836 26868
rect 33060 22460 33180 22488
rect 33244 23616 33364 23644
rect 33428 26574 33640 26602
rect 32956 22228 33008 22234
rect 32956 22170 33008 22176
rect 32862 22128 32918 22137
rect 33060 22094 33088 22460
rect 33138 22400 33194 22409
rect 33138 22335 33194 22344
rect 32862 22063 32864 22072
rect 32916 22063 32918 22072
rect 32968 22066 33088 22094
rect 32864 22034 32916 22040
rect 32864 21956 32916 21962
rect 32864 21898 32916 21904
rect 32876 16658 32904 21898
rect 32968 18358 32996 22066
rect 33152 22012 33180 22335
rect 33060 21984 33180 22012
rect 33060 21010 33088 21984
rect 33244 21622 33272 23616
rect 33324 23180 33376 23186
rect 33324 23122 33376 23128
rect 33336 22574 33364 23122
rect 33324 22568 33376 22574
rect 33324 22510 33376 22516
rect 33324 22228 33376 22234
rect 33324 22170 33376 22176
rect 33336 21962 33364 22170
rect 33324 21956 33376 21962
rect 33324 21898 33376 21904
rect 33232 21616 33284 21622
rect 33232 21558 33284 21564
rect 33048 21004 33100 21010
rect 33048 20946 33100 20952
rect 33140 20936 33192 20942
rect 33140 20878 33192 20884
rect 33152 19360 33180 20878
rect 33324 20800 33376 20806
rect 33324 20742 33376 20748
rect 33336 20534 33364 20742
rect 33324 20528 33376 20534
rect 33324 20470 33376 20476
rect 33232 19780 33284 19786
rect 33232 19722 33284 19728
rect 33244 19514 33272 19722
rect 33428 19514 33456 26574
rect 33888 26466 33916 29106
rect 33612 26438 33916 26466
rect 33508 24812 33560 24818
rect 33508 24754 33560 24760
rect 33520 23633 33548 24754
rect 33506 23624 33562 23633
rect 33506 23559 33562 23568
rect 33232 19508 33284 19514
rect 33232 19450 33284 19456
rect 33416 19508 33468 19514
rect 33416 19450 33468 19456
rect 33152 19332 33272 19360
rect 32956 18352 33008 18358
rect 32956 18294 33008 18300
rect 33140 17128 33192 17134
rect 33140 17070 33192 17076
rect 32956 17060 33008 17066
rect 32956 17002 33008 17008
rect 32968 16658 32996 17002
rect 32864 16652 32916 16658
rect 32864 16594 32916 16600
rect 32956 16652 33008 16658
rect 32956 16594 33008 16600
rect 32968 15026 32996 16594
rect 33152 16590 33180 17070
rect 33140 16584 33192 16590
rect 33140 16526 33192 16532
rect 32956 15020 33008 15026
rect 32956 14962 33008 14968
rect 33140 14816 33192 14822
rect 33140 14758 33192 14764
rect 33152 14482 33180 14758
rect 33140 14476 33192 14482
rect 33140 14418 33192 14424
rect 33140 13320 33192 13326
rect 33140 13262 33192 13268
rect 33152 12306 33180 13262
rect 33140 12300 33192 12306
rect 33140 12242 33192 12248
rect 32772 11824 32824 11830
rect 32772 11766 32824 11772
rect 32680 11688 32732 11694
rect 32680 11630 32732 11636
rect 32128 10056 32180 10062
rect 32128 9998 32180 10004
rect 32588 7880 32640 7886
rect 32588 7822 32640 7828
rect 31668 6792 31720 6798
rect 31668 6734 31720 6740
rect 31680 5778 31708 6734
rect 32496 6112 32548 6118
rect 32496 6054 32548 6060
rect 32312 5908 32364 5914
rect 32312 5850 32364 5856
rect 31668 5772 31720 5778
rect 31668 5714 31720 5720
rect 31484 5704 31536 5710
rect 31484 5646 31536 5652
rect 31392 5228 31444 5234
rect 31392 5170 31444 5176
rect 31404 5098 31432 5170
rect 31392 5092 31444 5098
rect 31392 5034 31444 5040
rect 30840 5024 30892 5030
rect 30840 4966 30892 4972
rect 30748 4072 30800 4078
rect 30748 4014 30800 4020
rect 30656 3460 30708 3466
rect 30656 3402 30708 3408
rect 30668 3194 30696 3402
rect 30656 3188 30708 3194
rect 30656 3130 30708 3136
rect 30472 2576 30524 2582
rect 30472 2518 30524 2524
rect 30852 2378 30880 4966
rect 30932 4684 30984 4690
rect 30932 4626 30984 4632
rect 30840 2372 30892 2378
rect 30840 2314 30892 2320
rect 30944 800 30972 4626
rect 31496 4146 31524 5646
rect 31852 5636 31904 5642
rect 31852 5578 31904 5584
rect 31484 4140 31536 4146
rect 31484 4082 31536 4088
rect 31864 2650 31892 5578
rect 32220 5160 32272 5166
rect 32220 5102 32272 5108
rect 32036 4072 32088 4078
rect 32036 4014 32088 4020
rect 31852 2644 31904 2650
rect 31852 2586 31904 2592
rect 32048 2145 32076 4014
rect 32232 3534 32260 5102
rect 32324 4690 32352 5850
rect 32312 4684 32364 4690
rect 32312 4626 32364 4632
rect 32312 4072 32364 4078
rect 32312 4014 32364 4020
rect 32324 3738 32352 4014
rect 32312 3732 32364 3738
rect 32312 3674 32364 3680
rect 32220 3528 32272 3534
rect 32220 3470 32272 3476
rect 32508 2990 32536 6054
rect 32600 5166 32628 7822
rect 32588 5160 32640 5166
rect 32588 5102 32640 5108
rect 32496 2984 32548 2990
rect 32496 2926 32548 2932
rect 32220 2848 32272 2854
rect 32220 2790 32272 2796
rect 32034 2136 32090 2145
rect 32034 2071 32090 2080
rect 32232 800 32260 2790
rect -10 0 102 800
rect 634 0 746 800
rect 1278 0 1390 800
rect 1922 0 2034 800
rect 2566 0 2678 800
rect 3210 0 3322 800
rect 3854 0 3966 800
rect 4498 0 4610 800
rect 5142 0 5254 800
rect 6430 0 6542 800
rect 7074 0 7186 800
rect 7718 0 7830 800
rect 8362 0 8474 800
rect 9006 0 9118 800
rect 9650 0 9762 800
rect 10294 0 10406 800
rect 10938 0 11050 800
rect 11582 0 11694 800
rect 12870 0 12982 800
rect 13514 0 13626 800
rect 14158 0 14270 800
rect 14802 0 14914 800
rect 15446 0 15558 800
rect 16090 0 16202 800
rect 16734 0 16846 800
rect 17378 0 17490 800
rect 18022 0 18134 800
rect 19310 0 19422 800
rect 19954 0 20066 800
rect 20598 0 20710 800
rect 21242 0 21354 800
rect 21886 0 21998 800
rect 22530 0 22642 800
rect 23174 0 23286 800
rect 23818 0 23930 800
rect 24462 0 24574 800
rect 25750 0 25862 800
rect 26394 0 26506 800
rect 27038 0 27150 800
rect 27682 0 27794 800
rect 28326 0 28438 800
rect 28970 0 29082 800
rect 29614 0 29726 800
rect 30258 0 30370 800
rect 30902 0 31014 800
rect 32190 0 32302 800
rect 32586 96 32642 105
rect 32692 82 32720 11630
rect 32956 6316 33008 6322
rect 32956 6258 33008 6264
rect 32968 5370 32996 6258
rect 33048 6112 33100 6118
rect 33048 6054 33100 6060
rect 32956 5364 33008 5370
rect 32956 5306 33008 5312
rect 33060 4690 33088 6054
rect 33140 5772 33192 5778
rect 33140 5714 33192 5720
rect 33048 4684 33100 4690
rect 33048 4626 33100 4632
rect 33048 4072 33100 4078
rect 33048 4014 33100 4020
rect 33060 3505 33088 4014
rect 33046 3496 33102 3505
rect 33046 3431 33102 3440
rect 33152 2854 33180 5714
rect 33244 2922 33272 19332
rect 33416 16992 33468 16998
rect 33416 16934 33468 16940
rect 33428 16658 33456 16934
rect 33416 16652 33468 16658
rect 33416 16594 33468 16600
rect 33428 13326 33456 16594
rect 33416 13320 33468 13326
rect 33416 13262 33468 13268
rect 33520 12434 33548 23559
rect 33612 22030 33640 26438
rect 33980 26042 34008 30670
rect 34072 29306 34100 31214
rect 34244 30796 34296 30802
rect 34244 30738 34296 30744
rect 34152 29640 34204 29646
rect 34152 29582 34204 29588
rect 34060 29300 34112 29306
rect 34060 29242 34112 29248
rect 34164 28994 34192 29582
rect 34072 28966 34192 28994
rect 33968 26036 34020 26042
rect 33968 25978 34020 25984
rect 34072 25922 34100 28966
rect 34152 28008 34204 28014
rect 34150 27976 34152 27985
rect 34204 27976 34206 27985
rect 34150 27911 34206 27920
rect 33888 25894 34100 25922
rect 34150 25936 34206 25945
rect 33692 23044 33744 23050
rect 33692 22986 33744 22992
rect 33704 22098 33732 22986
rect 33888 22642 33916 25894
rect 34150 25871 34152 25880
rect 34204 25871 34206 25880
rect 34152 25842 34204 25848
rect 34060 25832 34112 25838
rect 34060 25774 34112 25780
rect 33968 25220 34020 25226
rect 33968 25162 34020 25168
rect 33876 22636 33928 22642
rect 33876 22578 33928 22584
rect 33692 22092 33744 22098
rect 33888 22094 33916 22578
rect 33692 22034 33744 22040
rect 33796 22066 33916 22094
rect 33600 22024 33652 22030
rect 33600 21966 33652 21972
rect 33796 21554 33824 22066
rect 33980 21690 34008 25162
rect 34072 24818 34100 25774
rect 34152 25288 34204 25294
rect 34150 25256 34152 25265
rect 34204 25256 34206 25265
rect 34150 25191 34206 25200
rect 34060 24812 34112 24818
rect 34060 24754 34112 24760
rect 34060 24676 34112 24682
rect 34060 24618 34112 24624
rect 33968 21684 34020 21690
rect 33968 21626 34020 21632
rect 33784 21548 33836 21554
rect 33784 21490 33836 21496
rect 33876 21548 33928 21554
rect 33876 21490 33928 21496
rect 33692 18692 33744 18698
rect 33692 18634 33744 18640
rect 33704 18426 33732 18634
rect 33692 18420 33744 18426
rect 33692 18362 33744 18368
rect 33600 18284 33652 18290
rect 33600 18226 33652 18232
rect 33612 15586 33640 18226
rect 33784 17604 33836 17610
rect 33784 17546 33836 17552
rect 33796 16590 33824 17546
rect 33784 16584 33836 16590
rect 33784 16526 33836 16532
rect 33692 16040 33744 16046
rect 33692 15982 33744 15988
rect 33704 15706 33732 15982
rect 33692 15700 33744 15706
rect 33692 15642 33744 15648
rect 33612 15558 33732 15586
rect 33600 15496 33652 15502
rect 33600 15438 33652 15444
rect 33428 12406 33548 12434
rect 33324 9920 33376 9926
rect 33324 9862 33376 9868
rect 33336 9654 33364 9862
rect 33324 9648 33376 9654
rect 33324 9590 33376 9596
rect 33428 6322 33456 12406
rect 33612 11150 33640 15438
rect 33704 12434 33732 15558
rect 33784 14816 33836 14822
rect 33784 14758 33836 14764
rect 33796 14006 33824 14758
rect 33784 14000 33836 14006
rect 33784 13942 33836 13948
rect 33704 12406 33824 12434
rect 33692 12164 33744 12170
rect 33692 12106 33744 12112
rect 33704 11354 33732 12106
rect 33692 11348 33744 11354
rect 33692 11290 33744 11296
rect 33600 11144 33652 11150
rect 33600 11086 33652 11092
rect 33416 6316 33468 6322
rect 33416 6258 33468 6264
rect 33232 2916 33284 2922
rect 33232 2858 33284 2864
rect 33140 2848 33192 2854
rect 33140 2790 33192 2796
rect 32864 2508 32916 2514
rect 32864 2450 32916 2456
rect 32876 800 32904 2450
rect 33612 2310 33640 11086
rect 33692 6724 33744 6730
rect 33692 6666 33744 6672
rect 33704 6458 33732 6666
rect 33692 6452 33744 6458
rect 33692 6394 33744 6400
rect 33796 3466 33824 12406
rect 33888 5098 33916 21490
rect 34072 19378 34100 24618
rect 34150 24576 34206 24585
rect 34150 24511 34206 24520
rect 34164 24274 34192 24511
rect 34152 24268 34204 24274
rect 34152 24210 34204 24216
rect 34150 23896 34206 23905
rect 34150 23831 34206 23840
rect 34164 23798 34192 23831
rect 34152 23792 34204 23798
rect 34152 23734 34204 23740
rect 34150 23216 34206 23225
rect 34150 23151 34152 23160
rect 34204 23151 34206 23160
rect 34152 23122 34204 23128
rect 34150 20496 34206 20505
rect 34150 20431 34152 20440
rect 34204 20431 34206 20440
rect 34152 20402 34204 20408
rect 34150 19816 34206 19825
rect 34150 19751 34152 19760
rect 34204 19751 34206 19760
rect 34152 19722 34204 19728
rect 34060 19372 34112 19378
rect 34060 19314 34112 19320
rect 34150 19136 34206 19145
rect 34150 19071 34206 19080
rect 34164 18834 34192 19071
rect 34256 18902 34284 30738
rect 34348 20874 34376 36518
rect 34520 25356 34572 25362
rect 34520 25298 34572 25304
rect 34428 24132 34480 24138
rect 34428 24074 34480 24080
rect 34336 20868 34388 20874
rect 34336 20810 34388 20816
rect 34244 18896 34296 18902
rect 34244 18838 34296 18844
rect 34152 18828 34204 18834
rect 34152 18770 34204 18776
rect 34150 17776 34206 17785
rect 34150 17711 34152 17720
rect 34204 17711 34206 17720
rect 34152 17682 34204 17688
rect 34152 17128 34204 17134
rect 34150 17096 34152 17105
rect 34204 17096 34206 17105
rect 34150 17031 34206 17040
rect 34150 16416 34206 16425
rect 34150 16351 34206 16360
rect 34164 16182 34192 16351
rect 34152 16176 34204 16182
rect 34152 16118 34204 16124
rect 34440 15638 34468 24074
rect 34532 16726 34560 25298
rect 34520 16720 34572 16726
rect 34520 16662 34572 16668
rect 34428 15632 34480 15638
rect 34428 15574 34480 15580
rect 34150 14376 34206 14385
rect 34150 14311 34152 14320
rect 34204 14311 34206 14320
rect 34152 14282 34204 14288
rect 34152 13864 34204 13870
rect 34152 13806 34204 13812
rect 34164 13705 34192 13806
rect 34150 13696 34206 13705
rect 34150 13631 34206 13640
rect 34150 13016 34206 13025
rect 34150 12951 34206 12960
rect 34164 12918 34192 12951
rect 34152 12912 34204 12918
rect 34152 12854 34204 12860
rect 34150 12336 34206 12345
rect 34150 12271 34152 12280
rect 34204 12271 34206 12280
rect 34152 12242 34204 12248
rect 33968 11620 34020 11626
rect 33968 11562 34020 11568
rect 33980 10674 34008 11562
rect 33968 10668 34020 10674
rect 33968 10610 34020 10616
rect 33968 9988 34020 9994
rect 33968 9930 34020 9936
rect 33980 9625 34008 9930
rect 33966 9616 34022 9625
rect 33966 9551 34022 9560
rect 33968 9512 34020 9518
rect 33968 9454 34020 9460
rect 34152 9512 34204 9518
rect 34152 9454 34204 9460
rect 33980 9178 34008 9454
rect 33968 9172 34020 9178
rect 33968 9114 34020 9120
rect 34164 8945 34192 9454
rect 34150 8936 34206 8945
rect 34150 8871 34206 8880
rect 33968 7200 34020 7206
rect 33968 7142 34020 7148
rect 33980 6866 34008 7142
rect 34150 6896 34206 6905
rect 33968 6860 34020 6866
rect 34150 6831 34152 6840
rect 33968 6802 34020 6808
rect 34204 6831 34206 6840
rect 34152 6802 34204 6808
rect 34060 5568 34112 5574
rect 34060 5510 34112 5516
rect 33876 5092 33928 5098
rect 33876 5034 33928 5040
rect 33784 3460 33836 3466
rect 33784 3402 33836 3408
rect 34072 3126 34100 5510
rect 34152 5160 34204 5166
rect 34152 5102 34204 5108
rect 34164 4865 34192 5102
rect 34150 4856 34206 4865
rect 34150 4791 34206 4800
rect 34152 4548 34204 4554
rect 34152 4490 34204 4496
rect 34164 4185 34192 4490
rect 34150 4176 34206 4185
rect 34150 4111 34206 4120
rect 35440 3596 35492 3602
rect 35440 3538 35492 3544
rect 34060 3120 34112 3126
rect 34060 3062 34112 3068
rect 34796 2984 34848 2990
rect 34796 2926 34848 2932
rect 34428 2372 34480 2378
rect 34428 2314 34480 2320
rect 33600 2304 33652 2310
rect 33600 2246 33652 2252
rect 32642 54 32720 82
rect 32586 31 32642 40
rect 32834 0 32946 800
rect 33478 0 33590 800
rect 34122 0 34234 800
rect 34440 785 34468 2314
rect 34808 800 34836 2926
rect 35452 800 35480 3538
rect 34426 776 34482 785
rect 34426 711 34482 720
rect 34766 0 34878 800
rect 35410 0 35522 800
<< via2 >>
rect 2962 41520 3018 41576
rect 1398 38800 1454 38856
rect 4158 40840 4214 40896
rect 2778 36760 2834 36816
rect 1398 36080 1454 36136
rect 1950 31320 2006 31376
rect 1858 25200 1914 25256
rect 1950 17076 1952 17096
rect 1952 17076 2004 17096
rect 2004 17076 2006 17096
rect 1950 17040 2006 17076
rect 1950 14320 2006 14376
rect 1858 10920 1914 10976
rect 2226 19080 2282 19136
rect 1858 5480 1914 5536
rect 2778 35400 2834 35456
rect 2778 34060 2834 34096
rect 2778 34040 2780 34060
rect 2780 34040 2832 34060
rect 2832 34040 2834 34060
rect 2870 18400 2926 18456
rect 2778 15680 2834 15736
rect 3974 37440 4030 37496
rect 3422 32000 3478 32056
rect 3422 24792 3478 24848
rect 2778 13640 2834 13696
rect 2778 11636 2780 11656
rect 2780 11636 2832 11656
rect 2832 11636 2834 11656
rect 2778 11600 2834 11636
rect 2870 8880 2926 8936
rect 2778 8200 2834 8256
rect 2778 7520 2834 7576
rect 3054 4800 3110 4856
rect 2962 4120 3018 4176
rect 2778 2760 2834 2816
rect 3238 3440 3294 3496
rect 6588 39738 6644 39740
rect 6668 39738 6724 39740
rect 6748 39738 6804 39740
rect 6828 39738 6884 39740
rect 6588 39686 6634 39738
rect 6634 39686 6644 39738
rect 6668 39686 6698 39738
rect 6698 39686 6710 39738
rect 6710 39686 6724 39738
rect 6748 39686 6762 39738
rect 6762 39686 6774 39738
rect 6774 39686 6804 39738
rect 6828 39686 6838 39738
rect 6838 39686 6884 39738
rect 6588 39684 6644 39686
rect 6668 39684 6724 39686
rect 6748 39684 6804 39686
rect 6828 39684 6884 39686
rect 6588 38650 6644 38652
rect 6668 38650 6724 38652
rect 6748 38650 6804 38652
rect 6828 38650 6884 38652
rect 6588 38598 6634 38650
rect 6634 38598 6644 38650
rect 6668 38598 6698 38650
rect 6698 38598 6710 38650
rect 6710 38598 6724 38650
rect 6748 38598 6762 38650
rect 6762 38598 6774 38650
rect 6774 38598 6804 38650
rect 6828 38598 6838 38650
rect 6838 38598 6884 38650
rect 6588 38596 6644 38598
rect 6668 38596 6724 38598
rect 6748 38596 6804 38598
rect 6828 38596 6884 38598
rect 6588 37562 6644 37564
rect 6668 37562 6724 37564
rect 6748 37562 6804 37564
rect 6828 37562 6884 37564
rect 6588 37510 6634 37562
rect 6634 37510 6644 37562
rect 6668 37510 6698 37562
rect 6698 37510 6710 37562
rect 6710 37510 6724 37562
rect 6748 37510 6762 37562
rect 6762 37510 6774 37562
rect 6774 37510 6804 37562
rect 6828 37510 6838 37562
rect 6838 37510 6884 37562
rect 6588 37508 6644 37510
rect 6668 37508 6724 37510
rect 6748 37508 6804 37510
rect 6828 37508 6884 37510
rect 11058 40568 11114 40624
rect 9770 40160 9826 40216
rect 9586 39516 9588 39536
rect 9588 39516 9640 39536
rect 9640 39516 9642 39536
rect 9586 39480 9642 39516
rect 6588 36474 6644 36476
rect 6668 36474 6724 36476
rect 6748 36474 6804 36476
rect 6828 36474 6884 36476
rect 6588 36422 6634 36474
rect 6634 36422 6644 36474
rect 6668 36422 6698 36474
rect 6698 36422 6710 36474
rect 6710 36422 6724 36474
rect 6748 36422 6762 36474
rect 6762 36422 6774 36474
rect 6774 36422 6804 36474
rect 6828 36422 6838 36474
rect 6838 36422 6884 36474
rect 6588 36420 6644 36422
rect 6668 36420 6724 36422
rect 6748 36420 6804 36422
rect 6828 36420 6884 36422
rect 6588 35386 6644 35388
rect 6668 35386 6724 35388
rect 6748 35386 6804 35388
rect 6828 35386 6884 35388
rect 6588 35334 6634 35386
rect 6634 35334 6644 35386
rect 6668 35334 6698 35386
rect 6698 35334 6710 35386
rect 6710 35334 6724 35386
rect 6748 35334 6762 35386
rect 6762 35334 6774 35386
rect 6774 35334 6804 35386
rect 6828 35334 6838 35386
rect 6838 35334 6884 35386
rect 6588 35332 6644 35334
rect 6668 35332 6724 35334
rect 6748 35332 6804 35334
rect 6828 35332 6884 35334
rect 6588 34298 6644 34300
rect 6668 34298 6724 34300
rect 6748 34298 6804 34300
rect 6828 34298 6884 34300
rect 6588 34246 6634 34298
rect 6634 34246 6644 34298
rect 6668 34246 6698 34298
rect 6698 34246 6710 34298
rect 6710 34246 6724 34298
rect 6748 34246 6762 34298
rect 6762 34246 6774 34298
rect 6774 34246 6804 34298
rect 6828 34246 6838 34298
rect 6838 34246 6884 34298
rect 6588 34244 6644 34246
rect 6668 34244 6724 34246
rect 6748 34244 6804 34246
rect 6828 34244 6884 34246
rect 6588 33210 6644 33212
rect 6668 33210 6724 33212
rect 6748 33210 6804 33212
rect 6828 33210 6884 33212
rect 6588 33158 6634 33210
rect 6634 33158 6644 33210
rect 6668 33158 6698 33210
rect 6698 33158 6710 33210
rect 6710 33158 6724 33210
rect 6748 33158 6762 33210
rect 6762 33158 6774 33210
rect 6774 33158 6804 33210
rect 6828 33158 6838 33210
rect 6838 33158 6884 33210
rect 6588 33156 6644 33158
rect 6668 33156 6724 33158
rect 6748 33156 6804 33158
rect 6828 33156 6884 33158
rect 6588 32122 6644 32124
rect 6668 32122 6724 32124
rect 6748 32122 6804 32124
rect 6828 32122 6884 32124
rect 6588 32070 6634 32122
rect 6634 32070 6644 32122
rect 6668 32070 6698 32122
rect 6698 32070 6710 32122
rect 6710 32070 6724 32122
rect 6748 32070 6762 32122
rect 6762 32070 6774 32122
rect 6774 32070 6804 32122
rect 6828 32070 6838 32122
rect 6838 32070 6884 32122
rect 6588 32068 6644 32070
rect 6668 32068 6724 32070
rect 6748 32068 6804 32070
rect 6828 32068 6884 32070
rect 6588 31034 6644 31036
rect 6668 31034 6724 31036
rect 6748 31034 6804 31036
rect 6828 31034 6884 31036
rect 6588 30982 6634 31034
rect 6634 30982 6644 31034
rect 6668 30982 6698 31034
rect 6698 30982 6710 31034
rect 6710 30982 6724 31034
rect 6748 30982 6762 31034
rect 6762 30982 6774 31034
rect 6774 30982 6804 31034
rect 6828 30982 6838 31034
rect 6838 30982 6884 31034
rect 6588 30980 6644 30982
rect 6668 30980 6724 30982
rect 6748 30980 6804 30982
rect 6828 30980 6884 30982
rect 6588 29946 6644 29948
rect 6668 29946 6724 29948
rect 6748 29946 6804 29948
rect 6828 29946 6884 29948
rect 6588 29894 6634 29946
rect 6634 29894 6644 29946
rect 6668 29894 6698 29946
rect 6698 29894 6710 29946
rect 6710 29894 6724 29946
rect 6748 29894 6762 29946
rect 6762 29894 6774 29946
rect 6774 29894 6804 29946
rect 6828 29894 6838 29946
rect 6838 29894 6884 29946
rect 6588 29892 6644 29894
rect 6668 29892 6724 29894
rect 6748 29892 6804 29894
rect 6828 29892 6884 29894
rect 6588 28858 6644 28860
rect 6668 28858 6724 28860
rect 6748 28858 6804 28860
rect 6828 28858 6884 28860
rect 6588 28806 6634 28858
rect 6634 28806 6644 28858
rect 6668 28806 6698 28858
rect 6698 28806 6710 28858
rect 6710 28806 6724 28858
rect 6748 28806 6762 28858
rect 6762 28806 6774 28858
rect 6774 28806 6804 28858
rect 6828 28806 6838 28858
rect 6838 28806 6884 28858
rect 6588 28804 6644 28806
rect 6668 28804 6724 28806
rect 6748 28804 6804 28806
rect 6828 28804 6884 28806
rect 6588 27770 6644 27772
rect 6668 27770 6724 27772
rect 6748 27770 6804 27772
rect 6828 27770 6884 27772
rect 6588 27718 6634 27770
rect 6634 27718 6644 27770
rect 6668 27718 6698 27770
rect 6698 27718 6710 27770
rect 6710 27718 6724 27770
rect 6748 27718 6762 27770
rect 6762 27718 6774 27770
rect 6774 27718 6804 27770
rect 6828 27718 6838 27770
rect 6838 27718 6884 27770
rect 6588 27716 6644 27718
rect 6668 27716 6724 27718
rect 6748 27716 6804 27718
rect 6828 27716 6884 27718
rect 6588 26682 6644 26684
rect 6668 26682 6724 26684
rect 6748 26682 6804 26684
rect 6828 26682 6884 26684
rect 6588 26630 6634 26682
rect 6634 26630 6644 26682
rect 6668 26630 6698 26682
rect 6698 26630 6710 26682
rect 6710 26630 6724 26682
rect 6748 26630 6762 26682
rect 6762 26630 6774 26682
rect 6774 26630 6804 26682
rect 6828 26630 6838 26682
rect 6838 26630 6884 26682
rect 6588 26628 6644 26630
rect 6668 26628 6724 26630
rect 6748 26628 6804 26630
rect 6828 26628 6884 26630
rect 9678 37732 9734 37768
rect 9678 37712 9680 37732
rect 9680 37712 9732 37732
rect 9732 37712 9734 37732
rect 10322 39888 10378 39944
rect 10966 39380 10968 39400
rect 10968 39380 11020 39400
rect 11020 39380 11022 39400
rect 10966 39344 11022 39380
rect 10322 38936 10378 38992
rect 10874 38256 10930 38312
rect 10230 37324 10286 37360
rect 10230 37304 10232 37324
rect 10232 37304 10284 37324
rect 10284 37304 10286 37324
rect 10782 37848 10838 37904
rect 13174 40704 13230 40760
rect 12220 39194 12276 39196
rect 12300 39194 12356 39196
rect 12380 39194 12436 39196
rect 12460 39194 12516 39196
rect 12220 39142 12266 39194
rect 12266 39142 12276 39194
rect 12300 39142 12330 39194
rect 12330 39142 12342 39194
rect 12342 39142 12356 39194
rect 12380 39142 12394 39194
rect 12394 39142 12406 39194
rect 12406 39142 12436 39194
rect 12460 39142 12470 39194
rect 12470 39142 12516 39194
rect 12220 39140 12276 39142
rect 12300 39140 12356 39142
rect 12380 39140 12436 39142
rect 12460 39140 12516 39142
rect 12254 38528 12310 38584
rect 12220 38106 12276 38108
rect 12300 38106 12356 38108
rect 12380 38106 12436 38108
rect 12460 38106 12516 38108
rect 12220 38054 12266 38106
rect 12266 38054 12276 38106
rect 12300 38054 12330 38106
rect 12330 38054 12342 38106
rect 12342 38054 12356 38106
rect 12380 38054 12394 38106
rect 12394 38054 12406 38106
rect 12406 38054 12436 38106
rect 12460 38054 12470 38106
rect 12470 38054 12516 38106
rect 12220 38052 12276 38054
rect 12300 38052 12356 38054
rect 12380 38052 12436 38054
rect 12460 38052 12516 38054
rect 11426 37440 11482 37496
rect 12346 37576 12402 37632
rect 12898 38120 12954 38176
rect 11978 37168 12034 37224
rect 12622 37068 12624 37088
rect 12624 37068 12676 37088
rect 12676 37068 12678 37088
rect 12622 37032 12678 37068
rect 12220 37018 12276 37020
rect 12300 37018 12356 37020
rect 12380 37018 12436 37020
rect 12460 37018 12516 37020
rect 12220 36966 12266 37018
rect 12266 36966 12276 37018
rect 12300 36966 12330 37018
rect 12330 36966 12342 37018
rect 12342 36966 12356 37018
rect 12380 36966 12394 37018
rect 12394 36966 12406 37018
rect 12406 36966 12436 37018
rect 12460 36966 12470 37018
rect 12470 36966 12516 37018
rect 12220 36964 12276 36966
rect 12300 36964 12356 36966
rect 12380 36964 12436 36966
rect 12460 36964 12516 36966
rect 12070 36644 12126 36680
rect 12070 36624 12072 36644
rect 12072 36624 12124 36644
rect 12124 36624 12126 36644
rect 11610 36252 11612 36272
rect 11612 36252 11664 36272
rect 11664 36252 11666 36272
rect 11610 36216 11666 36252
rect 12346 36352 12402 36408
rect 12806 36896 12862 36952
rect 12162 36080 12218 36136
rect 12714 35980 12716 36000
rect 12716 35980 12768 36000
rect 12768 35980 12770 36000
rect 12714 35944 12770 35980
rect 12220 35930 12276 35932
rect 12300 35930 12356 35932
rect 12380 35930 12436 35932
rect 12460 35930 12516 35932
rect 12220 35878 12266 35930
rect 12266 35878 12276 35930
rect 12300 35878 12330 35930
rect 12330 35878 12342 35930
rect 12342 35878 12356 35930
rect 12380 35878 12394 35930
rect 12394 35878 12406 35930
rect 12406 35878 12436 35930
rect 12460 35878 12470 35930
rect 12470 35878 12516 35930
rect 12220 35876 12276 35878
rect 12300 35876 12356 35878
rect 12380 35876 12436 35878
rect 12460 35876 12516 35878
rect 12530 35556 12586 35592
rect 12530 35536 12532 35556
rect 12532 35536 12584 35556
rect 12584 35536 12586 35556
rect 12220 34842 12276 34844
rect 12300 34842 12356 34844
rect 12380 34842 12436 34844
rect 12460 34842 12516 34844
rect 12220 34790 12266 34842
rect 12266 34790 12276 34842
rect 12300 34790 12330 34842
rect 12330 34790 12342 34842
rect 12342 34790 12356 34842
rect 12380 34790 12394 34842
rect 12394 34790 12406 34842
rect 12406 34790 12436 34842
rect 12460 34790 12470 34842
rect 12470 34790 12516 34842
rect 12220 34788 12276 34790
rect 12300 34788 12356 34790
rect 12380 34788 12436 34790
rect 12460 34788 12516 34790
rect 12714 34740 12770 34776
rect 12714 34720 12716 34740
rect 12716 34720 12768 34740
rect 12768 34720 12770 34740
rect 13082 38412 13138 38448
rect 13082 38392 13084 38412
rect 13084 38392 13136 38412
rect 13136 38392 13138 38412
rect 13082 37984 13138 38040
rect 14278 40296 14334 40352
rect 14002 40024 14058 40080
rect 13450 39208 13506 39264
rect 13266 39072 13322 39128
rect 13450 38664 13506 38720
rect 13358 38528 13414 38584
rect 13082 36624 13138 36680
rect 13174 36488 13230 36544
rect 13450 36624 13506 36680
rect 13726 37984 13782 38040
rect 13818 36760 13874 36816
rect 13266 35264 13322 35320
rect 13174 34856 13230 34912
rect 13358 34740 13414 34776
rect 13358 34720 13360 34740
rect 13360 34720 13412 34740
rect 13412 34720 13414 34740
rect 12254 34468 12310 34504
rect 12254 34448 12256 34468
rect 12256 34448 12308 34468
rect 12308 34448 12310 34468
rect 11794 32308 11796 32328
rect 11796 32308 11848 32328
rect 11848 32308 11850 32328
rect 11794 32272 11850 32308
rect 12220 33754 12276 33756
rect 12300 33754 12356 33756
rect 12380 33754 12436 33756
rect 12460 33754 12516 33756
rect 12220 33702 12266 33754
rect 12266 33702 12276 33754
rect 12300 33702 12330 33754
rect 12330 33702 12342 33754
rect 12342 33702 12356 33754
rect 12380 33702 12394 33754
rect 12394 33702 12406 33754
rect 12406 33702 12436 33754
rect 12460 33702 12470 33754
rect 12470 33702 12516 33754
rect 12220 33700 12276 33702
rect 12300 33700 12356 33702
rect 12380 33700 12436 33702
rect 12460 33700 12516 33702
rect 12898 34312 12954 34368
rect 12714 34176 12770 34232
rect 12622 33496 12678 33552
rect 13266 34060 13322 34096
rect 13266 34040 13268 34060
rect 13268 34040 13320 34060
rect 13320 34040 13322 34060
rect 13450 33904 13506 33960
rect 12220 32666 12276 32668
rect 12300 32666 12356 32668
rect 12380 32666 12436 32668
rect 12460 32666 12516 32668
rect 12220 32614 12266 32666
rect 12266 32614 12276 32666
rect 12300 32614 12330 32666
rect 12330 32614 12342 32666
rect 12342 32614 12356 32666
rect 12380 32614 12394 32666
rect 12394 32614 12406 32666
rect 12406 32614 12436 32666
rect 12460 32614 12470 32666
rect 12470 32614 12516 32666
rect 12220 32612 12276 32614
rect 12300 32612 12356 32614
rect 12380 32612 12436 32614
rect 12460 32612 12516 32614
rect 12806 33260 12808 33280
rect 12808 33260 12860 33280
rect 12860 33260 12862 33280
rect 12806 33224 12862 33260
rect 12990 32680 13046 32736
rect 12806 32408 12862 32464
rect 12220 31578 12276 31580
rect 12300 31578 12356 31580
rect 12380 31578 12436 31580
rect 12460 31578 12516 31580
rect 12220 31526 12266 31578
rect 12266 31526 12276 31578
rect 12300 31526 12330 31578
rect 12330 31526 12342 31578
rect 12342 31526 12356 31578
rect 12380 31526 12394 31578
rect 12394 31526 12406 31578
rect 12406 31526 12436 31578
rect 12460 31526 12470 31578
rect 12470 31526 12516 31578
rect 12220 31524 12276 31526
rect 12300 31524 12356 31526
rect 12380 31524 12436 31526
rect 12460 31524 12516 31526
rect 12070 31048 12126 31104
rect 12898 31728 12954 31784
rect 12714 31456 12770 31512
rect 12806 30796 12862 30832
rect 12806 30776 12808 30796
rect 12808 30776 12860 30796
rect 12860 30776 12862 30796
rect 13910 35808 13966 35864
rect 14094 39616 14150 39672
rect 14278 37984 14334 38040
rect 14002 35128 14058 35184
rect 13634 33088 13690 33144
rect 13358 32952 13414 33008
rect 13910 33396 13912 33416
rect 13912 33396 13964 33416
rect 13964 33396 13966 33416
rect 13910 33360 13966 33396
rect 13266 32136 13322 32192
rect 13634 31864 13690 31920
rect 13634 31320 13690 31376
rect 13266 30912 13322 30968
rect 13174 30660 13230 30696
rect 13174 30640 13176 30660
rect 13176 30640 13228 30660
rect 13228 30640 13230 30660
rect 12220 30490 12276 30492
rect 12300 30490 12356 30492
rect 12380 30490 12436 30492
rect 12460 30490 12516 30492
rect 12220 30438 12266 30490
rect 12266 30438 12276 30490
rect 12300 30438 12330 30490
rect 12330 30438 12342 30490
rect 12342 30438 12356 30490
rect 12380 30438 12394 30490
rect 12394 30438 12406 30490
rect 12406 30438 12436 30490
rect 12460 30438 12470 30490
rect 12470 30438 12516 30490
rect 12220 30436 12276 30438
rect 12300 30436 12356 30438
rect 12380 30436 12436 30438
rect 12460 30436 12516 30438
rect 12714 29824 12770 29880
rect 12220 29402 12276 29404
rect 12300 29402 12356 29404
rect 12380 29402 12436 29404
rect 12460 29402 12516 29404
rect 12220 29350 12266 29402
rect 12266 29350 12276 29402
rect 12300 29350 12330 29402
rect 12330 29350 12342 29402
rect 12342 29350 12356 29402
rect 12380 29350 12394 29402
rect 12394 29350 12406 29402
rect 12406 29350 12436 29402
rect 12460 29350 12470 29402
rect 12470 29350 12516 29402
rect 12220 29348 12276 29350
rect 12300 29348 12356 29350
rect 12380 29348 12436 29350
rect 12460 29348 12516 29350
rect 11978 28736 12034 28792
rect 12220 28314 12276 28316
rect 12300 28314 12356 28316
rect 12380 28314 12436 28316
rect 12460 28314 12516 28316
rect 12220 28262 12266 28314
rect 12266 28262 12276 28314
rect 12300 28262 12330 28314
rect 12330 28262 12342 28314
rect 12342 28262 12356 28314
rect 12380 28262 12394 28314
rect 12394 28262 12406 28314
rect 12406 28262 12436 28314
rect 12460 28262 12470 28314
rect 12470 28262 12516 28314
rect 12220 28260 12276 28262
rect 12300 28260 12356 28262
rect 12380 28260 12436 28262
rect 12460 28260 12516 28262
rect 12220 27226 12276 27228
rect 12300 27226 12356 27228
rect 12380 27226 12436 27228
rect 12460 27226 12516 27228
rect 12220 27174 12266 27226
rect 12266 27174 12276 27226
rect 12300 27174 12330 27226
rect 12330 27174 12342 27226
rect 12342 27174 12356 27226
rect 12380 27174 12394 27226
rect 12394 27174 12406 27226
rect 12406 27174 12436 27226
rect 12460 27174 12470 27226
rect 12470 27174 12516 27226
rect 12220 27172 12276 27174
rect 12300 27172 12356 27174
rect 12380 27172 12436 27174
rect 12460 27172 12516 27174
rect 6588 25594 6644 25596
rect 6668 25594 6724 25596
rect 6748 25594 6804 25596
rect 6828 25594 6884 25596
rect 6588 25542 6634 25594
rect 6634 25542 6644 25594
rect 6668 25542 6698 25594
rect 6698 25542 6710 25594
rect 6710 25542 6724 25594
rect 6748 25542 6762 25594
rect 6762 25542 6774 25594
rect 6774 25542 6804 25594
rect 6828 25542 6838 25594
rect 6838 25542 6884 25594
rect 6588 25540 6644 25542
rect 6668 25540 6724 25542
rect 6748 25540 6804 25542
rect 6828 25540 6884 25542
rect 6588 24506 6644 24508
rect 6668 24506 6724 24508
rect 6748 24506 6804 24508
rect 6828 24506 6884 24508
rect 6588 24454 6634 24506
rect 6634 24454 6644 24506
rect 6668 24454 6698 24506
rect 6698 24454 6710 24506
rect 6710 24454 6724 24506
rect 6748 24454 6762 24506
rect 6762 24454 6774 24506
rect 6774 24454 6804 24506
rect 6828 24454 6838 24506
rect 6838 24454 6884 24506
rect 6588 24452 6644 24454
rect 6668 24452 6724 24454
rect 6748 24452 6804 24454
rect 6828 24452 6884 24454
rect 6588 23418 6644 23420
rect 6668 23418 6724 23420
rect 6748 23418 6804 23420
rect 6828 23418 6884 23420
rect 6588 23366 6634 23418
rect 6634 23366 6644 23418
rect 6668 23366 6698 23418
rect 6698 23366 6710 23418
rect 6710 23366 6724 23418
rect 6748 23366 6762 23418
rect 6762 23366 6774 23418
rect 6774 23366 6804 23418
rect 6828 23366 6838 23418
rect 6838 23366 6884 23418
rect 6588 23364 6644 23366
rect 6668 23364 6724 23366
rect 6748 23364 6804 23366
rect 6828 23364 6884 23366
rect 6588 22330 6644 22332
rect 6668 22330 6724 22332
rect 6748 22330 6804 22332
rect 6828 22330 6884 22332
rect 6588 22278 6634 22330
rect 6634 22278 6644 22330
rect 6668 22278 6698 22330
rect 6698 22278 6710 22330
rect 6710 22278 6724 22330
rect 6748 22278 6762 22330
rect 6762 22278 6774 22330
rect 6774 22278 6804 22330
rect 6828 22278 6838 22330
rect 6838 22278 6884 22330
rect 6588 22276 6644 22278
rect 6668 22276 6724 22278
rect 6748 22276 6804 22278
rect 6828 22276 6884 22278
rect 6588 21242 6644 21244
rect 6668 21242 6724 21244
rect 6748 21242 6804 21244
rect 6828 21242 6884 21244
rect 6588 21190 6634 21242
rect 6634 21190 6644 21242
rect 6668 21190 6698 21242
rect 6698 21190 6710 21242
rect 6710 21190 6724 21242
rect 6748 21190 6762 21242
rect 6762 21190 6774 21242
rect 6774 21190 6804 21242
rect 6828 21190 6838 21242
rect 6838 21190 6884 21242
rect 6588 21188 6644 21190
rect 6668 21188 6724 21190
rect 6748 21188 6804 21190
rect 6828 21188 6884 21190
rect 6588 20154 6644 20156
rect 6668 20154 6724 20156
rect 6748 20154 6804 20156
rect 6828 20154 6884 20156
rect 6588 20102 6634 20154
rect 6634 20102 6644 20154
rect 6668 20102 6698 20154
rect 6698 20102 6710 20154
rect 6710 20102 6724 20154
rect 6748 20102 6762 20154
rect 6762 20102 6774 20154
rect 6774 20102 6804 20154
rect 6828 20102 6838 20154
rect 6838 20102 6884 20154
rect 6588 20100 6644 20102
rect 6668 20100 6724 20102
rect 6748 20100 6804 20102
rect 6828 20100 6884 20102
rect 6588 19066 6644 19068
rect 6668 19066 6724 19068
rect 6748 19066 6804 19068
rect 6828 19066 6884 19068
rect 6588 19014 6634 19066
rect 6634 19014 6644 19066
rect 6668 19014 6698 19066
rect 6698 19014 6710 19066
rect 6710 19014 6724 19066
rect 6748 19014 6762 19066
rect 6762 19014 6774 19066
rect 6774 19014 6804 19066
rect 6828 19014 6838 19066
rect 6838 19014 6884 19066
rect 6588 19012 6644 19014
rect 6668 19012 6724 19014
rect 6748 19012 6804 19014
rect 6828 19012 6884 19014
rect 6588 17978 6644 17980
rect 6668 17978 6724 17980
rect 6748 17978 6804 17980
rect 6828 17978 6884 17980
rect 6588 17926 6634 17978
rect 6634 17926 6644 17978
rect 6668 17926 6698 17978
rect 6698 17926 6710 17978
rect 6710 17926 6724 17978
rect 6748 17926 6762 17978
rect 6762 17926 6774 17978
rect 6774 17926 6804 17978
rect 6828 17926 6838 17978
rect 6838 17926 6884 17978
rect 6588 17924 6644 17926
rect 6668 17924 6724 17926
rect 6748 17924 6804 17926
rect 6828 17924 6884 17926
rect 6588 16890 6644 16892
rect 6668 16890 6724 16892
rect 6748 16890 6804 16892
rect 6828 16890 6884 16892
rect 6588 16838 6634 16890
rect 6634 16838 6644 16890
rect 6668 16838 6698 16890
rect 6698 16838 6710 16890
rect 6710 16838 6724 16890
rect 6748 16838 6762 16890
rect 6762 16838 6774 16890
rect 6774 16838 6804 16890
rect 6828 16838 6838 16890
rect 6838 16838 6884 16890
rect 6588 16836 6644 16838
rect 6668 16836 6724 16838
rect 6748 16836 6804 16838
rect 6828 16836 6884 16838
rect 6588 15802 6644 15804
rect 6668 15802 6724 15804
rect 6748 15802 6804 15804
rect 6828 15802 6884 15804
rect 6588 15750 6634 15802
rect 6634 15750 6644 15802
rect 6668 15750 6698 15802
rect 6698 15750 6710 15802
rect 6710 15750 6724 15802
rect 6748 15750 6762 15802
rect 6762 15750 6774 15802
rect 6774 15750 6804 15802
rect 6828 15750 6838 15802
rect 6838 15750 6884 15802
rect 6588 15748 6644 15750
rect 6668 15748 6724 15750
rect 6748 15748 6804 15750
rect 6828 15748 6884 15750
rect 6588 14714 6644 14716
rect 6668 14714 6724 14716
rect 6748 14714 6804 14716
rect 6828 14714 6884 14716
rect 6588 14662 6634 14714
rect 6634 14662 6644 14714
rect 6668 14662 6698 14714
rect 6698 14662 6710 14714
rect 6710 14662 6724 14714
rect 6748 14662 6762 14714
rect 6762 14662 6774 14714
rect 6774 14662 6804 14714
rect 6828 14662 6838 14714
rect 6838 14662 6884 14714
rect 6588 14660 6644 14662
rect 6668 14660 6724 14662
rect 6748 14660 6804 14662
rect 6828 14660 6884 14662
rect 6588 13626 6644 13628
rect 6668 13626 6724 13628
rect 6748 13626 6804 13628
rect 6828 13626 6884 13628
rect 6588 13574 6634 13626
rect 6634 13574 6644 13626
rect 6668 13574 6698 13626
rect 6698 13574 6710 13626
rect 6710 13574 6724 13626
rect 6748 13574 6762 13626
rect 6762 13574 6774 13626
rect 6774 13574 6804 13626
rect 6828 13574 6838 13626
rect 6838 13574 6884 13626
rect 6588 13572 6644 13574
rect 6668 13572 6724 13574
rect 6748 13572 6804 13574
rect 6828 13572 6884 13574
rect 6588 12538 6644 12540
rect 6668 12538 6724 12540
rect 6748 12538 6804 12540
rect 6828 12538 6884 12540
rect 6588 12486 6634 12538
rect 6634 12486 6644 12538
rect 6668 12486 6698 12538
rect 6698 12486 6710 12538
rect 6710 12486 6724 12538
rect 6748 12486 6762 12538
rect 6762 12486 6774 12538
rect 6774 12486 6804 12538
rect 6828 12486 6838 12538
rect 6838 12486 6884 12538
rect 6588 12484 6644 12486
rect 6668 12484 6724 12486
rect 6748 12484 6804 12486
rect 6828 12484 6884 12486
rect 6588 11450 6644 11452
rect 6668 11450 6724 11452
rect 6748 11450 6804 11452
rect 6828 11450 6884 11452
rect 6588 11398 6634 11450
rect 6634 11398 6644 11450
rect 6668 11398 6698 11450
rect 6698 11398 6710 11450
rect 6710 11398 6724 11450
rect 6748 11398 6762 11450
rect 6762 11398 6774 11450
rect 6774 11398 6804 11450
rect 6828 11398 6838 11450
rect 6838 11398 6884 11450
rect 6588 11396 6644 11398
rect 6668 11396 6724 11398
rect 6748 11396 6804 11398
rect 6828 11396 6884 11398
rect 6588 10362 6644 10364
rect 6668 10362 6724 10364
rect 6748 10362 6804 10364
rect 6828 10362 6884 10364
rect 6588 10310 6634 10362
rect 6634 10310 6644 10362
rect 6668 10310 6698 10362
rect 6698 10310 6710 10362
rect 6710 10310 6724 10362
rect 6748 10310 6762 10362
rect 6762 10310 6774 10362
rect 6774 10310 6804 10362
rect 6828 10310 6838 10362
rect 6838 10310 6884 10362
rect 6588 10308 6644 10310
rect 6668 10308 6724 10310
rect 6748 10308 6804 10310
rect 6828 10308 6884 10310
rect 6588 9274 6644 9276
rect 6668 9274 6724 9276
rect 6748 9274 6804 9276
rect 6828 9274 6884 9276
rect 6588 9222 6634 9274
rect 6634 9222 6644 9274
rect 6668 9222 6698 9274
rect 6698 9222 6710 9274
rect 6710 9222 6724 9274
rect 6748 9222 6762 9274
rect 6762 9222 6774 9274
rect 6774 9222 6804 9274
rect 6828 9222 6838 9274
rect 6838 9222 6884 9274
rect 6588 9220 6644 9222
rect 6668 9220 6724 9222
rect 6748 9220 6804 9222
rect 6828 9220 6884 9222
rect 6588 8186 6644 8188
rect 6668 8186 6724 8188
rect 6748 8186 6804 8188
rect 6828 8186 6884 8188
rect 6588 8134 6634 8186
rect 6634 8134 6644 8186
rect 6668 8134 6698 8186
rect 6698 8134 6710 8186
rect 6710 8134 6724 8186
rect 6748 8134 6762 8186
rect 6762 8134 6774 8186
rect 6774 8134 6804 8186
rect 6828 8134 6838 8186
rect 6838 8134 6884 8186
rect 6588 8132 6644 8134
rect 6668 8132 6724 8134
rect 6748 8132 6804 8134
rect 6828 8132 6884 8134
rect 6588 7098 6644 7100
rect 6668 7098 6724 7100
rect 6748 7098 6804 7100
rect 6828 7098 6884 7100
rect 6588 7046 6634 7098
rect 6634 7046 6644 7098
rect 6668 7046 6698 7098
rect 6698 7046 6710 7098
rect 6710 7046 6724 7098
rect 6748 7046 6762 7098
rect 6762 7046 6774 7098
rect 6774 7046 6804 7098
rect 6828 7046 6838 7098
rect 6838 7046 6884 7098
rect 6588 7044 6644 7046
rect 6668 7044 6724 7046
rect 6748 7044 6804 7046
rect 6828 7044 6884 7046
rect 2870 2080 2926 2136
rect 3422 1400 3478 1456
rect 6588 6010 6644 6012
rect 6668 6010 6724 6012
rect 6748 6010 6804 6012
rect 6828 6010 6884 6012
rect 6588 5958 6634 6010
rect 6634 5958 6644 6010
rect 6668 5958 6698 6010
rect 6698 5958 6710 6010
rect 6710 5958 6724 6010
rect 6748 5958 6762 6010
rect 6762 5958 6774 6010
rect 6774 5958 6804 6010
rect 6828 5958 6838 6010
rect 6838 5958 6884 6010
rect 6588 5956 6644 5958
rect 6668 5956 6724 5958
rect 6748 5956 6804 5958
rect 6828 5956 6884 5958
rect 6588 4922 6644 4924
rect 6668 4922 6724 4924
rect 6748 4922 6804 4924
rect 6828 4922 6884 4924
rect 6588 4870 6634 4922
rect 6634 4870 6644 4922
rect 6668 4870 6698 4922
rect 6698 4870 6710 4922
rect 6710 4870 6724 4922
rect 6748 4870 6762 4922
rect 6762 4870 6774 4922
rect 6774 4870 6804 4922
rect 6828 4870 6838 4922
rect 6838 4870 6884 4922
rect 6588 4868 6644 4870
rect 6668 4868 6724 4870
rect 6748 4868 6804 4870
rect 6828 4868 6884 4870
rect 6588 3834 6644 3836
rect 6668 3834 6724 3836
rect 6748 3834 6804 3836
rect 6828 3834 6884 3836
rect 6588 3782 6634 3834
rect 6634 3782 6644 3834
rect 6668 3782 6698 3834
rect 6698 3782 6710 3834
rect 6710 3782 6724 3834
rect 6748 3782 6762 3834
rect 6762 3782 6774 3834
rect 6774 3782 6804 3834
rect 6828 3782 6838 3834
rect 6838 3782 6884 3834
rect 6588 3780 6644 3782
rect 6668 3780 6724 3782
rect 6748 3780 6804 3782
rect 6828 3780 6884 3782
rect 6588 2746 6644 2748
rect 6668 2746 6724 2748
rect 6748 2746 6804 2748
rect 6828 2746 6884 2748
rect 6588 2694 6634 2746
rect 6634 2694 6644 2746
rect 6668 2694 6698 2746
rect 6698 2694 6710 2746
rect 6710 2694 6724 2746
rect 6748 2694 6762 2746
rect 6762 2694 6774 2746
rect 6774 2694 6804 2746
rect 6828 2694 6838 2746
rect 6838 2694 6884 2746
rect 6588 2692 6644 2694
rect 6668 2692 6724 2694
rect 6748 2692 6804 2694
rect 6828 2692 6884 2694
rect 12220 26138 12276 26140
rect 12300 26138 12356 26140
rect 12380 26138 12436 26140
rect 12460 26138 12516 26140
rect 12220 26086 12266 26138
rect 12266 26086 12276 26138
rect 12300 26086 12330 26138
rect 12330 26086 12342 26138
rect 12342 26086 12356 26138
rect 12380 26086 12394 26138
rect 12394 26086 12406 26138
rect 12406 26086 12436 26138
rect 12460 26086 12470 26138
rect 12470 26086 12516 26138
rect 12220 26084 12276 26086
rect 12300 26084 12356 26086
rect 12380 26084 12436 26086
rect 12460 26084 12516 26086
rect 12220 25050 12276 25052
rect 12300 25050 12356 25052
rect 12380 25050 12436 25052
rect 12460 25050 12516 25052
rect 12220 24998 12266 25050
rect 12266 24998 12276 25050
rect 12300 24998 12330 25050
rect 12330 24998 12342 25050
rect 12342 24998 12356 25050
rect 12380 24998 12394 25050
rect 12394 24998 12406 25050
rect 12406 24998 12436 25050
rect 12460 24998 12470 25050
rect 12470 24998 12516 25050
rect 12220 24996 12276 24998
rect 12300 24996 12356 24998
rect 12380 24996 12436 24998
rect 12460 24996 12516 24998
rect 12990 30096 13046 30152
rect 12806 24656 12862 24712
rect 12220 23962 12276 23964
rect 12300 23962 12356 23964
rect 12380 23962 12436 23964
rect 12460 23962 12516 23964
rect 12220 23910 12266 23962
rect 12266 23910 12276 23962
rect 12300 23910 12330 23962
rect 12330 23910 12342 23962
rect 12342 23910 12356 23962
rect 12380 23910 12394 23962
rect 12394 23910 12406 23962
rect 12406 23910 12436 23962
rect 12460 23910 12470 23962
rect 12470 23910 12516 23962
rect 12220 23908 12276 23910
rect 12300 23908 12356 23910
rect 12380 23908 12436 23910
rect 12460 23908 12516 23910
rect 12220 22874 12276 22876
rect 12300 22874 12356 22876
rect 12380 22874 12436 22876
rect 12460 22874 12516 22876
rect 12220 22822 12266 22874
rect 12266 22822 12276 22874
rect 12300 22822 12330 22874
rect 12330 22822 12342 22874
rect 12342 22822 12356 22874
rect 12380 22822 12394 22874
rect 12394 22822 12406 22874
rect 12406 22822 12436 22874
rect 12460 22822 12470 22874
rect 12470 22822 12516 22874
rect 12220 22820 12276 22822
rect 12300 22820 12356 22822
rect 12380 22820 12436 22822
rect 12460 22820 12516 22822
rect 12220 21786 12276 21788
rect 12300 21786 12356 21788
rect 12380 21786 12436 21788
rect 12460 21786 12516 21788
rect 12220 21734 12266 21786
rect 12266 21734 12276 21786
rect 12300 21734 12330 21786
rect 12330 21734 12342 21786
rect 12342 21734 12356 21786
rect 12380 21734 12394 21786
rect 12394 21734 12406 21786
rect 12406 21734 12436 21786
rect 12460 21734 12470 21786
rect 12470 21734 12516 21786
rect 12220 21732 12276 21734
rect 12300 21732 12356 21734
rect 12380 21732 12436 21734
rect 12460 21732 12516 21734
rect 12220 20698 12276 20700
rect 12300 20698 12356 20700
rect 12380 20698 12436 20700
rect 12460 20698 12516 20700
rect 12220 20646 12266 20698
rect 12266 20646 12276 20698
rect 12300 20646 12330 20698
rect 12330 20646 12342 20698
rect 12342 20646 12356 20698
rect 12380 20646 12394 20698
rect 12394 20646 12406 20698
rect 12406 20646 12436 20698
rect 12460 20646 12470 20698
rect 12470 20646 12516 20698
rect 12220 20644 12276 20646
rect 12300 20644 12356 20646
rect 12380 20644 12436 20646
rect 12460 20644 12516 20646
rect 12220 19610 12276 19612
rect 12300 19610 12356 19612
rect 12380 19610 12436 19612
rect 12460 19610 12516 19612
rect 12220 19558 12266 19610
rect 12266 19558 12276 19610
rect 12300 19558 12330 19610
rect 12330 19558 12342 19610
rect 12342 19558 12356 19610
rect 12380 19558 12394 19610
rect 12394 19558 12406 19610
rect 12406 19558 12436 19610
rect 12460 19558 12470 19610
rect 12470 19558 12516 19610
rect 12220 19556 12276 19558
rect 12300 19556 12356 19558
rect 12380 19556 12436 19558
rect 12460 19556 12516 19558
rect 12220 18522 12276 18524
rect 12300 18522 12356 18524
rect 12380 18522 12436 18524
rect 12460 18522 12516 18524
rect 12220 18470 12266 18522
rect 12266 18470 12276 18522
rect 12300 18470 12330 18522
rect 12330 18470 12342 18522
rect 12342 18470 12356 18522
rect 12380 18470 12394 18522
rect 12394 18470 12406 18522
rect 12406 18470 12436 18522
rect 12460 18470 12470 18522
rect 12470 18470 12516 18522
rect 12220 18468 12276 18470
rect 12300 18468 12356 18470
rect 12380 18468 12436 18470
rect 12460 18468 12516 18470
rect 12220 17434 12276 17436
rect 12300 17434 12356 17436
rect 12380 17434 12436 17436
rect 12460 17434 12516 17436
rect 12220 17382 12266 17434
rect 12266 17382 12276 17434
rect 12300 17382 12330 17434
rect 12330 17382 12342 17434
rect 12342 17382 12356 17434
rect 12380 17382 12394 17434
rect 12394 17382 12406 17434
rect 12406 17382 12436 17434
rect 12460 17382 12470 17434
rect 12470 17382 12516 17434
rect 12220 17380 12276 17382
rect 12300 17380 12356 17382
rect 12380 17380 12436 17382
rect 12460 17380 12516 17382
rect 13082 28736 13138 28792
rect 13082 25744 13138 25800
rect 13450 30368 13506 30424
rect 13450 27920 13506 27976
rect 13358 27648 13414 27704
rect 13726 29280 13782 29336
rect 13542 27104 13598 27160
rect 13542 26988 13598 27024
rect 13542 26968 13544 26988
rect 13544 26968 13596 26988
rect 13596 26968 13598 26988
rect 13174 22752 13230 22808
rect 14002 32816 14058 32872
rect 14094 32544 14150 32600
rect 14002 29144 14058 29200
rect 14002 29044 14004 29064
rect 14004 29044 14056 29064
rect 14056 29044 14058 29064
rect 14002 29008 14058 29044
rect 12220 16346 12276 16348
rect 12300 16346 12356 16348
rect 12380 16346 12436 16348
rect 12460 16346 12516 16348
rect 12220 16294 12266 16346
rect 12266 16294 12276 16346
rect 12300 16294 12330 16346
rect 12330 16294 12342 16346
rect 12342 16294 12356 16346
rect 12380 16294 12394 16346
rect 12394 16294 12406 16346
rect 12406 16294 12436 16346
rect 12460 16294 12470 16346
rect 12470 16294 12516 16346
rect 12220 16292 12276 16294
rect 12300 16292 12356 16294
rect 12380 16292 12436 16294
rect 12460 16292 12516 16294
rect 12220 15258 12276 15260
rect 12300 15258 12356 15260
rect 12380 15258 12436 15260
rect 12460 15258 12516 15260
rect 12220 15206 12266 15258
rect 12266 15206 12276 15258
rect 12300 15206 12330 15258
rect 12330 15206 12342 15258
rect 12342 15206 12356 15258
rect 12380 15206 12394 15258
rect 12394 15206 12406 15258
rect 12406 15206 12436 15258
rect 12460 15206 12470 15258
rect 12470 15206 12516 15258
rect 12220 15204 12276 15206
rect 12300 15204 12356 15206
rect 12380 15204 12436 15206
rect 12460 15204 12516 15206
rect 12220 14170 12276 14172
rect 12300 14170 12356 14172
rect 12380 14170 12436 14172
rect 12460 14170 12516 14172
rect 12220 14118 12266 14170
rect 12266 14118 12276 14170
rect 12300 14118 12330 14170
rect 12330 14118 12342 14170
rect 12342 14118 12356 14170
rect 12380 14118 12394 14170
rect 12394 14118 12406 14170
rect 12406 14118 12436 14170
rect 12460 14118 12470 14170
rect 12470 14118 12516 14170
rect 12220 14116 12276 14118
rect 12300 14116 12356 14118
rect 12380 14116 12436 14118
rect 12460 14116 12516 14118
rect 12220 13082 12276 13084
rect 12300 13082 12356 13084
rect 12380 13082 12436 13084
rect 12460 13082 12516 13084
rect 12220 13030 12266 13082
rect 12266 13030 12276 13082
rect 12300 13030 12330 13082
rect 12330 13030 12342 13082
rect 12342 13030 12356 13082
rect 12380 13030 12394 13082
rect 12394 13030 12406 13082
rect 12406 13030 12436 13082
rect 12460 13030 12470 13082
rect 12470 13030 12516 13082
rect 12220 13028 12276 13030
rect 12300 13028 12356 13030
rect 12380 13028 12436 13030
rect 12460 13028 12516 13030
rect 12220 11994 12276 11996
rect 12300 11994 12356 11996
rect 12380 11994 12436 11996
rect 12460 11994 12516 11996
rect 12220 11942 12266 11994
rect 12266 11942 12276 11994
rect 12300 11942 12330 11994
rect 12330 11942 12342 11994
rect 12342 11942 12356 11994
rect 12380 11942 12394 11994
rect 12394 11942 12406 11994
rect 12406 11942 12436 11994
rect 12460 11942 12470 11994
rect 12470 11942 12516 11994
rect 12220 11940 12276 11942
rect 12300 11940 12356 11942
rect 12380 11940 12436 11942
rect 12460 11940 12516 11942
rect 12220 10906 12276 10908
rect 12300 10906 12356 10908
rect 12380 10906 12436 10908
rect 12460 10906 12516 10908
rect 12220 10854 12266 10906
rect 12266 10854 12276 10906
rect 12300 10854 12330 10906
rect 12330 10854 12342 10906
rect 12342 10854 12356 10906
rect 12380 10854 12394 10906
rect 12394 10854 12406 10906
rect 12406 10854 12436 10906
rect 12460 10854 12470 10906
rect 12470 10854 12516 10906
rect 12220 10852 12276 10854
rect 12300 10852 12356 10854
rect 12380 10852 12436 10854
rect 12460 10852 12516 10854
rect 12220 9818 12276 9820
rect 12300 9818 12356 9820
rect 12380 9818 12436 9820
rect 12460 9818 12516 9820
rect 12220 9766 12266 9818
rect 12266 9766 12276 9818
rect 12300 9766 12330 9818
rect 12330 9766 12342 9818
rect 12342 9766 12356 9818
rect 12380 9766 12394 9818
rect 12394 9766 12406 9818
rect 12406 9766 12436 9818
rect 12460 9766 12470 9818
rect 12470 9766 12516 9818
rect 12220 9764 12276 9766
rect 12300 9764 12356 9766
rect 12380 9764 12436 9766
rect 12460 9764 12516 9766
rect 12220 8730 12276 8732
rect 12300 8730 12356 8732
rect 12380 8730 12436 8732
rect 12460 8730 12516 8732
rect 12220 8678 12266 8730
rect 12266 8678 12276 8730
rect 12300 8678 12330 8730
rect 12330 8678 12342 8730
rect 12342 8678 12356 8730
rect 12380 8678 12394 8730
rect 12394 8678 12406 8730
rect 12406 8678 12436 8730
rect 12460 8678 12470 8730
rect 12470 8678 12516 8730
rect 12220 8676 12276 8678
rect 12300 8676 12356 8678
rect 12380 8676 12436 8678
rect 12460 8676 12516 8678
rect 12220 7642 12276 7644
rect 12300 7642 12356 7644
rect 12380 7642 12436 7644
rect 12460 7642 12516 7644
rect 12220 7590 12266 7642
rect 12266 7590 12276 7642
rect 12300 7590 12330 7642
rect 12330 7590 12342 7642
rect 12342 7590 12356 7642
rect 12380 7590 12394 7642
rect 12394 7590 12406 7642
rect 12406 7590 12436 7642
rect 12460 7590 12470 7642
rect 12470 7590 12516 7642
rect 12220 7588 12276 7590
rect 12300 7588 12356 7590
rect 12380 7588 12436 7590
rect 12460 7588 12516 7590
rect 12220 6554 12276 6556
rect 12300 6554 12356 6556
rect 12380 6554 12436 6556
rect 12460 6554 12516 6556
rect 12220 6502 12266 6554
rect 12266 6502 12276 6554
rect 12300 6502 12330 6554
rect 12330 6502 12342 6554
rect 12342 6502 12356 6554
rect 12380 6502 12394 6554
rect 12394 6502 12406 6554
rect 12406 6502 12436 6554
rect 12460 6502 12470 6554
rect 12470 6502 12516 6554
rect 12220 6500 12276 6502
rect 12300 6500 12356 6502
rect 12380 6500 12436 6502
rect 12460 6500 12516 6502
rect 12220 5466 12276 5468
rect 12300 5466 12356 5468
rect 12380 5466 12436 5468
rect 12460 5466 12516 5468
rect 12220 5414 12266 5466
rect 12266 5414 12276 5466
rect 12300 5414 12330 5466
rect 12330 5414 12342 5466
rect 12342 5414 12356 5466
rect 12380 5414 12394 5466
rect 12394 5414 12406 5466
rect 12406 5414 12436 5466
rect 12460 5414 12470 5466
rect 12470 5414 12516 5466
rect 12220 5412 12276 5414
rect 12300 5412 12356 5414
rect 12380 5412 12436 5414
rect 12460 5412 12516 5414
rect 12220 4378 12276 4380
rect 12300 4378 12356 4380
rect 12380 4378 12436 4380
rect 12460 4378 12516 4380
rect 12220 4326 12266 4378
rect 12266 4326 12276 4378
rect 12300 4326 12330 4378
rect 12330 4326 12342 4378
rect 12342 4326 12356 4378
rect 12380 4326 12394 4378
rect 12394 4326 12406 4378
rect 12406 4326 12436 4378
rect 12460 4326 12470 4378
rect 12470 4326 12516 4378
rect 12220 4324 12276 4326
rect 12300 4324 12356 4326
rect 12380 4324 12436 4326
rect 12460 4324 12516 4326
rect 12220 3290 12276 3292
rect 12300 3290 12356 3292
rect 12380 3290 12436 3292
rect 12460 3290 12516 3292
rect 12220 3238 12266 3290
rect 12266 3238 12276 3290
rect 12300 3238 12330 3290
rect 12330 3238 12342 3290
rect 12342 3238 12356 3290
rect 12380 3238 12394 3290
rect 12394 3238 12406 3290
rect 12406 3238 12436 3290
rect 12460 3238 12470 3290
rect 12470 3238 12516 3290
rect 12220 3236 12276 3238
rect 12300 3236 12356 3238
rect 12380 3236 12436 3238
rect 12460 3236 12516 3238
rect 12220 2202 12276 2204
rect 12300 2202 12356 2204
rect 12380 2202 12436 2204
rect 12460 2202 12516 2204
rect 12220 2150 12266 2202
rect 12266 2150 12276 2202
rect 12300 2150 12330 2202
rect 12330 2150 12342 2202
rect 12342 2150 12356 2202
rect 12380 2150 12394 2202
rect 12394 2150 12406 2202
rect 12406 2150 12436 2202
rect 12460 2150 12470 2202
rect 12470 2150 12516 2202
rect 12220 2148 12276 2150
rect 12300 2148 12356 2150
rect 12380 2148 12436 2150
rect 12460 2148 12516 2150
rect 14462 35436 14464 35456
rect 14464 35436 14516 35456
rect 14516 35436 14518 35456
rect 14462 35400 14518 35436
rect 14554 34992 14610 35048
rect 14462 34584 14518 34640
rect 15290 40432 15346 40488
rect 14554 34060 14610 34096
rect 14554 34040 14556 34060
rect 14556 34040 14608 34060
rect 14608 34040 14610 34060
rect 14554 33768 14610 33824
rect 14462 33632 14518 33688
rect 14462 33360 14518 33416
rect 14646 33360 14702 33416
rect 14278 32544 14334 32600
rect 14554 32544 14610 32600
rect 15014 36352 15070 36408
rect 15014 34992 15070 35048
rect 14922 34040 14978 34096
rect 15198 36624 15254 36680
rect 15290 34040 15346 34096
rect 15750 37440 15806 37496
rect 16670 40160 16726 40216
rect 17038 39888 17094 39944
rect 16854 39480 16910 39536
rect 17038 39480 17094 39536
rect 17682 40160 17738 40216
rect 17498 39616 17554 39672
rect 16670 39208 16726 39264
rect 16854 39208 16910 39264
rect 16578 38664 16634 38720
rect 17038 38800 17094 38856
rect 16302 37984 16358 38040
rect 15842 36896 15898 36952
rect 16302 37440 16358 37496
rect 16486 37984 16542 38040
rect 16118 36896 16174 36952
rect 15658 36624 15714 36680
rect 15658 36352 15714 36408
rect 15934 36352 15990 36408
rect 16302 36624 16358 36680
rect 18510 40568 18566 40624
rect 17852 39738 17908 39740
rect 17932 39738 17988 39740
rect 18012 39738 18068 39740
rect 18092 39738 18148 39740
rect 17852 39686 17898 39738
rect 17898 39686 17908 39738
rect 17932 39686 17962 39738
rect 17962 39686 17974 39738
rect 17974 39686 17988 39738
rect 18012 39686 18026 39738
rect 18026 39686 18038 39738
rect 18038 39686 18068 39738
rect 18092 39686 18102 39738
rect 18102 39686 18148 39738
rect 17852 39684 17908 39686
rect 17932 39684 17988 39686
rect 18012 39684 18068 39686
rect 18092 39684 18148 39686
rect 18326 39752 18382 39808
rect 18326 39072 18382 39128
rect 18326 38836 18328 38856
rect 18328 38836 18380 38856
rect 18380 38836 18382 38856
rect 18326 38800 18382 38836
rect 18510 38800 18566 38856
rect 16854 37460 16910 37496
rect 16854 37440 16856 37460
rect 16856 37440 16908 37460
rect 16908 37440 16910 37460
rect 17038 37440 17094 37496
rect 16486 36644 16542 36680
rect 17406 38664 17462 38720
rect 17314 37440 17370 37496
rect 17682 38664 17738 38720
rect 17852 38650 17908 38652
rect 17932 38650 17988 38652
rect 18012 38650 18068 38652
rect 18092 38650 18148 38652
rect 17852 38598 17898 38650
rect 17898 38598 17908 38650
rect 17932 38598 17962 38650
rect 17962 38598 17974 38650
rect 17974 38598 17988 38650
rect 18012 38598 18026 38650
rect 18026 38598 18038 38650
rect 18038 38598 18068 38650
rect 18092 38598 18102 38650
rect 18102 38598 18148 38650
rect 17852 38596 17908 38598
rect 17932 38596 17988 38598
rect 18012 38596 18068 38598
rect 18092 38596 18148 38598
rect 17682 37576 17738 37632
rect 17590 37440 17646 37496
rect 16486 36624 16488 36644
rect 16488 36624 16540 36644
rect 16540 36624 16542 36644
rect 16210 36372 16266 36408
rect 16210 36352 16212 36372
rect 16212 36352 16264 36372
rect 16264 36352 16266 36372
rect 16394 36352 16450 36408
rect 15474 34992 15530 35048
rect 15474 34740 15530 34776
rect 15474 34720 15476 34740
rect 15476 34720 15528 34740
rect 15528 34720 15530 34740
rect 15934 35400 15990 35456
rect 15750 34040 15806 34096
rect 16302 35672 16358 35728
rect 18326 37576 18382 37632
rect 17852 37562 17908 37564
rect 17932 37562 17988 37564
rect 18012 37562 18068 37564
rect 18092 37562 18148 37564
rect 17852 37510 17898 37562
rect 17898 37510 17908 37562
rect 17932 37510 17962 37562
rect 17962 37510 17974 37562
rect 17974 37510 17988 37562
rect 18012 37510 18026 37562
rect 18026 37510 18038 37562
rect 18038 37510 18068 37562
rect 18092 37510 18102 37562
rect 18102 37510 18148 37562
rect 17852 37508 17908 37510
rect 17932 37508 17988 37510
rect 18012 37508 18068 37510
rect 18092 37508 18148 37510
rect 18234 37460 18290 37496
rect 18234 37440 18236 37460
rect 18236 37440 18288 37460
rect 18288 37440 18290 37460
rect 17682 36488 17738 36544
rect 18234 36488 18290 36544
rect 17852 36474 17908 36476
rect 17932 36474 17988 36476
rect 18012 36474 18068 36476
rect 18092 36474 18148 36476
rect 17852 36422 17898 36474
rect 17898 36422 17908 36474
rect 17932 36422 17962 36474
rect 17962 36422 17974 36474
rect 17974 36422 17988 36474
rect 18012 36422 18026 36474
rect 18026 36422 18038 36474
rect 18038 36422 18068 36474
rect 18092 36422 18102 36474
rect 18102 36422 18148 36474
rect 17852 36420 17908 36422
rect 17932 36420 17988 36422
rect 18012 36420 18068 36422
rect 18092 36420 18148 36422
rect 17682 36352 17738 36408
rect 19154 40296 19210 40352
rect 18786 38936 18842 38992
rect 18786 38664 18842 38720
rect 18694 38392 18750 38448
rect 19338 39616 19394 39672
rect 16762 35400 16818 35456
rect 16302 33940 16304 33960
rect 16304 33940 16356 33960
rect 16356 33940 16358 33960
rect 16302 33904 16358 33940
rect 15566 33496 15622 33552
rect 14738 32020 14794 32056
rect 14738 32000 14740 32020
rect 14740 32000 14792 32020
rect 14792 32000 14794 32020
rect 14922 32136 14978 32192
rect 14186 31592 14242 31648
rect 14646 31456 14702 31512
rect 14554 31184 14610 31240
rect 14186 29688 14242 29744
rect 14186 29144 14242 29200
rect 14278 28464 14334 28520
rect 14278 28328 14334 28384
rect 14186 26560 14242 26616
rect 14462 29552 14518 29608
rect 14462 29280 14518 29336
rect 14646 29280 14702 29336
rect 14646 29180 14648 29200
rect 14648 29180 14700 29200
rect 14700 29180 14702 29200
rect 14646 29144 14702 29180
rect 14646 28600 14702 28656
rect 14830 31456 14886 31512
rect 14830 30504 14886 30560
rect 14830 29960 14886 30016
rect 15198 30232 15254 30288
rect 15290 29688 15346 29744
rect 14922 28736 14978 28792
rect 15658 33360 15714 33416
rect 15658 29824 15714 29880
rect 15198 28872 15254 28928
rect 14738 26696 14794 26752
rect 14922 28328 14978 28384
rect 15198 28328 15254 28384
rect 15014 28192 15070 28248
rect 14462 25880 14518 25936
rect 14830 25472 14886 25528
rect 14738 25200 14794 25256
rect 15290 28056 15346 28112
rect 15198 27784 15254 27840
rect 15106 27240 15162 27296
rect 15014 26424 15070 26480
rect 15290 27376 15346 27432
rect 15198 26288 15254 26344
rect 15290 26016 15346 26072
rect 14922 24928 14978 24984
rect 14922 24248 14978 24304
rect 14646 24112 14702 24168
rect 15106 23840 15162 23896
rect 14738 23704 14794 23760
rect 15934 33360 15990 33416
rect 17038 35400 17094 35456
rect 17130 35284 17186 35320
rect 17130 35264 17132 35284
rect 17132 35264 17184 35284
rect 17184 35264 17186 35284
rect 18326 36352 18382 36408
rect 17590 35264 17646 35320
rect 18786 36624 18842 36680
rect 18786 36080 18842 36136
rect 18326 35536 18382 35592
rect 18510 35536 18566 35592
rect 17852 35386 17908 35388
rect 17932 35386 17988 35388
rect 18012 35386 18068 35388
rect 18092 35386 18148 35388
rect 17852 35334 17898 35386
rect 17898 35334 17908 35386
rect 17932 35334 17962 35386
rect 17962 35334 17974 35386
rect 17974 35334 17988 35386
rect 18012 35334 18026 35386
rect 18026 35334 18038 35386
rect 18038 35334 18068 35386
rect 18092 35334 18102 35386
rect 18102 35334 18148 35386
rect 17852 35332 17908 35334
rect 17932 35332 17988 35334
rect 18012 35332 18068 35334
rect 18092 35332 18148 35334
rect 18326 35284 18382 35320
rect 18326 35264 18328 35284
rect 18328 35264 18380 35284
rect 18380 35264 18382 35284
rect 16946 34176 17002 34232
rect 18234 34992 18290 35048
rect 17682 34312 17738 34368
rect 17852 34298 17908 34300
rect 17932 34298 17988 34300
rect 18012 34298 18068 34300
rect 18092 34298 18148 34300
rect 17852 34246 17898 34298
rect 17898 34246 17908 34298
rect 17932 34246 17962 34298
rect 17962 34246 17974 34298
rect 17974 34246 17988 34298
rect 18012 34246 18026 34298
rect 18026 34246 18038 34298
rect 18038 34246 18068 34298
rect 18092 34246 18102 34298
rect 18102 34246 18148 34298
rect 17852 34244 17908 34246
rect 17932 34244 17988 34246
rect 18012 34244 18068 34246
rect 18092 34244 18148 34246
rect 18326 34312 18382 34368
rect 15842 31320 15898 31376
rect 16118 31320 16174 31376
rect 16026 30368 16082 30424
rect 15474 28872 15530 28928
rect 15566 28600 15622 28656
rect 15750 28872 15806 28928
rect 15750 28600 15806 28656
rect 15474 27920 15530 27976
rect 15934 29824 15990 29880
rect 18510 34992 18566 35048
rect 19062 36624 19118 36680
rect 18970 36116 18972 36136
rect 18972 36116 19024 36136
rect 19024 36116 19026 36136
rect 18970 36080 19026 36116
rect 17498 33360 17554 33416
rect 20074 40024 20130 40080
rect 19798 38392 19854 38448
rect 19982 38528 20038 38584
rect 19430 36896 19486 36952
rect 19614 36896 19670 36952
rect 19614 35808 19670 35864
rect 20534 40160 20590 40216
rect 20166 38936 20222 38992
rect 19706 34720 19762 34776
rect 20074 35128 20130 35184
rect 19982 34720 20038 34776
rect 18694 33632 18750 33688
rect 17852 33210 17908 33212
rect 17932 33210 17988 33212
rect 18012 33210 18068 33212
rect 18092 33210 18148 33212
rect 17852 33158 17898 33210
rect 17898 33158 17908 33210
rect 17932 33158 17962 33210
rect 17962 33158 17974 33210
rect 17974 33158 17988 33210
rect 18012 33158 18026 33210
rect 18026 33158 18038 33210
rect 18038 33158 18068 33210
rect 18092 33158 18102 33210
rect 18102 33158 18148 33210
rect 17852 33156 17908 33158
rect 17932 33156 17988 33158
rect 18012 33156 18068 33158
rect 18092 33156 18148 33158
rect 16762 32020 16818 32056
rect 16762 32000 16764 32020
rect 16764 32000 16816 32020
rect 16816 32000 16818 32020
rect 17222 32544 17278 32600
rect 17406 33088 17462 33144
rect 17682 32836 17738 32872
rect 17682 32816 17684 32836
rect 17684 32816 17736 32836
rect 17736 32816 17738 32836
rect 17958 32816 18014 32872
rect 18602 33108 18658 33144
rect 18602 33088 18604 33108
rect 18604 33088 18656 33108
rect 18656 33088 18658 33108
rect 17222 32136 17278 32192
rect 17130 32000 17186 32056
rect 16394 31456 16450 31512
rect 16210 30368 16266 30424
rect 16578 29280 16634 29336
rect 18418 32680 18474 32736
rect 17682 32172 17684 32192
rect 17684 32172 17736 32192
rect 17736 32172 17738 32192
rect 17682 32136 17738 32172
rect 17406 31456 17462 31512
rect 17682 32000 17738 32056
rect 18234 32136 18290 32192
rect 17852 32122 17908 32124
rect 17932 32122 17988 32124
rect 18012 32122 18068 32124
rect 18092 32122 18148 32124
rect 17852 32070 17898 32122
rect 17898 32070 17908 32122
rect 17932 32070 17962 32122
rect 17962 32070 17974 32122
rect 17974 32070 17988 32122
rect 18012 32070 18026 32122
rect 18026 32070 18038 32122
rect 18038 32070 18068 32122
rect 18092 32070 18102 32122
rect 18102 32070 18148 32122
rect 17852 32068 17908 32070
rect 17932 32068 17988 32070
rect 18012 32068 18068 32070
rect 18092 32068 18148 32070
rect 18970 32408 19026 32464
rect 19430 33224 19486 33280
rect 19614 33224 19670 33280
rect 19154 32408 19210 32464
rect 17222 31048 17278 31104
rect 17682 31048 17738 31104
rect 17852 31034 17908 31036
rect 17932 31034 17988 31036
rect 18012 31034 18068 31036
rect 18092 31034 18148 31036
rect 17852 30982 17898 31034
rect 17898 30982 17908 31034
rect 17932 30982 17962 31034
rect 17962 30982 17974 31034
rect 17974 30982 17988 31034
rect 18012 30982 18026 31034
rect 18026 30982 18038 31034
rect 18038 30982 18068 31034
rect 18092 30982 18102 31034
rect 18102 30982 18148 31034
rect 17852 30980 17908 30982
rect 17932 30980 17988 30982
rect 18012 30980 18068 30982
rect 18092 30980 18148 30982
rect 18326 30912 18382 30968
rect 17038 29960 17094 30016
rect 17314 30096 17370 30152
rect 17222 29960 17278 30016
rect 17958 30096 18014 30152
rect 18234 30232 18290 30288
rect 17406 29824 17462 29880
rect 17038 29280 17094 29336
rect 16670 29144 16726 29200
rect 16854 29144 16910 29200
rect 16670 28600 16726 28656
rect 15842 27512 15898 27568
rect 15566 27104 15622 27160
rect 15474 26152 15530 26208
rect 15750 25064 15806 25120
rect 15934 27104 15990 27160
rect 15934 25608 15990 25664
rect 15842 23976 15898 24032
rect 16210 27512 16266 27568
rect 16302 27104 16358 27160
rect 16302 26832 16358 26888
rect 16118 26696 16174 26752
rect 16854 27240 16910 27296
rect 16670 26732 16672 26752
rect 16672 26732 16724 26752
rect 16724 26732 16726 26752
rect 16670 26696 16726 26732
rect 16670 25336 16726 25392
rect 17852 29946 17908 29948
rect 17932 29946 17988 29948
rect 18012 29946 18068 29948
rect 18092 29946 18148 29948
rect 17852 29894 17898 29946
rect 17898 29894 17908 29946
rect 17932 29894 17962 29946
rect 17962 29894 17974 29946
rect 17974 29894 17988 29946
rect 18012 29894 18026 29946
rect 18026 29894 18038 29946
rect 18038 29894 18068 29946
rect 18092 29894 18102 29946
rect 18102 29894 18148 29946
rect 17852 29892 17908 29894
rect 17932 29892 17988 29894
rect 18012 29892 18068 29894
rect 18092 29892 18148 29894
rect 17682 29824 17738 29880
rect 18234 29824 18290 29880
rect 17682 28872 17738 28928
rect 17498 28636 17500 28656
rect 17500 28636 17552 28656
rect 17552 28636 17554 28656
rect 17498 28600 17554 28636
rect 17852 28858 17908 28860
rect 17932 28858 17988 28860
rect 18012 28858 18068 28860
rect 18092 28858 18148 28860
rect 17852 28806 17898 28858
rect 17898 28806 17908 28858
rect 17932 28806 17962 28858
rect 17962 28806 17974 28858
rect 17974 28806 17988 28858
rect 18012 28806 18026 28858
rect 18026 28806 18038 28858
rect 18038 28806 18068 28858
rect 18092 28806 18102 28858
rect 18102 28806 18148 28858
rect 17852 28804 17908 28806
rect 17932 28804 17988 28806
rect 18012 28804 18068 28806
rect 18092 28804 18148 28806
rect 18326 28872 18382 28928
rect 18786 31084 18788 31104
rect 18788 31084 18840 31104
rect 18840 31084 18842 31104
rect 18786 31048 18842 31084
rect 19062 31592 19118 31648
rect 18510 29824 18566 29880
rect 21638 40840 21694 40896
rect 20718 37984 20774 38040
rect 20810 37440 20866 37496
rect 20994 37440 21050 37496
rect 20718 37032 20774 37088
rect 20810 36760 20866 36816
rect 20534 35944 20590 36000
rect 20902 36352 20958 36408
rect 20810 35944 20866 36000
rect 20442 35672 20498 35728
rect 20350 35536 20406 35592
rect 21454 38120 21510 38176
rect 21086 36352 21142 36408
rect 21086 36080 21142 36136
rect 21086 35536 21142 35592
rect 20994 35400 21050 35456
rect 20258 34060 20314 34096
rect 20258 34040 20260 34060
rect 20260 34040 20312 34060
rect 20312 34040 20314 34060
rect 20074 33632 20130 33688
rect 19982 32680 20038 32736
rect 19890 32408 19946 32464
rect 19430 31592 19486 31648
rect 19338 31340 19394 31376
rect 19338 31320 19340 31340
rect 19340 31320 19392 31340
rect 19392 31320 19394 31340
rect 19614 31320 19670 31376
rect 17590 27784 17646 27840
rect 17852 27770 17908 27772
rect 17932 27770 17988 27772
rect 18012 27770 18068 27772
rect 18092 27770 18148 27772
rect 17852 27718 17898 27770
rect 17898 27718 17908 27770
rect 17932 27718 17962 27770
rect 17962 27718 17974 27770
rect 17974 27718 17988 27770
rect 18012 27718 18026 27770
rect 18026 27718 18038 27770
rect 18038 27718 18068 27770
rect 18092 27718 18102 27770
rect 18102 27718 18148 27770
rect 17852 27716 17908 27718
rect 17932 27716 17988 27718
rect 18012 27716 18068 27718
rect 18092 27716 18148 27718
rect 17682 27648 17738 27704
rect 18326 27784 18382 27840
rect 18234 27648 18290 27704
rect 17222 27240 17278 27296
rect 17406 26696 17462 26752
rect 18326 27512 18382 27568
rect 18510 27548 18512 27568
rect 18512 27548 18564 27568
rect 18564 27548 18566 27568
rect 18510 27512 18566 27548
rect 17590 26696 17646 26752
rect 17852 26682 17908 26684
rect 17932 26682 17988 26684
rect 18012 26682 18068 26684
rect 18092 26682 18148 26684
rect 17852 26630 17898 26682
rect 17898 26630 17908 26682
rect 17932 26630 17962 26682
rect 17962 26630 17974 26682
rect 17974 26630 17988 26682
rect 18012 26630 18026 26682
rect 18026 26630 18038 26682
rect 18038 26630 18068 26682
rect 18092 26630 18102 26682
rect 18102 26630 18148 26682
rect 17852 26628 17908 26630
rect 17932 26628 17988 26630
rect 18012 26628 18068 26630
rect 18092 26628 18148 26630
rect 17682 25608 17738 25664
rect 18234 25608 18290 25664
rect 17852 25594 17908 25596
rect 17932 25594 17988 25596
rect 18012 25594 18068 25596
rect 18092 25594 18148 25596
rect 17852 25542 17898 25594
rect 17898 25542 17908 25594
rect 17932 25542 17962 25594
rect 17962 25542 17974 25594
rect 17974 25542 17988 25594
rect 18012 25542 18026 25594
rect 18026 25542 18038 25594
rect 18038 25542 18068 25594
rect 18092 25542 18102 25594
rect 18102 25542 18148 25594
rect 17852 25540 17908 25542
rect 17932 25540 17988 25542
rect 18012 25540 18068 25542
rect 18092 25540 18148 25542
rect 17682 25472 17738 25528
rect 17852 24506 17908 24508
rect 17932 24506 17988 24508
rect 18012 24506 18068 24508
rect 18092 24506 18148 24508
rect 17852 24454 17898 24506
rect 17898 24454 17908 24506
rect 17932 24454 17962 24506
rect 17962 24454 17974 24506
rect 17974 24454 17988 24506
rect 18012 24454 18026 24506
rect 18026 24454 18038 24506
rect 18038 24454 18068 24506
rect 18092 24454 18102 24506
rect 18102 24454 18148 24506
rect 17852 24452 17908 24454
rect 17932 24452 17988 24454
rect 18012 24452 18068 24454
rect 18092 24452 18148 24454
rect 18510 25064 18566 25120
rect 18418 24248 18474 24304
rect 17852 23418 17908 23420
rect 17932 23418 17988 23420
rect 18012 23418 18068 23420
rect 18092 23418 18148 23420
rect 17852 23366 17898 23418
rect 17898 23366 17908 23418
rect 17932 23366 17962 23418
rect 17962 23366 17974 23418
rect 17974 23366 17988 23418
rect 18012 23366 18026 23418
rect 18026 23366 18038 23418
rect 18038 23366 18068 23418
rect 18092 23366 18102 23418
rect 18102 23366 18148 23418
rect 17852 23364 17908 23366
rect 17932 23364 17988 23366
rect 18012 23364 18068 23366
rect 18092 23364 18148 23366
rect 18418 23976 18474 24032
rect 18510 23860 18566 23896
rect 18510 23840 18512 23860
rect 18512 23840 18564 23860
rect 18564 23840 18566 23860
rect 17852 22330 17908 22332
rect 17932 22330 17988 22332
rect 18012 22330 18068 22332
rect 18092 22330 18148 22332
rect 17852 22278 17898 22330
rect 17898 22278 17908 22330
rect 17932 22278 17962 22330
rect 17962 22278 17974 22330
rect 17974 22278 17988 22330
rect 18012 22278 18026 22330
rect 18026 22278 18038 22330
rect 18038 22278 18068 22330
rect 18092 22278 18102 22330
rect 18102 22278 18148 22330
rect 17852 22276 17908 22278
rect 17932 22276 17988 22278
rect 18012 22276 18068 22278
rect 18092 22276 18148 22278
rect 19890 31184 19946 31240
rect 19430 30504 19486 30560
rect 19706 30368 19762 30424
rect 19890 30368 19946 30424
rect 19062 28600 19118 28656
rect 18786 26560 18842 26616
rect 18694 26424 18750 26480
rect 19706 28192 19762 28248
rect 19890 28192 19946 28248
rect 19890 27512 19946 27568
rect 19246 27376 19302 27432
rect 18970 26696 19026 26752
rect 18878 25744 18934 25800
rect 18786 25336 18842 25392
rect 18970 24656 19026 24712
rect 20074 32408 20130 32464
rect 20166 32000 20222 32056
rect 20074 31728 20130 31784
rect 19614 26016 19670 26072
rect 19338 24384 19394 24440
rect 19246 24112 19302 24168
rect 18694 23740 18696 23760
rect 18696 23740 18748 23760
rect 18748 23740 18750 23760
rect 18694 23704 18750 23740
rect 17852 21242 17908 21244
rect 17932 21242 17988 21244
rect 18012 21242 18068 21244
rect 18092 21242 18148 21244
rect 17852 21190 17898 21242
rect 17898 21190 17908 21242
rect 17932 21190 17962 21242
rect 17962 21190 17974 21242
rect 17974 21190 17988 21242
rect 18012 21190 18026 21242
rect 18026 21190 18038 21242
rect 18038 21190 18068 21242
rect 18092 21190 18102 21242
rect 18102 21190 18148 21242
rect 17852 21188 17908 21190
rect 17932 21188 17988 21190
rect 18012 21188 18068 21190
rect 18092 21188 18148 21190
rect 17852 20154 17908 20156
rect 17932 20154 17988 20156
rect 18012 20154 18068 20156
rect 18092 20154 18148 20156
rect 17852 20102 17898 20154
rect 17898 20102 17908 20154
rect 17932 20102 17962 20154
rect 17962 20102 17974 20154
rect 17974 20102 17988 20154
rect 18012 20102 18026 20154
rect 18026 20102 18038 20154
rect 18038 20102 18068 20154
rect 18092 20102 18102 20154
rect 18102 20102 18148 20154
rect 17852 20100 17908 20102
rect 17932 20100 17988 20102
rect 18012 20100 18068 20102
rect 18092 20100 18148 20102
rect 17852 19066 17908 19068
rect 17932 19066 17988 19068
rect 18012 19066 18068 19068
rect 18092 19066 18148 19068
rect 17852 19014 17898 19066
rect 17898 19014 17908 19066
rect 17932 19014 17962 19066
rect 17962 19014 17974 19066
rect 17974 19014 17988 19066
rect 18012 19014 18026 19066
rect 18026 19014 18038 19066
rect 18038 19014 18068 19066
rect 18092 19014 18102 19066
rect 18102 19014 18148 19066
rect 17852 19012 17908 19014
rect 17932 19012 17988 19014
rect 18012 19012 18068 19014
rect 18092 19012 18148 19014
rect 17852 17978 17908 17980
rect 17932 17978 17988 17980
rect 18012 17978 18068 17980
rect 18092 17978 18148 17980
rect 17852 17926 17898 17978
rect 17898 17926 17908 17978
rect 17932 17926 17962 17978
rect 17962 17926 17974 17978
rect 17974 17926 17988 17978
rect 18012 17926 18026 17978
rect 18026 17926 18038 17978
rect 18038 17926 18068 17978
rect 18092 17926 18102 17978
rect 18102 17926 18148 17978
rect 17852 17924 17908 17926
rect 17932 17924 17988 17926
rect 18012 17924 18068 17926
rect 18092 17924 18148 17926
rect 17852 16890 17908 16892
rect 17932 16890 17988 16892
rect 18012 16890 18068 16892
rect 18092 16890 18148 16892
rect 17852 16838 17898 16890
rect 17898 16838 17908 16890
rect 17932 16838 17962 16890
rect 17962 16838 17974 16890
rect 17974 16838 17988 16890
rect 18012 16838 18026 16890
rect 18026 16838 18038 16890
rect 18038 16838 18068 16890
rect 18092 16838 18102 16890
rect 18102 16838 18148 16890
rect 17852 16836 17908 16838
rect 17932 16836 17988 16838
rect 18012 16836 18068 16838
rect 18092 16836 18148 16838
rect 17852 15802 17908 15804
rect 17932 15802 17988 15804
rect 18012 15802 18068 15804
rect 18092 15802 18148 15804
rect 17852 15750 17898 15802
rect 17898 15750 17908 15802
rect 17932 15750 17962 15802
rect 17962 15750 17974 15802
rect 17974 15750 17988 15802
rect 18012 15750 18026 15802
rect 18026 15750 18038 15802
rect 18038 15750 18068 15802
rect 18092 15750 18102 15802
rect 18102 15750 18148 15802
rect 17852 15748 17908 15750
rect 17932 15748 17988 15750
rect 18012 15748 18068 15750
rect 18092 15748 18148 15750
rect 17852 14714 17908 14716
rect 17932 14714 17988 14716
rect 18012 14714 18068 14716
rect 18092 14714 18148 14716
rect 17852 14662 17898 14714
rect 17898 14662 17908 14714
rect 17932 14662 17962 14714
rect 17962 14662 17974 14714
rect 17974 14662 17988 14714
rect 18012 14662 18026 14714
rect 18026 14662 18038 14714
rect 18038 14662 18068 14714
rect 18092 14662 18102 14714
rect 18102 14662 18148 14714
rect 17852 14660 17908 14662
rect 17932 14660 17988 14662
rect 18012 14660 18068 14662
rect 18092 14660 18148 14662
rect 17852 13626 17908 13628
rect 17932 13626 17988 13628
rect 18012 13626 18068 13628
rect 18092 13626 18148 13628
rect 17852 13574 17898 13626
rect 17898 13574 17908 13626
rect 17932 13574 17962 13626
rect 17962 13574 17974 13626
rect 17974 13574 17988 13626
rect 18012 13574 18026 13626
rect 18026 13574 18038 13626
rect 18038 13574 18068 13626
rect 18092 13574 18102 13626
rect 18102 13574 18148 13626
rect 17852 13572 17908 13574
rect 17932 13572 17988 13574
rect 18012 13572 18068 13574
rect 18092 13572 18148 13574
rect 17852 12538 17908 12540
rect 17932 12538 17988 12540
rect 18012 12538 18068 12540
rect 18092 12538 18148 12540
rect 17852 12486 17898 12538
rect 17898 12486 17908 12538
rect 17932 12486 17962 12538
rect 17962 12486 17974 12538
rect 17974 12486 17988 12538
rect 18012 12486 18026 12538
rect 18026 12486 18038 12538
rect 18038 12486 18068 12538
rect 18092 12486 18102 12538
rect 18102 12486 18148 12538
rect 17852 12484 17908 12486
rect 17932 12484 17988 12486
rect 18012 12484 18068 12486
rect 18092 12484 18148 12486
rect 17852 11450 17908 11452
rect 17932 11450 17988 11452
rect 18012 11450 18068 11452
rect 18092 11450 18148 11452
rect 17852 11398 17898 11450
rect 17898 11398 17908 11450
rect 17932 11398 17962 11450
rect 17962 11398 17974 11450
rect 17974 11398 17988 11450
rect 18012 11398 18026 11450
rect 18026 11398 18038 11450
rect 18038 11398 18068 11450
rect 18092 11398 18102 11450
rect 18102 11398 18148 11450
rect 17852 11396 17908 11398
rect 17932 11396 17988 11398
rect 18012 11396 18068 11398
rect 18092 11396 18148 11398
rect 17852 10362 17908 10364
rect 17932 10362 17988 10364
rect 18012 10362 18068 10364
rect 18092 10362 18148 10364
rect 17852 10310 17898 10362
rect 17898 10310 17908 10362
rect 17932 10310 17962 10362
rect 17962 10310 17974 10362
rect 17974 10310 17988 10362
rect 18012 10310 18026 10362
rect 18026 10310 18038 10362
rect 18038 10310 18068 10362
rect 18092 10310 18102 10362
rect 18102 10310 18148 10362
rect 17852 10308 17908 10310
rect 17932 10308 17988 10310
rect 18012 10308 18068 10310
rect 18092 10308 18148 10310
rect 17852 9274 17908 9276
rect 17932 9274 17988 9276
rect 18012 9274 18068 9276
rect 18092 9274 18148 9276
rect 17852 9222 17898 9274
rect 17898 9222 17908 9274
rect 17932 9222 17962 9274
rect 17962 9222 17974 9274
rect 17974 9222 17988 9274
rect 18012 9222 18026 9274
rect 18026 9222 18038 9274
rect 18038 9222 18068 9274
rect 18092 9222 18102 9274
rect 18102 9222 18148 9274
rect 17852 9220 17908 9222
rect 17932 9220 17988 9222
rect 18012 9220 18068 9222
rect 18092 9220 18148 9222
rect 17852 8186 17908 8188
rect 17932 8186 17988 8188
rect 18012 8186 18068 8188
rect 18092 8186 18148 8188
rect 17852 8134 17898 8186
rect 17898 8134 17908 8186
rect 17932 8134 17962 8186
rect 17962 8134 17974 8186
rect 17974 8134 17988 8186
rect 18012 8134 18026 8186
rect 18026 8134 18038 8186
rect 18038 8134 18068 8186
rect 18092 8134 18102 8186
rect 18102 8134 18148 8186
rect 17852 8132 17908 8134
rect 17932 8132 17988 8134
rect 18012 8132 18068 8134
rect 18092 8132 18148 8134
rect 17852 7098 17908 7100
rect 17932 7098 17988 7100
rect 18012 7098 18068 7100
rect 18092 7098 18148 7100
rect 17852 7046 17898 7098
rect 17898 7046 17908 7098
rect 17932 7046 17962 7098
rect 17962 7046 17974 7098
rect 17974 7046 17988 7098
rect 18012 7046 18026 7098
rect 18026 7046 18038 7098
rect 18038 7046 18068 7098
rect 18092 7046 18102 7098
rect 18102 7046 18148 7098
rect 17852 7044 17908 7046
rect 17932 7044 17988 7046
rect 18012 7044 18068 7046
rect 18092 7044 18148 7046
rect 17852 6010 17908 6012
rect 17932 6010 17988 6012
rect 18012 6010 18068 6012
rect 18092 6010 18148 6012
rect 17852 5958 17898 6010
rect 17898 5958 17908 6010
rect 17932 5958 17962 6010
rect 17962 5958 17974 6010
rect 17974 5958 17988 6010
rect 18012 5958 18026 6010
rect 18026 5958 18038 6010
rect 18038 5958 18068 6010
rect 18092 5958 18102 6010
rect 18102 5958 18148 6010
rect 17852 5956 17908 5958
rect 17932 5956 17988 5958
rect 18012 5956 18068 5958
rect 18092 5956 18148 5958
rect 17852 4922 17908 4924
rect 17932 4922 17988 4924
rect 18012 4922 18068 4924
rect 18092 4922 18148 4924
rect 17852 4870 17898 4922
rect 17898 4870 17908 4922
rect 17932 4870 17962 4922
rect 17962 4870 17974 4922
rect 17974 4870 17988 4922
rect 18012 4870 18026 4922
rect 18026 4870 18038 4922
rect 18038 4870 18068 4922
rect 18092 4870 18102 4922
rect 18102 4870 18148 4922
rect 17852 4868 17908 4870
rect 17932 4868 17988 4870
rect 18012 4868 18068 4870
rect 18092 4868 18148 4870
rect 17852 3834 17908 3836
rect 17932 3834 17988 3836
rect 18012 3834 18068 3836
rect 18092 3834 18148 3836
rect 17852 3782 17898 3834
rect 17898 3782 17908 3834
rect 17932 3782 17962 3834
rect 17962 3782 17974 3834
rect 17974 3782 17988 3834
rect 18012 3782 18026 3834
rect 18026 3782 18038 3834
rect 18038 3782 18068 3834
rect 18092 3782 18102 3834
rect 18102 3782 18148 3834
rect 17852 3780 17908 3782
rect 17932 3780 17988 3782
rect 18012 3780 18068 3782
rect 18092 3780 18148 3782
rect 20534 34040 20590 34096
rect 21086 34620 21088 34640
rect 21088 34620 21140 34640
rect 21140 34620 21142 34640
rect 21086 34584 21142 34620
rect 20350 33088 20406 33144
rect 20350 31728 20406 31784
rect 20718 33768 20774 33824
rect 20902 33632 20958 33688
rect 20902 32952 20958 33008
rect 21362 36488 21418 36544
rect 22006 40160 22062 40216
rect 22926 40704 22982 40760
rect 22650 39072 22706 39128
rect 22834 38936 22890 38992
rect 22098 38528 22154 38584
rect 21730 38412 21786 38448
rect 21730 38392 21732 38412
rect 21732 38392 21784 38412
rect 21784 38392 21786 38412
rect 21914 38428 21916 38448
rect 21916 38428 21968 38448
rect 21968 38428 21970 38448
rect 21914 38392 21970 38428
rect 22282 38528 22338 38584
rect 22190 37576 22246 37632
rect 21822 36624 21878 36680
rect 22098 35944 22154 36000
rect 23662 39616 23718 39672
rect 23484 39194 23540 39196
rect 23564 39194 23620 39196
rect 23644 39194 23700 39196
rect 23724 39194 23780 39196
rect 23484 39142 23530 39194
rect 23530 39142 23540 39194
rect 23564 39142 23594 39194
rect 23594 39142 23606 39194
rect 23606 39142 23620 39194
rect 23644 39142 23658 39194
rect 23658 39142 23670 39194
rect 23670 39142 23700 39194
rect 23724 39142 23734 39194
rect 23734 39142 23780 39194
rect 23484 39140 23540 39142
rect 23564 39140 23620 39142
rect 23644 39140 23700 39142
rect 23724 39140 23780 39142
rect 23484 38106 23540 38108
rect 23564 38106 23620 38108
rect 23644 38106 23700 38108
rect 23724 38106 23780 38108
rect 23484 38054 23530 38106
rect 23530 38054 23540 38106
rect 23564 38054 23594 38106
rect 23594 38054 23606 38106
rect 23606 38054 23620 38106
rect 23644 38054 23658 38106
rect 23658 38054 23670 38106
rect 23670 38054 23700 38106
rect 23724 38054 23734 38106
rect 23734 38054 23780 38106
rect 23484 38052 23540 38054
rect 23564 38052 23620 38054
rect 23644 38052 23700 38054
rect 23724 38052 23780 38054
rect 22742 36760 22798 36816
rect 21638 35128 21694 35184
rect 22558 34720 22614 34776
rect 21362 34176 21418 34232
rect 21546 34176 21602 34232
rect 21178 33768 21234 33824
rect 21086 32952 21142 33008
rect 21362 32852 21364 32872
rect 21364 32852 21416 32872
rect 21416 32852 21418 32872
rect 21362 32816 21418 32852
rect 20718 32020 20774 32056
rect 20718 32000 20720 32020
rect 20720 32000 20772 32020
rect 20772 32000 20774 32020
rect 21546 33632 21602 33688
rect 21822 33768 21878 33824
rect 21730 33632 21786 33688
rect 21914 32544 21970 32600
rect 20258 31184 20314 31240
rect 20258 29008 20314 29064
rect 20166 27512 20222 27568
rect 20626 28464 20682 28520
rect 20810 29960 20866 30016
rect 20902 29008 20958 29064
rect 20810 28464 20866 28520
rect 20534 28056 20590 28112
rect 20718 28056 20774 28112
rect 20718 26968 20774 27024
rect 20442 25880 20498 25936
rect 20350 25472 20406 25528
rect 20718 24656 20774 24712
rect 20074 24248 20130 24304
rect 20442 23296 20498 23352
rect 20350 23160 20406 23216
rect 20074 22344 20130 22400
rect 19982 22072 20038 22128
rect 20534 21392 20590 21448
rect 20442 21256 20498 21312
rect 20810 19372 20866 19408
rect 20810 19352 20812 19372
rect 20812 19352 20864 19372
rect 20864 19352 20866 19372
rect 21362 30640 21418 30696
rect 22282 33768 22338 33824
rect 22282 32816 22338 32872
rect 22190 32544 22246 32600
rect 23018 34720 23074 34776
rect 23484 37018 23540 37020
rect 23564 37018 23620 37020
rect 23644 37018 23700 37020
rect 23724 37018 23780 37020
rect 23484 36966 23530 37018
rect 23530 36966 23540 37018
rect 23564 36966 23594 37018
rect 23594 36966 23606 37018
rect 23606 36966 23620 37018
rect 23644 36966 23658 37018
rect 23658 36966 23670 37018
rect 23670 36966 23700 37018
rect 23724 36966 23734 37018
rect 23734 36966 23780 37018
rect 23484 36964 23540 36966
rect 23564 36964 23620 36966
rect 23644 36964 23700 36966
rect 23724 36964 23780 36966
rect 23662 36352 23718 36408
rect 23484 35930 23540 35932
rect 23564 35930 23620 35932
rect 23644 35930 23700 35932
rect 23724 35930 23780 35932
rect 23484 35878 23530 35930
rect 23530 35878 23540 35930
rect 23564 35878 23594 35930
rect 23594 35878 23606 35930
rect 23606 35878 23620 35930
rect 23644 35878 23658 35930
rect 23658 35878 23670 35930
rect 23670 35878 23700 35930
rect 23724 35878 23734 35930
rect 23734 35878 23780 35930
rect 23484 35876 23540 35878
rect 23564 35876 23620 35878
rect 23644 35876 23700 35878
rect 23724 35876 23780 35878
rect 24490 38956 24546 38992
rect 24490 38936 24492 38956
rect 24492 38936 24544 38956
rect 24544 38936 24546 38956
rect 23938 36760 23994 36816
rect 22374 32680 22430 32736
rect 23570 34992 23626 35048
rect 23484 34842 23540 34844
rect 23564 34842 23620 34844
rect 23644 34842 23700 34844
rect 23724 34842 23780 34844
rect 23484 34790 23530 34842
rect 23530 34790 23540 34842
rect 23564 34790 23594 34842
rect 23594 34790 23606 34842
rect 23606 34790 23620 34842
rect 23644 34790 23658 34842
rect 23658 34790 23670 34842
rect 23670 34790 23700 34842
rect 23724 34790 23734 34842
rect 23734 34790 23780 34842
rect 23484 34788 23540 34790
rect 23564 34788 23620 34790
rect 23644 34788 23700 34790
rect 23724 34788 23780 34790
rect 23484 33754 23540 33756
rect 23564 33754 23620 33756
rect 23644 33754 23700 33756
rect 23724 33754 23780 33756
rect 23484 33702 23530 33754
rect 23530 33702 23540 33754
rect 23564 33702 23594 33754
rect 23594 33702 23606 33754
rect 23606 33702 23620 33754
rect 23644 33702 23658 33754
rect 23658 33702 23670 33754
rect 23670 33702 23700 33754
rect 23724 33702 23734 33754
rect 23734 33702 23780 33754
rect 23484 33700 23540 33702
rect 23564 33700 23620 33702
rect 23644 33700 23700 33702
rect 23724 33700 23780 33702
rect 23294 33632 23350 33688
rect 23386 33360 23442 33416
rect 23110 33260 23112 33280
rect 23112 33260 23164 33280
rect 23164 33260 23166 33280
rect 23110 33224 23166 33260
rect 22926 33088 22982 33144
rect 22650 32544 22706 32600
rect 23202 32544 23258 32600
rect 21730 29960 21786 30016
rect 21914 29824 21970 29880
rect 21822 29180 21824 29200
rect 21824 29180 21876 29200
rect 21876 29180 21878 29200
rect 21822 29144 21878 29180
rect 21270 27784 21326 27840
rect 20994 27240 21050 27296
rect 21546 27376 21602 27432
rect 21730 28736 21786 28792
rect 21914 28872 21970 28928
rect 22466 29960 22522 30016
rect 22742 31048 22798 31104
rect 22834 30640 22890 30696
rect 22650 29824 22706 29880
rect 22374 29416 22430 29472
rect 22190 29144 22246 29200
rect 22558 28872 22614 28928
rect 21914 27956 21916 27976
rect 21916 27956 21968 27976
rect 21968 27956 21970 27976
rect 21914 27920 21970 27956
rect 22006 27512 22062 27568
rect 21638 26152 21694 26208
rect 22190 27512 22246 27568
rect 21730 25336 21786 25392
rect 22834 29164 22890 29200
rect 22834 29144 22836 29164
rect 22836 29144 22888 29164
rect 22888 29144 22890 29164
rect 22650 28328 22706 28384
rect 23484 32666 23540 32668
rect 23564 32666 23620 32668
rect 23644 32666 23700 32668
rect 23724 32666 23780 32668
rect 23484 32614 23530 32666
rect 23530 32614 23540 32666
rect 23564 32614 23594 32666
rect 23594 32614 23606 32666
rect 23606 32614 23620 32666
rect 23644 32614 23658 32666
rect 23658 32614 23670 32666
rect 23670 32614 23700 32666
rect 23724 32614 23734 32666
rect 23734 32614 23780 32666
rect 23484 32612 23540 32614
rect 23564 32612 23620 32614
rect 23644 32612 23700 32614
rect 23724 32612 23780 32614
rect 23484 31578 23540 31580
rect 23564 31578 23620 31580
rect 23644 31578 23700 31580
rect 23724 31578 23780 31580
rect 23484 31526 23530 31578
rect 23530 31526 23540 31578
rect 23564 31526 23594 31578
rect 23594 31526 23606 31578
rect 23606 31526 23620 31578
rect 23644 31526 23658 31578
rect 23658 31526 23670 31578
rect 23670 31526 23700 31578
rect 23724 31526 23734 31578
rect 23734 31526 23780 31578
rect 23484 31524 23540 31526
rect 23564 31524 23620 31526
rect 23644 31524 23700 31526
rect 23724 31524 23780 31526
rect 23110 31456 23166 31512
rect 23110 31340 23166 31376
rect 23110 31320 23112 31340
rect 23112 31320 23164 31340
rect 23164 31320 23166 31340
rect 23110 30096 23166 30152
rect 23484 30490 23540 30492
rect 23564 30490 23620 30492
rect 23644 30490 23700 30492
rect 23724 30490 23780 30492
rect 23484 30438 23530 30490
rect 23530 30438 23540 30490
rect 23564 30438 23594 30490
rect 23594 30438 23606 30490
rect 23606 30438 23620 30490
rect 23644 30438 23658 30490
rect 23658 30438 23670 30490
rect 23670 30438 23700 30490
rect 23724 30438 23734 30490
rect 23734 30438 23780 30490
rect 23484 30436 23540 30438
rect 23564 30436 23620 30438
rect 23644 30436 23700 30438
rect 23724 30436 23780 30438
rect 23570 30232 23626 30288
rect 23478 29824 23534 29880
rect 25134 38292 25136 38312
rect 25136 38292 25188 38312
rect 25188 38292 25190 38312
rect 25134 38256 25190 38292
rect 24214 35808 24270 35864
rect 24122 33768 24178 33824
rect 24766 37440 24822 37496
rect 24858 37188 24914 37224
rect 24858 37168 24860 37188
rect 24860 37168 24912 37188
rect 24912 37168 24914 37188
rect 24674 35128 24730 35184
rect 24766 34856 24822 34912
rect 24766 34312 24822 34368
rect 24858 34040 24914 34096
rect 25134 33768 25190 33824
rect 23938 29996 23940 30016
rect 23940 29996 23992 30016
rect 23992 29996 23994 30016
rect 23938 29960 23994 29996
rect 23938 29416 23994 29472
rect 23484 29402 23540 29404
rect 23564 29402 23620 29404
rect 23644 29402 23700 29404
rect 23724 29402 23780 29404
rect 23484 29350 23530 29402
rect 23530 29350 23540 29402
rect 23564 29350 23594 29402
rect 23594 29350 23606 29402
rect 23606 29350 23620 29402
rect 23644 29350 23658 29402
rect 23658 29350 23670 29402
rect 23670 29350 23700 29402
rect 23724 29350 23734 29402
rect 23734 29350 23780 29402
rect 23484 29348 23540 29350
rect 23564 29348 23620 29350
rect 23644 29348 23700 29350
rect 23724 29348 23780 29350
rect 23294 29280 23350 29336
rect 23018 28484 23074 28520
rect 23018 28464 23020 28484
rect 23020 28464 23072 28484
rect 23072 28464 23074 28484
rect 22834 27784 22890 27840
rect 23018 27784 23074 27840
rect 22926 26988 22982 27024
rect 22926 26968 22928 26988
rect 22928 26968 22980 26988
rect 22980 26968 22982 26988
rect 22558 25608 22614 25664
rect 23484 28314 23540 28316
rect 23564 28314 23620 28316
rect 23644 28314 23700 28316
rect 23724 28314 23780 28316
rect 23484 28262 23530 28314
rect 23530 28262 23540 28314
rect 23564 28262 23594 28314
rect 23594 28262 23606 28314
rect 23606 28262 23620 28314
rect 23644 28262 23658 28314
rect 23658 28262 23670 28314
rect 23670 28262 23700 28314
rect 23724 28262 23734 28314
rect 23734 28262 23780 28314
rect 23484 28260 23540 28262
rect 23564 28260 23620 28262
rect 23644 28260 23700 28262
rect 23724 28260 23780 28262
rect 23938 27920 23994 27976
rect 23754 27784 23810 27840
rect 23484 27226 23540 27228
rect 23564 27226 23620 27228
rect 23644 27226 23700 27228
rect 23724 27226 23780 27228
rect 23484 27174 23530 27226
rect 23530 27174 23540 27226
rect 23564 27174 23594 27226
rect 23594 27174 23606 27226
rect 23606 27174 23620 27226
rect 23644 27174 23658 27226
rect 23658 27174 23670 27226
rect 23670 27174 23700 27226
rect 23724 27174 23734 27226
rect 23734 27174 23780 27226
rect 23484 27172 23540 27174
rect 23564 27172 23620 27174
rect 23644 27172 23700 27174
rect 23724 27172 23780 27174
rect 23478 26424 23534 26480
rect 23484 26138 23540 26140
rect 23564 26138 23620 26140
rect 23644 26138 23700 26140
rect 23724 26138 23780 26140
rect 23484 26086 23530 26138
rect 23530 26086 23540 26138
rect 23564 26086 23594 26138
rect 23594 26086 23606 26138
rect 23606 26086 23620 26138
rect 23644 26086 23658 26138
rect 23658 26086 23670 26138
rect 23670 26086 23700 26138
rect 23724 26086 23734 26138
rect 23734 26086 23780 26138
rect 23484 26084 23540 26086
rect 23564 26084 23620 26086
rect 23644 26084 23700 26086
rect 23724 26084 23780 26086
rect 23938 26832 23994 26888
rect 21730 24928 21786 24984
rect 21454 23568 21510 23624
rect 21822 24520 21878 24576
rect 21546 23044 21602 23080
rect 21546 23024 21548 23044
rect 21548 23024 21600 23044
rect 21600 23024 21602 23044
rect 21822 22888 21878 22944
rect 21914 22616 21970 22672
rect 22098 22752 22154 22808
rect 23484 25050 23540 25052
rect 23564 25050 23620 25052
rect 23644 25050 23700 25052
rect 23724 25050 23780 25052
rect 23484 24998 23530 25050
rect 23530 24998 23540 25050
rect 23564 24998 23594 25050
rect 23594 24998 23606 25050
rect 23606 24998 23620 25050
rect 23644 24998 23658 25050
rect 23658 24998 23670 25050
rect 23670 24998 23700 25050
rect 23724 24998 23734 25050
rect 23734 24998 23780 25050
rect 23484 24996 23540 24998
rect 23564 24996 23620 24998
rect 23644 24996 23700 24998
rect 23724 24996 23780 24998
rect 23662 24692 23664 24712
rect 23664 24692 23716 24712
rect 23716 24692 23718 24712
rect 23662 24656 23718 24692
rect 23938 24520 23994 24576
rect 22926 23160 22982 23216
rect 23202 22888 23258 22944
rect 23018 22616 23074 22672
rect 23018 22208 23074 22264
rect 23110 22072 23166 22128
rect 23294 22616 23350 22672
rect 21822 20340 21824 20360
rect 21824 20340 21876 20360
rect 21876 20340 21878 20360
rect 21822 20304 21878 20340
rect 22190 19488 22246 19544
rect 22374 19760 22430 19816
rect 22374 19508 22430 19544
rect 22374 19488 22376 19508
rect 22376 19488 22428 19508
rect 22428 19488 22430 19508
rect 22834 20848 22890 20904
rect 23484 23962 23540 23964
rect 23564 23962 23620 23964
rect 23644 23962 23700 23964
rect 23724 23962 23780 23964
rect 23484 23910 23530 23962
rect 23530 23910 23540 23962
rect 23564 23910 23594 23962
rect 23594 23910 23606 23962
rect 23606 23910 23620 23962
rect 23644 23910 23658 23962
rect 23658 23910 23670 23962
rect 23670 23910 23700 23962
rect 23724 23910 23734 23962
rect 23734 23910 23780 23962
rect 23484 23908 23540 23910
rect 23564 23908 23620 23910
rect 23644 23908 23700 23910
rect 23724 23908 23780 23910
rect 23484 22874 23540 22876
rect 23564 22874 23620 22876
rect 23644 22874 23700 22876
rect 23724 22874 23780 22876
rect 23484 22822 23530 22874
rect 23530 22822 23540 22874
rect 23564 22822 23594 22874
rect 23594 22822 23606 22874
rect 23606 22822 23620 22874
rect 23644 22822 23658 22874
rect 23658 22822 23670 22874
rect 23670 22822 23700 22874
rect 23724 22822 23734 22874
rect 23734 22822 23780 22874
rect 23484 22820 23540 22822
rect 23564 22820 23620 22822
rect 23644 22820 23700 22822
rect 23724 22820 23780 22822
rect 23484 21786 23540 21788
rect 23564 21786 23620 21788
rect 23644 21786 23700 21788
rect 23724 21786 23780 21788
rect 23484 21734 23530 21786
rect 23530 21734 23540 21786
rect 23564 21734 23594 21786
rect 23594 21734 23606 21786
rect 23606 21734 23620 21786
rect 23644 21734 23658 21786
rect 23658 21734 23670 21786
rect 23670 21734 23700 21786
rect 23724 21734 23734 21786
rect 23734 21734 23780 21786
rect 23484 21732 23540 21734
rect 23564 21732 23620 21734
rect 23644 21732 23700 21734
rect 23724 21732 23780 21734
rect 23570 21548 23626 21584
rect 23570 21528 23572 21548
rect 23572 21528 23624 21548
rect 23624 21528 23626 21548
rect 23202 20884 23204 20904
rect 23204 20884 23256 20904
rect 23256 20884 23258 20904
rect 23202 20848 23258 20884
rect 23484 20698 23540 20700
rect 23564 20698 23620 20700
rect 23644 20698 23700 20700
rect 23724 20698 23780 20700
rect 23484 20646 23530 20698
rect 23530 20646 23540 20698
rect 23564 20646 23594 20698
rect 23594 20646 23606 20698
rect 23606 20646 23620 20698
rect 23644 20646 23658 20698
rect 23658 20646 23670 20698
rect 23670 20646 23700 20698
rect 23724 20646 23734 20698
rect 23734 20646 23780 20698
rect 23484 20644 23540 20646
rect 23564 20644 23620 20646
rect 23644 20644 23700 20646
rect 23724 20644 23780 20646
rect 23110 20460 23166 20496
rect 23110 20440 23112 20460
rect 23112 20440 23164 20460
rect 23164 20440 23166 20460
rect 23484 19610 23540 19612
rect 23564 19610 23620 19612
rect 23644 19610 23700 19612
rect 23724 19610 23780 19612
rect 23484 19558 23530 19610
rect 23530 19558 23540 19610
rect 23564 19558 23594 19610
rect 23594 19558 23606 19610
rect 23606 19558 23620 19610
rect 23644 19558 23658 19610
rect 23658 19558 23670 19610
rect 23670 19558 23700 19610
rect 23724 19558 23734 19610
rect 23734 19558 23780 19610
rect 23484 19556 23540 19558
rect 23564 19556 23620 19558
rect 23644 19556 23700 19558
rect 23724 19556 23780 19558
rect 23938 19352 23994 19408
rect 23484 18522 23540 18524
rect 23564 18522 23620 18524
rect 23644 18522 23700 18524
rect 23724 18522 23780 18524
rect 23484 18470 23530 18522
rect 23530 18470 23540 18522
rect 23564 18470 23594 18522
rect 23594 18470 23606 18522
rect 23606 18470 23620 18522
rect 23644 18470 23658 18522
rect 23658 18470 23670 18522
rect 23670 18470 23700 18522
rect 23724 18470 23734 18522
rect 23734 18470 23780 18522
rect 23484 18468 23540 18470
rect 23564 18468 23620 18470
rect 23644 18468 23700 18470
rect 23724 18468 23780 18470
rect 23484 17434 23540 17436
rect 23564 17434 23620 17436
rect 23644 17434 23700 17436
rect 23724 17434 23780 17436
rect 23484 17382 23530 17434
rect 23530 17382 23540 17434
rect 23564 17382 23594 17434
rect 23594 17382 23606 17434
rect 23606 17382 23620 17434
rect 23644 17382 23658 17434
rect 23658 17382 23670 17434
rect 23670 17382 23700 17434
rect 23724 17382 23734 17434
rect 23734 17382 23780 17434
rect 23484 17380 23540 17382
rect 23564 17380 23620 17382
rect 23644 17380 23700 17382
rect 23724 17380 23780 17382
rect 23294 17176 23350 17232
rect 23484 16346 23540 16348
rect 23564 16346 23620 16348
rect 23644 16346 23700 16348
rect 23724 16346 23780 16348
rect 23484 16294 23530 16346
rect 23530 16294 23540 16346
rect 23564 16294 23594 16346
rect 23594 16294 23606 16346
rect 23606 16294 23620 16346
rect 23644 16294 23658 16346
rect 23658 16294 23670 16346
rect 23670 16294 23700 16346
rect 23724 16294 23734 16346
rect 23734 16294 23780 16346
rect 23484 16292 23540 16294
rect 23564 16292 23620 16294
rect 23644 16292 23700 16294
rect 23724 16292 23780 16294
rect 23484 15258 23540 15260
rect 23564 15258 23620 15260
rect 23644 15258 23700 15260
rect 23724 15258 23780 15260
rect 23484 15206 23530 15258
rect 23530 15206 23540 15258
rect 23564 15206 23594 15258
rect 23594 15206 23606 15258
rect 23606 15206 23620 15258
rect 23644 15206 23658 15258
rect 23658 15206 23670 15258
rect 23670 15206 23700 15258
rect 23724 15206 23734 15258
rect 23734 15206 23780 15258
rect 23484 15204 23540 15206
rect 23564 15204 23620 15206
rect 23644 15204 23700 15206
rect 23724 15204 23780 15206
rect 23484 14170 23540 14172
rect 23564 14170 23620 14172
rect 23644 14170 23700 14172
rect 23724 14170 23780 14172
rect 23484 14118 23530 14170
rect 23530 14118 23540 14170
rect 23564 14118 23594 14170
rect 23594 14118 23606 14170
rect 23606 14118 23620 14170
rect 23644 14118 23658 14170
rect 23658 14118 23670 14170
rect 23670 14118 23700 14170
rect 23724 14118 23734 14170
rect 23734 14118 23780 14170
rect 23484 14116 23540 14118
rect 23564 14116 23620 14118
rect 23644 14116 23700 14118
rect 23724 14116 23780 14118
rect 23484 13082 23540 13084
rect 23564 13082 23620 13084
rect 23644 13082 23700 13084
rect 23724 13082 23780 13084
rect 23484 13030 23530 13082
rect 23530 13030 23540 13082
rect 23564 13030 23594 13082
rect 23594 13030 23606 13082
rect 23606 13030 23620 13082
rect 23644 13030 23658 13082
rect 23658 13030 23670 13082
rect 23670 13030 23700 13082
rect 23724 13030 23734 13082
rect 23734 13030 23780 13082
rect 23484 13028 23540 13030
rect 23564 13028 23620 13030
rect 23644 13028 23700 13030
rect 23724 13028 23780 13030
rect 23484 11994 23540 11996
rect 23564 11994 23620 11996
rect 23644 11994 23700 11996
rect 23724 11994 23780 11996
rect 23484 11942 23530 11994
rect 23530 11942 23540 11994
rect 23564 11942 23594 11994
rect 23594 11942 23606 11994
rect 23606 11942 23620 11994
rect 23644 11942 23658 11994
rect 23658 11942 23670 11994
rect 23670 11942 23700 11994
rect 23724 11942 23734 11994
rect 23734 11942 23780 11994
rect 23484 11940 23540 11942
rect 23564 11940 23620 11942
rect 23644 11940 23700 11942
rect 23724 11940 23780 11942
rect 23484 10906 23540 10908
rect 23564 10906 23620 10908
rect 23644 10906 23700 10908
rect 23724 10906 23780 10908
rect 23484 10854 23530 10906
rect 23530 10854 23540 10906
rect 23564 10854 23594 10906
rect 23594 10854 23606 10906
rect 23606 10854 23620 10906
rect 23644 10854 23658 10906
rect 23658 10854 23670 10906
rect 23670 10854 23700 10906
rect 23724 10854 23734 10906
rect 23734 10854 23780 10906
rect 23484 10852 23540 10854
rect 23564 10852 23620 10854
rect 23644 10852 23700 10854
rect 23724 10852 23780 10854
rect 23484 9818 23540 9820
rect 23564 9818 23620 9820
rect 23644 9818 23700 9820
rect 23724 9818 23780 9820
rect 23484 9766 23530 9818
rect 23530 9766 23540 9818
rect 23564 9766 23594 9818
rect 23594 9766 23606 9818
rect 23606 9766 23620 9818
rect 23644 9766 23658 9818
rect 23658 9766 23670 9818
rect 23670 9766 23700 9818
rect 23724 9766 23734 9818
rect 23734 9766 23780 9818
rect 23484 9764 23540 9766
rect 23564 9764 23620 9766
rect 23644 9764 23700 9766
rect 23724 9764 23780 9766
rect 23484 8730 23540 8732
rect 23564 8730 23620 8732
rect 23644 8730 23700 8732
rect 23724 8730 23780 8732
rect 23484 8678 23530 8730
rect 23530 8678 23540 8730
rect 23564 8678 23594 8730
rect 23594 8678 23606 8730
rect 23606 8678 23620 8730
rect 23644 8678 23658 8730
rect 23658 8678 23670 8730
rect 23670 8678 23700 8730
rect 23724 8678 23734 8730
rect 23734 8678 23780 8730
rect 23484 8676 23540 8678
rect 23564 8676 23620 8678
rect 23644 8676 23700 8678
rect 23724 8676 23780 8678
rect 23484 7642 23540 7644
rect 23564 7642 23620 7644
rect 23644 7642 23700 7644
rect 23724 7642 23780 7644
rect 23484 7590 23530 7642
rect 23530 7590 23540 7642
rect 23564 7590 23594 7642
rect 23594 7590 23606 7642
rect 23606 7590 23620 7642
rect 23644 7590 23658 7642
rect 23658 7590 23670 7642
rect 23670 7590 23700 7642
rect 23724 7590 23734 7642
rect 23734 7590 23780 7642
rect 23484 7588 23540 7590
rect 23564 7588 23620 7590
rect 23644 7588 23700 7590
rect 23724 7588 23780 7590
rect 23484 6554 23540 6556
rect 23564 6554 23620 6556
rect 23644 6554 23700 6556
rect 23724 6554 23780 6556
rect 23484 6502 23530 6554
rect 23530 6502 23540 6554
rect 23564 6502 23594 6554
rect 23594 6502 23606 6554
rect 23606 6502 23620 6554
rect 23644 6502 23658 6554
rect 23658 6502 23670 6554
rect 23670 6502 23700 6554
rect 23724 6502 23734 6554
rect 23734 6502 23780 6554
rect 23484 6500 23540 6502
rect 23564 6500 23620 6502
rect 23644 6500 23700 6502
rect 23724 6500 23780 6502
rect 24122 31592 24178 31648
rect 24122 29824 24178 29880
rect 24398 30540 24400 30560
rect 24400 30540 24452 30560
rect 24452 30540 24454 30560
rect 24398 30504 24454 30540
rect 24306 27784 24362 27840
rect 26882 39888 26938 39944
rect 26514 39636 26570 39672
rect 26514 39616 26516 39636
rect 26516 39616 26568 39636
rect 26568 39616 26570 39636
rect 25318 35672 25374 35728
rect 25502 34176 25558 34232
rect 25226 32816 25282 32872
rect 25318 32544 25374 32600
rect 24950 32136 25006 32192
rect 26882 38936 26938 38992
rect 26974 38664 27030 38720
rect 26238 35692 26294 35728
rect 26238 35672 26240 35692
rect 26240 35672 26292 35692
rect 26292 35672 26294 35692
rect 26238 35264 26294 35320
rect 26054 34040 26110 34096
rect 25962 33224 26018 33280
rect 26146 33224 26202 33280
rect 25410 31456 25466 31512
rect 24950 28736 25006 28792
rect 24306 27376 24362 27432
rect 24214 25472 24270 25528
rect 24674 24384 24730 24440
rect 24214 23024 24270 23080
rect 24122 20340 24124 20360
rect 24124 20340 24176 20360
rect 24176 20340 24178 20360
rect 24122 20304 24178 20340
rect 24582 22480 24638 22536
rect 24306 21548 24362 21584
rect 24306 21528 24308 21548
rect 24308 21528 24360 21548
rect 24360 21528 24362 21548
rect 25686 31048 25742 31104
rect 25318 27648 25374 27704
rect 25318 25336 25374 25392
rect 26330 32000 26386 32056
rect 25778 30096 25834 30152
rect 26054 30640 26110 30696
rect 26238 31456 26294 31512
rect 27710 38836 27712 38856
rect 27712 38836 27764 38856
rect 27764 38836 27766 38856
rect 27710 38800 27766 38836
rect 28262 38528 28318 38584
rect 27710 38392 27766 38448
rect 27342 33496 27398 33552
rect 26330 29688 26386 29744
rect 26330 28464 26386 28520
rect 26606 28464 26662 28520
rect 25502 26560 25558 26616
rect 25502 25492 25558 25528
rect 25502 25472 25504 25492
rect 25504 25472 25556 25492
rect 25556 25472 25558 25492
rect 25962 27648 26018 27704
rect 26606 27784 26662 27840
rect 27158 31592 27214 31648
rect 26882 29688 26938 29744
rect 26882 29572 26938 29608
rect 26882 29552 26884 29572
rect 26884 29552 26936 29572
rect 26936 29552 26938 29572
rect 27066 29688 27122 29744
rect 28170 36660 28172 36680
rect 28172 36660 28224 36680
rect 28224 36660 28226 36680
rect 28170 36624 28226 36660
rect 27894 36080 27950 36136
rect 28630 38528 28686 38584
rect 28538 38392 28594 38448
rect 29116 39738 29172 39740
rect 29196 39738 29252 39740
rect 29276 39738 29332 39740
rect 29356 39738 29412 39740
rect 29116 39686 29162 39738
rect 29162 39686 29172 39738
rect 29196 39686 29226 39738
rect 29226 39686 29238 39738
rect 29238 39686 29252 39738
rect 29276 39686 29290 39738
rect 29290 39686 29302 39738
rect 29302 39686 29332 39738
rect 29356 39686 29366 39738
rect 29366 39686 29412 39738
rect 29116 39684 29172 39686
rect 29196 39684 29252 39686
rect 29276 39684 29332 39686
rect 29356 39684 29412 39686
rect 29116 38650 29172 38652
rect 29196 38650 29252 38652
rect 29276 38650 29332 38652
rect 29356 38650 29412 38652
rect 29116 38598 29162 38650
rect 29162 38598 29172 38650
rect 29196 38598 29226 38650
rect 29226 38598 29238 38650
rect 29238 38598 29252 38650
rect 29276 38598 29290 38650
rect 29290 38598 29302 38650
rect 29302 38598 29332 38650
rect 29356 38598 29366 38650
rect 29366 38598 29412 38650
rect 29116 38596 29172 38598
rect 29196 38596 29252 38598
rect 29276 38596 29332 38598
rect 29356 38596 29412 38598
rect 29116 37562 29172 37564
rect 29196 37562 29252 37564
rect 29276 37562 29332 37564
rect 29356 37562 29412 37564
rect 29116 37510 29162 37562
rect 29162 37510 29172 37562
rect 29196 37510 29226 37562
rect 29226 37510 29238 37562
rect 29238 37510 29252 37562
rect 29276 37510 29290 37562
rect 29290 37510 29302 37562
rect 29302 37510 29332 37562
rect 29356 37510 29366 37562
rect 29366 37510 29412 37562
rect 29116 37508 29172 37510
rect 29196 37508 29252 37510
rect 29276 37508 29332 37510
rect 29356 37508 29412 37510
rect 27802 33496 27858 33552
rect 27894 32680 27950 32736
rect 28078 32136 28134 32192
rect 28078 31764 28080 31784
rect 28080 31764 28132 31784
rect 28132 31764 28134 31784
rect 28078 31728 28134 31764
rect 27986 31048 28042 31104
rect 27802 29960 27858 30016
rect 27526 27920 27582 27976
rect 27342 27512 27398 27568
rect 26974 27396 27030 27432
rect 26974 27376 26976 27396
rect 26976 27376 27028 27396
rect 27028 27376 27030 27396
rect 25226 23296 25282 23352
rect 24766 21800 24822 21856
rect 24582 20984 24638 21040
rect 24950 22344 25006 22400
rect 24766 20848 24822 20904
rect 25134 21936 25190 21992
rect 25502 22636 25558 22672
rect 25502 22616 25504 22636
rect 25504 22616 25556 22636
rect 25556 22616 25558 22636
rect 25410 22072 25466 22128
rect 25410 21936 25466 21992
rect 25318 21120 25374 21176
rect 25594 21936 25650 21992
rect 25962 22344 26018 22400
rect 25778 21548 25834 21584
rect 25778 21528 25780 21548
rect 25780 21528 25832 21548
rect 25832 21528 25834 21548
rect 27250 26968 27306 27024
rect 26790 23704 26846 23760
rect 25686 20712 25742 20768
rect 25410 17196 25466 17232
rect 26238 21664 26294 21720
rect 25962 20460 26018 20496
rect 27250 22616 27306 22672
rect 27342 22516 27344 22536
rect 27344 22516 27396 22536
rect 27396 22516 27398 22536
rect 27066 22208 27122 22264
rect 27342 22480 27398 22516
rect 27066 21936 27122 21992
rect 26974 20712 27030 20768
rect 25962 20440 25964 20460
rect 25964 20440 26016 20460
rect 26016 20440 26018 20460
rect 26422 19624 26478 19680
rect 25410 17176 25412 17196
rect 25412 17176 25464 17196
rect 25464 17176 25466 17196
rect 23484 5466 23540 5468
rect 23564 5466 23620 5468
rect 23644 5466 23700 5468
rect 23724 5466 23780 5468
rect 23484 5414 23530 5466
rect 23530 5414 23540 5466
rect 23564 5414 23594 5466
rect 23594 5414 23606 5466
rect 23606 5414 23620 5466
rect 23644 5414 23658 5466
rect 23658 5414 23670 5466
rect 23670 5414 23700 5466
rect 23724 5414 23734 5466
rect 23734 5414 23780 5466
rect 23484 5412 23540 5414
rect 23564 5412 23620 5414
rect 23644 5412 23700 5414
rect 23724 5412 23780 5414
rect 27802 27920 27858 27976
rect 29116 36474 29172 36476
rect 29196 36474 29252 36476
rect 29276 36474 29332 36476
rect 29356 36474 29412 36476
rect 29116 36422 29162 36474
rect 29162 36422 29172 36474
rect 29196 36422 29226 36474
rect 29226 36422 29238 36474
rect 29238 36422 29252 36474
rect 29276 36422 29290 36474
rect 29290 36422 29302 36474
rect 29302 36422 29332 36474
rect 29356 36422 29366 36474
rect 29366 36422 29412 36474
rect 29116 36420 29172 36422
rect 29196 36420 29252 36422
rect 29276 36420 29332 36422
rect 29356 36420 29412 36422
rect 29550 37712 29606 37768
rect 29734 37304 29790 37360
rect 29458 35672 29514 35728
rect 28906 35400 28962 35456
rect 29116 35386 29172 35388
rect 29196 35386 29252 35388
rect 29276 35386 29332 35388
rect 29356 35386 29412 35388
rect 29116 35334 29162 35386
rect 29162 35334 29172 35386
rect 29196 35334 29226 35386
rect 29226 35334 29238 35386
rect 29238 35334 29252 35386
rect 29276 35334 29290 35386
rect 29290 35334 29302 35386
rect 29302 35334 29332 35386
rect 29356 35334 29366 35386
rect 29366 35334 29412 35386
rect 29116 35332 29172 35334
rect 29196 35332 29252 35334
rect 29276 35332 29332 35334
rect 29356 35332 29412 35334
rect 29366 34720 29422 34776
rect 28722 33224 28778 33280
rect 28630 33088 28686 33144
rect 29116 34298 29172 34300
rect 29196 34298 29252 34300
rect 29276 34298 29332 34300
rect 29356 34298 29412 34300
rect 29116 34246 29162 34298
rect 29162 34246 29172 34298
rect 29196 34246 29226 34298
rect 29226 34246 29238 34298
rect 29238 34246 29252 34298
rect 29276 34246 29290 34298
rect 29290 34246 29302 34298
rect 29302 34246 29332 34298
rect 29356 34246 29366 34298
rect 29366 34246 29412 34298
rect 29116 34244 29172 34246
rect 29196 34244 29252 34246
rect 29276 34244 29332 34246
rect 29356 34244 29412 34246
rect 29274 34040 29330 34096
rect 29458 33516 29514 33552
rect 29458 33496 29460 33516
rect 29460 33496 29512 33516
rect 29512 33496 29514 33516
rect 29116 33210 29172 33212
rect 29196 33210 29252 33212
rect 29276 33210 29332 33212
rect 29356 33210 29412 33212
rect 29116 33158 29162 33210
rect 29162 33158 29172 33210
rect 29196 33158 29226 33210
rect 29226 33158 29238 33210
rect 29238 33158 29252 33210
rect 29276 33158 29290 33210
rect 29290 33158 29302 33210
rect 29302 33158 29332 33210
rect 29356 33158 29366 33210
rect 29366 33158 29412 33210
rect 29116 33156 29172 33158
rect 29196 33156 29252 33158
rect 29276 33156 29332 33158
rect 29356 33156 29412 33158
rect 28814 32136 28870 32192
rect 28446 31184 28502 31240
rect 28354 30504 28410 30560
rect 28262 28464 28318 28520
rect 28538 30796 28594 30832
rect 28538 30776 28540 30796
rect 28540 30776 28592 30796
rect 28592 30776 28594 30796
rect 28722 30912 28778 30968
rect 29116 32122 29172 32124
rect 29196 32122 29252 32124
rect 29276 32122 29332 32124
rect 29356 32122 29412 32124
rect 29116 32070 29162 32122
rect 29162 32070 29172 32122
rect 29196 32070 29226 32122
rect 29226 32070 29238 32122
rect 29238 32070 29252 32122
rect 29276 32070 29290 32122
rect 29290 32070 29302 32122
rect 29302 32070 29332 32122
rect 29356 32070 29366 32122
rect 29366 32070 29412 32122
rect 29116 32068 29172 32070
rect 29196 32068 29252 32070
rect 29276 32068 29332 32070
rect 29356 32068 29412 32070
rect 29550 32000 29606 32056
rect 29366 31864 29422 31920
rect 29274 31592 29330 31648
rect 29116 31034 29172 31036
rect 29196 31034 29252 31036
rect 29276 31034 29332 31036
rect 29356 31034 29412 31036
rect 29116 30982 29162 31034
rect 29162 30982 29172 31034
rect 29196 30982 29226 31034
rect 29226 30982 29238 31034
rect 29238 30982 29252 31034
rect 29276 30982 29290 31034
rect 29290 30982 29302 31034
rect 29302 30982 29332 31034
rect 29356 30982 29366 31034
rect 29366 30982 29412 31034
rect 29116 30980 29172 30982
rect 29196 30980 29252 30982
rect 29276 30980 29332 30982
rect 29356 30980 29412 30982
rect 28446 29960 28502 30016
rect 28538 29824 28594 29880
rect 28446 29416 28502 29472
rect 28446 29144 28502 29200
rect 28446 27376 28502 27432
rect 28446 27276 28448 27296
rect 28448 27276 28500 27296
rect 28500 27276 28502 27296
rect 28446 27240 28502 27276
rect 28906 29960 28962 30016
rect 29116 29946 29172 29948
rect 29196 29946 29252 29948
rect 29276 29946 29332 29948
rect 29356 29946 29412 29948
rect 29116 29894 29162 29946
rect 29162 29894 29172 29946
rect 29196 29894 29226 29946
rect 29226 29894 29238 29946
rect 29238 29894 29252 29946
rect 29276 29894 29290 29946
rect 29290 29894 29302 29946
rect 29302 29894 29332 29946
rect 29356 29894 29366 29946
rect 29366 29894 29412 29946
rect 29116 29892 29172 29894
rect 29196 29892 29252 29894
rect 29276 29892 29332 29894
rect 29356 29892 29412 29894
rect 29366 29588 29368 29608
rect 29368 29588 29420 29608
rect 29420 29588 29422 29608
rect 29366 29552 29422 29588
rect 29274 29280 29330 29336
rect 28814 28872 28870 28928
rect 29116 28858 29172 28860
rect 29196 28858 29252 28860
rect 29276 28858 29332 28860
rect 29356 28858 29412 28860
rect 29116 28806 29162 28858
rect 29162 28806 29172 28858
rect 29196 28806 29226 28858
rect 29226 28806 29238 28858
rect 29238 28806 29252 28858
rect 29276 28806 29290 28858
rect 29290 28806 29302 28858
rect 29302 28806 29332 28858
rect 29356 28806 29366 28858
rect 29366 28806 29412 28858
rect 29116 28804 29172 28806
rect 29196 28804 29252 28806
rect 29276 28804 29332 28806
rect 29356 28804 29412 28806
rect 29918 34856 29974 34912
rect 31390 39888 31446 39944
rect 29734 32816 29790 32872
rect 29918 32816 29974 32872
rect 29734 30912 29790 30968
rect 29642 29960 29698 30016
rect 29550 28872 29606 28928
rect 29734 29416 29790 29472
rect 29642 28736 29698 28792
rect 28630 26696 28686 26752
rect 28078 25200 28134 25256
rect 27710 24248 27766 24304
rect 27894 21392 27950 21448
rect 28354 23976 28410 24032
rect 28262 22616 28318 22672
rect 28262 21800 28318 21856
rect 28078 21256 28134 21312
rect 28446 23160 28502 23216
rect 28446 21392 28502 21448
rect 27986 19624 28042 19680
rect 28722 23976 28778 24032
rect 28722 23568 28778 23624
rect 28630 19760 28686 19816
rect 29116 27770 29172 27772
rect 29196 27770 29252 27772
rect 29276 27770 29332 27772
rect 29356 27770 29412 27772
rect 29116 27718 29162 27770
rect 29162 27718 29172 27770
rect 29196 27718 29226 27770
rect 29226 27718 29238 27770
rect 29238 27718 29252 27770
rect 29276 27718 29290 27770
rect 29290 27718 29302 27770
rect 29302 27718 29332 27770
rect 29356 27718 29366 27770
rect 29366 27718 29412 27770
rect 29116 27716 29172 27718
rect 29196 27716 29252 27718
rect 29276 27716 29332 27718
rect 29356 27716 29412 27718
rect 29550 28192 29606 28248
rect 29550 26832 29606 26888
rect 29116 26682 29172 26684
rect 29196 26682 29252 26684
rect 29276 26682 29332 26684
rect 29356 26682 29412 26684
rect 29116 26630 29162 26682
rect 29162 26630 29172 26682
rect 29196 26630 29226 26682
rect 29226 26630 29238 26682
rect 29238 26630 29252 26682
rect 29276 26630 29290 26682
rect 29290 26630 29302 26682
rect 29302 26630 29332 26682
rect 29356 26630 29366 26682
rect 29366 26630 29412 26682
rect 29116 26628 29172 26630
rect 29196 26628 29252 26630
rect 29276 26628 29332 26630
rect 29356 26628 29412 26630
rect 29116 25594 29172 25596
rect 29196 25594 29252 25596
rect 29276 25594 29332 25596
rect 29356 25594 29412 25596
rect 29116 25542 29162 25594
rect 29162 25542 29172 25594
rect 29196 25542 29226 25594
rect 29226 25542 29238 25594
rect 29238 25542 29252 25594
rect 29276 25542 29290 25594
rect 29290 25542 29302 25594
rect 29302 25542 29332 25594
rect 29356 25542 29366 25594
rect 29366 25542 29412 25594
rect 29116 25540 29172 25542
rect 29196 25540 29252 25542
rect 29276 25540 29332 25542
rect 29356 25540 29412 25542
rect 29458 24656 29514 24712
rect 29734 24556 29736 24576
rect 29736 24556 29788 24576
rect 29788 24556 29790 24576
rect 29734 24520 29790 24556
rect 29116 24506 29172 24508
rect 29196 24506 29252 24508
rect 29276 24506 29332 24508
rect 29356 24506 29412 24508
rect 29116 24454 29162 24506
rect 29162 24454 29172 24506
rect 29196 24454 29226 24506
rect 29226 24454 29238 24506
rect 29238 24454 29252 24506
rect 29276 24454 29290 24506
rect 29290 24454 29302 24506
rect 29302 24454 29332 24506
rect 29356 24454 29366 24506
rect 29366 24454 29412 24506
rect 29116 24452 29172 24454
rect 29196 24452 29252 24454
rect 29276 24452 29332 24454
rect 29356 24452 29412 24454
rect 28998 23568 29054 23624
rect 29116 23418 29172 23420
rect 29196 23418 29252 23420
rect 29276 23418 29332 23420
rect 29356 23418 29412 23420
rect 29116 23366 29162 23418
rect 29162 23366 29172 23418
rect 29196 23366 29226 23418
rect 29226 23366 29238 23418
rect 29238 23366 29252 23418
rect 29276 23366 29290 23418
rect 29290 23366 29302 23418
rect 29302 23366 29332 23418
rect 29356 23366 29366 23418
rect 29366 23366 29412 23418
rect 29116 23364 29172 23366
rect 29196 23364 29252 23366
rect 29276 23364 29332 23366
rect 29356 23364 29412 23366
rect 28906 23180 28962 23216
rect 28906 23160 28908 23180
rect 28908 23160 28960 23180
rect 28960 23160 28962 23180
rect 29116 22330 29172 22332
rect 29196 22330 29252 22332
rect 29276 22330 29332 22332
rect 29356 22330 29412 22332
rect 29116 22278 29162 22330
rect 29162 22278 29172 22330
rect 29196 22278 29226 22330
rect 29226 22278 29238 22330
rect 29238 22278 29252 22330
rect 29276 22278 29290 22330
rect 29290 22278 29302 22330
rect 29302 22278 29332 22330
rect 29356 22278 29366 22330
rect 29366 22278 29412 22330
rect 29116 22276 29172 22278
rect 29196 22276 29252 22278
rect 29276 22276 29332 22278
rect 29356 22276 29412 22278
rect 29182 21800 29238 21856
rect 29274 21528 29330 21584
rect 29116 21242 29172 21244
rect 29196 21242 29252 21244
rect 29276 21242 29332 21244
rect 29356 21242 29412 21244
rect 29116 21190 29162 21242
rect 29162 21190 29172 21242
rect 29196 21190 29226 21242
rect 29226 21190 29238 21242
rect 29238 21190 29252 21242
rect 29276 21190 29290 21242
rect 29290 21190 29302 21242
rect 29302 21190 29332 21242
rect 29356 21190 29366 21242
rect 29366 21190 29412 21242
rect 29116 21188 29172 21190
rect 29196 21188 29252 21190
rect 29276 21188 29332 21190
rect 29356 21188 29412 21190
rect 29116 20154 29172 20156
rect 29196 20154 29252 20156
rect 29276 20154 29332 20156
rect 29356 20154 29412 20156
rect 29116 20102 29162 20154
rect 29162 20102 29172 20154
rect 29196 20102 29226 20154
rect 29226 20102 29238 20154
rect 29238 20102 29252 20154
rect 29276 20102 29290 20154
rect 29290 20102 29302 20154
rect 29302 20102 29332 20154
rect 29356 20102 29366 20154
rect 29366 20102 29412 20154
rect 29116 20100 29172 20102
rect 29196 20100 29252 20102
rect 29276 20100 29332 20102
rect 29356 20100 29412 20102
rect 29550 19760 29606 19816
rect 29274 19508 29330 19544
rect 29274 19488 29276 19508
rect 29276 19488 29328 19508
rect 29328 19488 29330 19508
rect 29458 19624 29514 19680
rect 29116 19066 29172 19068
rect 29196 19066 29252 19068
rect 29276 19066 29332 19068
rect 29356 19066 29412 19068
rect 29116 19014 29162 19066
rect 29162 19014 29172 19066
rect 29196 19014 29226 19066
rect 29226 19014 29238 19066
rect 29238 19014 29252 19066
rect 29276 19014 29290 19066
rect 29290 19014 29302 19066
rect 29302 19014 29332 19066
rect 29356 19014 29366 19066
rect 29366 19014 29412 19066
rect 29116 19012 29172 19014
rect 29196 19012 29252 19014
rect 29276 19012 29332 19014
rect 29356 19012 29412 19014
rect 29116 17978 29172 17980
rect 29196 17978 29252 17980
rect 29276 17978 29332 17980
rect 29356 17978 29412 17980
rect 29116 17926 29162 17978
rect 29162 17926 29172 17978
rect 29196 17926 29226 17978
rect 29226 17926 29238 17978
rect 29238 17926 29252 17978
rect 29276 17926 29290 17978
rect 29290 17926 29302 17978
rect 29302 17926 29332 17978
rect 29356 17926 29366 17978
rect 29366 17926 29412 17978
rect 29116 17924 29172 17926
rect 29196 17924 29252 17926
rect 29276 17924 29332 17926
rect 29356 17924 29412 17926
rect 29550 19352 29606 19408
rect 29116 16890 29172 16892
rect 29196 16890 29252 16892
rect 29276 16890 29332 16892
rect 29356 16890 29412 16892
rect 29116 16838 29162 16890
rect 29162 16838 29172 16890
rect 29196 16838 29226 16890
rect 29226 16838 29238 16890
rect 29238 16838 29252 16890
rect 29276 16838 29290 16890
rect 29290 16838 29302 16890
rect 29302 16838 29332 16890
rect 29356 16838 29366 16890
rect 29366 16838 29412 16890
rect 29116 16836 29172 16838
rect 29196 16836 29252 16838
rect 29276 16836 29332 16838
rect 29356 16836 29412 16838
rect 29116 15802 29172 15804
rect 29196 15802 29252 15804
rect 29276 15802 29332 15804
rect 29356 15802 29412 15804
rect 29116 15750 29162 15802
rect 29162 15750 29172 15802
rect 29196 15750 29226 15802
rect 29226 15750 29238 15802
rect 29238 15750 29252 15802
rect 29276 15750 29290 15802
rect 29290 15750 29302 15802
rect 29302 15750 29332 15802
rect 29356 15750 29366 15802
rect 29366 15750 29412 15802
rect 29116 15748 29172 15750
rect 29196 15748 29252 15750
rect 29276 15748 29332 15750
rect 29356 15748 29412 15750
rect 29116 14714 29172 14716
rect 29196 14714 29252 14716
rect 29276 14714 29332 14716
rect 29356 14714 29412 14716
rect 29116 14662 29162 14714
rect 29162 14662 29172 14714
rect 29196 14662 29226 14714
rect 29226 14662 29238 14714
rect 29238 14662 29252 14714
rect 29276 14662 29290 14714
rect 29290 14662 29302 14714
rect 29302 14662 29332 14714
rect 29356 14662 29366 14714
rect 29366 14662 29412 14714
rect 29116 14660 29172 14662
rect 29196 14660 29252 14662
rect 29276 14660 29332 14662
rect 29356 14660 29412 14662
rect 29116 13626 29172 13628
rect 29196 13626 29252 13628
rect 29276 13626 29332 13628
rect 29356 13626 29412 13628
rect 29116 13574 29162 13626
rect 29162 13574 29172 13626
rect 29196 13574 29226 13626
rect 29226 13574 29238 13626
rect 29238 13574 29252 13626
rect 29276 13574 29290 13626
rect 29290 13574 29302 13626
rect 29302 13574 29332 13626
rect 29356 13574 29366 13626
rect 29366 13574 29412 13626
rect 29116 13572 29172 13574
rect 29196 13572 29252 13574
rect 29276 13572 29332 13574
rect 29356 13572 29412 13574
rect 29116 12538 29172 12540
rect 29196 12538 29252 12540
rect 29276 12538 29332 12540
rect 29356 12538 29412 12540
rect 29116 12486 29162 12538
rect 29162 12486 29172 12538
rect 29196 12486 29226 12538
rect 29226 12486 29238 12538
rect 29238 12486 29252 12538
rect 29276 12486 29290 12538
rect 29290 12486 29302 12538
rect 29302 12486 29332 12538
rect 29356 12486 29366 12538
rect 29366 12486 29412 12538
rect 29116 12484 29172 12486
rect 29196 12484 29252 12486
rect 29276 12484 29332 12486
rect 29356 12484 29412 12486
rect 29116 11450 29172 11452
rect 29196 11450 29252 11452
rect 29276 11450 29332 11452
rect 29356 11450 29412 11452
rect 29116 11398 29162 11450
rect 29162 11398 29172 11450
rect 29196 11398 29226 11450
rect 29226 11398 29238 11450
rect 29238 11398 29252 11450
rect 29276 11398 29290 11450
rect 29290 11398 29302 11450
rect 29302 11398 29332 11450
rect 29356 11398 29366 11450
rect 29366 11398 29412 11450
rect 29116 11396 29172 11398
rect 29196 11396 29252 11398
rect 29276 11396 29332 11398
rect 29356 11396 29412 11398
rect 29116 10362 29172 10364
rect 29196 10362 29252 10364
rect 29276 10362 29332 10364
rect 29356 10362 29412 10364
rect 29116 10310 29162 10362
rect 29162 10310 29172 10362
rect 29196 10310 29226 10362
rect 29226 10310 29238 10362
rect 29238 10310 29252 10362
rect 29276 10310 29290 10362
rect 29290 10310 29302 10362
rect 29302 10310 29332 10362
rect 29356 10310 29366 10362
rect 29366 10310 29412 10362
rect 29116 10308 29172 10310
rect 29196 10308 29252 10310
rect 29276 10308 29332 10310
rect 29356 10308 29412 10310
rect 29116 9274 29172 9276
rect 29196 9274 29252 9276
rect 29276 9274 29332 9276
rect 29356 9274 29412 9276
rect 29116 9222 29162 9274
rect 29162 9222 29172 9274
rect 29196 9222 29226 9274
rect 29226 9222 29238 9274
rect 29238 9222 29252 9274
rect 29276 9222 29290 9274
rect 29290 9222 29302 9274
rect 29302 9222 29332 9274
rect 29356 9222 29366 9274
rect 29366 9222 29412 9274
rect 29116 9220 29172 9222
rect 29196 9220 29252 9222
rect 29276 9220 29332 9222
rect 29356 9220 29412 9222
rect 29116 8186 29172 8188
rect 29196 8186 29252 8188
rect 29276 8186 29332 8188
rect 29356 8186 29412 8188
rect 29116 8134 29162 8186
rect 29162 8134 29172 8186
rect 29196 8134 29226 8186
rect 29226 8134 29238 8186
rect 29238 8134 29252 8186
rect 29276 8134 29290 8186
rect 29290 8134 29302 8186
rect 29302 8134 29332 8186
rect 29356 8134 29366 8186
rect 29366 8134 29412 8186
rect 29116 8132 29172 8134
rect 29196 8132 29252 8134
rect 29276 8132 29332 8134
rect 29356 8132 29412 8134
rect 29116 7098 29172 7100
rect 29196 7098 29252 7100
rect 29276 7098 29332 7100
rect 29356 7098 29412 7100
rect 29116 7046 29162 7098
rect 29162 7046 29172 7098
rect 29196 7046 29226 7098
rect 29226 7046 29238 7098
rect 29238 7046 29252 7098
rect 29276 7046 29290 7098
rect 29290 7046 29302 7098
rect 29302 7046 29332 7098
rect 29356 7046 29366 7098
rect 29366 7046 29412 7098
rect 29116 7044 29172 7046
rect 29196 7044 29252 7046
rect 29276 7044 29332 7046
rect 29356 7044 29412 7046
rect 29116 6010 29172 6012
rect 29196 6010 29252 6012
rect 29276 6010 29332 6012
rect 29356 6010 29412 6012
rect 29116 5958 29162 6010
rect 29162 5958 29172 6010
rect 29196 5958 29226 6010
rect 29226 5958 29238 6010
rect 29238 5958 29252 6010
rect 29276 5958 29290 6010
rect 29290 5958 29302 6010
rect 29302 5958 29332 6010
rect 29356 5958 29366 6010
rect 29366 5958 29412 6010
rect 29116 5956 29172 5958
rect 29196 5956 29252 5958
rect 29276 5956 29332 5958
rect 29356 5956 29412 5958
rect 29116 4922 29172 4924
rect 29196 4922 29252 4924
rect 29276 4922 29332 4924
rect 29356 4922 29412 4924
rect 29116 4870 29162 4922
rect 29162 4870 29172 4922
rect 29196 4870 29226 4922
rect 29226 4870 29238 4922
rect 29238 4870 29252 4922
rect 29276 4870 29290 4922
rect 29290 4870 29302 4922
rect 29302 4870 29332 4922
rect 29356 4870 29366 4922
rect 29366 4870 29412 4922
rect 29116 4868 29172 4870
rect 29196 4868 29252 4870
rect 29276 4868 29332 4870
rect 29356 4868 29412 4870
rect 23484 4378 23540 4380
rect 23564 4378 23620 4380
rect 23644 4378 23700 4380
rect 23724 4378 23780 4380
rect 23484 4326 23530 4378
rect 23530 4326 23540 4378
rect 23564 4326 23594 4378
rect 23594 4326 23606 4378
rect 23606 4326 23620 4378
rect 23644 4326 23658 4378
rect 23658 4326 23670 4378
rect 23670 4326 23700 4378
rect 23724 4326 23734 4378
rect 23734 4326 23780 4378
rect 23484 4324 23540 4326
rect 23564 4324 23620 4326
rect 23644 4324 23700 4326
rect 23724 4324 23780 4326
rect 17852 2746 17908 2748
rect 17932 2746 17988 2748
rect 18012 2746 18068 2748
rect 18092 2746 18148 2748
rect 17852 2694 17898 2746
rect 17898 2694 17908 2746
rect 17932 2694 17962 2746
rect 17962 2694 17974 2746
rect 17974 2694 17988 2746
rect 18012 2694 18026 2746
rect 18026 2694 18038 2746
rect 18038 2694 18068 2746
rect 18092 2694 18102 2746
rect 18102 2694 18148 2746
rect 17852 2692 17908 2694
rect 17932 2692 17988 2694
rect 18012 2692 18068 2694
rect 18092 2692 18148 2694
rect 23484 3290 23540 3292
rect 23564 3290 23620 3292
rect 23644 3290 23700 3292
rect 23724 3290 23780 3292
rect 23484 3238 23530 3290
rect 23530 3238 23540 3290
rect 23564 3238 23594 3290
rect 23594 3238 23606 3290
rect 23606 3238 23620 3290
rect 23644 3238 23658 3290
rect 23658 3238 23670 3290
rect 23670 3238 23700 3290
rect 23724 3238 23734 3290
rect 23734 3238 23780 3290
rect 23484 3236 23540 3238
rect 23564 3236 23620 3238
rect 23644 3236 23700 3238
rect 23724 3236 23780 3238
rect 23484 2202 23540 2204
rect 23564 2202 23620 2204
rect 23644 2202 23700 2204
rect 23724 2202 23780 2204
rect 23484 2150 23530 2202
rect 23530 2150 23540 2202
rect 23564 2150 23594 2202
rect 23594 2150 23606 2202
rect 23606 2150 23620 2202
rect 23644 2150 23658 2202
rect 23658 2150 23670 2202
rect 23670 2150 23700 2202
rect 23724 2150 23734 2202
rect 23734 2150 23780 2202
rect 23484 2148 23540 2150
rect 23564 2148 23620 2150
rect 23644 2148 23700 2150
rect 23724 2148 23780 2150
rect 29116 3834 29172 3836
rect 29196 3834 29252 3836
rect 29276 3834 29332 3836
rect 29356 3834 29412 3836
rect 29116 3782 29162 3834
rect 29162 3782 29172 3834
rect 29196 3782 29226 3834
rect 29226 3782 29238 3834
rect 29238 3782 29252 3834
rect 29276 3782 29290 3834
rect 29290 3782 29302 3834
rect 29302 3782 29332 3834
rect 29356 3782 29366 3834
rect 29366 3782 29412 3834
rect 29116 3780 29172 3782
rect 29196 3780 29252 3782
rect 29276 3780 29332 3782
rect 29356 3780 29412 3782
rect 30470 35808 30526 35864
rect 30378 32816 30434 32872
rect 30654 32680 30710 32736
rect 30470 32136 30526 32192
rect 30838 32136 30894 32192
rect 30194 30776 30250 30832
rect 30010 30232 30066 30288
rect 30286 30504 30342 30560
rect 30746 31864 30802 31920
rect 30378 30368 30434 30424
rect 30654 30388 30710 30424
rect 30654 30368 30656 30388
rect 30656 30368 30708 30388
rect 30708 30368 30710 30388
rect 30654 30252 30710 30288
rect 30654 30232 30656 30252
rect 30656 30232 30708 30252
rect 30708 30232 30710 30252
rect 30746 30096 30802 30152
rect 30838 29996 30840 30016
rect 30840 29996 30892 30016
rect 30892 29996 30894 30016
rect 30838 29960 30894 29996
rect 30838 29824 30894 29880
rect 30286 28600 30342 28656
rect 30562 29552 30618 29608
rect 30654 29416 30710 29472
rect 30838 27104 30894 27160
rect 31022 31592 31078 31648
rect 31022 27240 31078 27296
rect 31298 35536 31354 35592
rect 32126 39480 32182 39536
rect 32034 39344 32090 39400
rect 31942 37848 31998 37904
rect 31574 35128 31630 35184
rect 31574 33360 31630 33416
rect 31390 31864 31446 31920
rect 31482 31764 31484 31784
rect 31484 31764 31536 31784
rect 31536 31764 31538 31784
rect 31482 31728 31538 31764
rect 32310 38936 32366 38992
rect 32954 39480 33010 39536
rect 32310 36236 32366 36272
rect 33046 38120 33102 38176
rect 34150 40840 34206 40896
rect 34150 38800 34206 38856
rect 32310 36216 32312 36236
rect 32312 36216 32364 36236
rect 32364 36216 32366 36236
rect 33322 36080 33378 36136
rect 31482 30676 31484 30696
rect 31484 30676 31536 30696
rect 31536 30676 31538 30696
rect 31482 30640 31538 30676
rect 31390 29008 31446 29064
rect 31666 29688 31722 29744
rect 31666 29164 31722 29200
rect 31666 29144 31668 29164
rect 31668 29144 31720 29164
rect 31720 29144 31722 29164
rect 30654 25916 30656 25936
rect 30656 25916 30708 25936
rect 30708 25916 30710 25936
rect 30654 25880 30710 25916
rect 30010 22480 30066 22536
rect 30102 22380 30104 22400
rect 30104 22380 30156 22400
rect 30156 22380 30158 22400
rect 30102 22344 30158 22380
rect 30102 22208 30158 22264
rect 30562 22616 30618 22672
rect 30378 22500 30434 22536
rect 30378 22480 30380 22500
rect 30380 22480 30432 22500
rect 30432 22480 30434 22500
rect 30286 21956 30342 21992
rect 30286 21936 30288 21956
rect 30288 21936 30340 21956
rect 30340 21936 30342 21956
rect 30010 20032 30066 20088
rect 30010 19760 30066 19816
rect 30194 19896 30250 19952
rect 30102 18536 30158 18592
rect 30470 21256 30526 21312
rect 30654 19352 30710 19408
rect 30930 22344 30986 22400
rect 30930 21392 30986 21448
rect 31022 20748 31024 20768
rect 31024 20748 31076 20768
rect 31076 20748 31078 20768
rect 31022 20712 31078 20748
rect 31850 33904 31906 33960
rect 32034 32952 32090 33008
rect 31850 29688 31906 29744
rect 32310 34448 32366 34504
rect 32310 32428 32366 32464
rect 32310 32408 32312 32428
rect 32312 32408 32364 32428
rect 32364 32408 32366 32428
rect 32310 32272 32366 32328
rect 32310 31220 32312 31240
rect 32312 31220 32364 31240
rect 32364 31220 32366 31240
rect 32310 31184 32366 31220
rect 32310 30776 32366 30832
rect 31482 25336 31538 25392
rect 31298 23704 31354 23760
rect 31298 23024 31354 23080
rect 31666 24656 31722 24712
rect 31666 22616 31722 22672
rect 31850 22516 31852 22536
rect 31852 22516 31904 22536
rect 31904 22516 31906 22536
rect 31850 22480 31906 22516
rect 31758 22380 31760 22400
rect 31760 22380 31812 22400
rect 31812 22380 31814 22400
rect 31758 22344 31814 22380
rect 31666 21800 31722 21856
rect 32310 28076 32366 28112
rect 32310 28056 32312 28076
rect 32312 28056 32364 28076
rect 32364 28056 32366 28076
rect 33230 34720 33286 34776
rect 34150 36780 34206 36816
rect 34150 36760 34152 36780
rect 34152 36760 34204 36780
rect 34204 36760 34206 36780
rect 32586 33224 32642 33280
rect 33138 32544 33194 32600
rect 31850 20460 31906 20496
rect 31850 20440 31852 20460
rect 31852 20440 31904 20460
rect 31904 20440 31906 20460
rect 31574 19508 31630 19544
rect 31574 19488 31576 19508
rect 31576 19488 31628 19508
rect 31628 19488 31630 19508
rect 29116 2746 29172 2748
rect 29196 2746 29252 2748
rect 29276 2746 29332 2748
rect 29356 2746 29412 2748
rect 29116 2694 29162 2746
rect 29162 2694 29172 2746
rect 29196 2694 29226 2746
rect 29226 2694 29238 2746
rect 29238 2694 29252 2746
rect 29276 2694 29290 2746
rect 29290 2694 29302 2746
rect 29302 2694 29332 2746
rect 29356 2694 29366 2746
rect 29366 2694 29412 2746
rect 29116 2692 29172 2694
rect 29196 2692 29252 2694
rect 29276 2692 29332 2694
rect 29356 2692 29412 2694
rect 32402 23840 32458 23896
rect 32218 22208 32274 22264
rect 32218 22072 32274 22128
rect 32402 22888 32458 22944
rect 32402 22752 32458 22808
rect 32402 21800 32458 21856
rect 32678 22480 32734 22536
rect 32954 25336 33010 25392
rect 34150 34720 34206 34776
rect 34150 34060 34206 34096
rect 34150 34040 34152 34060
rect 34152 34040 34204 34060
rect 34204 34040 34206 34060
rect 34150 33396 34152 33416
rect 34152 33396 34204 33416
rect 34204 33396 34206 33416
rect 34150 33360 34206 33396
rect 34150 32680 34206 32736
rect 34150 32000 34206 32056
rect 34150 31340 34206 31376
rect 34150 31320 34152 31340
rect 34152 31320 34204 31340
rect 34204 31320 34206 31340
rect 33874 30912 33930 30968
rect 33506 30096 33562 30152
rect 33414 26832 33470 26888
rect 33046 22616 33102 22672
rect 32862 22092 32918 22128
rect 33138 22344 33194 22400
rect 32862 22072 32864 22092
rect 32864 22072 32916 22092
rect 32916 22072 32918 22092
rect 33506 23568 33562 23624
rect 32034 2080 32090 2136
rect 32586 40 32642 96
rect 33046 3440 33102 3496
rect 34150 27956 34152 27976
rect 34152 27956 34204 27976
rect 34204 27956 34206 27976
rect 34150 27920 34206 27956
rect 34150 25900 34206 25936
rect 34150 25880 34152 25900
rect 34152 25880 34204 25900
rect 34204 25880 34206 25900
rect 34150 25236 34152 25256
rect 34152 25236 34204 25256
rect 34204 25236 34206 25256
rect 34150 25200 34206 25236
rect 34150 24520 34206 24576
rect 34150 23840 34206 23896
rect 34150 23180 34206 23216
rect 34150 23160 34152 23180
rect 34152 23160 34204 23180
rect 34204 23160 34206 23180
rect 34150 20460 34206 20496
rect 34150 20440 34152 20460
rect 34152 20440 34204 20460
rect 34204 20440 34206 20460
rect 34150 19780 34206 19816
rect 34150 19760 34152 19780
rect 34152 19760 34204 19780
rect 34204 19760 34206 19780
rect 34150 19080 34206 19136
rect 34150 17740 34206 17776
rect 34150 17720 34152 17740
rect 34152 17720 34204 17740
rect 34204 17720 34206 17740
rect 34150 17076 34152 17096
rect 34152 17076 34204 17096
rect 34204 17076 34206 17096
rect 34150 17040 34206 17076
rect 34150 16360 34206 16416
rect 34150 14340 34206 14376
rect 34150 14320 34152 14340
rect 34152 14320 34204 14340
rect 34204 14320 34206 14340
rect 34150 13640 34206 13696
rect 34150 12960 34206 13016
rect 34150 12300 34206 12336
rect 34150 12280 34152 12300
rect 34152 12280 34204 12300
rect 34204 12280 34206 12300
rect 33966 9560 34022 9616
rect 34150 8880 34206 8936
rect 34150 6860 34206 6896
rect 34150 6840 34152 6860
rect 34152 6840 34204 6860
rect 34204 6840 34206 6860
rect 34150 4800 34206 4856
rect 34150 4120 34206 4176
rect 34426 720 34482 776
<< metal3 >>
rect 0 41578 800 41668
rect 2957 41578 3023 41581
rect 0 41576 3023 41578
rect 0 41520 2962 41576
rect 3018 41520 3023 41576
rect 0 41518 3023 41520
rect 0 41428 800 41518
rect 2957 41515 3023 41518
rect 0 40898 800 40988
rect 4153 40898 4219 40901
rect 0 40896 4219 40898
rect 0 40840 4158 40896
rect 4214 40840 4219 40896
rect 0 40838 4219 40840
rect 0 40748 800 40838
rect 4153 40835 4219 40838
rect 14590 40836 14596 40900
rect 14660 40898 14666 40900
rect 21633 40898 21699 40901
rect 14660 40896 21699 40898
rect 14660 40840 21638 40896
rect 21694 40840 21699 40896
rect 14660 40838 21699 40840
rect 14660 40836 14666 40838
rect 21633 40835 21699 40838
rect 34145 40898 34211 40901
rect 35200 40898 36000 40988
rect 34145 40896 36000 40898
rect 34145 40840 34150 40896
rect 34206 40840 36000 40896
rect 34145 40838 36000 40840
rect 34145 40835 34211 40838
rect 13169 40762 13235 40765
rect 22921 40762 22987 40765
rect 13169 40760 22987 40762
rect 13169 40704 13174 40760
rect 13230 40704 22926 40760
rect 22982 40704 22987 40760
rect 35200 40748 36000 40838
rect 13169 40702 22987 40704
rect 13169 40699 13235 40702
rect 22921 40699 22987 40702
rect 11053 40626 11119 40629
rect 18505 40626 18571 40629
rect 11053 40624 18571 40626
rect 11053 40568 11058 40624
rect 11114 40568 18510 40624
rect 18566 40568 18571 40624
rect 11053 40566 18571 40568
rect 11053 40563 11119 40566
rect 18505 40563 18571 40566
rect 15285 40490 15351 40493
rect 18454 40490 18460 40492
rect 15285 40488 18460 40490
rect 15285 40432 15290 40488
rect 15346 40432 18460 40488
rect 15285 40430 18460 40432
rect 15285 40427 15351 40430
rect 18454 40428 18460 40430
rect 18524 40428 18530 40492
rect 14273 40354 14339 40357
rect 19149 40354 19215 40357
rect 14273 40352 19215 40354
rect 14273 40296 14278 40352
rect 14334 40296 19154 40352
rect 19210 40296 19215 40352
rect 14273 40294 19215 40296
rect 14273 40291 14339 40294
rect 19149 40291 19215 40294
rect 9765 40218 9831 40221
rect 16665 40218 16731 40221
rect 9765 40216 16731 40218
rect 9765 40160 9770 40216
rect 9826 40160 16670 40216
rect 16726 40160 16731 40216
rect 9765 40158 16731 40160
rect 9765 40155 9831 40158
rect 16665 40155 16731 40158
rect 17677 40218 17743 40221
rect 20529 40218 20595 40221
rect 22001 40218 22067 40221
rect 17677 40216 22067 40218
rect 17677 40160 17682 40216
rect 17738 40160 20534 40216
rect 20590 40160 22006 40216
rect 22062 40160 22067 40216
rect 17677 40158 22067 40160
rect 17677 40155 17743 40158
rect 20529 40155 20595 40158
rect 22001 40155 22067 40158
rect 13997 40082 14063 40085
rect 20069 40082 20135 40085
rect 13997 40080 20135 40082
rect 13997 40024 14002 40080
rect 14058 40024 20074 40080
rect 20130 40024 20135 40080
rect 35200 40068 36000 40308
rect 13997 40022 20135 40024
rect 13997 40019 14063 40022
rect 20069 40019 20135 40022
rect 10317 39946 10383 39949
rect 17033 39946 17099 39949
rect 26877 39946 26943 39949
rect 31385 39946 31451 39949
rect 10317 39944 17099 39946
rect 10317 39888 10322 39944
rect 10378 39888 17038 39944
rect 17094 39888 17099 39944
rect 10317 39886 17099 39888
rect 10317 39883 10383 39886
rect 17033 39883 17099 39886
rect 17174 39944 26943 39946
rect 17174 39888 26882 39944
rect 26938 39888 26943 39944
rect 17174 39886 26943 39888
rect 12014 39748 12020 39812
rect 12084 39810 12090 39812
rect 17174 39810 17234 39886
rect 26877 39883 26943 39886
rect 28950 39944 31451 39946
rect 28950 39888 31390 39944
rect 31446 39888 31451 39944
rect 28950 39886 31451 39888
rect 12084 39750 17234 39810
rect 18321 39810 18387 39813
rect 28950 39810 29010 39886
rect 31385 39883 31451 39886
rect 18321 39808 29010 39810
rect 18321 39752 18326 39808
rect 18382 39752 29010 39808
rect 18321 39750 29010 39752
rect 12084 39748 12090 39750
rect 18321 39747 18387 39750
rect 6576 39744 6896 39745
rect 6576 39680 6584 39744
rect 6648 39680 6664 39744
rect 6728 39680 6744 39744
rect 6808 39680 6824 39744
rect 6888 39680 6896 39744
rect 6576 39679 6896 39680
rect 17840 39744 18160 39745
rect 17840 39680 17848 39744
rect 17912 39680 17928 39744
rect 17992 39680 18008 39744
rect 18072 39680 18088 39744
rect 18152 39680 18160 39744
rect 17840 39679 18160 39680
rect 29104 39744 29424 39745
rect 29104 39680 29112 39744
rect 29176 39680 29192 39744
rect 29256 39680 29272 39744
rect 29336 39680 29352 39744
rect 29416 39680 29424 39744
rect 29104 39679 29424 39680
rect 14089 39674 14155 39677
rect 17493 39674 17559 39677
rect 14089 39672 17559 39674
rect 0 39388 800 39628
rect 14089 39616 14094 39672
rect 14150 39616 17498 39672
rect 17554 39616 17559 39672
rect 14089 39614 17559 39616
rect 14089 39611 14155 39614
rect 17493 39611 17559 39614
rect 19333 39674 19399 39677
rect 23657 39674 23723 39677
rect 26509 39674 26575 39677
rect 19333 39672 26575 39674
rect 19333 39616 19338 39672
rect 19394 39616 23662 39672
rect 23718 39616 26514 39672
rect 26570 39616 26575 39672
rect 19333 39614 26575 39616
rect 19333 39611 19399 39614
rect 23657 39611 23723 39614
rect 26509 39611 26575 39614
rect 9581 39538 9647 39541
rect 16849 39538 16915 39541
rect 9581 39536 16915 39538
rect 9581 39480 9586 39536
rect 9642 39480 16854 39536
rect 16910 39480 16915 39536
rect 9581 39478 16915 39480
rect 9581 39475 9647 39478
rect 16849 39475 16915 39478
rect 17033 39538 17099 39541
rect 32121 39538 32187 39541
rect 17033 39536 32187 39538
rect 17033 39480 17038 39536
rect 17094 39480 32126 39536
rect 32182 39480 32187 39536
rect 17033 39478 32187 39480
rect 17033 39475 17099 39478
rect 32121 39475 32187 39478
rect 32949 39538 33015 39541
rect 35200 39538 36000 39628
rect 32949 39536 36000 39538
rect 32949 39480 32954 39536
rect 33010 39480 36000 39536
rect 32949 39478 36000 39480
rect 32949 39475 33015 39478
rect 10961 39402 11027 39405
rect 32029 39402 32095 39405
rect 10961 39400 32095 39402
rect 10961 39344 10966 39400
rect 11022 39344 32034 39400
rect 32090 39344 32095 39400
rect 35200 39388 36000 39478
rect 10961 39342 32095 39344
rect 10961 39339 11027 39342
rect 32029 39339 32095 39342
rect 13445 39266 13511 39269
rect 16665 39266 16731 39269
rect 13445 39264 16731 39266
rect 13445 39208 13450 39264
rect 13506 39208 16670 39264
rect 16726 39208 16731 39264
rect 13445 39206 16731 39208
rect 13445 39203 13511 39206
rect 16665 39203 16731 39206
rect 16849 39266 16915 39269
rect 16849 39264 23306 39266
rect 16849 39208 16854 39264
rect 16910 39208 23306 39264
rect 16849 39206 23306 39208
rect 16849 39203 16915 39206
rect 12208 39200 12528 39201
rect 12208 39136 12216 39200
rect 12280 39136 12296 39200
rect 12360 39136 12376 39200
rect 12440 39136 12456 39200
rect 12520 39136 12528 39200
rect 12208 39135 12528 39136
rect 13261 39130 13327 39133
rect 18321 39130 18387 39133
rect 13261 39128 18387 39130
rect 13261 39072 13266 39128
rect 13322 39072 18326 39128
rect 18382 39072 18387 39128
rect 13261 39070 18387 39072
rect 13261 39067 13327 39070
rect 18321 39067 18387 39070
rect 18454 39068 18460 39132
rect 18524 39130 18530 39132
rect 22645 39130 22711 39133
rect 18524 39128 22711 39130
rect 18524 39072 22650 39128
rect 22706 39072 22711 39128
rect 18524 39070 22711 39072
rect 18524 39068 18530 39070
rect 22645 39067 22711 39070
rect 10317 38994 10383 38997
rect 18781 38994 18847 38997
rect 10317 38992 18847 38994
rect 0 38858 800 38948
rect 10317 38936 10322 38992
rect 10378 38936 18786 38992
rect 18842 38936 18847 38992
rect 10317 38934 18847 38936
rect 10317 38931 10383 38934
rect 18781 38931 18847 38934
rect 20161 38994 20227 38997
rect 22829 38994 22895 38997
rect 20161 38992 22895 38994
rect 20161 38936 20166 38992
rect 20222 38936 22834 38992
rect 22890 38936 22895 38992
rect 20161 38934 22895 38936
rect 23246 38994 23306 39206
rect 23472 39200 23792 39201
rect 23472 39136 23480 39200
rect 23544 39136 23560 39200
rect 23624 39136 23640 39200
rect 23704 39136 23720 39200
rect 23784 39136 23792 39200
rect 23472 39135 23792 39136
rect 24485 38994 24551 38997
rect 23246 38992 24551 38994
rect 23246 38936 24490 38992
rect 24546 38936 24551 38992
rect 23246 38934 24551 38936
rect 20161 38931 20227 38934
rect 22829 38931 22895 38934
rect 24485 38931 24551 38934
rect 26877 38994 26943 38997
rect 32305 38994 32371 38997
rect 26877 38992 32371 38994
rect 26877 38936 26882 38992
rect 26938 38936 32310 38992
rect 32366 38936 32371 38992
rect 26877 38934 32371 38936
rect 26877 38931 26943 38934
rect 32305 38931 32371 38934
rect 1393 38858 1459 38861
rect 0 38856 1459 38858
rect 0 38800 1398 38856
rect 1454 38800 1459 38856
rect 0 38798 1459 38800
rect 0 38708 800 38798
rect 1393 38795 1459 38798
rect 12750 38796 12756 38860
rect 12820 38858 12826 38860
rect 17033 38858 17099 38861
rect 18321 38858 18387 38861
rect 12820 38798 16820 38858
rect 12820 38796 12826 38798
rect 13445 38722 13511 38725
rect 16573 38722 16639 38725
rect 13445 38720 16639 38722
rect 13445 38664 13450 38720
rect 13506 38664 16578 38720
rect 16634 38664 16639 38720
rect 13445 38662 16639 38664
rect 16760 38722 16820 38798
rect 17033 38856 18387 38858
rect 17033 38800 17038 38856
rect 17094 38800 18326 38856
rect 18382 38800 18387 38856
rect 17033 38798 18387 38800
rect 17033 38795 17099 38798
rect 18321 38795 18387 38798
rect 18505 38858 18571 38861
rect 27705 38858 27771 38861
rect 18505 38856 27771 38858
rect 18505 38800 18510 38856
rect 18566 38800 27710 38856
rect 27766 38800 27771 38856
rect 18505 38798 27771 38800
rect 18505 38795 18571 38798
rect 27705 38795 27771 38798
rect 34145 38858 34211 38861
rect 35200 38858 36000 38948
rect 34145 38856 36000 38858
rect 34145 38800 34150 38856
rect 34206 38800 36000 38856
rect 34145 38798 36000 38800
rect 34145 38795 34211 38798
rect 17401 38722 17467 38725
rect 17677 38722 17743 38725
rect 16760 38720 17467 38722
rect 16760 38664 17406 38720
rect 17462 38664 17467 38720
rect 16760 38662 17467 38664
rect 13445 38659 13511 38662
rect 16573 38659 16639 38662
rect 17401 38659 17467 38662
rect 17542 38720 17743 38722
rect 17542 38664 17682 38720
rect 17738 38664 17743 38720
rect 17542 38662 17743 38664
rect 6576 38656 6896 38657
rect 6576 38592 6584 38656
rect 6648 38592 6664 38656
rect 6728 38592 6744 38656
rect 6808 38592 6824 38656
rect 6888 38592 6896 38656
rect 6576 38591 6896 38592
rect 12014 38524 12020 38588
rect 12084 38586 12090 38588
rect 12249 38586 12315 38589
rect 12084 38584 12315 38586
rect 12084 38528 12254 38584
rect 12310 38528 12315 38584
rect 12084 38526 12315 38528
rect 12084 38524 12090 38526
rect 12249 38523 12315 38526
rect 13353 38586 13419 38589
rect 17542 38586 17602 38662
rect 17677 38659 17743 38662
rect 18781 38722 18847 38725
rect 26969 38722 27035 38725
rect 18781 38720 27035 38722
rect 18781 38664 18786 38720
rect 18842 38664 26974 38720
rect 27030 38664 27035 38720
rect 35200 38708 36000 38798
rect 18781 38662 27035 38664
rect 18781 38659 18847 38662
rect 26969 38659 27035 38662
rect 17840 38656 18160 38657
rect 17840 38592 17848 38656
rect 17912 38592 17928 38656
rect 17992 38592 18008 38656
rect 18072 38592 18088 38656
rect 18152 38592 18160 38656
rect 17840 38591 18160 38592
rect 29104 38656 29424 38657
rect 29104 38592 29112 38656
rect 29176 38592 29192 38656
rect 29256 38592 29272 38656
rect 29336 38592 29352 38656
rect 29416 38592 29424 38656
rect 29104 38591 29424 38592
rect 13353 38584 17602 38586
rect 13353 38528 13358 38584
rect 13414 38528 17602 38584
rect 13353 38526 17602 38528
rect 19977 38586 20043 38589
rect 22093 38586 22159 38589
rect 19977 38584 22159 38586
rect 19977 38528 19982 38584
rect 20038 38528 22098 38584
rect 22154 38528 22159 38584
rect 19977 38526 22159 38528
rect 13353 38523 13419 38526
rect 19977 38523 20043 38526
rect 22093 38523 22159 38526
rect 22277 38586 22343 38589
rect 28257 38586 28323 38589
rect 28625 38586 28691 38589
rect 22277 38584 28691 38586
rect 22277 38528 22282 38584
rect 22338 38528 28262 38584
rect 28318 38528 28630 38584
rect 28686 38528 28691 38584
rect 22277 38526 28691 38528
rect 22277 38523 22343 38526
rect 28257 38523 28323 38526
rect 28625 38523 28691 38526
rect 13077 38450 13143 38453
rect 18689 38450 18755 38453
rect 13077 38448 18755 38450
rect 13077 38392 13082 38448
rect 13138 38392 18694 38448
rect 18750 38392 18755 38448
rect 13077 38390 18755 38392
rect 13077 38387 13143 38390
rect 18689 38387 18755 38390
rect 19793 38450 19859 38453
rect 21725 38450 21791 38453
rect 19793 38448 21791 38450
rect 19793 38392 19798 38448
rect 19854 38392 21730 38448
rect 21786 38392 21791 38448
rect 19793 38390 21791 38392
rect 19793 38387 19859 38390
rect 21725 38387 21791 38390
rect 21909 38450 21975 38453
rect 27705 38450 27771 38453
rect 28533 38450 28599 38453
rect 21909 38448 28599 38450
rect 21909 38392 21914 38448
rect 21970 38392 27710 38448
rect 27766 38392 28538 38448
rect 28594 38392 28599 38448
rect 21909 38390 28599 38392
rect 21909 38387 21975 38390
rect 27705 38387 27771 38390
rect 28533 38387 28599 38390
rect 10869 38314 10935 38317
rect 25129 38314 25195 38317
rect 10869 38312 25195 38314
rect 0 38028 800 38268
rect 10869 38256 10874 38312
rect 10930 38256 25134 38312
rect 25190 38256 25195 38312
rect 10869 38254 25195 38256
rect 10869 38251 10935 38254
rect 25129 38251 25195 38254
rect 12893 38178 12959 38181
rect 21449 38178 21515 38181
rect 12893 38176 21515 38178
rect 12893 38120 12898 38176
rect 12954 38120 21454 38176
rect 21510 38120 21515 38176
rect 12893 38118 21515 38120
rect 12893 38115 12959 38118
rect 21449 38115 21515 38118
rect 33041 38178 33107 38181
rect 35200 38178 36000 38268
rect 33041 38176 36000 38178
rect 33041 38120 33046 38176
rect 33102 38120 36000 38176
rect 33041 38118 36000 38120
rect 33041 38115 33107 38118
rect 12208 38112 12528 38113
rect 12208 38048 12216 38112
rect 12280 38048 12296 38112
rect 12360 38048 12376 38112
rect 12440 38048 12456 38112
rect 12520 38048 12528 38112
rect 12208 38047 12528 38048
rect 23472 38112 23792 38113
rect 23472 38048 23480 38112
rect 23544 38048 23560 38112
rect 23624 38048 23640 38112
rect 23704 38048 23720 38112
rect 23784 38048 23792 38112
rect 23472 38047 23792 38048
rect 13077 38042 13143 38045
rect 13721 38042 13787 38045
rect 13077 38040 13787 38042
rect 13077 37984 13082 38040
rect 13138 37984 13726 38040
rect 13782 37984 13787 38040
rect 13077 37982 13787 37984
rect 13077 37979 13143 37982
rect 13721 37979 13787 37982
rect 14273 38042 14339 38045
rect 16297 38042 16363 38045
rect 14273 38040 16363 38042
rect 14273 37984 14278 38040
rect 14334 37984 16302 38040
rect 16358 37984 16363 38040
rect 14273 37982 16363 37984
rect 14273 37979 14339 37982
rect 16297 37979 16363 37982
rect 16481 38042 16547 38045
rect 20713 38042 20779 38045
rect 16481 38040 20779 38042
rect 16481 37984 16486 38040
rect 16542 37984 20718 38040
rect 20774 37984 20779 38040
rect 35200 38028 36000 38118
rect 16481 37982 20779 37984
rect 16481 37979 16547 37982
rect 20713 37979 20779 37982
rect 10777 37906 10843 37909
rect 31937 37906 32003 37909
rect 10777 37904 32003 37906
rect 10777 37848 10782 37904
rect 10838 37848 31942 37904
rect 31998 37848 32003 37904
rect 10777 37846 32003 37848
rect 10777 37843 10843 37846
rect 31937 37843 32003 37846
rect 9673 37770 9739 37773
rect 29545 37770 29611 37773
rect 9673 37768 29611 37770
rect 9673 37712 9678 37768
rect 9734 37712 29550 37768
rect 29606 37712 29611 37768
rect 9673 37710 29611 37712
rect 9673 37707 9739 37710
rect 29545 37707 29611 37710
rect 12341 37634 12407 37637
rect 17677 37634 17743 37637
rect 12341 37632 17743 37634
rect 0 37498 800 37588
rect 12341 37576 12346 37632
rect 12402 37576 17682 37632
rect 17738 37576 17743 37632
rect 12341 37574 17743 37576
rect 12341 37571 12407 37574
rect 17677 37571 17743 37574
rect 18321 37634 18387 37637
rect 22185 37634 22251 37637
rect 18321 37632 22251 37634
rect 18321 37576 18326 37632
rect 18382 37576 22190 37632
rect 22246 37576 22251 37632
rect 18321 37574 22251 37576
rect 18321 37571 18387 37574
rect 22185 37571 22251 37574
rect 6576 37568 6896 37569
rect 6576 37504 6584 37568
rect 6648 37504 6664 37568
rect 6728 37504 6744 37568
rect 6808 37504 6824 37568
rect 6888 37504 6896 37568
rect 6576 37503 6896 37504
rect 17840 37568 18160 37569
rect 17840 37504 17848 37568
rect 17912 37504 17928 37568
rect 17992 37504 18008 37568
rect 18072 37504 18088 37568
rect 18152 37504 18160 37568
rect 17840 37503 18160 37504
rect 29104 37568 29424 37569
rect 29104 37504 29112 37568
rect 29176 37504 29192 37568
rect 29256 37504 29272 37568
rect 29336 37504 29352 37568
rect 29416 37504 29424 37568
rect 29104 37503 29424 37504
rect 3969 37498 4035 37501
rect 0 37496 4035 37498
rect 0 37440 3974 37496
rect 4030 37440 4035 37496
rect 0 37438 4035 37440
rect 0 37348 800 37438
rect 3969 37435 4035 37438
rect 11421 37498 11487 37501
rect 15745 37498 15811 37501
rect 11421 37496 15811 37498
rect 11421 37440 11426 37496
rect 11482 37440 15750 37496
rect 15806 37440 15811 37496
rect 11421 37438 15811 37440
rect 11421 37435 11487 37438
rect 15745 37435 15811 37438
rect 16297 37498 16363 37501
rect 16849 37498 16915 37501
rect 16297 37496 16915 37498
rect 16297 37440 16302 37496
rect 16358 37440 16854 37496
rect 16910 37440 16915 37496
rect 16297 37438 16915 37440
rect 16297 37435 16363 37438
rect 16849 37435 16915 37438
rect 17033 37498 17099 37501
rect 17309 37498 17375 37501
rect 17585 37500 17651 37501
rect 17033 37496 17375 37498
rect 17033 37440 17038 37496
rect 17094 37440 17314 37496
rect 17370 37440 17375 37496
rect 17033 37438 17375 37440
rect 17033 37435 17099 37438
rect 17309 37435 17375 37438
rect 17534 37436 17540 37500
rect 17604 37498 17651 37500
rect 18229 37498 18295 37501
rect 20805 37498 20871 37501
rect 17604 37496 17696 37498
rect 17646 37440 17696 37496
rect 17604 37438 17696 37440
rect 18229 37496 20871 37498
rect 18229 37440 18234 37496
rect 18290 37440 20810 37496
rect 20866 37440 20871 37496
rect 18229 37438 20871 37440
rect 17604 37436 17651 37438
rect 17585 37435 17651 37436
rect 18229 37435 18295 37438
rect 20805 37435 20871 37438
rect 20989 37498 21055 37501
rect 24761 37498 24827 37501
rect 20989 37496 24827 37498
rect 20989 37440 20994 37496
rect 21050 37440 24766 37496
rect 24822 37440 24827 37496
rect 20989 37438 24827 37440
rect 20989 37435 21055 37438
rect 24761 37435 24827 37438
rect 10225 37362 10291 37365
rect 29729 37362 29795 37365
rect 10225 37360 29795 37362
rect 10225 37304 10230 37360
rect 10286 37304 29734 37360
rect 29790 37304 29795 37360
rect 35200 37348 36000 37588
rect 10225 37302 29795 37304
rect 10225 37299 10291 37302
rect 29729 37299 29795 37302
rect 11973 37226 12039 37229
rect 24853 37226 24919 37229
rect 11973 37224 24919 37226
rect 11973 37168 11978 37224
rect 12034 37168 24858 37224
rect 24914 37168 24919 37224
rect 11973 37166 24919 37168
rect 11973 37163 12039 37166
rect 24853 37163 24919 37166
rect 12617 37090 12683 37093
rect 20713 37090 20779 37093
rect 12617 37088 20779 37090
rect 12617 37032 12622 37088
rect 12678 37032 20718 37088
rect 20774 37032 20779 37088
rect 12617 37030 20779 37032
rect 12617 37027 12683 37030
rect 20713 37027 20779 37030
rect 12208 37024 12528 37025
rect 12208 36960 12216 37024
rect 12280 36960 12296 37024
rect 12360 36960 12376 37024
rect 12440 36960 12456 37024
rect 12520 36960 12528 37024
rect 12208 36959 12528 36960
rect 23472 37024 23792 37025
rect 23472 36960 23480 37024
rect 23544 36960 23560 37024
rect 23624 36960 23640 37024
rect 23704 36960 23720 37024
rect 23784 36960 23792 37024
rect 23472 36959 23792 36960
rect 12801 36954 12867 36957
rect 15837 36954 15903 36957
rect 12801 36952 15903 36954
rect 0 36818 800 36908
rect 12801 36896 12806 36952
rect 12862 36896 15842 36952
rect 15898 36896 15903 36952
rect 12801 36894 15903 36896
rect 12801 36891 12867 36894
rect 15837 36891 15903 36894
rect 16113 36954 16179 36957
rect 19425 36954 19491 36957
rect 16113 36952 19491 36954
rect 16113 36896 16118 36952
rect 16174 36896 19430 36952
rect 19486 36896 19491 36952
rect 16113 36894 19491 36896
rect 16113 36891 16179 36894
rect 19425 36891 19491 36894
rect 19609 36954 19675 36957
rect 19609 36952 23122 36954
rect 19609 36896 19614 36952
rect 19670 36896 23122 36952
rect 19609 36894 23122 36896
rect 19609 36891 19675 36894
rect 2773 36818 2839 36821
rect 0 36816 2839 36818
rect 0 36760 2778 36816
rect 2834 36760 2839 36816
rect 0 36758 2839 36760
rect 0 36668 800 36758
rect 2773 36755 2839 36758
rect 13813 36818 13879 36821
rect 20805 36818 20871 36821
rect 22737 36818 22803 36821
rect 13813 36816 20871 36818
rect 13813 36760 13818 36816
rect 13874 36760 20810 36816
rect 20866 36760 20871 36816
rect 13813 36758 20871 36760
rect 13813 36755 13879 36758
rect 20805 36755 20871 36758
rect 20992 36816 22803 36818
rect 20992 36760 22742 36816
rect 22798 36760 22803 36816
rect 20992 36758 22803 36760
rect 23062 36818 23122 36894
rect 23933 36818 23999 36821
rect 23062 36816 23999 36818
rect 23062 36760 23938 36816
rect 23994 36760 23999 36816
rect 23062 36758 23999 36760
rect 12065 36682 12131 36685
rect 13077 36682 13143 36685
rect 12065 36680 13143 36682
rect 12065 36624 12070 36680
rect 12126 36624 13082 36680
rect 13138 36624 13143 36680
rect 12065 36622 13143 36624
rect 12065 36619 12131 36622
rect 13077 36619 13143 36622
rect 13445 36682 13511 36685
rect 15193 36682 15259 36685
rect 13445 36680 15259 36682
rect 13445 36624 13450 36680
rect 13506 36624 15198 36680
rect 15254 36624 15259 36680
rect 13445 36622 15259 36624
rect 13445 36619 13511 36622
rect 15193 36619 15259 36622
rect 15653 36682 15719 36685
rect 16297 36682 16363 36685
rect 15653 36680 16363 36682
rect 15653 36624 15658 36680
rect 15714 36624 16302 36680
rect 16358 36624 16363 36680
rect 15653 36622 16363 36624
rect 15653 36619 15719 36622
rect 16297 36619 16363 36622
rect 16481 36682 16547 36685
rect 18781 36682 18847 36685
rect 16481 36680 18847 36682
rect 16481 36624 16486 36680
rect 16542 36624 18786 36680
rect 18842 36624 18847 36680
rect 16481 36622 18847 36624
rect 16481 36619 16547 36622
rect 18781 36619 18847 36622
rect 19057 36682 19123 36685
rect 20992 36682 21052 36758
rect 22737 36755 22803 36758
rect 23933 36755 23999 36758
rect 34145 36818 34211 36821
rect 35200 36818 36000 36908
rect 34145 36816 36000 36818
rect 34145 36760 34150 36816
rect 34206 36760 36000 36816
rect 34145 36758 36000 36760
rect 34145 36755 34211 36758
rect 19057 36680 21052 36682
rect 19057 36624 19062 36680
rect 19118 36624 21052 36680
rect 19057 36622 21052 36624
rect 21817 36682 21883 36685
rect 28165 36682 28231 36685
rect 21817 36680 28231 36682
rect 21817 36624 21822 36680
rect 21878 36624 28170 36680
rect 28226 36624 28231 36680
rect 35200 36668 36000 36758
rect 21817 36622 28231 36624
rect 19057 36619 19123 36622
rect 21817 36619 21883 36622
rect 28165 36619 28231 36622
rect 13169 36546 13235 36549
rect 17677 36546 17743 36549
rect 13169 36544 17743 36546
rect 13169 36488 13174 36544
rect 13230 36488 17682 36544
rect 17738 36488 17743 36544
rect 13169 36486 17743 36488
rect 13169 36483 13235 36486
rect 17677 36483 17743 36486
rect 18229 36546 18295 36549
rect 21357 36546 21423 36549
rect 18229 36544 21423 36546
rect 18229 36488 18234 36544
rect 18290 36488 21362 36544
rect 21418 36488 21423 36544
rect 18229 36486 21423 36488
rect 18229 36483 18295 36486
rect 21357 36483 21423 36486
rect 6576 36480 6896 36481
rect 6576 36416 6584 36480
rect 6648 36416 6664 36480
rect 6728 36416 6744 36480
rect 6808 36416 6824 36480
rect 6888 36416 6896 36480
rect 6576 36415 6896 36416
rect 17840 36480 18160 36481
rect 17840 36416 17848 36480
rect 17912 36416 17928 36480
rect 17992 36416 18008 36480
rect 18072 36416 18088 36480
rect 18152 36416 18160 36480
rect 17840 36415 18160 36416
rect 29104 36480 29424 36481
rect 29104 36416 29112 36480
rect 29176 36416 29192 36480
rect 29256 36416 29272 36480
rect 29336 36416 29352 36480
rect 29416 36416 29424 36480
rect 29104 36415 29424 36416
rect 12341 36410 12407 36413
rect 15009 36410 15075 36413
rect 15653 36410 15719 36413
rect 12341 36408 15719 36410
rect 12341 36352 12346 36408
rect 12402 36352 15014 36408
rect 15070 36352 15658 36408
rect 15714 36352 15719 36408
rect 12341 36350 15719 36352
rect 12341 36347 12407 36350
rect 15009 36347 15075 36350
rect 15653 36347 15719 36350
rect 15929 36410 15995 36413
rect 16205 36410 16271 36413
rect 15929 36408 16271 36410
rect 15929 36352 15934 36408
rect 15990 36352 16210 36408
rect 16266 36352 16271 36408
rect 15929 36350 16271 36352
rect 15929 36347 15995 36350
rect 16205 36347 16271 36350
rect 16389 36410 16455 36413
rect 17677 36410 17743 36413
rect 16389 36408 17743 36410
rect 16389 36352 16394 36408
rect 16450 36352 17682 36408
rect 17738 36352 17743 36408
rect 16389 36350 17743 36352
rect 16389 36347 16455 36350
rect 17677 36347 17743 36350
rect 18321 36410 18387 36413
rect 20897 36410 20963 36413
rect 18321 36408 20963 36410
rect 18321 36352 18326 36408
rect 18382 36352 20902 36408
rect 20958 36352 20963 36408
rect 18321 36350 20963 36352
rect 18321 36347 18387 36350
rect 20897 36347 20963 36350
rect 21081 36410 21147 36413
rect 23657 36410 23723 36413
rect 21081 36408 23723 36410
rect 21081 36352 21086 36408
rect 21142 36352 23662 36408
rect 23718 36352 23723 36408
rect 21081 36350 23723 36352
rect 21081 36347 21147 36350
rect 23657 36347 23723 36350
rect 11605 36274 11671 36277
rect 32305 36274 32371 36277
rect 11605 36272 32371 36274
rect 0 36138 800 36228
rect 11605 36216 11610 36272
rect 11666 36216 32310 36272
rect 32366 36216 32371 36272
rect 11605 36214 32371 36216
rect 11605 36211 11671 36214
rect 32305 36211 32371 36214
rect 1393 36138 1459 36141
rect 0 36136 1459 36138
rect 0 36080 1398 36136
rect 1454 36080 1459 36136
rect 0 36078 1459 36080
rect 0 35988 800 36078
rect 1393 36075 1459 36078
rect 12157 36138 12223 36141
rect 18781 36138 18847 36141
rect 12157 36136 18847 36138
rect 12157 36080 12162 36136
rect 12218 36080 18786 36136
rect 18842 36080 18847 36136
rect 12157 36078 18847 36080
rect 12157 36075 12223 36078
rect 18781 36075 18847 36078
rect 18965 36138 19031 36141
rect 21081 36138 21147 36141
rect 27889 36138 27955 36141
rect 18965 36136 21147 36138
rect 18965 36080 18970 36136
rect 19026 36080 21086 36136
rect 21142 36080 21147 36136
rect 18965 36078 21147 36080
rect 18965 36075 19031 36078
rect 21081 36075 21147 36078
rect 22280 36136 27955 36138
rect 22280 36080 27894 36136
rect 27950 36080 27955 36136
rect 22280 36078 27955 36080
rect 12709 36002 12775 36005
rect 20529 36002 20595 36005
rect 12709 36000 20595 36002
rect 12709 35944 12714 36000
rect 12770 35944 20534 36000
rect 20590 35944 20595 36000
rect 12709 35942 20595 35944
rect 12709 35939 12775 35942
rect 20529 35939 20595 35942
rect 20805 36002 20871 36005
rect 22093 36002 22159 36005
rect 20805 36000 22159 36002
rect 20805 35944 20810 36000
rect 20866 35944 22098 36000
rect 22154 35944 22159 36000
rect 20805 35942 22159 35944
rect 20805 35939 20871 35942
rect 22093 35939 22159 35942
rect 12208 35936 12528 35937
rect 12208 35872 12216 35936
rect 12280 35872 12296 35936
rect 12360 35872 12376 35936
rect 12440 35872 12456 35936
rect 12520 35872 12528 35936
rect 12208 35871 12528 35872
rect 13905 35866 13971 35869
rect 19609 35866 19675 35869
rect 22280 35866 22340 36078
rect 27889 36075 27955 36078
rect 33317 36138 33383 36141
rect 35200 36138 36000 36228
rect 33317 36136 36000 36138
rect 33317 36080 33322 36136
rect 33378 36080 36000 36136
rect 33317 36078 36000 36080
rect 33317 36075 33383 36078
rect 35200 35988 36000 36078
rect 23472 35936 23792 35937
rect 23472 35872 23480 35936
rect 23544 35872 23560 35936
rect 23624 35872 23640 35936
rect 23704 35872 23720 35936
rect 23784 35872 23792 35936
rect 23472 35871 23792 35872
rect 13905 35864 19675 35866
rect 13905 35808 13910 35864
rect 13966 35808 19614 35864
rect 19670 35808 19675 35864
rect 13905 35806 19675 35808
rect 13905 35803 13971 35806
rect 19609 35803 19675 35806
rect 19750 35806 22340 35866
rect 24209 35866 24275 35869
rect 30465 35866 30531 35869
rect 24209 35864 30531 35866
rect 24209 35808 24214 35864
rect 24270 35808 30470 35864
rect 30526 35808 30531 35864
rect 24209 35806 30531 35808
rect 16297 35730 16363 35733
rect 19750 35730 19810 35806
rect 24209 35803 24275 35806
rect 30465 35803 30531 35806
rect 16297 35728 19810 35730
rect 16297 35672 16302 35728
rect 16358 35672 19810 35728
rect 16297 35670 19810 35672
rect 20437 35730 20503 35733
rect 25313 35730 25379 35733
rect 20437 35728 25379 35730
rect 20437 35672 20442 35728
rect 20498 35672 25318 35728
rect 25374 35672 25379 35728
rect 20437 35670 25379 35672
rect 16297 35667 16363 35670
rect 20437 35667 20503 35670
rect 25313 35667 25379 35670
rect 26233 35730 26299 35733
rect 29453 35730 29519 35733
rect 26233 35728 29519 35730
rect 26233 35672 26238 35728
rect 26294 35672 29458 35728
rect 29514 35672 29519 35728
rect 26233 35670 29519 35672
rect 26233 35667 26299 35670
rect 29453 35667 29519 35670
rect 12525 35594 12591 35597
rect 17350 35594 17356 35596
rect 12525 35592 17356 35594
rect 0 35458 800 35548
rect 12525 35536 12530 35592
rect 12586 35536 17356 35592
rect 12525 35534 17356 35536
rect 12525 35531 12591 35534
rect 17350 35532 17356 35534
rect 17420 35532 17426 35596
rect 18321 35594 18387 35597
rect 17496 35592 18387 35594
rect 17496 35536 18326 35592
rect 18382 35536 18387 35592
rect 17496 35534 18387 35536
rect 2773 35458 2839 35461
rect 0 35456 2839 35458
rect 0 35400 2778 35456
rect 2834 35400 2839 35456
rect 0 35398 2839 35400
rect 0 35308 800 35398
rect 2773 35395 2839 35398
rect 14457 35458 14523 35461
rect 15929 35458 15995 35461
rect 16757 35458 16823 35461
rect 14457 35456 16823 35458
rect 14457 35400 14462 35456
rect 14518 35400 15934 35456
rect 15990 35400 16762 35456
rect 16818 35400 16823 35456
rect 14457 35398 16823 35400
rect 14457 35395 14523 35398
rect 15929 35395 15995 35398
rect 16757 35395 16823 35398
rect 17033 35458 17099 35461
rect 17496 35458 17556 35534
rect 18321 35531 18387 35534
rect 18505 35594 18571 35597
rect 20345 35594 20411 35597
rect 18505 35592 20411 35594
rect 18505 35536 18510 35592
rect 18566 35536 20350 35592
rect 20406 35536 20411 35592
rect 18505 35534 20411 35536
rect 18505 35531 18571 35534
rect 20345 35531 20411 35534
rect 21081 35594 21147 35597
rect 31293 35594 31359 35597
rect 21081 35592 31359 35594
rect 21081 35536 21086 35592
rect 21142 35536 31298 35592
rect 31354 35536 31359 35592
rect 21081 35534 31359 35536
rect 21081 35531 21147 35534
rect 31293 35531 31359 35534
rect 17033 35456 17556 35458
rect 17033 35400 17038 35456
rect 17094 35400 17556 35456
rect 17033 35398 17556 35400
rect 20989 35458 21055 35461
rect 28901 35458 28967 35461
rect 20989 35456 28967 35458
rect 20989 35400 20994 35456
rect 21050 35400 28906 35456
rect 28962 35400 28967 35456
rect 20989 35398 28967 35400
rect 17033 35395 17099 35398
rect 20989 35395 21055 35398
rect 28901 35395 28967 35398
rect 6576 35392 6896 35393
rect 6576 35328 6584 35392
rect 6648 35328 6664 35392
rect 6728 35328 6744 35392
rect 6808 35328 6824 35392
rect 6888 35328 6896 35392
rect 6576 35327 6896 35328
rect 17840 35392 18160 35393
rect 17840 35328 17848 35392
rect 17912 35328 17928 35392
rect 17992 35328 18008 35392
rect 18072 35328 18088 35392
rect 18152 35328 18160 35392
rect 17840 35327 18160 35328
rect 29104 35392 29424 35393
rect 29104 35328 29112 35392
rect 29176 35328 29192 35392
rect 29256 35328 29272 35392
rect 29336 35328 29352 35392
rect 29416 35328 29424 35392
rect 29104 35327 29424 35328
rect 13261 35322 13327 35325
rect 17125 35322 17191 35325
rect 13261 35320 17191 35322
rect 13261 35264 13266 35320
rect 13322 35264 17130 35320
rect 17186 35264 17191 35320
rect 13261 35262 17191 35264
rect 13261 35259 13327 35262
rect 17125 35259 17191 35262
rect 17350 35260 17356 35324
rect 17420 35322 17426 35324
rect 17585 35322 17651 35325
rect 17420 35320 17651 35322
rect 17420 35264 17590 35320
rect 17646 35264 17651 35320
rect 17420 35262 17651 35264
rect 17420 35260 17426 35262
rect 17585 35259 17651 35262
rect 18321 35322 18387 35325
rect 26233 35322 26299 35325
rect 18321 35320 26299 35322
rect 18321 35264 18326 35320
rect 18382 35264 26238 35320
rect 26294 35264 26299 35320
rect 18321 35262 26299 35264
rect 18321 35259 18387 35262
rect 26233 35259 26299 35262
rect 13997 35186 14063 35189
rect 20069 35186 20135 35189
rect 13997 35184 20135 35186
rect 13997 35128 14002 35184
rect 14058 35128 20074 35184
rect 20130 35128 20135 35184
rect 13997 35126 20135 35128
rect 13997 35123 14063 35126
rect 20069 35123 20135 35126
rect 21633 35186 21699 35189
rect 24669 35186 24735 35189
rect 31569 35188 31635 35189
rect 21633 35184 24735 35186
rect 21633 35128 21638 35184
rect 21694 35128 24674 35184
rect 24730 35128 24735 35184
rect 21633 35126 24735 35128
rect 21633 35123 21699 35126
rect 24669 35123 24735 35126
rect 31518 35124 31524 35188
rect 31588 35186 31635 35188
rect 31588 35184 31680 35186
rect 31630 35128 31680 35184
rect 31588 35126 31680 35128
rect 31588 35124 31635 35126
rect 31569 35123 31635 35124
rect 14222 34988 14228 35052
rect 14292 35050 14298 35052
rect 14549 35050 14615 35053
rect 14292 35048 14615 35050
rect 14292 34992 14554 35048
rect 14610 34992 14615 35048
rect 14292 34990 14615 34992
rect 14292 34988 14298 34990
rect 14549 34987 14615 34990
rect 15009 35050 15075 35053
rect 15326 35050 15332 35052
rect 15009 35048 15332 35050
rect 15009 34992 15014 35048
rect 15070 34992 15332 35048
rect 15009 34990 15332 34992
rect 15009 34987 15075 34990
rect 15326 34988 15332 34990
rect 15396 34988 15402 35052
rect 15469 35050 15535 35053
rect 18229 35050 18295 35053
rect 15469 35048 18295 35050
rect 15469 34992 15474 35048
rect 15530 34992 18234 35048
rect 18290 34992 18295 35048
rect 15469 34990 18295 34992
rect 15469 34987 15535 34990
rect 18229 34987 18295 34990
rect 18505 35050 18571 35053
rect 23565 35050 23631 35053
rect 18505 35048 23631 35050
rect 18505 34992 18510 35048
rect 18566 34992 23570 35048
rect 23626 34992 23631 35048
rect 18505 34990 23631 34992
rect 18505 34987 18571 34990
rect 23565 34987 23631 34990
rect 13169 34914 13235 34917
rect 24761 34914 24827 34917
rect 29913 34914 29979 34917
rect 13169 34912 23076 34914
rect 0 34628 800 34868
rect 13169 34856 13174 34912
rect 13230 34856 23076 34912
rect 13169 34854 23076 34856
rect 13169 34851 13235 34854
rect 12208 34848 12528 34849
rect 12208 34784 12216 34848
rect 12280 34784 12296 34848
rect 12360 34784 12376 34848
rect 12440 34784 12456 34848
rect 12520 34784 12528 34848
rect 12208 34783 12528 34784
rect 23016 34781 23076 34854
rect 24761 34912 29979 34914
rect 24761 34856 24766 34912
rect 24822 34856 29918 34912
rect 29974 34856 29979 34912
rect 24761 34854 29979 34856
rect 24761 34851 24827 34854
rect 29913 34851 29979 34854
rect 23472 34848 23792 34849
rect 23472 34784 23480 34848
rect 23544 34784 23560 34848
rect 23624 34784 23640 34848
rect 23704 34784 23720 34848
rect 23784 34784 23792 34848
rect 23472 34783 23792 34784
rect 12709 34780 12775 34781
rect 12709 34778 12756 34780
rect 12664 34776 12756 34778
rect 12664 34720 12714 34776
rect 12664 34718 12756 34720
rect 12709 34716 12756 34718
rect 12820 34716 12826 34780
rect 13353 34778 13419 34781
rect 15469 34778 15535 34781
rect 19701 34778 19767 34781
rect 13353 34776 15394 34778
rect 13353 34720 13358 34776
rect 13414 34720 15394 34776
rect 13353 34718 15394 34720
rect 12709 34715 12775 34716
rect 13353 34715 13419 34718
rect 14457 34642 14523 34645
rect 14590 34642 14596 34644
rect 14457 34640 14596 34642
rect 14457 34584 14462 34640
rect 14518 34584 14596 34640
rect 14457 34582 14596 34584
rect 14457 34579 14523 34582
rect 14590 34580 14596 34582
rect 14660 34580 14666 34644
rect 15334 34642 15394 34718
rect 15469 34776 19767 34778
rect 15469 34720 15474 34776
rect 15530 34720 19706 34776
rect 19762 34720 19767 34776
rect 15469 34718 19767 34720
rect 15469 34715 15535 34718
rect 19701 34715 19767 34718
rect 19977 34778 20043 34781
rect 22553 34778 22619 34781
rect 19977 34776 22619 34778
rect 19977 34720 19982 34776
rect 20038 34720 22558 34776
rect 22614 34720 22619 34776
rect 19977 34718 22619 34720
rect 19977 34715 20043 34718
rect 22553 34715 22619 34718
rect 23013 34776 23079 34781
rect 23013 34720 23018 34776
rect 23074 34720 23079 34776
rect 23013 34715 23079 34720
rect 29361 34778 29427 34781
rect 33225 34778 33291 34781
rect 29361 34776 33291 34778
rect 29361 34720 29366 34776
rect 29422 34720 33230 34776
rect 33286 34720 33291 34776
rect 29361 34718 33291 34720
rect 29361 34715 29427 34718
rect 33225 34715 33291 34718
rect 34145 34778 34211 34781
rect 35200 34778 36000 34868
rect 34145 34776 36000 34778
rect 34145 34720 34150 34776
rect 34206 34720 36000 34776
rect 34145 34718 36000 34720
rect 34145 34715 34211 34718
rect 21081 34642 21147 34645
rect 15334 34640 21147 34642
rect 15334 34584 21086 34640
rect 21142 34584 21147 34640
rect 35200 34628 36000 34718
rect 15334 34582 21147 34584
rect 21081 34579 21147 34582
rect 12249 34506 12315 34509
rect 32305 34506 32371 34509
rect 12249 34504 32371 34506
rect 12249 34448 12254 34504
rect 12310 34448 32310 34504
rect 32366 34448 32371 34504
rect 12249 34446 32371 34448
rect 12249 34443 12315 34446
rect 32305 34443 32371 34446
rect 12893 34370 12959 34373
rect 17677 34370 17743 34373
rect 12893 34368 17743 34370
rect 12893 34312 12898 34368
rect 12954 34312 17682 34368
rect 17738 34312 17743 34368
rect 12893 34310 17743 34312
rect 12893 34307 12959 34310
rect 17677 34307 17743 34310
rect 18321 34370 18387 34373
rect 24761 34370 24827 34373
rect 18321 34368 24827 34370
rect 18321 34312 18326 34368
rect 18382 34312 24766 34368
rect 24822 34312 24827 34368
rect 18321 34310 24827 34312
rect 18321 34307 18387 34310
rect 24761 34307 24827 34310
rect 6576 34304 6896 34305
rect 6576 34240 6584 34304
rect 6648 34240 6664 34304
rect 6728 34240 6744 34304
rect 6808 34240 6824 34304
rect 6888 34240 6896 34304
rect 6576 34239 6896 34240
rect 17840 34304 18160 34305
rect 17840 34240 17848 34304
rect 17912 34240 17928 34304
rect 17992 34240 18008 34304
rect 18072 34240 18088 34304
rect 18152 34240 18160 34304
rect 17840 34239 18160 34240
rect 29104 34304 29424 34305
rect 29104 34240 29112 34304
rect 29176 34240 29192 34304
rect 29256 34240 29272 34304
rect 29336 34240 29352 34304
rect 29416 34240 29424 34304
rect 29104 34239 29424 34240
rect 12709 34234 12775 34237
rect 16941 34234 17007 34237
rect 12709 34232 17007 34234
rect 0 34098 800 34188
rect 12709 34176 12714 34232
rect 12770 34176 16946 34232
rect 17002 34176 17007 34232
rect 12709 34174 17007 34176
rect 12709 34171 12775 34174
rect 16941 34171 17007 34174
rect 18454 34172 18460 34236
rect 18524 34234 18530 34236
rect 21357 34234 21423 34237
rect 18524 34232 21423 34234
rect 18524 34176 21362 34232
rect 21418 34176 21423 34232
rect 18524 34174 21423 34176
rect 18524 34172 18530 34174
rect 21357 34171 21423 34174
rect 21541 34234 21607 34237
rect 25497 34234 25563 34237
rect 21541 34232 25563 34234
rect 21541 34176 21546 34232
rect 21602 34176 25502 34232
rect 25558 34176 25563 34232
rect 21541 34174 25563 34176
rect 21541 34171 21607 34174
rect 25497 34171 25563 34174
rect 2773 34098 2839 34101
rect 0 34096 2839 34098
rect 0 34040 2778 34096
rect 2834 34040 2839 34096
rect 0 34038 2839 34040
rect 0 33948 800 34038
rect 2773 34035 2839 34038
rect 13261 34098 13327 34101
rect 14549 34100 14615 34101
rect 14222 34098 14228 34100
rect 13261 34096 14228 34098
rect 13261 34040 13266 34096
rect 13322 34040 14228 34096
rect 13261 34038 14228 34040
rect 13261 34035 13327 34038
rect 14222 34036 14228 34038
rect 14292 34036 14298 34100
rect 14549 34098 14596 34100
rect 14504 34096 14596 34098
rect 14504 34040 14554 34096
rect 14504 34038 14596 34040
rect 14549 34036 14596 34038
rect 14660 34036 14666 34100
rect 14917 34098 14983 34101
rect 15285 34098 15351 34101
rect 14917 34096 15351 34098
rect 14917 34040 14922 34096
rect 14978 34040 15290 34096
rect 15346 34040 15351 34096
rect 14917 34038 15351 34040
rect 14549 34035 14615 34036
rect 14917 34035 14983 34038
rect 15285 34035 15351 34038
rect 15745 34098 15811 34101
rect 20253 34098 20319 34101
rect 15745 34096 20319 34098
rect 15745 34040 15750 34096
rect 15806 34040 20258 34096
rect 20314 34040 20319 34096
rect 15745 34038 20319 34040
rect 15745 34035 15811 34038
rect 20253 34035 20319 34038
rect 20529 34098 20595 34101
rect 24853 34098 24919 34101
rect 20529 34096 24919 34098
rect 20529 34040 20534 34096
rect 20590 34040 24858 34096
rect 24914 34040 24919 34096
rect 20529 34038 24919 34040
rect 20529 34035 20595 34038
rect 24853 34035 24919 34038
rect 26049 34098 26115 34101
rect 29269 34098 29335 34101
rect 26049 34096 29335 34098
rect 26049 34040 26054 34096
rect 26110 34040 29274 34096
rect 29330 34040 29335 34096
rect 26049 34038 29335 34040
rect 26049 34035 26115 34038
rect 29269 34035 29335 34038
rect 34145 34098 34211 34101
rect 35200 34098 36000 34188
rect 34145 34096 36000 34098
rect 34145 34040 34150 34096
rect 34206 34040 36000 34096
rect 34145 34038 36000 34040
rect 34145 34035 34211 34038
rect 13445 33962 13511 33965
rect 15878 33962 15884 33964
rect 13445 33960 15884 33962
rect 13445 33904 13450 33960
rect 13506 33904 15884 33960
rect 13445 33902 15884 33904
rect 13445 33899 13511 33902
rect 15878 33900 15884 33902
rect 15948 33900 15954 33964
rect 16297 33962 16363 33965
rect 31845 33962 31911 33965
rect 16297 33960 31911 33962
rect 16297 33904 16302 33960
rect 16358 33904 31850 33960
rect 31906 33904 31911 33960
rect 35200 33948 36000 34038
rect 16297 33902 31911 33904
rect 16297 33899 16363 33902
rect 31845 33899 31911 33902
rect 14549 33826 14615 33829
rect 20713 33826 20779 33829
rect 14549 33824 20779 33826
rect 14549 33768 14554 33824
rect 14610 33768 20718 33824
rect 20774 33768 20779 33824
rect 14549 33766 20779 33768
rect 14549 33763 14615 33766
rect 20713 33763 20779 33766
rect 20846 33764 20852 33828
rect 20916 33826 20922 33828
rect 21173 33826 21239 33829
rect 20916 33824 21239 33826
rect 20916 33768 21178 33824
rect 21234 33768 21239 33824
rect 20916 33766 21239 33768
rect 20916 33764 20922 33766
rect 21173 33763 21239 33766
rect 21817 33826 21883 33829
rect 22277 33826 22343 33829
rect 21817 33824 22343 33826
rect 21817 33768 21822 33824
rect 21878 33768 22282 33824
rect 22338 33768 22343 33824
rect 21817 33766 22343 33768
rect 21817 33763 21883 33766
rect 22277 33763 22343 33766
rect 24117 33826 24183 33829
rect 25129 33826 25195 33829
rect 24117 33824 25195 33826
rect 24117 33768 24122 33824
rect 24178 33768 25134 33824
rect 25190 33768 25195 33824
rect 24117 33766 25195 33768
rect 24117 33763 24183 33766
rect 25129 33763 25195 33766
rect 12208 33760 12528 33761
rect 12208 33696 12216 33760
rect 12280 33696 12296 33760
rect 12360 33696 12376 33760
rect 12440 33696 12456 33760
rect 12520 33696 12528 33760
rect 12208 33695 12528 33696
rect 23472 33760 23792 33761
rect 23472 33696 23480 33760
rect 23544 33696 23560 33760
rect 23624 33696 23640 33760
rect 23704 33696 23720 33760
rect 23784 33696 23792 33760
rect 23472 33695 23792 33696
rect 14457 33690 14523 33693
rect 18454 33690 18460 33692
rect 14457 33688 18460 33690
rect 14457 33632 14462 33688
rect 14518 33632 18460 33688
rect 14457 33630 18460 33632
rect 14457 33627 14523 33630
rect 18454 33628 18460 33630
rect 18524 33628 18530 33692
rect 18689 33690 18755 33693
rect 20069 33690 20135 33693
rect 18689 33688 20135 33690
rect 18689 33632 18694 33688
rect 18750 33632 20074 33688
rect 20130 33632 20135 33688
rect 18689 33630 20135 33632
rect 18689 33627 18755 33630
rect 20069 33627 20135 33630
rect 20897 33690 20963 33693
rect 21541 33690 21607 33693
rect 20897 33688 21607 33690
rect 20897 33632 20902 33688
rect 20958 33632 21546 33688
rect 21602 33632 21607 33688
rect 20897 33630 21607 33632
rect 20897 33627 20963 33630
rect 21541 33627 21607 33630
rect 21725 33690 21791 33693
rect 23289 33690 23355 33693
rect 21725 33688 23355 33690
rect 21725 33632 21730 33688
rect 21786 33632 23294 33688
rect 23350 33632 23355 33688
rect 21725 33630 23355 33632
rect 21725 33627 21791 33630
rect 23289 33627 23355 33630
rect 12617 33554 12683 33557
rect 15561 33554 15627 33557
rect 12617 33552 15627 33554
rect 12617 33496 12622 33552
rect 12678 33496 15566 33552
rect 15622 33496 15627 33552
rect 12617 33494 15627 33496
rect 12617 33491 12683 33494
rect 15561 33491 15627 33494
rect 15878 33492 15884 33556
rect 15948 33554 15954 33556
rect 27337 33554 27403 33557
rect 15948 33552 27403 33554
rect 15948 33496 27342 33552
rect 27398 33496 27403 33552
rect 15948 33494 27403 33496
rect 15948 33492 15954 33494
rect 27337 33491 27403 33494
rect 27797 33554 27863 33557
rect 29453 33554 29519 33557
rect 27797 33552 29519 33554
rect 27797 33496 27802 33552
rect 27858 33496 29458 33552
rect 29514 33496 29519 33552
rect 27797 33494 29519 33496
rect 27797 33491 27863 33494
rect 29453 33491 29519 33494
rect 13905 33418 13971 33421
rect 14457 33418 14523 33421
rect 13905 33416 14523 33418
rect 13905 33360 13910 33416
rect 13966 33360 14462 33416
rect 14518 33360 14523 33416
rect 13905 33358 14523 33360
rect 13905 33355 13971 33358
rect 14457 33355 14523 33358
rect 14641 33418 14707 33421
rect 15653 33418 15719 33421
rect 14641 33416 15719 33418
rect 14641 33360 14646 33416
rect 14702 33360 15658 33416
rect 15714 33360 15719 33416
rect 14641 33358 15719 33360
rect 14641 33355 14707 33358
rect 15653 33355 15719 33358
rect 15929 33418 15995 33421
rect 17493 33418 17559 33421
rect 18270 33418 18276 33420
rect 15929 33416 17559 33418
rect 15929 33360 15934 33416
rect 15990 33360 17498 33416
rect 17554 33360 17559 33416
rect 15929 33358 17559 33360
rect 15929 33355 15995 33358
rect 17493 33355 17559 33358
rect 17680 33358 18276 33418
rect 12801 33282 12867 33285
rect 17680 33282 17740 33358
rect 18270 33356 18276 33358
rect 18340 33356 18346 33420
rect 18454 33356 18460 33420
rect 18524 33418 18530 33420
rect 23381 33418 23447 33421
rect 31569 33420 31635 33421
rect 31518 33418 31524 33420
rect 18524 33358 23306 33418
rect 18524 33356 18530 33358
rect 12801 33280 17740 33282
rect 12801 33224 12806 33280
rect 12862 33224 17740 33280
rect 12801 33222 17740 33224
rect 12801 33219 12867 33222
rect 18270 33220 18276 33284
rect 18340 33282 18346 33284
rect 19425 33282 19491 33285
rect 18340 33280 19491 33282
rect 18340 33224 19430 33280
rect 19486 33224 19491 33280
rect 18340 33222 19491 33224
rect 18340 33220 18346 33222
rect 19425 33219 19491 33222
rect 19609 33282 19675 33285
rect 23105 33282 23171 33285
rect 19609 33280 23171 33282
rect 19609 33224 19614 33280
rect 19670 33224 23110 33280
rect 23166 33224 23171 33280
rect 19609 33222 23171 33224
rect 23246 33282 23306 33358
rect 23381 33416 30804 33418
rect 23381 33360 23386 33416
rect 23442 33360 30804 33416
rect 23381 33358 30804 33360
rect 31478 33358 31524 33418
rect 31588 33416 31635 33420
rect 31630 33360 31635 33416
rect 23381 33355 23447 33358
rect 25957 33282 26023 33285
rect 23246 33280 26023 33282
rect 23246 33224 25962 33280
rect 26018 33224 26023 33280
rect 23246 33222 26023 33224
rect 19609 33219 19675 33222
rect 23105 33219 23171 33222
rect 25957 33219 26023 33222
rect 26141 33282 26207 33285
rect 28717 33282 28783 33285
rect 26141 33280 28783 33282
rect 26141 33224 26146 33280
rect 26202 33224 28722 33280
rect 28778 33224 28783 33280
rect 26141 33222 28783 33224
rect 30744 33282 30804 33358
rect 31518 33356 31524 33358
rect 31588 33356 31635 33360
rect 31569 33355 31635 33356
rect 34145 33418 34211 33421
rect 35200 33418 36000 33508
rect 34145 33416 36000 33418
rect 34145 33360 34150 33416
rect 34206 33360 36000 33416
rect 34145 33358 36000 33360
rect 34145 33355 34211 33358
rect 32581 33282 32647 33285
rect 30744 33280 32647 33282
rect 30744 33224 32586 33280
rect 32642 33224 32647 33280
rect 35200 33268 36000 33358
rect 30744 33222 32647 33224
rect 26141 33219 26207 33222
rect 28717 33219 28783 33222
rect 32581 33219 32647 33222
rect 6576 33216 6896 33217
rect 6576 33152 6584 33216
rect 6648 33152 6664 33216
rect 6728 33152 6744 33216
rect 6808 33152 6824 33216
rect 6888 33152 6896 33216
rect 6576 33151 6896 33152
rect 17840 33216 18160 33217
rect 17840 33152 17848 33216
rect 17912 33152 17928 33216
rect 17992 33152 18008 33216
rect 18072 33152 18088 33216
rect 18152 33152 18160 33216
rect 17840 33151 18160 33152
rect 29104 33216 29424 33217
rect 29104 33152 29112 33216
rect 29176 33152 29192 33216
rect 29256 33152 29272 33216
rect 29336 33152 29352 33216
rect 29416 33152 29424 33216
rect 29104 33151 29424 33152
rect 13629 33146 13695 33149
rect 13629 33144 16268 33146
rect 13629 33088 13634 33144
rect 13690 33088 16268 33144
rect 13629 33086 16268 33088
rect 13629 33083 13695 33086
rect 13353 33010 13419 33013
rect 16062 33010 16068 33012
rect 13353 33008 16068 33010
rect 13353 32952 13358 33008
rect 13414 32952 16068 33008
rect 13353 32950 16068 32952
rect 13353 32947 13419 32950
rect 16062 32948 16068 32950
rect 16132 32948 16138 33012
rect 16208 33010 16268 33086
rect 16430 33084 16436 33148
rect 16500 33146 16506 33148
rect 17401 33146 17467 33149
rect 16500 33144 17467 33146
rect 16500 33088 17406 33144
rect 17462 33088 17467 33144
rect 16500 33086 17467 33088
rect 16500 33084 16506 33086
rect 17401 33083 17467 33086
rect 18597 33146 18663 33149
rect 20345 33146 20411 33149
rect 18597 33144 20411 33146
rect 18597 33088 18602 33144
rect 18658 33088 20350 33144
rect 20406 33088 20411 33144
rect 18597 33086 20411 33088
rect 18597 33083 18663 33086
rect 20345 33083 20411 33086
rect 22921 33146 22987 33149
rect 28625 33146 28691 33149
rect 22921 33144 28691 33146
rect 22921 33088 22926 33144
rect 22982 33088 28630 33144
rect 28686 33088 28691 33144
rect 22921 33086 28691 33088
rect 22921 33083 22987 33086
rect 28625 33083 28691 33086
rect 17588 33010 17970 33044
rect 20897 33010 20963 33013
rect 16208 33008 20963 33010
rect 16208 32984 20902 33008
rect 16208 32950 17648 32984
rect 17910 32952 20902 32984
rect 20958 32952 20963 33008
rect 17910 32950 20963 32952
rect 20897 32947 20963 32950
rect 21081 33010 21147 33013
rect 32029 33010 32095 33013
rect 21081 33008 32095 33010
rect 21081 32952 21086 33008
rect 21142 32952 32034 33008
rect 32090 32952 32095 33008
rect 21081 32950 32095 32952
rect 21081 32947 21147 32950
rect 32029 32947 32095 32950
rect 13997 32874 14063 32877
rect 17677 32874 17743 32877
rect 13997 32872 17743 32874
rect 0 32588 800 32828
rect 13997 32816 14002 32872
rect 14058 32816 17682 32872
rect 17738 32816 17743 32872
rect 13997 32814 17743 32816
rect 13997 32811 14063 32814
rect 17677 32811 17743 32814
rect 17953 32874 18019 32877
rect 21357 32874 21423 32877
rect 22277 32874 22343 32877
rect 25221 32874 25287 32877
rect 29729 32874 29795 32877
rect 17953 32872 20730 32874
rect 17953 32816 17958 32872
rect 18014 32816 20730 32872
rect 17953 32814 20730 32816
rect 17953 32811 18019 32814
rect 12985 32738 13051 32741
rect 12985 32736 17418 32738
rect 12985 32680 12990 32736
rect 13046 32680 17418 32736
rect 12985 32678 17418 32680
rect 12985 32675 13051 32678
rect 12208 32672 12528 32673
rect 12208 32608 12216 32672
rect 12280 32608 12296 32672
rect 12360 32608 12376 32672
rect 12440 32608 12456 32672
rect 12520 32608 12528 32672
rect 12208 32607 12528 32608
rect 14089 32602 14155 32605
rect 14273 32602 14339 32605
rect 14089 32600 14339 32602
rect 14089 32544 14094 32600
rect 14150 32544 14278 32600
rect 14334 32544 14339 32600
rect 14089 32542 14339 32544
rect 14089 32539 14155 32542
rect 14273 32539 14339 32542
rect 14549 32602 14615 32605
rect 17217 32602 17283 32605
rect 14549 32600 17283 32602
rect 14549 32544 14554 32600
rect 14610 32544 17222 32600
rect 17278 32544 17283 32600
rect 14549 32542 17283 32544
rect 17358 32602 17418 32678
rect 17534 32676 17540 32740
rect 17604 32738 17610 32740
rect 18270 32738 18276 32740
rect 17604 32678 18276 32738
rect 17604 32676 17610 32678
rect 18270 32676 18276 32678
rect 18340 32676 18346 32740
rect 18413 32738 18479 32741
rect 19977 32738 20043 32741
rect 18413 32736 20043 32738
rect 18413 32680 18418 32736
rect 18474 32680 19982 32736
rect 20038 32680 20043 32736
rect 18413 32678 20043 32680
rect 20670 32738 20730 32814
rect 21357 32872 22343 32874
rect 21357 32816 21362 32872
rect 21418 32816 22282 32872
rect 22338 32816 22343 32872
rect 21357 32814 22343 32816
rect 21357 32811 21423 32814
rect 22277 32811 22343 32814
rect 22510 32814 24870 32874
rect 22369 32738 22435 32741
rect 20670 32736 22435 32738
rect 20670 32680 22374 32736
rect 22430 32680 22435 32736
rect 20670 32678 22435 32680
rect 18413 32675 18479 32678
rect 19977 32675 20043 32678
rect 22369 32675 22435 32678
rect 21909 32602 21975 32605
rect 17358 32600 21975 32602
rect 17358 32544 21914 32600
rect 21970 32544 21975 32600
rect 17358 32542 21975 32544
rect 14549 32539 14615 32542
rect 17217 32539 17283 32542
rect 21909 32539 21975 32542
rect 22185 32602 22251 32605
rect 22510 32602 22570 32814
rect 24810 32738 24870 32814
rect 25221 32872 29795 32874
rect 25221 32816 25226 32872
rect 25282 32816 29734 32872
rect 29790 32816 29795 32872
rect 25221 32814 29795 32816
rect 25221 32811 25287 32814
rect 29729 32811 29795 32814
rect 29913 32874 29979 32877
rect 30373 32874 30439 32877
rect 29913 32872 30439 32874
rect 29913 32816 29918 32872
rect 29974 32816 30378 32872
rect 30434 32816 30439 32872
rect 29913 32814 30439 32816
rect 29913 32811 29979 32814
rect 30373 32811 30439 32814
rect 27889 32738 27955 32741
rect 30649 32738 30715 32741
rect 24810 32736 30715 32738
rect 24810 32680 27894 32736
rect 27950 32680 30654 32736
rect 30710 32680 30715 32736
rect 24810 32678 30715 32680
rect 27889 32675 27955 32678
rect 30649 32675 30715 32678
rect 34145 32738 34211 32741
rect 35200 32738 36000 32828
rect 34145 32736 36000 32738
rect 34145 32680 34150 32736
rect 34206 32680 36000 32736
rect 34145 32678 36000 32680
rect 34145 32675 34211 32678
rect 23472 32672 23792 32673
rect 23472 32608 23480 32672
rect 23544 32608 23560 32672
rect 23624 32608 23640 32672
rect 23704 32608 23720 32672
rect 23784 32608 23792 32672
rect 23472 32607 23792 32608
rect 22185 32600 22570 32602
rect 22185 32544 22190 32600
rect 22246 32544 22570 32600
rect 22185 32542 22570 32544
rect 22645 32602 22711 32605
rect 23197 32602 23263 32605
rect 22645 32600 23263 32602
rect 22645 32544 22650 32600
rect 22706 32544 23202 32600
rect 23258 32544 23263 32600
rect 22645 32542 23263 32544
rect 22185 32539 22251 32542
rect 22645 32539 22711 32542
rect 23197 32539 23263 32542
rect 25313 32602 25379 32605
rect 33133 32602 33199 32605
rect 25313 32600 33199 32602
rect 25313 32544 25318 32600
rect 25374 32544 33138 32600
rect 33194 32544 33199 32600
rect 35200 32588 36000 32678
rect 25313 32542 33199 32544
rect 25313 32539 25379 32542
rect 33133 32539 33199 32542
rect 12801 32466 12867 32469
rect 18454 32466 18460 32468
rect 12801 32464 18460 32466
rect 12801 32408 12806 32464
rect 12862 32408 18460 32464
rect 12801 32406 18460 32408
rect 12801 32403 12867 32406
rect 18454 32404 18460 32406
rect 18524 32404 18530 32468
rect 18638 32404 18644 32468
rect 18708 32466 18714 32468
rect 18965 32466 19031 32469
rect 18708 32464 19031 32466
rect 18708 32408 18970 32464
rect 19026 32408 19031 32464
rect 18708 32406 19031 32408
rect 18708 32404 18714 32406
rect 18965 32403 19031 32406
rect 19149 32466 19215 32469
rect 19885 32466 19951 32469
rect 19149 32464 19951 32466
rect 19149 32408 19154 32464
rect 19210 32408 19890 32464
rect 19946 32408 19951 32464
rect 19149 32406 19951 32408
rect 19149 32403 19215 32406
rect 19885 32403 19951 32406
rect 20069 32466 20135 32469
rect 32305 32466 32371 32469
rect 20069 32464 32371 32466
rect 20069 32408 20074 32464
rect 20130 32408 32310 32464
rect 32366 32408 32371 32464
rect 20069 32406 32371 32408
rect 20069 32403 20135 32406
rect 32305 32403 32371 32406
rect 11789 32330 11855 32333
rect 32305 32330 32371 32333
rect 11789 32328 32371 32330
rect 11789 32272 11794 32328
rect 11850 32272 32310 32328
rect 32366 32272 32371 32328
rect 11789 32270 32371 32272
rect 11789 32267 11855 32270
rect 32305 32267 32371 32270
rect 13261 32194 13327 32197
rect 14774 32194 14780 32196
rect 13261 32192 14780 32194
rect 0 32058 800 32148
rect 13261 32136 13266 32192
rect 13322 32136 14780 32192
rect 13261 32134 14780 32136
rect 13261 32131 13327 32134
rect 14774 32132 14780 32134
rect 14844 32132 14850 32196
rect 14917 32194 14983 32197
rect 17217 32194 17283 32197
rect 14917 32192 17283 32194
rect 14917 32136 14922 32192
rect 14978 32136 17222 32192
rect 17278 32136 17283 32192
rect 14917 32134 17283 32136
rect 14917 32131 14983 32134
rect 17217 32131 17283 32134
rect 17350 32132 17356 32196
rect 17420 32194 17426 32196
rect 17677 32194 17743 32197
rect 17420 32192 17743 32194
rect 17420 32136 17682 32192
rect 17738 32136 17743 32192
rect 17420 32134 17743 32136
rect 17420 32132 17426 32134
rect 17677 32131 17743 32134
rect 18229 32196 18295 32197
rect 18229 32192 18276 32196
rect 18340 32194 18346 32196
rect 18229 32136 18234 32192
rect 18229 32132 18276 32136
rect 18340 32134 18386 32194
rect 18340 32132 18346 32134
rect 18454 32132 18460 32196
rect 18524 32194 18530 32196
rect 24945 32194 25011 32197
rect 18524 32192 25011 32194
rect 18524 32136 24950 32192
rect 25006 32136 25011 32192
rect 18524 32134 25011 32136
rect 18524 32132 18530 32134
rect 18229 32131 18295 32132
rect 24945 32131 25011 32134
rect 28073 32194 28139 32197
rect 28809 32194 28875 32197
rect 30465 32196 30531 32197
rect 30833 32196 30899 32197
rect 30414 32194 30420 32196
rect 28073 32192 28875 32194
rect 28073 32136 28078 32192
rect 28134 32136 28814 32192
rect 28870 32136 28875 32192
rect 28073 32134 28875 32136
rect 30374 32134 30420 32194
rect 30484 32192 30531 32196
rect 30782 32194 30788 32196
rect 30526 32136 30531 32192
rect 28073 32131 28139 32134
rect 28809 32131 28875 32134
rect 30414 32132 30420 32134
rect 30484 32132 30531 32136
rect 30742 32134 30788 32194
rect 30852 32192 30899 32196
rect 30894 32136 30899 32192
rect 30782 32132 30788 32134
rect 30852 32132 30899 32136
rect 30465 32131 30531 32132
rect 30833 32131 30899 32132
rect 6576 32128 6896 32129
rect 6576 32064 6584 32128
rect 6648 32064 6664 32128
rect 6728 32064 6744 32128
rect 6808 32064 6824 32128
rect 6888 32064 6896 32128
rect 6576 32063 6896 32064
rect 17840 32128 18160 32129
rect 17840 32064 17848 32128
rect 17912 32064 17928 32128
rect 17992 32064 18008 32128
rect 18072 32064 18088 32128
rect 18152 32064 18160 32128
rect 17840 32063 18160 32064
rect 29104 32128 29424 32129
rect 29104 32064 29112 32128
rect 29176 32064 29192 32128
rect 29256 32064 29272 32128
rect 29336 32064 29352 32128
rect 29416 32064 29424 32128
rect 29104 32063 29424 32064
rect 3417 32058 3483 32061
rect 0 32056 3483 32058
rect 0 32000 3422 32056
rect 3478 32000 3483 32056
rect 0 31998 3483 32000
rect 0 31908 800 31998
rect 3417 31995 3483 31998
rect 14733 32058 14799 32061
rect 16757 32058 16823 32061
rect 14733 32056 16823 32058
rect 14733 32000 14738 32056
rect 14794 32000 16762 32056
rect 16818 32000 16823 32056
rect 14733 31998 16823 32000
rect 14733 31995 14799 31998
rect 16757 31995 16823 31998
rect 17125 32058 17191 32061
rect 17677 32058 17743 32061
rect 17125 32056 17743 32058
rect 17125 32000 17130 32056
rect 17186 32000 17682 32056
rect 17738 32000 17743 32056
rect 17125 31998 17743 32000
rect 17125 31995 17191 31998
rect 17677 31995 17743 31998
rect 18822 31996 18828 32060
rect 18892 32058 18898 32060
rect 20161 32058 20227 32061
rect 18892 32056 20227 32058
rect 18892 32000 20166 32056
rect 20222 32000 20227 32056
rect 18892 31998 20227 32000
rect 18892 31996 18898 31998
rect 20161 31995 20227 31998
rect 20713 32058 20779 32061
rect 26325 32058 26391 32061
rect 20713 32056 26391 32058
rect 20713 32000 20718 32056
rect 20774 32000 26330 32056
rect 26386 32000 26391 32056
rect 20713 31998 26391 32000
rect 20713 31995 20779 31998
rect 26325 31995 26391 31998
rect 29545 32056 29611 32061
rect 29545 32000 29550 32056
rect 29606 32000 29611 32056
rect 29545 31995 29611 32000
rect 34145 32058 34211 32061
rect 35200 32058 36000 32148
rect 34145 32056 36000 32058
rect 34145 32000 34150 32056
rect 34206 32000 36000 32056
rect 34145 31998 36000 32000
rect 34145 31995 34211 31998
rect 13629 31922 13695 31925
rect 29361 31922 29427 31925
rect 29548 31922 29608 31995
rect 13629 31920 29010 31922
rect 13629 31864 13634 31920
rect 13690 31864 29010 31920
rect 13629 31862 29010 31864
rect 13629 31859 13695 31862
rect 12893 31786 12959 31789
rect 16246 31786 16252 31788
rect 12893 31784 16252 31786
rect 12893 31728 12898 31784
rect 12954 31728 16252 31784
rect 12893 31726 16252 31728
rect 12893 31723 12959 31726
rect 16246 31724 16252 31726
rect 16316 31724 16322 31788
rect 16430 31724 16436 31788
rect 16500 31786 16506 31788
rect 20069 31786 20135 31789
rect 16500 31784 20135 31786
rect 16500 31728 20074 31784
rect 20130 31728 20135 31784
rect 16500 31726 20135 31728
rect 16500 31724 16506 31726
rect 20069 31723 20135 31726
rect 20345 31786 20411 31789
rect 28073 31786 28139 31789
rect 20345 31784 28139 31786
rect 20345 31728 20350 31784
rect 20406 31728 28078 31784
rect 28134 31728 28139 31784
rect 20345 31726 28139 31728
rect 28950 31786 29010 31862
rect 29361 31920 29608 31922
rect 29361 31864 29366 31920
rect 29422 31864 29608 31920
rect 29361 31862 29608 31864
rect 30741 31922 30807 31925
rect 31385 31922 31451 31925
rect 30741 31920 31451 31922
rect 30741 31864 30746 31920
rect 30802 31864 31390 31920
rect 31446 31864 31451 31920
rect 35200 31908 36000 31998
rect 30741 31862 31451 31864
rect 29361 31859 29427 31862
rect 30741 31859 30807 31862
rect 31385 31859 31451 31862
rect 31477 31786 31543 31789
rect 28950 31784 31543 31786
rect 28950 31728 31482 31784
rect 31538 31728 31543 31784
rect 28950 31726 31543 31728
rect 20345 31723 20411 31726
rect 28073 31723 28139 31726
rect 31477 31723 31543 31726
rect 14181 31650 14247 31653
rect 19057 31650 19123 31653
rect 14181 31648 19123 31650
rect 14181 31592 14186 31648
rect 14242 31592 19062 31648
rect 19118 31592 19123 31648
rect 14181 31590 19123 31592
rect 14181 31587 14247 31590
rect 19057 31587 19123 31590
rect 19425 31650 19491 31653
rect 24117 31650 24183 31653
rect 27153 31650 27219 31653
rect 19425 31648 23306 31650
rect 19425 31592 19430 31648
rect 19486 31592 23306 31648
rect 19425 31590 23306 31592
rect 19425 31587 19491 31590
rect 12208 31584 12528 31585
rect 12208 31520 12216 31584
rect 12280 31520 12296 31584
rect 12360 31520 12376 31584
rect 12440 31520 12456 31584
rect 12520 31520 12528 31584
rect 12208 31519 12528 31520
rect 12709 31514 12775 31517
rect 14641 31514 14707 31517
rect 12709 31512 14707 31514
rect 0 31378 800 31468
rect 12709 31456 12714 31512
rect 12770 31456 14646 31512
rect 14702 31456 14707 31512
rect 12709 31454 14707 31456
rect 12709 31451 12775 31454
rect 14641 31451 14707 31454
rect 14825 31514 14891 31517
rect 16389 31514 16455 31517
rect 14825 31512 16455 31514
rect 14825 31456 14830 31512
rect 14886 31456 16394 31512
rect 16450 31456 16455 31512
rect 14825 31454 16455 31456
rect 14825 31451 14891 31454
rect 16389 31451 16455 31454
rect 17401 31514 17467 31517
rect 23105 31514 23171 31517
rect 17401 31512 23171 31514
rect 17401 31456 17406 31512
rect 17462 31456 23110 31512
rect 23166 31456 23171 31512
rect 17401 31454 23171 31456
rect 17401 31451 17467 31454
rect 23105 31451 23171 31454
rect 1945 31378 2011 31381
rect 0 31376 2011 31378
rect 0 31320 1950 31376
rect 2006 31320 2011 31376
rect 0 31318 2011 31320
rect 0 31228 800 31318
rect 1945 31315 2011 31318
rect 13629 31378 13695 31381
rect 15837 31378 15903 31381
rect 13629 31376 15903 31378
rect 13629 31320 13634 31376
rect 13690 31320 15842 31376
rect 15898 31320 15903 31376
rect 13629 31318 15903 31320
rect 13629 31315 13695 31318
rect 15837 31315 15903 31318
rect 16113 31378 16179 31381
rect 19333 31378 19399 31381
rect 16113 31376 19399 31378
rect 16113 31320 16118 31376
rect 16174 31320 19338 31376
rect 19394 31320 19399 31376
rect 16113 31318 19399 31320
rect 16113 31315 16179 31318
rect 19333 31315 19399 31318
rect 19609 31378 19675 31381
rect 23105 31378 23171 31381
rect 19609 31376 23171 31378
rect 19609 31320 19614 31376
rect 19670 31320 23110 31376
rect 23166 31320 23171 31376
rect 19609 31318 23171 31320
rect 23246 31378 23306 31590
rect 24117 31648 27219 31650
rect 24117 31592 24122 31648
rect 24178 31592 27158 31648
rect 27214 31592 27219 31648
rect 24117 31590 27219 31592
rect 24117 31587 24183 31590
rect 27153 31587 27219 31590
rect 29269 31650 29335 31653
rect 31017 31650 31083 31653
rect 29269 31648 31083 31650
rect 29269 31592 29274 31648
rect 29330 31592 31022 31648
rect 31078 31592 31083 31648
rect 29269 31590 31083 31592
rect 29269 31587 29335 31590
rect 31017 31587 31083 31590
rect 23472 31584 23792 31585
rect 23472 31520 23480 31584
rect 23544 31520 23560 31584
rect 23624 31520 23640 31584
rect 23704 31520 23720 31584
rect 23784 31520 23792 31584
rect 23472 31519 23792 31520
rect 25405 31514 25471 31517
rect 26233 31514 26299 31517
rect 25405 31512 26299 31514
rect 25405 31456 25410 31512
rect 25466 31456 26238 31512
rect 26294 31456 26299 31512
rect 25405 31454 26299 31456
rect 25405 31451 25471 31454
rect 26233 31451 26299 31454
rect 34145 31378 34211 31381
rect 35200 31378 36000 31468
rect 23246 31318 29562 31378
rect 19609 31315 19675 31318
rect 23105 31315 23171 31318
rect 14549 31242 14615 31245
rect 19885 31242 19951 31245
rect 14549 31240 19951 31242
rect 14549 31184 14554 31240
rect 14610 31184 19890 31240
rect 19946 31184 19951 31240
rect 14549 31182 19951 31184
rect 14549 31179 14615 31182
rect 19885 31179 19951 31182
rect 20253 31242 20319 31245
rect 28441 31242 28507 31245
rect 20253 31240 28507 31242
rect 20253 31184 20258 31240
rect 20314 31184 28446 31240
rect 28502 31184 28507 31240
rect 20253 31182 28507 31184
rect 20253 31179 20319 31182
rect 28441 31179 28507 31182
rect 12065 31106 12131 31109
rect 17217 31106 17283 31109
rect 17534 31106 17540 31108
rect 12065 31104 17540 31106
rect 12065 31048 12070 31104
rect 12126 31048 17222 31104
rect 17278 31048 17540 31104
rect 12065 31046 17540 31048
rect 12065 31043 12131 31046
rect 17217 31043 17283 31046
rect 17534 31044 17540 31046
rect 17604 31044 17610 31108
rect 17677 31104 17743 31109
rect 17677 31048 17682 31104
rect 17738 31048 17743 31104
rect 17677 31043 17743 31048
rect 18781 31106 18847 31109
rect 18781 31104 21604 31106
rect 18781 31048 18786 31104
rect 18842 31048 21604 31104
rect 18781 31046 21604 31048
rect 18781 31043 18847 31046
rect 6576 31040 6896 31041
rect 6576 30976 6584 31040
rect 6648 30976 6664 31040
rect 6728 30976 6744 31040
rect 6808 30976 6824 31040
rect 6888 30976 6896 31040
rect 6576 30975 6896 30976
rect 13261 30970 13327 30973
rect 17680 30970 17740 31043
rect 17840 31040 18160 31041
rect 17840 30976 17848 31040
rect 17912 30976 17928 31040
rect 17992 30976 18008 31040
rect 18072 30976 18088 31040
rect 18152 30976 18160 31040
rect 17840 30975 18160 30976
rect 13261 30968 17740 30970
rect 13261 30912 13266 30968
rect 13322 30912 17740 30968
rect 13261 30910 17740 30912
rect 18321 30970 18387 30973
rect 18454 30970 18460 30972
rect 18321 30968 18460 30970
rect 18321 30912 18326 30968
rect 18382 30912 18460 30968
rect 18321 30910 18460 30912
rect 13261 30907 13327 30910
rect 18321 30907 18387 30910
rect 18454 30908 18460 30910
rect 18524 30908 18530 30972
rect 18638 30908 18644 30972
rect 18708 30970 18714 30972
rect 21544 30970 21604 31046
rect 21766 31044 21772 31108
rect 21836 31106 21842 31108
rect 22737 31106 22803 31109
rect 21836 31104 22803 31106
rect 21836 31048 22742 31104
rect 22798 31048 22803 31104
rect 21836 31046 22803 31048
rect 21836 31044 21842 31046
rect 22737 31043 22803 31046
rect 23054 31044 23060 31108
rect 23124 31106 23130 31108
rect 25681 31106 25747 31109
rect 23124 31104 25747 31106
rect 23124 31048 25686 31104
rect 25742 31048 25747 31104
rect 23124 31046 25747 31048
rect 23124 31044 23130 31046
rect 25681 31043 25747 31046
rect 27654 31044 27660 31108
rect 27724 31106 27730 31108
rect 27981 31106 28047 31109
rect 27724 31104 28047 31106
rect 27724 31048 27986 31104
rect 28042 31048 28047 31104
rect 27724 31046 28047 31048
rect 29502 31106 29562 31318
rect 34145 31376 36000 31378
rect 34145 31320 34150 31376
rect 34206 31320 36000 31376
rect 34145 31318 36000 31320
rect 34145 31315 34211 31318
rect 32305 31242 32371 31245
rect 31710 31240 32371 31242
rect 31710 31184 32310 31240
rect 32366 31184 32371 31240
rect 35200 31228 36000 31318
rect 31710 31182 32371 31184
rect 31710 31106 31770 31182
rect 32305 31179 32371 31182
rect 29502 31046 31770 31106
rect 27724 31044 27730 31046
rect 27981 31043 28047 31046
rect 29104 31040 29424 31041
rect 29104 30976 29112 31040
rect 29176 30976 29192 31040
rect 29256 30976 29272 31040
rect 29336 30976 29352 31040
rect 29416 30976 29424 31040
rect 29104 30975 29424 30976
rect 28717 30970 28783 30973
rect 18708 30910 21420 30970
rect 21544 30968 28783 30970
rect 21544 30912 28722 30968
rect 28778 30912 28783 30968
rect 21544 30910 28783 30912
rect 18708 30908 18714 30910
rect 12801 30834 12867 30837
rect 21214 30834 21220 30836
rect 12801 30832 21220 30834
rect 0 30548 800 30788
rect 12801 30776 12806 30832
rect 12862 30776 21220 30832
rect 12801 30774 21220 30776
rect 12801 30771 12867 30774
rect 21214 30772 21220 30774
rect 21284 30772 21290 30836
rect 21360 30834 21420 30910
rect 28717 30907 28783 30910
rect 29729 30970 29795 30973
rect 33869 30970 33935 30973
rect 29729 30968 33935 30970
rect 29729 30912 29734 30968
rect 29790 30912 33874 30968
rect 33930 30912 33935 30968
rect 29729 30910 33935 30912
rect 29729 30907 29795 30910
rect 33869 30907 33935 30910
rect 28533 30834 28599 30837
rect 21360 30832 28599 30834
rect 21360 30776 28538 30832
rect 28594 30776 28599 30832
rect 21360 30774 28599 30776
rect 28533 30771 28599 30774
rect 30189 30834 30255 30837
rect 32305 30834 32371 30837
rect 30189 30832 32371 30834
rect 30189 30776 30194 30832
rect 30250 30776 32310 30832
rect 32366 30776 32371 30832
rect 30189 30774 32371 30776
rect 30189 30771 30255 30774
rect 32305 30771 32371 30774
rect 13169 30698 13235 30701
rect 21214 30698 21220 30700
rect 13169 30696 21220 30698
rect 13169 30640 13174 30696
rect 13230 30640 21220 30696
rect 13169 30638 21220 30640
rect 13169 30635 13235 30638
rect 21214 30636 21220 30638
rect 21284 30636 21290 30700
rect 21357 30698 21423 30701
rect 22829 30698 22895 30701
rect 26049 30698 26115 30701
rect 21357 30696 22895 30698
rect 21357 30640 21362 30696
rect 21418 30640 22834 30696
rect 22890 30640 22895 30696
rect 21357 30638 22895 30640
rect 21357 30635 21423 30638
rect 22829 30635 22895 30638
rect 23292 30696 26115 30698
rect 23292 30640 26054 30696
rect 26110 30640 26115 30696
rect 23292 30638 26115 30640
rect 14825 30562 14891 30565
rect 19425 30562 19491 30565
rect 23054 30562 23060 30564
rect 14825 30560 19304 30562
rect 14825 30504 14830 30560
rect 14886 30504 19304 30560
rect 14825 30502 19304 30504
rect 14825 30499 14891 30502
rect 12208 30496 12528 30497
rect 12208 30432 12216 30496
rect 12280 30432 12296 30496
rect 12360 30432 12376 30496
rect 12440 30432 12456 30496
rect 12520 30432 12528 30496
rect 12208 30431 12528 30432
rect 13445 30426 13511 30429
rect 16021 30426 16087 30429
rect 13445 30424 16087 30426
rect 13445 30368 13450 30424
rect 13506 30368 16026 30424
rect 16082 30368 16087 30424
rect 13445 30366 16087 30368
rect 13445 30363 13511 30366
rect 16021 30363 16087 30366
rect 16205 30426 16271 30429
rect 18822 30426 18828 30428
rect 16205 30424 18828 30426
rect 16205 30368 16210 30424
rect 16266 30368 18828 30424
rect 16205 30366 18828 30368
rect 16205 30363 16271 30366
rect 18822 30364 18828 30366
rect 18892 30364 18898 30428
rect 19244 30426 19304 30502
rect 19425 30560 23060 30562
rect 19425 30504 19430 30560
rect 19486 30504 23060 30560
rect 19425 30502 23060 30504
rect 19425 30499 19491 30502
rect 23054 30500 23060 30502
rect 23124 30500 23130 30564
rect 19701 30426 19767 30429
rect 19244 30424 19767 30426
rect 19244 30368 19706 30424
rect 19762 30368 19767 30424
rect 19244 30366 19767 30368
rect 19701 30363 19767 30366
rect 19885 30426 19951 30429
rect 23292 30426 23352 30638
rect 26049 30635 26115 30638
rect 28574 30636 28580 30700
rect 28644 30698 28650 30700
rect 31477 30698 31543 30701
rect 28644 30696 31543 30698
rect 28644 30640 31482 30696
rect 31538 30640 31543 30696
rect 28644 30638 31543 30640
rect 28644 30636 28650 30638
rect 31477 30635 31543 30638
rect 24393 30562 24459 30565
rect 28349 30562 28415 30565
rect 24393 30560 28415 30562
rect 24393 30504 24398 30560
rect 24454 30504 28354 30560
rect 28410 30504 28415 30560
rect 24393 30502 28415 30504
rect 24393 30499 24459 30502
rect 28349 30499 28415 30502
rect 30281 30562 30347 30565
rect 30414 30562 30420 30564
rect 30281 30560 30420 30562
rect 30281 30504 30286 30560
rect 30342 30504 30420 30560
rect 30281 30502 30420 30504
rect 30281 30499 30347 30502
rect 30414 30500 30420 30502
rect 30484 30500 30490 30564
rect 35200 30548 36000 30788
rect 23472 30496 23792 30497
rect 23472 30432 23480 30496
rect 23544 30432 23560 30496
rect 23624 30432 23640 30496
rect 23704 30432 23720 30496
rect 23784 30432 23792 30496
rect 23472 30431 23792 30432
rect 19885 30424 23352 30426
rect 19885 30368 19890 30424
rect 19946 30368 23352 30424
rect 19885 30366 23352 30368
rect 30373 30426 30439 30429
rect 30649 30426 30715 30429
rect 30373 30424 30715 30426
rect 30373 30368 30378 30424
rect 30434 30368 30654 30424
rect 30710 30368 30715 30424
rect 30373 30366 30715 30368
rect 19885 30363 19951 30366
rect 30373 30363 30439 30366
rect 30649 30363 30715 30366
rect 15193 30290 15259 30293
rect 18229 30290 18295 30293
rect 23565 30290 23631 30293
rect 15193 30288 18154 30290
rect 15193 30232 15198 30288
rect 15254 30232 18154 30288
rect 15193 30230 18154 30232
rect 15193 30227 15259 30230
rect 12985 30154 13051 30157
rect 17309 30154 17375 30157
rect 17953 30154 18019 30157
rect 12985 30152 17375 30154
rect 0 29868 800 30108
rect 12985 30096 12990 30152
rect 13046 30096 17314 30152
rect 17370 30096 17375 30152
rect 12985 30094 17375 30096
rect 12985 30091 13051 30094
rect 17309 30091 17375 30094
rect 17496 30152 18019 30154
rect 17496 30096 17958 30152
rect 18014 30096 18019 30152
rect 17496 30094 18019 30096
rect 18094 30154 18154 30230
rect 18229 30288 23631 30290
rect 18229 30232 18234 30288
rect 18290 30232 23570 30288
rect 23626 30232 23631 30288
rect 18229 30230 23631 30232
rect 18229 30227 18295 30230
rect 23565 30227 23631 30230
rect 30005 30290 30071 30293
rect 30649 30290 30715 30293
rect 30005 30288 30715 30290
rect 30005 30232 30010 30288
rect 30066 30232 30654 30288
rect 30710 30232 30715 30288
rect 30005 30230 30715 30232
rect 30005 30227 30071 30230
rect 30649 30227 30715 30230
rect 23105 30154 23171 30157
rect 18094 30152 23171 30154
rect 18094 30096 23110 30152
rect 23166 30096 23171 30152
rect 18094 30094 23171 30096
rect 14825 30018 14891 30021
rect 17033 30018 17099 30021
rect 14825 30016 17099 30018
rect 14825 29960 14830 30016
rect 14886 29960 17038 30016
rect 17094 29960 17099 30016
rect 14825 29958 17099 29960
rect 14825 29955 14891 29958
rect 17033 29955 17099 29958
rect 17217 30018 17283 30021
rect 17496 30018 17556 30094
rect 17953 30091 18019 30094
rect 23105 30091 23171 30094
rect 25773 30154 25839 30157
rect 30741 30154 30807 30157
rect 33501 30154 33567 30157
rect 25773 30152 33567 30154
rect 25773 30096 25778 30152
rect 25834 30096 30746 30152
rect 30802 30096 33506 30152
rect 33562 30096 33567 30152
rect 25773 30094 33567 30096
rect 25773 30091 25839 30094
rect 30741 30091 30807 30094
rect 33501 30091 33567 30094
rect 17217 30016 17556 30018
rect 17217 29960 17222 30016
rect 17278 29960 17556 30016
rect 17217 29958 17556 29960
rect 17217 29955 17283 29958
rect 18454 29956 18460 30020
rect 18524 30018 18530 30020
rect 20805 30018 20871 30021
rect 18524 30016 20871 30018
rect 18524 29960 20810 30016
rect 20866 29960 20871 30016
rect 18524 29958 20871 29960
rect 18524 29956 18530 29958
rect 20805 29955 20871 29958
rect 21725 30018 21791 30021
rect 22461 30018 22527 30021
rect 21725 30016 22527 30018
rect 21725 29960 21730 30016
rect 21786 29960 22466 30016
rect 22522 29960 22527 30016
rect 21725 29958 22527 29960
rect 21725 29955 21791 29958
rect 22461 29955 22527 29958
rect 22686 29956 22692 30020
rect 22756 30018 22762 30020
rect 23933 30018 23999 30021
rect 27797 30018 27863 30021
rect 22756 29958 23858 30018
rect 22756 29956 22762 29958
rect 6576 29952 6896 29953
rect 6576 29888 6584 29952
rect 6648 29888 6664 29952
rect 6728 29888 6744 29952
rect 6808 29888 6824 29952
rect 6888 29888 6896 29952
rect 6576 29887 6896 29888
rect 17840 29952 18160 29953
rect 17840 29888 17848 29952
rect 17912 29888 17928 29952
rect 17992 29888 18008 29952
rect 18072 29888 18088 29952
rect 18152 29888 18160 29952
rect 17840 29887 18160 29888
rect 12709 29882 12775 29885
rect 15653 29882 15719 29885
rect 12709 29880 15719 29882
rect 12709 29824 12714 29880
rect 12770 29824 15658 29880
rect 15714 29824 15719 29880
rect 12709 29822 15719 29824
rect 12709 29819 12775 29822
rect 15653 29819 15719 29822
rect 15929 29882 15995 29885
rect 17401 29882 17467 29885
rect 15929 29880 17467 29882
rect 15929 29824 15934 29880
rect 15990 29824 17406 29880
rect 17462 29824 17467 29880
rect 15929 29822 17467 29824
rect 15929 29819 15995 29822
rect 17401 29819 17467 29822
rect 17534 29820 17540 29884
rect 17604 29882 17610 29884
rect 17677 29882 17743 29885
rect 17604 29880 17743 29882
rect 17604 29824 17682 29880
rect 17738 29824 17743 29880
rect 17604 29822 17743 29824
rect 17604 29820 17610 29822
rect 17677 29819 17743 29822
rect 18229 29884 18295 29885
rect 18229 29880 18276 29884
rect 18340 29882 18346 29884
rect 18505 29882 18571 29885
rect 21909 29882 21975 29885
rect 22645 29882 22711 29885
rect 18229 29824 18234 29880
rect 18229 29820 18276 29824
rect 18340 29822 18386 29882
rect 18505 29880 22711 29882
rect 18505 29824 18510 29880
rect 18566 29824 21914 29880
rect 21970 29824 22650 29880
rect 22706 29824 22711 29880
rect 18505 29822 22711 29824
rect 18340 29820 18346 29822
rect 18229 29819 18295 29820
rect 18505 29819 18571 29822
rect 21909 29819 21975 29822
rect 22645 29819 22711 29822
rect 23238 29820 23244 29884
rect 23308 29882 23314 29884
rect 23473 29882 23539 29885
rect 23308 29880 23539 29882
rect 23308 29824 23478 29880
rect 23534 29824 23539 29880
rect 23308 29822 23539 29824
rect 23798 29882 23858 29958
rect 23933 30016 27863 30018
rect 23933 29960 23938 30016
rect 23994 29960 27802 30016
rect 27858 29960 27863 30016
rect 23933 29958 27863 29960
rect 23933 29955 23999 29958
rect 27797 29955 27863 29958
rect 28441 30018 28507 30021
rect 28901 30018 28967 30021
rect 28441 30016 28967 30018
rect 28441 29960 28446 30016
rect 28502 29960 28906 30016
rect 28962 29960 28967 30016
rect 28441 29958 28967 29960
rect 28441 29955 28507 29958
rect 28901 29955 28967 29958
rect 29637 30018 29703 30021
rect 30833 30018 30899 30021
rect 29637 30016 30899 30018
rect 29637 29960 29642 30016
rect 29698 29960 30838 30016
rect 30894 29960 30899 30016
rect 29637 29958 30899 29960
rect 29637 29955 29703 29958
rect 30833 29955 30899 29958
rect 29104 29952 29424 29953
rect 29104 29888 29112 29952
rect 29176 29888 29192 29952
rect 29256 29888 29272 29952
rect 29336 29888 29352 29952
rect 29416 29888 29424 29952
rect 29104 29887 29424 29888
rect 24117 29882 24183 29885
rect 28533 29884 28599 29885
rect 30833 29884 30899 29885
rect 28533 29882 28580 29884
rect 23798 29880 24183 29882
rect 23798 29824 24122 29880
rect 24178 29824 24183 29880
rect 23798 29822 24183 29824
rect 28488 29880 28580 29882
rect 28488 29824 28538 29880
rect 28488 29822 28580 29824
rect 23308 29820 23314 29822
rect 23473 29819 23539 29822
rect 24117 29819 24183 29822
rect 28533 29820 28580 29822
rect 28644 29820 28650 29884
rect 30782 29882 30788 29884
rect 30742 29822 30788 29882
rect 30852 29880 30899 29884
rect 30894 29824 30899 29880
rect 35200 29868 36000 30108
rect 30782 29820 30788 29822
rect 30852 29820 30899 29824
rect 28533 29819 28599 29820
rect 30790 29819 30899 29820
rect 14181 29744 14247 29749
rect 14181 29688 14186 29744
rect 14242 29688 14247 29744
rect 14181 29683 14247 29688
rect 15285 29746 15351 29749
rect 26325 29746 26391 29749
rect 26877 29746 26943 29749
rect 15285 29744 26943 29746
rect 15285 29688 15290 29744
rect 15346 29688 26330 29744
rect 26386 29688 26882 29744
rect 26938 29688 26943 29744
rect 15285 29686 26943 29688
rect 15285 29683 15351 29686
rect 26325 29683 26391 29686
rect 26877 29683 26943 29686
rect 27061 29746 27127 29749
rect 30790 29746 30850 29819
rect 27061 29744 30850 29746
rect 27061 29688 27066 29744
rect 27122 29688 30850 29744
rect 27061 29686 30850 29688
rect 31661 29746 31727 29749
rect 31845 29746 31911 29749
rect 31661 29744 31911 29746
rect 31661 29688 31666 29744
rect 31722 29688 31850 29744
rect 31906 29688 31911 29744
rect 31661 29686 31911 29688
rect 27061 29683 27127 29686
rect 31661 29683 31727 29686
rect 31845 29683 31911 29686
rect 14184 29474 14244 29683
rect 14457 29610 14523 29613
rect 26877 29610 26943 29613
rect 14457 29608 26943 29610
rect 14457 29552 14462 29608
rect 14518 29552 26882 29608
rect 26938 29552 26943 29608
rect 14457 29550 26943 29552
rect 14457 29547 14523 29550
rect 26877 29547 26943 29550
rect 29361 29610 29427 29613
rect 30557 29610 30623 29613
rect 29361 29608 30623 29610
rect 29361 29552 29366 29608
rect 29422 29552 30562 29608
rect 30618 29552 30623 29608
rect 29361 29550 30623 29552
rect 29361 29547 29427 29550
rect 30557 29547 30623 29550
rect 22369 29474 22435 29477
rect 23238 29474 23244 29476
rect 14184 29472 23244 29474
rect 0 29188 800 29428
rect 14184 29416 22374 29472
rect 22430 29416 23244 29472
rect 14184 29414 23244 29416
rect 22369 29411 22435 29414
rect 23238 29412 23244 29414
rect 23308 29412 23314 29476
rect 23933 29474 23999 29477
rect 28441 29474 28507 29477
rect 23933 29472 28507 29474
rect 23933 29416 23938 29472
rect 23994 29416 28446 29472
rect 28502 29416 28507 29472
rect 23933 29414 28507 29416
rect 23933 29411 23999 29414
rect 28441 29411 28507 29414
rect 29729 29474 29795 29477
rect 30649 29474 30715 29477
rect 29729 29472 30715 29474
rect 29729 29416 29734 29472
rect 29790 29416 30654 29472
rect 30710 29416 30715 29472
rect 29729 29414 30715 29416
rect 29729 29411 29795 29414
rect 30649 29411 30715 29414
rect 12208 29408 12528 29409
rect 12208 29344 12216 29408
rect 12280 29344 12296 29408
rect 12360 29344 12376 29408
rect 12440 29344 12456 29408
rect 12520 29344 12528 29408
rect 12208 29343 12528 29344
rect 23472 29408 23792 29409
rect 23472 29344 23480 29408
rect 23544 29344 23560 29408
rect 23624 29344 23640 29408
rect 23704 29344 23720 29408
rect 23784 29344 23792 29408
rect 23472 29343 23792 29344
rect 13721 29338 13787 29341
rect 14457 29338 14523 29341
rect 13721 29336 14523 29338
rect 13721 29280 13726 29336
rect 13782 29280 14462 29336
rect 14518 29280 14523 29336
rect 13721 29278 14523 29280
rect 13721 29275 13787 29278
rect 14457 29275 14523 29278
rect 14641 29338 14707 29341
rect 16573 29338 16639 29341
rect 14641 29336 16639 29338
rect 14641 29280 14646 29336
rect 14702 29280 16578 29336
rect 16634 29280 16639 29336
rect 14641 29278 16639 29280
rect 14641 29275 14707 29278
rect 16573 29275 16639 29278
rect 17033 29338 17099 29341
rect 23289 29338 23355 29341
rect 17033 29336 23355 29338
rect 17033 29280 17038 29336
rect 17094 29280 23294 29336
rect 23350 29280 23355 29336
rect 17033 29278 23355 29280
rect 17033 29275 17099 29278
rect 23289 29275 23355 29278
rect 29269 29338 29335 29341
rect 35200 29338 36000 29428
rect 29269 29336 36000 29338
rect 29269 29280 29274 29336
rect 29330 29280 36000 29336
rect 29269 29278 36000 29280
rect 29269 29275 29335 29278
rect 13997 29202 14063 29205
rect 14181 29202 14247 29205
rect 13997 29200 14247 29202
rect 13997 29144 14002 29200
rect 14058 29144 14186 29200
rect 14242 29144 14247 29200
rect 13997 29142 14247 29144
rect 13997 29139 14063 29142
rect 14181 29139 14247 29142
rect 14641 29202 14707 29205
rect 16665 29202 16731 29205
rect 14641 29200 16731 29202
rect 14641 29144 14646 29200
rect 14702 29144 16670 29200
rect 16726 29144 16731 29200
rect 14641 29142 16731 29144
rect 14641 29139 14707 29142
rect 16665 29139 16731 29142
rect 16849 29202 16915 29205
rect 21817 29202 21883 29205
rect 16849 29200 21883 29202
rect 16849 29144 16854 29200
rect 16910 29144 21822 29200
rect 21878 29144 21883 29200
rect 16849 29142 21883 29144
rect 16849 29139 16915 29142
rect 21817 29139 21883 29142
rect 22185 29202 22251 29205
rect 22829 29202 22895 29205
rect 22185 29200 22895 29202
rect 22185 29144 22190 29200
rect 22246 29144 22834 29200
rect 22890 29144 22895 29200
rect 22185 29142 22895 29144
rect 22185 29139 22251 29142
rect 22829 29139 22895 29142
rect 28441 29202 28507 29205
rect 31661 29202 31727 29205
rect 28441 29200 31727 29202
rect 28441 29144 28446 29200
rect 28502 29144 31666 29200
rect 31722 29144 31727 29200
rect 35200 29188 36000 29278
rect 28441 29142 31727 29144
rect 28441 29139 28507 29142
rect 31661 29139 31727 29142
rect 13997 29066 14063 29069
rect 20253 29066 20319 29069
rect 20897 29068 20963 29069
rect 20846 29066 20852 29068
rect 13997 29064 20319 29066
rect 13997 29008 14002 29064
rect 14058 29008 20258 29064
rect 20314 29008 20319 29064
rect 13997 29006 20319 29008
rect 20806 29006 20852 29066
rect 20916 29064 20963 29068
rect 31385 29066 31451 29069
rect 20958 29008 20963 29064
rect 13997 29003 14063 29006
rect 20253 29003 20319 29006
rect 20846 29004 20852 29006
rect 20916 29004 20963 29008
rect 20897 29003 20963 29004
rect 21038 29064 31451 29066
rect 21038 29008 31390 29064
rect 31446 29008 31451 29064
rect 21038 29006 31451 29008
rect 15193 28930 15259 28933
rect 15469 28930 15535 28933
rect 15193 28928 15535 28930
rect 15193 28872 15198 28928
rect 15254 28872 15474 28928
rect 15530 28872 15535 28928
rect 15193 28870 15535 28872
rect 15193 28867 15259 28870
rect 15469 28867 15535 28870
rect 15745 28930 15811 28933
rect 17677 28930 17743 28933
rect 15745 28928 17743 28930
rect 15745 28872 15750 28928
rect 15806 28872 17682 28928
rect 17738 28872 17743 28928
rect 15745 28870 17743 28872
rect 15745 28867 15811 28870
rect 17677 28867 17743 28870
rect 18321 28930 18387 28933
rect 21038 28930 21098 29006
rect 31385 29003 31451 29006
rect 21909 28930 21975 28933
rect 18321 28928 21098 28930
rect 18321 28872 18326 28928
rect 18382 28872 21098 28928
rect 18321 28870 21098 28872
rect 21590 28928 21975 28930
rect 21590 28872 21914 28928
rect 21970 28872 21975 28928
rect 21590 28870 21975 28872
rect 18321 28867 18387 28870
rect 6576 28864 6896 28865
rect 6576 28800 6584 28864
rect 6648 28800 6664 28864
rect 6728 28800 6744 28864
rect 6808 28800 6824 28864
rect 6888 28800 6896 28864
rect 6576 28799 6896 28800
rect 17840 28864 18160 28865
rect 17840 28800 17848 28864
rect 17912 28800 17928 28864
rect 17992 28800 18008 28864
rect 18072 28800 18088 28864
rect 18152 28800 18160 28864
rect 17840 28799 18160 28800
rect 11973 28794 12039 28797
rect 13077 28794 13143 28797
rect 11973 28792 13143 28794
rect 0 28508 800 28748
rect 11973 28736 11978 28792
rect 12034 28736 13082 28792
rect 13138 28736 13143 28792
rect 11973 28734 13143 28736
rect 11973 28731 12039 28734
rect 13077 28731 13143 28734
rect 14917 28794 14983 28797
rect 21590 28794 21650 28870
rect 21909 28867 21975 28870
rect 22553 28930 22619 28933
rect 28809 28930 28875 28933
rect 22553 28928 28875 28930
rect 22553 28872 22558 28928
rect 22614 28872 28814 28928
rect 28870 28872 28875 28928
rect 22553 28870 28875 28872
rect 22553 28867 22619 28870
rect 28809 28867 28875 28870
rect 29545 28930 29611 28933
rect 29862 28930 29868 28932
rect 29545 28928 29868 28930
rect 29545 28872 29550 28928
rect 29606 28872 29868 28928
rect 29545 28870 29868 28872
rect 29545 28867 29611 28870
rect 29862 28868 29868 28870
rect 29932 28868 29938 28932
rect 29104 28864 29424 28865
rect 29104 28800 29112 28864
rect 29176 28800 29192 28864
rect 29256 28800 29272 28864
rect 29336 28800 29352 28864
rect 29416 28800 29424 28864
rect 29104 28799 29424 28800
rect 14917 28792 17740 28794
rect 14917 28736 14922 28792
rect 14978 28736 17740 28792
rect 14917 28734 17740 28736
rect 14917 28731 14983 28734
rect 14641 28658 14707 28661
rect 15561 28658 15627 28661
rect 14641 28656 15627 28658
rect 14641 28600 14646 28656
rect 14702 28600 15566 28656
rect 15622 28600 15627 28656
rect 14641 28598 15627 28600
rect 14641 28595 14707 28598
rect 15561 28595 15627 28598
rect 15745 28658 15811 28661
rect 16665 28658 16731 28661
rect 15745 28656 16731 28658
rect 15745 28600 15750 28656
rect 15806 28600 16670 28656
rect 16726 28600 16731 28656
rect 15745 28598 16731 28600
rect 15745 28595 15811 28598
rect 16665 28595 16731 28598
rect 16798 28596 16804 28660
rect 16868 28658 16874 28660
rect 17493 28658 17559 28661
rect 16868 28656 17559 28658
rect 16868 28600 17498 28656
rect 17554 28600 17559 28656
rect 16868 28598 17559 28600
rect 17680 28658 17740 28734
rect 18278 28734 21650 28794
rect 21725 28794 21791 28797
rect 24945 28794 25011 28797
rect 21725 28792 25011 28794
rect 21725 28736 21730 28792
rect 21786 28736 24950 28792
rect 25006 28736 25011 28792
rect 21725 28734 25011 28736
rect 18278 28658 18338 28734
rect 21725 28731 21791 28734
rect 24945 28731 25011 28734
rect 29637 28794 29703 28797
rect 29637 28792 29746 28794
rect 29637 28736 29642 28792
rect 29698 28736 29746 28792
rect 29637 28731 29746 28736
rect 17680 28598 18338 28658
rect 19057 28658 19123 28661
rect 29686 28658 29746 28731
rect 30281 28658 30347 28661
rect 19057 28656 30347 28658
rect 19057 28600 19062 28656
rect 19118 28600 30286 28656
rect 30342 28600 30347 28656
rect 19057 28598 30347 28600
rect 16868 28596 16874 28598
rect 17493 28595 17559 28598
rect 19057 28595 19123 28598
rect 30281 28595 30347 28598
rect 14273 28522 14339 28525
rect 20621 28522 20687 28525
rect 14273 28520 20687 28522
rect 14273 28464 14278 28520
rect 14334 28464 20626 28520
rect 20682 28464 20687 28520
rect 14273 28462 20687 28464
rect 14273 28459 14339 28462
rect 20621 28459 20687 28462
rect 20805 28522 20871 28525
rect 23013 28522 23079 28525
rect 26325 28522 26391 28525
rect 20805 28520 23079 28522
rect 20805 28464 20810 28520
rect 20866 28464 23018 28520
rect 23074 28464 23079 28520
rect 20805 28462 23079 28464
rect 20805 28459 20871 28462
rect 23013 28459 23079 28462
rect 23200 28520 26391 28522
rect 23200 28464 26330 28520
rect 26386 28464 26391 28520
rect 23200 28462 26391 28464
rect 14273 28388 14339 28389
rect 14222 28386 14228 28388
rect 14182 28326 14228 28386
rect 14292 28384 14339 28388
rect 14334 28328 14339 28384
rect 14222 28324 14228 28326
rect 14292 28324 14339 28328
rect 14273 28323 14339 28324
rect 14917 28386 14983 28389
rect 15193 28386 15259 28389
rect 22645 28386 22711 28389
rect 14917 28384 22711 28386
rect 14917 28328 14922 28384
rect 14978 28328 15198 28384
rect 15254 28328 22650 28384
rect 22706 28328 22711 28384
rect 14917 28326 22711 28328
rect 14917 28323 14983 28326
rect 15193 28323 15259 28326
rect 22645 28323 22711 28326
rect 12208 28320 12528 28321
rect 12208 28256 12216 28320
rect 12280 28256 12296 28320
rect 12360 28256 12376 28320
rect 12440 28256 12456 28320
rect 12520 28256 12528 28320
rect 12208 28255 12528 28256
rect 15009 28250 15075 28253
rect 19701 28250 19767 28253
rect 15009 28248 19767 28250
rect 15009 28192 15014 28248
rect 15070 28192 19706 28248
rect 19762 28192 19767 28248
rect 15009 28190 19767 28192
rect 15009 28187 15075 28190
rect 19701 28187 19767 28190
rect 19885 28250 19951 28253
rect 23200 28250 23260 28462
rect 26325 28459 26391 28462
rect 26601 28522 26667 28525
rect 28257 28522 28323 28525
rect 26601 28520 28323 28522
rect 26601 28464 26606 28520
rect 26662 28464 28262 28520
rect 28318 28464 28323 28520
rect 26601 28462 28323 28464
rect 26601 28459 26667 28462
rect 28257 28459 28323 28462
rect 23472 28320 23792 28321
rect 23472 28256 23480 28320
rect 23544 28256 23560 28320
rect 23624 28256 23640 28320
rect 23704 28256 23720 28320
rect 23784 28256 23792 28320
rect 23472 28255 23792 28256
rect 19885 28248 23260 28250
rect 19885 28192 19890 28248
rect 19946 28192 23260 28248
rect 19885 28190 23260 28192
rect 29545 28250 29611 28253
rect 30046 28250 30052 28252
rect 29545 28248 30052 28250
rect 29545 28192 29550 28248
rect 29606 28192 30052 28248
rect 29545 28190 30052 28192
rect 19885 28187 19951 28190
rect 29545 28187 29611 28190
rect 30046 28188 30052 28190
rect 30116 28188 30122 28252
rect 15285 28114 15351 28117
rect 20529 28114 20595 28117
rect 15285 28112 20595 28114
rect 0 27828 800 28068
rect 15285 28056 15290 28112
rect 15346 28056 20534 28112
rect 20590 28056 20595 28112
rect 15285 28054 20595 28056
rect 15285 28051 15351 28054
rect 20529 28051 20595 28054
rect 20713 28114 20779 28117
rect 32305 28114 32371 28117
rect 20713 28112 32371 28114
rect 20713 28056 20718 28112
rect 20774 28056 32310 28112
rect 32366 28056 32371 28112
rect 20713 28054 32371 28056
rect 20713 28051 20779 28054
rect 32305 28051 32371 28054
rect 13445 27978 13511 27981
rect 15326 27978 15332 27980
rect 13445 27976 15332 27978
rect 13445 27920 13450 27976
rect 13506 27920 15332 27976
rect 13445 27918 15332 27920
rect 13445 27915 13511 27918
rect 15326 27916 15332 27918
rect 15396 27916 15402 27980
rect 15469 27978 15535 27981
rect 21909 27978 21975 27981
rect 23933 27978 23999 27981
rect 15469 27976 21834 27978
rect 15469 27920 15474 27976
rect 15530 27920 21834 27976
rect 15469 27918 21834 27920
rect 15469 27915 15535 27918
rect 15193 27842 15259 27845
rect 17585 27842 17651 27845
rect 15193 27840 17651 27842
rect 15193 27784 15198 27840
rect 15254 27784 17590 27840
rect 17646 27784 17651 27840
rect 15193 27782 17651 27784
rect 15193 27779 15259 27782
rect 17585 27779 17651 27782
rect 18321 27842 18387 27845
rect 21265 27842 21331 27845
rect 18321 27840 21331 27842
rect 18321 27784 18326 27840
rect 18382 27784 21270 27840
rect 21326 27784 21331 27840
rect 18321 27782 21331 27784
rect 21774 27842 21834 27918
rect 21909 27976 23999 27978
rect 21909 27920 21914 27976
rect 21970 27920 23938 27976
rect 23994 27920 23999 27976
rect 21909 27918 23999 27920
rect 21909 27915 21975 27918
rect 23933 27915 23999 27918
rect 27521 27978 27587 27981
rect 27797 27978 27863 27981
rect 27521 27976 27863 27978
rect 27521 27920 27526 27976
rect 27582 27920 27802 27976
rect 27858 27920 27863 27976
rect 27521 27918 27863 27920
rect 27521 27915 27587 27918
rect 27797 27915 27863 27918
rect 34145 27978 34211 27981
rect 35200 27978 36000 28068
rect 34145 27976 36000 27978
rect 34145 27920 34150 27976
rect 34206 27920 36000 27976
rect 34145 27918 36000 27920
rect 34145 27915 34211 27918
rect 22829 27842 22895 27845
rect 21774 27840 22895 27842
rect 21774 27784 22834 27840
rect 22890 27784 22895 27840
rect 21774 27782 22895 27784
rect 18321 27779 18387 27782
rect 21265 27779 21331 27782
rect 22829 27779 22895 27782
rect 23013 27842 23079 27845
rect 23749 27842 23815 27845
rect 23013 27840 23815 27842
rect 23013 27784 23018 27840
rect 23074 27784 23754 27840
rect 23810 27784 23815 27840
rect 23013 27782 23815 27784
rect 23013 27779 23079 27782
rect 23749 27779 23815 27782
rect 24301 27842 24367 27845
rect 26601 27842 26667 27845
rect 24301 27840 26667 27842
rect 24301 27784 24306 27840
rect 24362 27784 26606 27840
rect 26662 27784 26667 27840
rect 35200 27828 36000 27918
rect 24301 27782 26667 27784
rect 24301 27779 24367 27782
rect 26601 27779 26667 27782
rect 6576 27776 6896 27777
rect 6576 27712 6584 27776
rect 6648 27712 6664 27776
rect 6728 27712 6744 27776
rect 6808 27712 6824 27776
rect 6888 27712 6896 27776
rect 6576 27711 6896 27712
rect 17840 27776 18160 27777
rect 17840 27712 17848 27776
rect 17912 27712 17928 27776
rect 17992 27712 18008 27776
rect 18072 27712 18088 27776
rect 18152 27712 18160 27776
rect 17840 27711 18160 27712
rect 29104 27776 29424 27777
rect 29104 27712 29112 27776
rect 29176 27712 29192 27776
rect 29256 27712 29272 27776
rect 29336 27712 29352 27776
rect 29416 27712 29424 27776
rect 29104 27711 29424 27712
rect 13353 27706 13419 27709
rect 17677 27706 17743 27709
rect 13353 27704 17743 27706
rect 13353 27648 13358 27704
rect 13414 27648 17682 27704
rect 17738 27648 17743 27704
rect 13353 27646 17743 27648
rect 13353 27643 13419 27646
rect 17677 27643 17743 27646
rect 18229 27706 18295 27709
rect 25313 27706 25379 27709
rect 25957 27706 26023 27709
rect 18229 27704 26023 27706
rect 18229 27648 18234 27704
rect 18290 27648 25318 27704
rect 25374 27648 25962 27704
rect 26018 27648 26023 27704
rect 18229 27646 26023 27648
rect 18229 27643 18295 27646
rect 25313 27643 25379 27646
rect 25957 27643 26023 27646
rect 15837 27570 15903 27573
rect 16062 27570 16068 27572
rect 15837 27568 16068 27570
rect 15837 27512 15842 27568
rect 15898 27512 16068 27568
rect 15837 27510 16068 27512
rect 15837 27507 15903 27510
rect 16062 27508 16068 27510
rect 16132 27508 16138 27572
rect 16205 27570 16271 27573
rect 18321 27570 18387 27573
rect 16205 27568 18387 27570
rect 16205 27512 16210 27568
rect 16266 27512 18326 27568
rect 18382 27512 18387 27568
rect 16205 27510 18387 27512
rect 16205 27507 16271 27510
rect 18321 27507 18387 27510
rect 18505 27570 18571 27573
rect 19885 27570 19951 27573
rect 18505 27568 19951 27570
rect 18505 27512 18510 27568
rect 18566 27512 19890 27568
rect 19946 27512 19951 27568
rect 18505 27510 19951 27512
rect 18505 27507 18571 27510
rect 19885 27507 19951 27510
rect 20161 27570 20227 27573
rect 22001 27570 22067 27573
rect 20161 27568 22067 27570
rect 20161 27512 20166 27568
rect 20222 27512 22006 27568
rect 22062 27512 22067 27568
rect 20161 27510 22067 27512
rect 20161 27507 20227 27510
rect 22001 27507 22067 27510
rect 22185 27570 22251 27573
rect 27337 27570 27403 27573
rect 22185 27568 27403 27570
rect 22185 27512 22190 27568
rect 22246 27512 27342 27568
rect 27398 27512 27403 27568
rect 22185 27510 27403 27512
rect 22185 27507 22251 27510
rect 27337 27507 27403 27510
rect 15285 27434 15351 27437
rect 19241 27434 19307 27437
rect 15285 27432 19307 27434
rect 0 27148 800 27388
rect 15285 27376 15290 27432
rect 15346 27376 19246 27432
rect 19302 27376 19307 27432
rect 15285 27374 19307 27376
rect 15285 27371 15351 27374
rect 19241 27371 19307 27374
rect 21541 27434 21607 27437
rect 24301 27434 24367 27437
rect 21541 27432 24367 27434
rect 21541 27376 21546 27432
rect 21602 27376 24306 27432
rect 24362 27376 24367 27432
rect 21541 27374 24367 27376
rect 21541 27371 21607 27374
rect 24301 27371 24367 27374
rect 26969 27434 27035 27437
rect 28441 27434 28507 27437
rect 26969 27432 28507 27434
rect 26969 27376 26974 27432
rect 27030 27376 28446 27432
rect 28502 27376 28507 27432
rect 26969 27374 28507 27376
rect 26969 27371 27035 27374
rect 28441 27371 28507 27374
rect 15101 27298 15167 27301
rect 15101 27296 16498 27298
rect 15101 27240 15106 27296
rect 15162 27240 16498 27296
rect 15101 27238 16498 27240
rect 15101 27235 15167 27238
rect 12208 27232 12528 27233
rect 12208 27168 12216 27232
rect 12280 27168 12296 27232
rect 12360 27168 12376 27232
rect 12440 27168 12456 27232
rect 12520 27168 12528 27232
rect 12208 27167 12528 27168
rect 13537 27162 13603 27165
rect 15561 27162 15627 27165
rect 13537 27160 15627 27162
rect 13537 27104 13542 27160
rect 13598 27104 15566 27160
rect 15622 27104 15627 27160
rect 13537 27102 15627 27104
rect 13537 27099 13603 27102
rect 15561 27099 15627 27102
rect 15929 27162 15995 27165
rect 16297 27162 16363 27165
rect 15929 27160 16363 27162
rect 15929 27104 15934 27160
rect 15990 27104 16302 27160
rect 16358 27104 16363 27160
rect 15929 27102 16363 27104
rect 16438 27162 16498 27238
rect 16614 27236 16620 27300
rect 16684 27298 16690 27300
rect 16849 27298 16915 27301
rect 16684 27296 16915 27298
rect 16684 27240 16854 27296
rect 16910 27240 16915 27296
rect 16684 27238 16915 27240
rect 16684 27236 16690 27238
rect 16849 27235 16915 27238
rect 17217 27298 17283 27301
rect 20989 27298 21055 27301
rect 17217 27296 21055 27298
rect 17217 27240 17222 27296
rect 17278 27240 20994 27296
rect 21050 27240 21055 27296
rect 17217 27238 21055 27240
rect 17217 27235 17283 27238
rect 20989 27235 21055 27238
rect 28441 27298 28507 27301
rect 30414 27298 30420 27300
rect 28441 27296 30420 27298
rect 28441 27240 28446 27296
rect 28502 27240 30420 27296
rect 28441 27238 30420 27240
rect 28441 27235 28507 27238
rect 30414 27236 30420 27238
rect 30484 27298 30490 27300
rect 31017 27298 31083 27301
rect 30484 27296 31083 27298
rect 30484 27240 31022 27296
rect 31078 27240 31083 27296
rect 30484 27238 31083 27240
rect 30484 27236 30490 27238
rect 31017 27235 31083 27238
rect 23472 27232 23792 27233
rect 23472 27168 23480 27232
rect 23544 27168 23560 27232
rect 23624 27168 23640 27232
rect 23704 27168 23720 27232
rect 23784 27168 23792 27232
rect 23472 27167 23792 27168
rect 30833 27164 30899 27165
rect 16438 27102 22984 27162
rect 15929 27099 15995 27102
rect 16297 27099 16363 27102
rect 22924 27029 22984 27102
rect 30782 27100 30788 27164
rect 30852 27162 30899 27164
rect 30852 27160 30944 27162
rect 30894 27104 30944 27160
rect 35200 27148 36000 27388
rect 30852 27102 30944 27104
rect 30852 27100 30899 27102
rect 30833 27099 30899 27100
rect 13537 27026 13603 27029
rect 20713 27026 20779 27029
rect 13537 27024 20779 27026
rect 13537 26968 13542 27024
rect 13598 26968 20718 27024
rect 20774 26968 20779 27024
rect 13537 26966 20779 26968
rect 13537 26963 13603 26966
rect 20713 26963 20779 26966
rect 22921 27026 22987 27029
rect 27245 27026 27311 27029
rect 22921 27024 27311 27026
rect 22921 26968 22926 27024
rect 22982 26968 27250 27024
rect 27306 26968 27311 27024
rect 22921 26966 27311 26968
rect 22921 26963 22987 26966
rect 27245 26963 27311 26966
rect 16297 26890 16363 26893
rect 23933 26890 23999 26893
rect 29545 26892 29611 26893
rect 29494 26890 29500 26892
rect 16297 26888 23999 26890
rect 16297 26832 16302 26888
rect 16358 26832 23938 26888
rect 23994 26832 23999 26888
rect 16297 26830 23999 26832
rect 29418 26830 29500 26890
rect 29564 26890 29611 26892
rect 33409 26890 33475 26893
rect 29564 26888 33475 26890
rect 29606 26832 33414 26888
rect 33470 26832 33475 26888
rect 16297 26827 16363 26830
rect 23933 26827 23999 26830
rect 29494 26828 29500 26830
rect 29564 26830 33475 26832
rect 29564 26828 29611 26830
rect 29545 26827 29611 26828
rect 33409 26827 33475 26830
rect 14733 26754 14799 26757
rect 16113 26754 16179 26757
rect 14733 26752 16179 26754
rect 14733 26696 14738 26752
rect 14794 26696 16118 26752
rect 16174 26696 16179 26752
rect 14733 26694 16179 26696
rect 14733 26691 14799 26694
rect 16113 26691 16179 26694
rect 16665 26754 16731 26757
rect 17401 26754 17467 26757
rect 17585 26754 17651 26757
rect 16665 26752 17467 26754
rect 16665 26696 16670 26752
rect 16726 26696 17406 26752
rect 17462 26696 17467 26752
rect 16665 26694 17467 26696
rect 16665 26691 16731 26694
rect 17401 26691 17467 26694
rect 17542 26752 17651 26754
rect 17542 26696 17590 26752
rect 17646 26696 17651 26752
rect 17542 26691 17651 26696
rect 18965 26754 19031 26757
rect 28625 26754 28691 26757
rect 18965 26752 28691 26754
rect 18965 26696 18970 26752
rect 19026 26696 28630 26752
rect 28686 26696 28691 26752
rect 18965 26694 28691 26696
rect 18965 26691 19031 26694
rect 28625 26691 28691 26694
rect 6576 26688 6896 26689
rect 6576 26624 6584 26688
rect 6648 26624 6664 26688
rect 6728 26624 6744 26688
rect 6808 26624 6824 26688
rect 6888 26624 6896 26688
rect 6576 26623 6896 26624
rect 14181 26618 14247 26621
rect 17542 26618 17602 26691
rect 17840 26688 18160 26689
rect 17840 26624 17848 26688
rect 17912 26624 17928 26688
rect 17992 26624 18008 26688
rect 18072 26624 18088 26688
rect 18152 26624 18160 26688
rect 17840 26623 18160 26624
rect 29104 26688 29424 26689
rect 29104 26624 29112 26688
rect 29176 26624 29192 26688
rect 29256 26624 29272 26688
rect 29336 26624 29352 26688
rect 29416 26624 29424 26688
rect 29104 26623 29424 26624
rect 14181 26616 17602 26618
rect 14181 26560 14186 26616
rect 14242 26560 17602 26616
rect 14181 26558 17602 26560
rect 18781 26618 18847 26621
rect 25497 26618 25563 26621
rect 18781 26616 25563 26618
rect 18781 26560 18786 26616
rect 18842 26560 25502 26616
rect 25558 26560 25563 26616
rect 18781 26558 25563 26560
rect 14181 26555 14247 26558
rect 18781 26555 18847 26558
rect 25497 26555 25563 26558
rect 15009 26482 15075 26485
rect 18689 26482 18755 26485
rect 23473 26482 23539 26485
rect 15009 26480 18755 26482
rect 15009 26424 15014 26480
rect 15070 26424 18694 26480
rect 18750 26424 18755 26480
rect 15009 26422 18755 26424
rect 15009 26419 15075 26422
rect 18689 26419 18755 26422
rect 21038 26480 23539 26482
rect 21038 26424 23478 26480
rect 23534 26424 23539 26480
rect 35200 26468 36000 26708
rect 21038 26422 23539 26424
rect 15193 26346 15259 26349
rect 21038 26346 21098 26422
rect 23473 26419 23539 26422
rect 15193 26344 21098 26346
rect 15193 26288 15198 26344
rect 15254 26288 21098 26344
rect 15193 26286 21098 26288
rect 15193 26283 15259 26286
rect 15469 26210 15535 26213
rect 21633 26210 21699 26213
rect 15469 26208 21699 26210
rect 15469 26152 15474 26208
rect 15530 26152 21638 26208
rect 21694 26152 21699 26208
rect 15469 26150 21699 26152
rect 15469 26147 15535 26150
rect 21633 26147 21699 26150
rect 12208 26144 12528 26145
rect 12208 26080 12216 26144
rect 12280 26080 12296 26144
rect 12360 26080 12376 26144
rect 12440 26080 12456 26144
rect 12520 26080 12528 26144
rect 12208 26079 12528 26080
rect 23472 26144 23792 26145
rect 23472 26080 23480 26144
rect 23544 26080 23560 26144
rect 23624 26080 23640 26144
rect 23704 26080 23720 26144
rect 23784 26080 23792 26144
rect 23472 26079 23792 26080
rect 15285 26074 15351 26077
rect 19609 26074 19675 26077
rect 15285 26072 19675 26074
rect 0 25788 800 26028
rect 15285 26016 15290 26072
rect 15346 26016 19614 26072
rect 19670 26016 19675 26072
rect 15285 26014 19675 26016
rect 15285 26011 15351 26014
rect 19609 26011 19675 26014
rect 14457 25938 14523 25941
rect 20437 25938 20503 25941
rect 14457 25936 20503 25938
rect 14457 25880 14462 25936
rect 14518 25880 20442 25936
rect 20498 25880 20503 25936
rect 14457 25878 20503 25880
rect 14457 25875 14523 25878
rect 20437 25875 20503 25878
rect 30649 25938 30715 25941
rect 31702 25938 31708 25940
rect 30649 25936 31708 25938
rect 30649 25880 30654 25936
rect 30710 25880 31708 25936
rect 30649 25878 31708 25880
rect 30649 25875 30715 25878
rect 31702 25876 31708 25878
rect 31772 25876 31778 25940
rect 34145 25938 34211 25941
rect 35200 25938 36000 26028
rect 34145 25936 36000 25938
rect 34145 25880 34150 25936
rect 34206 25880 36000 25936
rect 34145 25878 36000 25880
rect 34145 25875 34211 25878
rect 13077 25802 13143 25805
rect 18873 25802 18939 25805
rect 13077 25800 18939 25802
rect 13077 25744 13082 25800
rect 13138 25744 18878 25800
rect 18934 25744 18939 25800
rect 35200 25788 36000 25878
rect 13077 25742 18939 25744
rect 13077 25739 13143 25742
rect 18873 25739 18939 25742
rect 15929 25666 15995 25669
rect 17677 25666 17743 25669
rect 15929 25664 17743 25666
rect 15929 25608 15934 25664
rect 15990 25608 17682 25664
rect 17738 25608 17743 25664
rect 15929 25606 17743 25608
rect 15929 25603 15995 25606
rect 17677 25603 17743 25606
rect 18229 25666 18295 25669
rect 22553 25666 22619 25669
rect 18229 25664 22619 25666
rect 18229 25608 18234 25664
rect 18290 25608 22558 25664
rect 22614 25608 22619 25664
rect 18229 25606 22619 25608
rect 18229 25603 18295 25606
rect 22553 25603 22619 25606
rect 6576 25600 6896 25601
rect 6576 25536 6584 25600
rect 6648 25536 6664 25600
rect 6728 25536 6744 25600
rect 6808 25536 6824 25600
rect 6888 25536 6896 25600
rect 6576 25535 6896 25536
rect 17840 25600 18160 25601
rect 17840 25536 17848 25600
rect 17912 25536 17928 25600
rect 17992 25536 18008 25600
rect 18072 25536 18088 25600
rect 18152 25536 18160 25600
rect 17840 25535 18160 25536
rect 29104 25600 29424 25601
rect 29104 25536 29112 25600
rect 29176 25536 29192 25600
rect 29256 25536 29272 25600
rect 29336 25536 29352 25600
rect 29416 25536 29424 25600
rect 29104 25535 29424 25536
rect 14825 25530 14891 25533
rect 17677 25530 17743 25533
rect 14825 25528 17743 25530
rect 14825 25472 14830 25528
rect 14886 25472 17682 25528
rect 17738 25472 17743 25528
rect 14825 25470 17743 25472
rect 14825 25467 14891 25470
rect 17677 25467 17743 25470
rect 20345 25530 20411 25533
rect 24209 25530 24275 25533
rect 25497 25530 25563 25533
rect 20345 25528 25563 25530
rect 20345 25472 20350 25528
rect 20406 25472 24214 25528
rect 24270 25472 25502 25528
rect 25558 25472 25563 25528
rect 20345 25470 25563 25472
rect 20345 25467 20411 25470
rect 24209 25467 24275 25470
rect 25497 25467 25563 25470
rect 16665 25394 16731 25397
rect 18781 25394 18847 25397
rect 16665 25392 18847 25394
rect 0 25258 800 25348
rect 16665 25336 16670 25392
rect 16726 25336 18786 25392
rect 18842 25336 18847 25392
rect 16665 25334 18847 25336
rect 16665 25331 16731 25334
rect 18781 25331 18847 25334
rect 21725 25394 21791 25397
rect 25313 25394 25379 25397
rect 21725 25392 25379 25394
rect 21725 25336 21730 25392
rect 21786 25336 25318 25392
rect 25374 25336 25379 25392
rect 21725 25334 25379 25336
rect 21725 25331 21791 25334
rect 25313 25331 25379 25334
rect 31477 25394 31543 25397
rect 32949 25394 33015 25397
rect 31477 25392 33015 25394
rect 31477 25336 31482 25392
rect 31538 25336 32954 25392
rect 33010 25336 33015 25392
rect 31477 25334 33015 25336
rect 31477 25331 31543 25334
rect 32949 25331 33015 25334
rect 1853 25258 1919 25261
rect 0 25256 1919 25258
rect 0 25200 1858 25256
rect 1914 25200 1919 25256
rect 0 25198 1919 25200
rect 0 25108 800 25198
rect 1853 25195 1919 25198
rect 14733 25258 14799 25261
rect 28073 25258 28139 25261
rect 14733 25256 28139 25258
rect 14733 25200 14738 25256
rect 14794 25200 28078 25256
rect 28134 25200 28139 25256
rect 14733 25198 28139 25200
rect 14733 25195 14799 25198
rect 28073 25195 28139 25198
rect 34145 25258 34211 25261
rect 35200 25258 36000 25348
rect 34145 25256 36000 25258
rect 34145 25200 34150 25256
rect 34206 25200 36000 25256
rect 34145 25198 36000 25200
rect 34145 25195 34211 25198
rect 15745 25122 15811 25125
rect 18505 25122 18571 25125
rect 15745 25120 18571 25122
rect 15745 25064 15750 25120
rect 15806 25064 18510 25120
rect 18566 25064 18571 25120
rect 35200 25108 36000 25198
rect 15745 25062 18571 25064
rect 15745 25059 15811 25062
rect 18505 25059 18571 25062
rect 12208 25056 12528 25057
rect 12208 24992 12216 25056
rect 12280 24992 12296 25056
rect 12360 24992 12376 25056
rect 12440 24992 12456 25056
rect 12520 24992 12528 25056
rect 12208 24991 12528 24992
rect 23472 25056 23792 25057
rect 23472 24992 23480 25056
rect 23544 24992 23560 25056
rect 23624 24992 23640 25056
rect 23704 24992 23720 25056
rect 23784 24992 23792 25056
rect 23472 24991 23792 24992
rect 14917 24986 14983 24989
rect 21725 24986 21791 24989
rect 14917 24984 21791 24986
rect 14917 24928 14922 24984
rect 14978 24928 21730 24984
rect 21786 24928 21791 24984
rect 14917 24926 21791 24928
rect 14917 24923 14983 24926
rect 21725 24923 21791 24926
rect 3417 24850 3483 24853
rect 27654 24850 27660 24852
rect 3417 24848 27660 24850
rect 3417 24792 3422 24848
rect 3478 24792 27660 24848
rect 3417 24790 27660 24792
rect 3417 24787 3483 24790
rect 27654 24788 27660 24790
rect 27724 24788 27730 24852
rect 12801 24714 12867 24717
rect 18965 24714 19031 24717
rect 12801 24712 19031 24714
rect 0 24428 800 24668
rect 12801 24656 12806 24712
rect 12862 24656 18970 24712
rect 19026 24656 19031 24712
rect 12801 24654 19031 24656
rect 12801 24651 12867 24654
rect 18965 24651 19031 24654
rect 20713 24714 20779 24717
rect 23657 24714 23723 24717
rect 20713 24712 23723 24714
rect 20713 24656 20718 24712
rect 20774 24656 23662 24712
rect 23718 24656 23723 24712
rect 20713 24654 23723 24656
rect 20713 24651 20779 24654
rect 23657 24651 23723 24654
rect 29453 24714 29519 24717
rect 31661 24714 31727 24717
rect 29453 24712 31727 24714
rect 29453 24656 29458 24712
rect 29514 24656 31666 24712
rect 31722 24656 31727 24712
rect 29453 24654 31727 24656
rect 29453 24651 29519 24654
rect 31661 24651 31727 24654
rect 21817 24578 21883 24581
rect 23933 24578 23999 24581
rect 29729 24580 29795 24581
rect 21817 24576 23999 24578
rect 21817 24520 21822 24576
rect 21878 24520 23938 24576
rect 23994 24520 23999 24576
rect 21817 24518 23999 24520
rect 21817 24515 21883 24518
rect 23933 24515 23999 24518
rect 29678 24516 29684 24580
rect 29748 24578 29795 24580
rect 34145 24578 34211 24581
rect 35200 24578 36000 24668
rect 29748 24576 29840 24578
rect 29790 24520 29840 24576
rect 29748 24518 29840 24520
rect 34145 24576 36000 24578
rect 34145 24520 34150 24576
rect 34206 24520 36000 24576
rect 34145 24518 36000 24520
rect 29748 24516 29795 24518
rect 29729 24515 29795 24516
rect 34145 24515 34211 24518
rect 6576 24512 6896 24513
rect 6576 24448 6584 24512
rect 6648 24448 6664 24512
rect 6728 24448 6744 24512
rect 6808 24448 6824 24512
rect 6888 24448 6896 24512
rect 6576 24447 6896 24448
rect 17840 24512 18160 24513
rect 17840 24448 17848 24512
rect 17912 24448 17928 24512
rect 17992 24448 18008 24512
rect 18072 24448 18088 24512
rect 18152 24448 18160 24512
rect 17840 24447 18160 24448
rect 29104 24512 29424 24513
rect 29104 24448 29112 24512
rect 29176 24448 29192 24512
rect 29256 24448 29272 24512
rect 29336 24448 29352 24512
rect 29416 24448 29424 24512
rect 29104 24447 29424 24448
rect 19333 24442 19399 24445
rect 24669 24442 24735 24445
rect 19333 24440 24735 24442
rect 19333 24384 19338 24440
rect 19394 24384 24674 24440
rect 24730 24384 24735 24440
rect 35200 24428 36000 24518
rect 19333 24382 24735 24384
rect 19333 24379 19399 24382
rect 24669 24379 24735 24382
rect 14917 24306 14983 24309
rect 18413 24306 18479 24309
rect 14917 24304 18479 24306
rect 14917 24248 14922 24304
rect 14978 24248 18418 24304
rect 18474 24248 18479 24304
rect 14917 24246 18479 24248
rect 14917 24243 14983 24246
rect 18413 24243 18479 24246
rect 20069 24306 20135 24309
rect 27705 24306 27771 24309
rect 20069 24304 27771 24306
rect 20069 24248 20074 24304
rect 20130 24248 27710 24304
rect 27766 24248 27771 24304
rect 20069 24246 27771 24248
rect 20069 24243 20135 24246
rect 27705 24243 27771 24246
rect 14641 24170 14707 24173
rect 19241 24170 19307 24173
rect 14641 24168 19307 24170
rect 14641 24112 14646 24168
rect 14702 24112 19246 24168
rect 19302 24112 19307 24168
rect 14641 24110 19307 24112
rect 14641 24107 14707 24110
rect 19241 24107 19307 24110
rect 15837 24034 15903 24037
rect 18413 24034 18479 24037
rect 15837 24032 18479 24034
rect 0 23748 800 23988
rect 15837 23976 15842 24032
rect 15898 23976 18418 24032
rect 18474 23976 18479 24032
rect 15837 23974 18479 23976
rect 15837 23971 15903 23974
rect 18413 23971 18479 23974
rect 28349 24034 28415 24037
rect 28717 24034 28783 24037
rect 28349 24032 28783 24034
rect 28349 23976 28354 24032
rect 28410 23976 28722 24032
rect 28778 23976 28783 24032
rect 28349 23974 28783 23976
rect 28349 23971 28415 23974
rect 28717 23971 28783 23974
rect 12208 23968 12528 23969
rect 12208 23904 12216 23968
rect 12280 23904 12296 23968
rect 12360 23904 12376 23968
rect 12440 23904 12456 23968
rect 12520 23904 12528 23968
rect 12208 23903 12528 23904
rect 23472 23968 23792 23969
rect 23472 23904 23480 23968
rect 23544 23904 23560 23968
rect 23624 23904 23640 23968
rect 23704 23904 23720 23968
rect 23784 23904 23792 23968
rect 23472 23903 23792 23904
rect 15101 23898 15167 23901
rect 18505 23898 18571 23901
rect 15101 23896 18571 23898
rect 15101 23840 15106 23896
rect 15162 23840 18510 23896
rect 18566 23840 18571 23896
rect 15101 23838 18571 23840
rect 15101 23835 15167 23838
rect 18505 23835 18571 23838
rect 32397 23898 32463 23901
rect 32622 23898 32628 23900
rect 32397 23896 32628 23898
rect 32397 23840 32402 23896
rect 32458 23840 32628 23896
rect 32397 23838 32628 23840
rect 32397 23835 32463 23838
rect 32622 23836 32628 23838
rect 32692 23836 32698 23900
rect 34145 23898 34211 23901
rect 35200 23898 36000 23988
rect 34145 23896 36000 23898
rect 34145 23840 34150 23896
rect 34206 23840 36000 23896
rect 34145 23838 36000 23840
rect 34145 23835 34211 23838
rect 14733 23762 14799 23765
rect 18689 23762 18755 23765
rect 14733 23760 18755 23762
rect 14733 23704 14738 23760
rect 14794 23704 18694 23760
rect 18750 23704 18755 23760
rect 14733 23702 18755 23704
rect 14733 23699 14799 23702
rect 18689 23699 18755 23702
rect 26785 23762 26851 23765
rect 31293 23762 31359 23765
rect 26785 23760 31359 23762
rect 26785 23704 26790 23760
rect 26846 23704 31298 23760
rect 31354 23704 31359 23760
rect 35200 23748 36000 23838
rect 26785 23702 31359 23704
rect 26785 23699 26851 23702
rect 31293 23699 31359 23702
rect 21449 23626 21515 23629
rect 28717 23626 28783 23629
rect 21449 23624 28783 23626
rect 21449 23568 21454 23624
rect 21510 23568 28722 23624
rect 28778 23568 28783 23624
rect 21449 23566 28783 23568
rect 21449 23563 21515 23566
rect 28717 23563 28783 23566
rect 28993 23626 29059 23629
rect 33501 23626 33567 23629
rect 28993 23624 33567 23626
rect 28993 23568 28998 23624
rect 29054 23568 33506 23624
rect 33562 23568 33567 23624
rect 28993 23566 33567 23568
rect 28993 23563 29059 23566
rect 33501 23563 33567 23566
rect 6576 23424 6896 23425
rect 6576 23360 6584 23424
rect 6648 23360 6664 23424
rect 6728 23360 6744 23424
rect 6808 23360 6824 23424
rect 6888 23360 6896 23424
rect 6576 23359 6896 23360
rect 17840 23424 18160 23425
rect 17840 23360 17848 23424
rect 17912 23360 17928 23424
rect 17992 23360 18008 23424
rect 18072 23360 18088 23424
rect 18152 23360 18160 23424
rect 17840 23359 18160 23360
rect 29104 23424 29424 23425
rect 29104 23360 29112 23424
rect 29176 23360 29192 23424
rect 29256 23360 29272 23424
rect 29336 23360 29352 23424
rect 29416 23360 29424 23424
rect 29104 23359 29424 23360
rect 20437 23354 20503 23357
rect 25221 23354 25287 23357
rect 20437 23352 25287 23354
rect 0 23068 800 23308
rect 20437 23296 20442 23352
rect 20498 23296 25226 23352
rect 25282 23296 25287 23352
rect 20437 23294 25287 23296
rect 20437 23291 20503 23294
rect 25221 23291 25287 23294
rect 20345 23218 20411 23221
rect 22921 23218 22987 23221
rect 20345 23216 22987 23218
rect 20345 23160 20350 23216
rect 20406 23160 22926 23216
rect 22982 23160 22987 23216
rect 20345 23158 22987 23160
rect 20345 23155 20411 23158
rect 22921 23155 22987 23158
rect 28441 23218 28507 23221
rect 28901 23218 28967 23221
rect 28441 23216 28967 23218
rect 28441 23160 28446 23216
rect 28502 23160 28906 23216
rect 28962 23160 28967 23216
rect 28441 23158 28967 23160
rect 28441 23155 28507 23158
rect 28901 23155 28967 23158
rect 34145 23218 34211 23221
rect 35200 23218 36000 23308
rect 34145 23216 36000 23218
rect 34145 23160 34150 23216
rect 34206 23160 36000 23216
rect 34145 23158 36000 23160
rect 34145 23155 34211 23158
rect 21541 23082 21607 23085
rect 24209 23082 24275 23085
rect 31293 23082 31359 23085
rect 21541 23080 31359 23082
rect 21541 23024 21546 23080
rect 21602 23024 24214 23080
rect 24270 23024 31298 23080
rect 31354 23024 31359 23080
rect 35200 23068 36000 23158
rect 21541 23022 31359 23024
rect 21541 23019 21607 23022
rect 24209 23019 24275 23022
rect 31293 23019 31359 23022
rect 21817 22946 21883 22949
rect 23197 22946 23263 22949
rect 21817 22944 23263 22946
rect 21817 22888 21822 22944
rect 21878 22888 23202 22944
rect 23258 22888 23263 22944
rect 21817 22886 23263 22888
rect 21817 22883 21883 22886
rect 23197 22883 23263 22886
rect 32397 22946 32463 22949
rect 32806 22946 32812 22948
rect 32397 22944 32812 22946
rect 32397 22888 32402 22944
rect 32458 22888 32812 22944
rect 32397 22886 32812 22888
rect 32397 22883 32463 22886
rect 32806 22884 32812 22886
rect 32876 22884 32882 22948
rect 12208 22880 12528 22881
rect 12208 22816 12216 22880
rect 12280 22816 12296 22880
rect 12360 22816 12376 22880
rect 12440 22816 12456 22880
rect 12520 22816 12528 22880
rect 12208 22815 12528 22816
rect 23472 22880 23792 22881
rect 23472 22816 23480 22880
rect 23544 22816 23560 22880
rect 23624 22816 23640 22880
rect 23704 22816 23720 22880
rect 23784 22816 23792 22880
rect 23472 22815 23792 22816
rect 13169 22810 13235 22813
rect 22093 22810 22159 22813
rect 13169 22808 22159 22810
rect 13169 22752 13174 22808
rect 13230 22752 22098 22808
rect 22154 22752 22159 22808
rect 13169 22750 22159 22752
rect 13169 22747 13235 22750
rect 22093 22747 22159 22750
rect 29862 22748 29868 22812
rect 29932 22810 29938 22812
rect 32397 22810 32463 22813
rect 29932 22808 32463 22810
rect 29932 22752 32402 22808
rect 32458 22752 32463 22808
rect 29932 22750 32463 22752
rect 29932 22748 29938 22750
rect 32397 22747 32463 22750
rect 21909 22674 21975 22677
rect 23013 22674 23079 22677
rect 21909 22672 23079 22674
rect 0 22388 800 22628
rect 21909 22616 21914 22672
rect 21970 22616 23018 22672
rect 23074 22616 23079 22672
rect 21909 22614 23079 22616
rect 21909 22611 21975 22614
rect 23013 22611 23079 22614
rect 23289 22674 23355 22677
rect 25497 22674 25563 22677
rect 23289 22672 25563 22674
rect 23289 22616 23294 22672
rect 23350 22616 25502 22672
rect 25558 22616 25563 22672
rect 23289 22614 25563 22616
rect 23289 22611 23355 22614
rect 25497 22611 25563 22614
rect 27245 22674 27311 22677
rect 28257 22674 28323 22677
rect 27245 22672 28323 22674
rect 27245 22616 27250 22672
rect 27306 22616 28262 22672
rect 28318 22616 28323 22672
rect 27245 22614 28323 22616
rect 27245 22611 27311 22614
rect 28257 22611 28323 22614
rect 30557 22674 30623 22677
rect 30782 22674 30788 22676
rect 30557 22672 30788 22674
rect 30557 22616 30562 22672
rect 30618 22616 30788 22672
rect 30557 22614 30788 22616
rect 30557 22611 30623 22614
rect 30782 22612 30788 22614
rect 30852 22612 30858 22676
rect 31661 22674 31727 22677
rect 31526 22672 31727 22674
rect 31526 22616 31666 22672
rect 31722 22616 31727 22672
rect 31526 22614 31727 22616
rect 24577 22538 24643 22541
rect 27337 22538 27403 22541
rect 24577 22536 27403 22538
rect 24577 22480 24582 22536
rect 24638 22480 27342 22536
rect 27398 22480 27403 22536
rect 24577 22478 27403 22480
rect 24577 22475 24643 22478
rect 27337 22475 27403 22478
rect 30005 22538 30071 22541
rect 30373 22538 30439 22541
rect 30005 22536 30439 22538
rect 30005 22480 30010 22536
rect 30066 22480 30378 22536
rect 30434 22480 30439 22536
rect 30005 22478 30439 22480
rect 30005 22475 30071 22478
rect 30373 22475 30439 22478
rect 20069 22402 20135 22405
rect 24945 22402 25011 22405
rect 25957 22402 26023 22405
rect 20069 22400 26023 22402
rect 20069 22344 20074 22400
rect 20130 22344 24950 22400
rect 25006 22344 25962 22400
rect 26018 22344 26023 22400
rect 20069 22342 26023 22344
rect 20069 22339 20135 22342
rect 24945 22339 25011 22342
rect 25957 22339 26023 22342
rect 30097 22402 30163 22405
rect 30230 22402 30236 22404
rect 30097 22400 30236 22402
rect 30097 22344 30102 22400
rect 30158 22344 30236 22400
rect 30097 22342 30236 22344
rect 30097 22339 30163 22342
rect 30230 22340 30236 22342
rect 30300 22340 30306 22404
rect 30925 22402 30991 22405
rect 31526 22402 31586 22614
rect 31661 22611 31727 22614
rect 33041 22674 33107 22677
rect 33041 22672 33242 22674
rect 33041 22616 33046 22672
rect 33102 22616 33242 22672
rect 33041 22614 33242 22616
rect 33041 22611 33107 22614
rect 31845 22540 31911 22541
rect 31845 22538 31892 22540
rect 31800 22536 31892 22538
rect 31800 22480 31850 22536
rect 31800 22478 31892 22480
rect 31845 22476 31892 22478
rect 31956 22476 31962 22540
rect 32673 22538 32739 22541
rect 32446 22536 32739 22538
rect 32446 22480 32678 22536
rect 32734 22480 32739 22536
rect 32446 22478 32739 22480
rect 31845 22475 31911 22476
rect 31753 22404 31819 22405
rect 30925 22400 31586 22402
rect 30925 22344 30930 22400
rect 30986 22344 31586 22400
rect 30925 22342 31586 22344
rect 30925 22339 30991 22342
rect 31702 22340 31708 22404
rect 31772 22402 31819 22404
rect 31772 22400 31864 22402
rect 31814 22344 31864 22400
rect 31772 22342 31864 22344
rect 31772 22340 31819 22342
rect 31753 22339 31819 22340
rect 6576 22336 6896 22337
rect 6576 22272 6584 22336
rect 6648 22272 6664 22336
rect 6728 22272 6744 22336
rect 6808 22272 6824 22336
rect 6888 22272 6896 22336
rect 6576 22271 6896 22272
rect 17840 22336 18160 22337
rect 17840 22272 17848 22336
rect 17912 22272 17928 22336
rect 17992 22272 18008 22336
rect 18072 22272 18088 22336
rect 18152 22272 18160 22336
rect 17840 22271 18160 22272
rect 29104 22336 29424 22337
rect 29104 22272 29112 22336
rect 29176 22272 29192 22336
rect 29256 22272 29272 22336
rect 29336 22272 29352 22336
rect 29416 22272 29424 22336
rect 29104 22271 29424 22272
rect 23013 22266 23079 22269
rect 27061 22266 27127 22269
rect 23013 22264 27127 22266
rect 23013 22208 23018 22264
rect 23074 22208 27066 22264
rect 27122 22208 27127 22264
rect 23013 22206 27127 22208
rect 23013 22203 23079 22206
rect 27061 22203 27127 22206
rect 30097 22266 30163 22269
rect 32213 22266 32279 22269
rect 30097 22264 32279 22266
rect 30097 22208 30102 22264
rect 30158 22208 32218 22264
rect 32274 22208 32279 22264
rect 30097 22206 32279 22208
rect 30097 22203 30163 22206
rect 32213 22203 32279 22206
rect 19977 22130 20043 22133
rect 23105 22130 23171 22133
rect 19977 22128 23171 22130
rect 19977 22072 19982 22128
rect 20038 22072 23110 22128
rect 23166 22072 23171 22128
rect 19977 22070 23171 22072
rect 19977 22067 20043 22070
rect 23105 22067 23171 22070
rect 25262 22068 25268 22132
rect 25332 22130 25338 22132
rect 25405 22130 25471 22133
rect 25332 22128 25471 22130
rect 25332 22072 25410 22128
rect 25466 22072 25471 22128
rect 25332 22070 25471 22072
rect 25332 22068 25338 22070
rect 25405 22067 25471 22070
rect 32213 22130 32279 22133
rect 32446 22130 32506 22478
rect 32673 22475 32739 22478
rect 33182 22405 33242 22614
rect 33133 22400 33242 22405
rect 33133 22344 33138 22400
rect 33194 22344 33242 22400
rect 35200 22388 36000 22628
rect 33133 22342 33242 22344
rect 33133 22339 33199 22342
rect 32213 22128 32506 22130
rect 32213 22072 32218 22128
rect 32274 22072 32506 22128
rect 32213 22070 32506 22072
rect 32213 22067 32279 22070
rect 32622 22068 32628 22132
rect 32692 22130 32698 22132
rect 32857 22130 32923 22133
rect 32692 22128 32923 22130
rect 32692 22072 32862 22128
rect 32918 22072 32923 22128
rect 32692 22070 32923 22072
rect 32692 22068 32698 22070
rect 32857 22067 32923 22070
rect 25129 21994 25195 21997
rect 25405 21994 25471 21997
rect 25129 21992 25471 21994
rect 0 21708 800 21948
rect 25129 21936 25134 21992
rect 25190 21936 25410 21992
rect 25466 21936 25471 21992
rect 25129 21934 25471 21936
rect 25129 21931 25195 21934
rect 25405 21931 25471 21934
rect 25589 21994 25655 21997
rect 27061 21994 27127 21997
rect 30281 21996 30347 21997
rect 25589 21992 27127 21994
rect 25589 21936 25594 21992
rect 25650 21936 27066 21992
rect 27122 21936 27127 21992
rect 25589 21934 27127 21936
rect 25589 21931 25655 21934
rect 27061 21931 27127 21934
rect 30230 21932 30236 21996
rect 30300 21994 30347 21996
rect 30300 21992 30392 21994
rect 30342 21936 30392 21992
rect 30300 21934 30392 21936
rect 30300 21932 30347 21934
rect 30281 21931 30347 21932
rect 24761 21858 24827 21861
rect 28257 21858 28323 21861
rect 24761 21856 28323 21858
rect 24761 21800 24766 21856
rect 24822 21800 28262 21856
rect 28318 21800 28323 21856
rect 24761 21798 28323 21800
rect 24761 21795 24827 21798
rect 28257 21795 28323 21798
rect 29177 21858 29243 21861
rect 31661 21858 31727 21861
rect 29177 21856 31727 21858
rect 29177 21800 29182 21856
rect 29238 21800 31666 21856
rect 31722 21800 31727 21856
rect 29177 21798 31727 21800
rect 29177 21795 29243 21798
rect 31661 21795 31727 21798
rect 32397 21858 32463 21861
rect 32806 21858 32812 21860
rect 32397 21856 32812 21858
rect 32397 21800 32402 21856
rect 32458 21800 32812 21856
rect 32397 21798 32812 21800
rect 32397 21795 32463 21798
rect 32806 21796 32812 21798
rect 32876 21796 32882 21860
rect 12208 21792 12528 21793
rect 12208 21728 12216 21792
rect 12280 21728 12296 21792
rect 12360 21728 12376 21792
rect 12440 21728 12456 21792
rect 12520 21728 12528 21792
rect 12208 21727 12528 21728
rect 23472 21792 23792 21793
rect 23472 21728 23480 21792
rect 23544 21728 23560 21792
rect 23624 21728 23640 21792
rect 23704 21728 23720 21792
rect 23784 21728 23792 21792
rect 23472 21727 23792 21728
rect 26233 21722 26299 21725
rect 24166 21720 26299 21722
rect 24166 21664 26238 21720
rect 26294 21664 26299 21720
rect 24166 21662 26299 21664
rect 23565 21586 23631 21589
rect 24166 21586 24226 21662
rect 26233 21659 26299 21662
rect 23565 21584 24226 21586
rect 23565 21528 23570 21584
rect 23626 21528 24226 21584
rect 23565 21526 24226 21528
rect 24301 21586 24367 21589
rect 25773 21586 25839 21589
rect 24301 21584 25839 21586
rect 24301 21528 24306 21584
rect 24362 21528 25778 21584
rect 25834 21528 25839 21584
rect 24301 21526 25839 21528
rect 23565 21523 23631 21526
rect 24301 21523 24367 21526
rect 25773 21523 25839 21526
rect 29269 21586 29335 21589
rect 29269 21584 35266 21586
rect 29269 21528 29274 21584
rect 29330 21528 35266 21584
rect 29269 21526 35266 21528
rect 29269 21523 29335 21526
rect 20529 21450 20595 21453
rect 27889 21450 27955 21453
rect 20529 21448 27955 21450
rect 20529 21392 20534 21448
rect 20590 21392 27894 21448
rect 27950 21392 27955 21448
rect 20529 21390 27955 21392
rect 20529 21387 20595 21390
rect 27889 21387 27955 21390
rect 28441 21450 28507 21453
rect 30925 21450 30991 21453
rect 28441 21448 30991 21450
rect 28441 21392 28446 21448
rect 28502 21392 30930 21448
rect 30986 21392 30991 21448
rect 28441 21390 30991 21392
rect 28441 21387 28507 21390
rect 30925 21387 30991 21390
rect 20437 21314 20503 21317
rect 28073 21314 28139 21317
rect 30465 21316 30531 21317
rect 20437 21312 28139 21314
rect 0 21028 800 21268
rect 20437 21256 20442 21312
rect 20498 21256 28078 21312
rect 28134 21256 28139 21312
rect 20437 21254 28139 21256
rect 20437 21251 20503 21254
rect 28073 21251 28139 21254
rect 30414 21252 30420 21316
rect 30484 21314 30531 21316
rect 35206 21314 35266 21526
rect 30484 21312 30576 21314
rect 30526 21256 30576 21312
rect 30484 21254 30576 21256
rect 35022 21268 35266 21314
rect 35022 21254 36000 21268
rect 30484 21252 30531 21254
rect 30465 21251 30531 21252
rect 6576 21248 6896 21249
rect 6576 21184 6584 21248
rect 6648 21184 6664 21248
rect 6728 21184 6744 21248
rect 6808 21184 6824 21248
rect 6888 21184 6896 21248
rect 6576 21183 6896 21184
rect 17840 21248 18160 21249
rect 17840 21184 17848 21248
rect 17912 21184 17928 21248
rect 17992 21184 18008 21248
rect 18072 21184 18088 21248
rect 18152 21184 18160 21248
rect 17840 21183 18160 21184
rect 29104 21248 29424 21249
rect 29104 21184 29112 21248
rect 29176 21184 29192 21248
rect 29256 21184 29272 21248
rect 29336 21184 29352 21248
rect 29416 21184 29424 21248
rect 29104 21183 29424 21184
rect 25313 21180 25379 21181
rect 25262 21116 25268 21180
rect 25332 21178 25379 21180
rect 35022 21178 35082 21254
rect 35200 21178 36000 21254
rect 25332 21176 25424 21178
rect 25374 21120 25424 21176
rect 25332 21118 25424 21120
rect 35022 21118 36000 21178
rect 25332 21116 25379 21118
rect 25313 21115 25379 21116
rect 24577 21042 24643 21045
rect 24577 21040 25698 21042
rect 24577 20984 24582 21040
rect 24638 20984 25698 21040
rect 35200 21028 36000 21118
rect 24577 20982 25698 20984
rect 24577 20979 24643 20982
rect 22829 20906 22895 20909
rect 23197 20906 23263 20909
rect 24761 20906 24827 20909
rect 22829 20904 24827 20906
rect 22829 20848 22834 20904
rect 22890 20848 23202 20904
rect 23258 20848 24766 20904
rect 24822 20848 24827 20904
rect 22829 20846 24827 20848
rect 22829 20843 22895 20846
rect 23197 20843 23263 20846
rect 24761 20843 24827 20846
rect 25638 20773 25698 20982
rect 25638 20768 25747 20773
rect 25638 20712 25686 20768
rect 25742 20712 25747 20768
rect 25638 20710 25747 20712
rect 25681 20707 25747 20710
rect 26969 20770 27035 20773
rect 31017 20770 31083 20773
rect 26969 20768 31083 20770
rect 26969 20712 26974 20768
rect 27030 20712 31022 20768
rect 31078 20712 31083 20768
rect 26969 20710 31083 20712
rect 26969 20707 27035 20710
rect 31017 20707 31083 20710
rect 12208 20704 12528 20705
rect 12208 20640 12216 20704
rect 12280 20640 12296 20704
rect 12360 20640 12376 20704
rect 12440 20640 12456 20704
rect 12520 20640 12528 20704
rect 12208 20639 12528 20640
rect 23472 20704 23792 20705
rect 23472 20640 23480 20704
rect 23544 20640 23560 20704
rect 23624 20640 23640 20704
rect 23704 20640 23720 20704
rect 23784 20640 23792 20704
rect 23472 20639 23792 20640
rect 0 20348 800 20588
rect 23105 20498 23171 20501
rect 25957 20498 26023 20501
rect 31845 20500 31911 20501
rect 31845 20498 31892 20500
rect 23105 20496 26023 20498
rect 23105 20440 23110 20496
rect 23166 20440 25962 20496
rect 26018 20440 26023 20496
rect 23105 20438 26023 20440
rect 31800 20496 31892 20498
rect 31800 20440 31850 20496
rect 31800 20438 31892 20440
rect 23105 20435 23171 20438
rect 25957 20435 26023 20438
rect 31845 20436 31892 20438
rect 31956 20436 31962 20500
rect 34145 20498 34211 20501
rect 35200 20498 36000 20588
rect 34145 20496 36000 20498
rect 34145 20440 34150 20496
rect 34206 20440 36000 20496
rect 34145 20438 36000 20440
rect 31845 20435 31911 20436
rect 34145 20435 34211 20438
rect 21817 20362 21883 20365
rect 24117 20362 24183 20365
rect 21817 20360 24183 20362
rect 21817 20304 21822 20360
rect 21878 20304 24122 20360
rect 24178 20304 24183 20360
rect 35200 20348 36000 20438
rect 21817 20302 24183 20304
rect 21817 20299 21883 20302
rect 24117 20299 24183 20302
rect 6576 20160 6896 20161
rect 6576 20096 6584 20160
rect 6648 20096 6664 20160
rect 6728 20096 6744 20160
rect 6808 20096 6824 20160
rect 6888 20096 6896 20160
rect 6576 20095 6896 20096
rect 17840 20160 18160 20161
rect 17840 20096 17848 20160
rect 17912 20096 17928 20160
rect 17992 20096 18008 20160
rect 18072 20096 18088 20160
rect 18152 20096 18160 20160
rect 17840 20095 18160 20096
rect 29104 20160 29424 20161
rect 29104 20096 29112 20160
rect 29176 20096 29192 20160
rect 29256 20096 29272 20160
rect 29336 20096 29352 20160
rect 29416 20096 29424 20160
rect 29104 20095 29424 20096
rect 30005 20090 30071 20093
rect 30005 20088 30252 20090
rect 30005 20032 30010 20088
rect 30066 20032 30252 20088
rect 30005 20030 30252 20032
rect 30005 20027 30071 20030
rect 30192 19957 30252 20030
rect 30189 19952 30255 19957
rect 30189 19896 30194 19952
rect 30250 19896 30255 19952
rect 30189 19891 30255 19896
rect 22369 19818 22435 19821
rect 28625 19818 28691 19821
rect 22369 19816 28691 19818
rect 22369 19760 22374 19816
rect 22430 19760 28630 19816
rect 28686 19760 28691 19816
rect 22369 19758 28691 19760
rect 22369 19755 22435 19758
rect 28625 19755 28691 19758
rect 29545 19818 29611 19821
rect 30005 19818 30071 19821
rect 29545 19816 30071 19818
rect 29545 19760 29550 19816
rect 29606 19760 30010 19816
rect 30066 19760 30071 19816
rect 29545 19758 30071 19760
rect 29545 19755 29611 19758
rect 30005 19755 30071 19758
rect 34145 19818 34211 19821
rect 35200 19818 36000 19908
rect 34145 19816 36000 19818
rect 34145 19760 34150 19816
rect 34206 19760 36000 19816
rect 34145 19758 36000 19760
rect 34145 19755 34211 19758
rect 26417 19682 26483 19685
rect 27981 19682 28047 19685
rect 26417 19680 28047 19682
rect 26417 19624 26422 19680
rect 26478 19624 27986 19680
rect 28042 19624 28047 19680
rect 26417 19622 28047 19624
rect 26417 19619 26483 19622
rect 27981 19619 28047 19622
rect 29453 19682 29519 19685
rect 29678 19682 29684 19684
rect 29453 19680 29684 19682
rect 29453 19624 29458 19680
rect 29514 19624 29684 19680
rect 29453 19622 29684 19624
rect 29453 19619 29519 19622
rect 29678 19620 29684 19622
rect 29748 19620 29754 19684
rect 30560 19622 31632 19682
rect 35200 19668 36000 19758
rect 12208 19616 12528 19617
rect 12208 19552 12216 19616
rect 12280 19552 12296 19616
rect 12360 19552 12376 19616
rect 12440 19552 12456 19616
rect 12520 19552 12528 19616
rect 12208 19551 12528 19552
rect 23472 19616 23792 19617
rect 23472 19552 23480 19616
rect 23544 19552 23560 19616
rect 23624 19552 23640 19616
rect 23704 19552 23720 19616
rect 23784 19552 23792 19616
rect 23472 19551 23792 19552
rect 22185 19546 22251 19549
rect 22369 19546 22435 19549
rect 22185 19544 22435 19546
rect 22185 19488 22190 19544
rect 22246 19488 22374 19544
rect 22430 19488 22435 19544
rect 22185 19486 22435 19488
rect 22185 19483 22251 19486
rect 22369 19483 22435 19486
rect 29269 19546 29335 19549
rect 30560 19546 30620 19622
rect 31572 19549 31632 19622
rect 29269 19544 30620 19546
rect 29269 19488 29274 19544
rect 29330 19488 30620 19544
rect 29269 19486 30620 19488
rect 31569 19544 31635 19549
rect 31569 19488 31574 19544
rect 31630 19488 31635 19544
rect 29269 19483 29335 19486
rect 31569 19483 31635 19488
rect 20805 19410 20871 19413
rect 23933 19410 23999 19413
rect 29545 19412 29611 19413
rect 20805 19408 23999 19410
rect 20805 19352 20810 19408
rect 20866 19352 23938 19408
rect 23994 19352 23999 19408
rect 20805 19350 23999 19352
rect 20805 19347 20871 19350
rect 23933 19347 23999 19350
rect 29494 19348 29500 19412
rect 29564 19410 29611 19412
rect 29564 19408 29656 19410
rect 29606 19352 29656 19408
rect 29564 19350 29656 19352
rect 29564 19348 29611 19350
rect 30414 19348 30420 19412
rect 30484 19410 30490 19412
rect 30649 19410 30715 19413
rect 30484 19408 30715 19410
rect 30484 19352 30654 19408
rect 30710 19352 30715 19408
rect 30484 19350 30715 19352
rect 30484 19348 30490 19350
rect 29545 19347 29611 19348
rect 30649 19347 30715 19350
rect 0 19138 800 19228
rect 2221 19138 2287 19141
rect 0 19136 2287 19138
rect 0 19080 2226 19136
rect 2282 19080 2287 19136
rect 0 19078 2287 19080
rect 0 18988 800 19078
rect 2221 19075 2287 19078
rect 34145 19138 34211 19141
rect 35200 19138 36000 19228
rect 34145 19136 36000 19138
rect 34145 19080 34150 19136
rect 34206 19080 36000 19136
rect 34145 19078 36000 19080
rect 34145 19075 34211 19078
rect 6576 19072 6896 19073
rect 6576 19008 6584 19072
rect 6648 19008 6664 19072
rect 6728 19008 6744 19072
rect 6808 19008 6824 19072
rect 6888 19008 6896 19072
rect 6576 19007 6896 19008
rect 17840 19072 18160 19073
rect 17840 19008 17848 19072
rect 17912 19008 17928 19072
rect 17992 19008 18008 19072
rect 18072 19008 18088 19072
rect 18152 19008 18160 19072
rect 17840 19007 18160 19008
rect 29104 19072 29424 19073
rect 29104 19008 29112 19072
rect 29176 19008 29192 19072
rect 29256 19008 29272 19072
rect 29336 19008 29352 19072
rect 29416 19008 29424 19072
rect 29104 19007 29424 19008
rect 35200 18988 36000 19078
rect 30097 18596 30163 18597
rect 30046 18594 30052 18596
rect 0 18458 800 18548
rect 30006 18534 30052 18594
rect 30116 18592 30163 18596
rect 30158 18536 30163 18592
rect 30046 18532 30052 18534
rect 30116 18532 30163 18536
rect 30097 18531 30163 18532
rect 12208 18528 12528 18529
rect 12208 18464 12216 18528
rect 12280 18464 12296 18528
rect 12360 18464 12376 18528
rect 12440 18464 12456 18528
rect 12520 18464 12528 18528
rect 12208 18463 12528 18464
rect 23472 18528 23792 18529
rect 23472 18464 23480 18528
rect 23544 18464 23560 18528
rect 23624 18464 23640 18528
rect 23704 18464 23720 18528
rect 23784 18464 23792 18528
rect 23472 18463 23792 18464
rect 2865 18458 2931 18461
rect 0 18456 2931 18458
rect 0 18400 2870 18456
rect 2926 18400 2931 18456
rect 0 18398 2931 18400
rect 0 18308 800 18398
rect 2865 18395 2931 18398
rect 35200 18308 36000 18548
rect 6576 17984 6896 17985
rect 6576 17920 6584 17984
rect 6648 17920 6664 17984
rect 6728 17920 6744 17984
rect 6808 17920 6824 17984
rect 6888 17920 6896 17984
rect 6576 17919 6896 17920
rect 17840 17984 18160 17985
rect 17840 17920 17848 17984
rect 17912 17920 17928 17984
rect 17992 17920 18008 17984
rect 18072 17920 18088 17984
rect 18152 17920 18160 17984
rect 17840 17919 18160 17920
rect 29104 17984 29424 17985
rect 29104 17920 29112 17984
rect 29176 17920 29192 17984
rect 29256 17920 29272 17984
rect 29336 17920 29352 17984
rect 29416 17920 29424 17984
rect 29104 17919 29424 17920
rect 0 17628 800 17868
rect 34145 17778 34211 17781
rect 35200 17778 36000 17868
rect 34145 17776 36000 17778
rect 34145 17720 34150 17776
rect 34206 17720 36000 17776
rect 34145 17718 36000 17720
rect 34145 17715 34211 17718
rect 35200 17628 36000 17718
rect 12208 17440 12528 17441
rect 12208 17376 12216 17440
rect 12280 17376 12296 17440
rect 12360 17376 12376 17440
rect 12440 17376 12456 17440
rect 12520 17376 12528 17440
rect 12208 17375 12528 17376
rect 23472 17440 23792 17441
rect 23472 17376 23480 17440
rect 23544 17376 23560 17440
rect 23624 17376 23640 17440
rect 23704 17376 23720 17440
rect 23784 17376 23792 17440
rect 23472 17375 23792 17376
rect 23289 17234 23355 17237
rect 25405 17234 25471 17237
rect 23289 17232 25471 17234
rect 0 17098 800 17188
rect 23289 17176 23294 17232
rect 23350 17176 25410 17232
rect 25466 17176 25471 17232
rect 23289 17174 25471 17176
rect 23289 17171 23355 17174
rect 25405 17171 25471 17174
rect 1945 17098 2011 17101
rect 0 17096 2011 17098
rect 0 17040 1950 17096
rect 2006 17040 2011 17096
rect 0 17038 2011 17040
rect 0 16948 800 17038
rect 1945 17035 2011 17038
rect 34145 17098 34211 17101
rect 35200 17098 36000 17188
rect 34145 17096 36000 17098
rect 34145 17040 34150 17096
rect 34206 17040 36000 17096
rect 34145 17038 36000 17040
rect 34145 17035 34211 17038
rect 35200 16948 36000 17038
rect 6576 16896 6896 16897
rect 6576 16832 6584 16896
rect 6648 16832 6664 16896
rect 6728 16832 6744 16896
rect 6808 16832 6824 16896
rect 6888 16832 6896 16896
rect 6576 16831 6896 16832
rect 17840 16896 18160 16897
rect 17840 16832 17848 16896
rect 17912 16832 17928 16896
rect 17992 16832 18008 16896
rect 18072 16832 18088 16896
rect 18152 16832 18160 16896
rect 17840 16831 18160 16832
rect 29104 16896 29424 16897
rect 29104 16832 29112 16896
rect 29176 16832 29192 16896
rect 29256 16832 29272 16896
rect 29336 16832 29352 16896
rect 29416 16832 29424 16896
rect 29104 16831 29424 16832
rect 0 16268 800 16508
rect 34145 16418 34211 16421
rect 35200 16418 36000 16508
rect 34145 16416 36000 16418
rect 34145 16360 34150 16416
rect 34206 16360 36000 16416
rect 34145 16358 36000 16360
rect 34145 16355 34211 16358
rect 12208 16352 12528 16353
rect 12208 16288 12216 16352
rect 12280 16288 12296 16352
rect 12360 16288 12376 16352
rect 12440 16288 12456 16352
rect 12520 16288 12528 16352
rect 12208 16287 12528 16288
rect 23472 16352 23792 16353
rect 23472 16288 23480 16352
rect 23544 16288 23560 16352
rect 23624 16288 23640 16352
rect 23704 16288 23720 16352
rect 23784 16288 23792 16352
rect 23472 16287 23792 16288
rect 35200 16268 36000 16358
rect 0 15738 800 15828
rect 6576 15808 6896 15809
rect 6576 15744 6584 15808
rect 6648 15744 6664 15808
rect 6728 15744 6744 15808
rect 6808 15744 6824 15808
rect 6888 15744 6896 15808
rect 6576 15743 6896 15744
rect 17840 15808 18160 15809
rect 17840 15744 17848 15808
rect 17912 15744 17928 15808
rect 17992 15744 18008 15808
rect 18072 15744 18088 15808
rect 18152 15744 18160 15808
rect 17840 15743 18160 15744
rect 29104 15808 29424 15809
rect 29104 15744 29112 15808
rect 29176 15744 29192 15808
rect 29256 15744 29272 15808
rect 29336 15744 29352 15808
rect 29416 15744 29424 15808
rect 29104 15743 29424 15744
rect 2773 15738 2839 15741
rect 0 15736 2839 15738
rect 0 15680 2778 15736
rect 2834 15680 2839 15736
rect 0 15678 2839 15680
rect 0 15588 800 15678
rect 2773 15675 2839 15678
rect 35200 15588 36000 15828
rect 12208 15264 12528 15265
rect 12208 15200 12216 15264
rect 12280 15200 12296 15264
rect 12360 15200 12376 15264
rect 12440 15200 12456 15264
rect 12520 15200 12528 15264
rect 12208 15199 12528 15200
rect 23472 15264 23792 15265
rect 23472 15200 23480 15264
rect 23544 15200 23560 15264
rect 23624 15200 23640 15264
rect 23704 15200 23720 15264
rect 23784 15200 23792 15264
rect 23472 15199 23792 15200
rect 0 14908 800 15148
rect 6576 14720 6896 14721
rect 6576 14656 6584 14720
rect 6648 14656 6664 14720
rect 6728 14656 6744 14720
rect 6808 14656 6824 14720
rect 6888 14656 6896 14720
rect 6576 14655 6896 14656
rect 17840 14720 18160 14721
rect 17840 14656 17848 14720
rect 17912 14656 17928 14720
rect 17992 14656 18008 14720
rect 18072 14656 18088 14720
rect 18152 14656 18160 14720
rect 17840 14655 18160 14656
rect 29104 14720 29424 14721
rect 29104 14656 29112 14720
rect 29176 14656 29192 14720
rect 29256 14656 29272 14720
rect 29336 14656 29352 14720
rect 29416 14656 29424 14720
rect 29104 14655 29424 14656
rect 0 14378 800 14468
rect 1945 14378 2011 14381
rect 0 14376 2011 14378
rect 0 14320 1950 14376
rect 2006 14320 2011 14376
rect 0 14318 2011 14320
rect 0 14228 800 14318
rect 1945 14315 2011 14318
rect 34145 14378 34211 14381
rect 35200 14378 36000 14468
rect 34145 14376 36000 14378
rect 34145 14320 34150 14376
rect 34206 14320 36000 14376
rect 34145 14318 36000 14320
rect 34145 14315 34211 14318
rect 35200 14228 36000 14318
rect 12208 14176 12528 14177
rect 12208 14112 12216 14176
rect 12280 14112 12296 14176
rect 12360 14112 12376 14176
rect 12440 14112 12456 14176
rect 12520 14112 12528 14176
rect 12208 14111 12528 14112
rect 23472 14176 23792 14177
rect 23472 14112 23480 14176
rect 23544 14112 23560 14176
rect 23624 14112 23640 14176
rect 23704 14112 23720 14176
rect 23784 14112 23792 14176
rect 23472 14111 23792 14112
rect 0 13698 800 13788
rect 2773 13698 2839 13701
rect 0 13696 2839 13698
rect 0 13640 2778 13696
rect 2834 13640 2839 13696
rect 0 13638 2839 13640
rect 0 13548 800 13638
rect 2773 13635 2839 13638
rect 34145 13698 34211 13701
rect 35200 13698 36000 13788
rect 34145 13696 36000 13698
rect 34145 13640 34150 13696
rect 34206 13640 36000 13696
rect 34145 13638 36000 13640
rect 34145 13635 34211 13638
rect 6576 13632 6896 13633
rect 6576 13568 6584 13632
rect 6648 13568 6664 13632
rect 6728 13568 6744 13632
rect 6808 13568 6824 13632
rect 6888 13568 6896 13632
rect 6576 13567 6896 13568
rect 17840 13632 18160 13633
rect 17840 13568 17848 13632
rect 17912 13568 17928 13632
rect 17992 13568 18008 13632
rect 18072 13568 18088 13632
rect 18152 13568 18160 13632
rect 17840 13567 18160 13568
rect 29104 13632 29424 13633
rect 29104 13568 29112 13632
rect 29176 13568 29192 13632
rect 29256 13568 29272 13632
rect 29336 13568 29352 13632
rect 29416 13568 29424 13632
rect 29104 13567 29424 13568
rect 35200 13548 36000 13638
rect 12208 13088 12528 13089
rect 12208 13024 12216 13088
rect 12280 13024 12296 13088
rect 12360 13024 12376 13088
rect 12440 13024 12456 13088
rect 12520 13024 12528 13088
rect 12208 13023 12528 13024
rect 23472 13088 23792 13089
rect 23472 13024 23480 13088
rect 23544 13024 23560 13088
rect 23624 13024 23640 13088
rect 23704 13024 23720 13088
rect 23784 13024 23792 13088
rect 23472 13023 23792 13024
rect 34145 13018 34211 13021
rect 35200 13018 36000 13108
rect 34145 13016 36000 13018
rect 34145 12960 34150 13016
rect 34206 12960 36000 13016
rect 34145 12958 36000 12960
rect 34145 12955 34211 12958
rect 35200 12868 36000 12958
rect 6576 12544 6896 12545
rect 6576 12480 6584 12544
rect 6648 12480 6664 12544
rect 6728 12480 6744 12544
rect 6808 12480 6824 12544
rect 6888 12480 6896 12544
rect 6576 12479 6896 12480
rect 17840 12544 18160 12545
rect 17840 12480 17848 12544
rect 17912 12480 17928 12544
rect 17992 12480 18008 12544
rect 18072 12480 18088 12544
rect 18152 12480 18160 12544
rect 17840 12479 18160 12480
rect 29104 12544 29424 12545
rect 29104 12480 29112 12544
rect 29176 12480 29192 12544
rect 29256 12480 29272 12544
rect 29336 12480 29352 12544
rect 29416 12480 29424 12544
rect 29104 12479 29424 12480
rect 0 12188 800 12428
rect 34145 12338 34211 12341
rect 35200 12338 36000 12428
rect 34145 12336 36000 12338
rect 34145 12280 34150 12336
rect 34206 12280 36000 12336
rect 34145 12278 36000 12280
rect 34145 12275 34211 12278
rect 35200 12188 36000 12278
rect 12208 12000 12528 12001
rect 12208 11936 12216 12000
rect 12280 11936 12296 12000
rect 12360 11936 12376 12000
rect 12440 11936 12456 12000
rect 12520 11936 12528 12000
rect 12208 11935 12528 11936
rect 23472 12000 23792 12001
rect 23472 11936 23480 12000
rect 23544 11936 23560 12000
rect 23624 11936 23640 12000
rect 23704 11936 23720 12000
rect 23784 11936 23792 12000
rect 23472 11935 23792 11936
rect 0 11658 800 11748
rect 2773 11658 2839 11661
rect 0 11656 2839 11658
rect 0 11600 2778 11656
rect 2834 11600 2839 11656
rect 0 11598 2839 11600
rect 0 11508 800 11598
rect 2773 11595 2839 11598
rect 35200 11508 36000 11748
rect 6576 11456 6896 11457
rect 6576 11392 6584 11456
rect 6648 11392 6664 11456
rect 6728 11392 6744 11456
rect 6808 11392 6824 11456
rect 6888 11392 6896 11456
rect 6576 11391 6896 11392
rect 17840 11456 18160 11457
rect 17840 11392 17848 11456
rect 17912 11392 17928 11456
rect 17992 11392 18008 11456
rect 18072 11392 18088 11456
rect 18152 11392 18160 11456
rect 17840 11391 18160 11392
rect 29104 11456 29424 11457
rect 29104 11392 29112 11456
rect 29176 11392 29192 11456
rect 29256 11392 29272 11456
rect 29336 11392 29352 11456
rect 29416 11392 29424 11456
rect 29104 11391 29424 11392
rect 0 10978 800 11068
rect 1853 10978 1919 10981
rect 0 10976 1919 10978
rect 0 10920 1858 10976
rect 1914 10920 1919 10976
rect 0 10918 1919 10920
rect 0 10828 800 10918
rect 1853 10915 1919 10918
rect 12208 10912 12528 10913
rect 12208 10848 12216 10912
rect 12280 10848 12296 10912
rect 12360 10848 12376 10912
rect 12440 10848 12456 10912
rect 12520 10848 12528 10912
rect 12208 10847 12528 10848
rect 23472 10912 23792 10913
rect 23472 10848 23480 10912
rect 23544 10848 23560 10912
rect 23624 10848 23640 10912
rect 23704 10848 23720 10912
rect 23784 10848 23792 10912
rect 23472 10847 23792 10848
rect 35200 10828 36000 11068
rect 0 10148 800 10388
rect 6576 10368 6896 10369
rect 6576 10304 6584 10368
rect 6648 10304 6664 10368
rect 6728 10304 6744 10368
rect 6808 10304 6824 10368
rect 6888 10304 6896 10368
rect 6576 10303 6896 10304
rect 17840 10368 18160 10369
rect 17840 10304 17848 10368
rect 17912 10304 17928 10368
rect 17992 10304 18008 10368
rect 18072 10304 18088 10368
rect 18152 10304 18160 10368
rect 17840 10303 18160 10304
rect 29104 10368 29424 10369
rect 29104 10304 29112 10368
rect 29176 10304 29192 10368
rect 29256 10304 29272 10368
rect 29336 10304 29352 10368
rect 29416 10304 29424 10368
rect 29104 10303 29424 10304
rect 35200 10148 36000 10388
rect 12208 9824 12528 9825
rect 12208 9760 12216 9824
rect 12280 9760 12296 9824
rect 12360 9760 12376 9824
rect 12440 9760 12456 9824
rect 12520 9760 12528 9824
rect 12208 9759 12528 9760
rect 23472 9824 23792 9825
rect 23472 9760 23480 9824
rect 23544 9760 23560 9824
rect 23624 9760 23640 9824
rect 23704 9760 23720 9824
rect 23784 9760 23792 9824
rect 23472 9759 23792 9760
rect 0 9468 800 9708
rect 33961 9618 34027 9621
rect 35200 9618 36000 9708
rect 33961 9616 36000 9618
rect 33961 9560 33966 9616
rect 34022 9560 36000 9616
rect 33961 9558 36000 9560
rect 33961 9555 34027 9558
rect 35200 9468 36000 9558
rect 6576 9280 6896 9281
rect 6576 9216 6584 9280
rect 6648 9216 6664 9280
rect 6728 9216 6744 9280
rect 6808 9216 6824 9280
rect 6888 9216 6896 9280
rect 6576 9215 6896 9216
rect 17840 9280 18160 9281
rect 17840 9216 17848 9280
rect 17912 9216 17928 9280
rect 17992 9216 18008 9280
rect 18072 9216 18088 9280
rect 18152 9216 18160 9280
rect 17840 9215 18160 9216
rect 29104 9280 29424 9281
rect 29104 9216 29112 9280
rect 29176 9216 29192 9280
rect 29256 9216 29272 9280
rect 29336 9216 29352 9280
rect 29416 9216 29424 9280
rect 29104 9215 29424 9216
rect 0 8938 800 9028
rect 2865 8938 2931 8941
rect 0 8936 2931 8938
rect 0 8880 2870 8936
rect 2926 8880 2931 8936
rect 0 8878 2931 8880
rect 0 8788 800 8878
rect 2865 8875 2931 8878
rect 34145 8938 34211 8941
rect 35200 8938 36000 9028
rect 34145 8936 36000 8938
rect 34145 8880 34150 8936
rect 34206 8880 36000 8936
rect 34145 8878 36000 8880
rect 34145 8875 34211 8878
rect 35200 8788 36000 8878
rect 12208 8736 12528 8737
rect 12208 8672 12216 8736
rect 12280 8672 12296 8736
rect 12360 8672 12376 8736
rect 12440 8672 12456 8736
rect 12520 8672 12528 8736
rect 12208 8671 12528 8672
rect 23472 8736 23792 8737
rect 23472 8672 23480 8736
rect 23544 8672 23560 8736
rect 23624 8672 23640 8736
rect 23704 8672 23720 8736
rect 23784 8672 23792 8736
rect 23472 8671 23792 8672
rect 0 8258 800 8348
rect 2773 8258 2839 8261
rect 0 8256 2839 8258
rect 0 8200 2778 8256
rect 2834 8200 2839 8256
rect 0 8198 2839 8200
rect 0 8108 800 8198
rect 2773 8195 2839 8198
rect 6576 8192 6896 8193
rect 6576 8128 6584 8192
rect 6648 8128 6664 8192
rect 6728 8128 6744 8192
rect 6808 8128 6824 8192
rect 6888 8128 6896 8192
rect 6576 8127 6896 8128
rect 17840 8192 18160 8193
rect 17840 8128 17848 8192
rect 17912 8128 17928 8192
rect 17992 8128 18008 8192
rect 18072 8128 18088 8192
rect 18152 8128 18160 8192
rect 17840 8127 18160 8128
rect 29104 8192 29424 8193
rect 29104 8128 29112 8192
rect 29176 8128 29192 8192
rect 29256 8128 29272 8192
rect 29336 8128 29352 8192
rect 29416 8128 29424 8192
rect 29104 8127 29424 8128
rect 0 7578 800 7668
rect 12208 7648 12528 7649
rect 12208 7584 12216 7648
rect 12280 7584 12296 7648
rect 12360 7584 12376 7648
rect 12440 7584 12456 7648
rect 12520 7584 12528 7648
rect 12208 7583 12528 7584
rect 23472 7648 23792 7649
rect 23472 7584 23480 7648
rect 23544 7584 23560 7648
rect 23624 7584 23640 7648
rect 23704 7584 23720 7648
rect 23784 7584 23792 7648
rect 23472 7583 23792 7584
rect 2773 7578 2839 7581
rect 0 7576 2839 7578
rect 0 7520 2778 7576
rect 2834 7520 2839 7576
rect 0 7518 2839 7520
rect 0 7428 800 7518
rect 2773 7515 2839 7518
rect 35200 7428 36000 7668
rect 6576 7104 6896 7105
rect 6576 7040 6584 7104
rect 6648 7040 6664 7104
rect 6728 7040 6744 7104
rect 6808 7040 6824 7104
rect 6888 7040 6896 7104
rect 6576 7039 6896 7040
rect 17840 7104 18160 7105
rect 17840 7040 17848 7104
rect 17912 7040 17928 7104
rect 17992 7040 18008 7104
rect 18072 7040 18088 7104
rect 18152 7040 18160 7104
rect 17840 7039 18160 7040
rect 29104 7104 29424 7105
rect 29104 7040 29112 7104
rect 29176 7040 29192 7104
rect 29256 7040 29272 7104
rect 29336 7040 29352 7104
rect 29416 7040 29424 7104
rect 29104 7039 29424 7040
rect 0 6748 800 6988
rect 34145 6898 34211 6901
rect 35200 6898 36000 6988
rect 34145 6896 36000 6898
rect 34145 6840 34150 6896
rect 34206 6840 36000 6896
rect 34145 6838 36000 6840
rect 34145 6835 34211 6838
rect 35200 6748 36000 6838
rect 12208 6560 12528 6561
rect 12208 6496 12216 6560
rect 12280 6496 12296 6560
rect 12360 6496 12376 6560
rect 12440 6496 12456 6560
rect 12520 6496 12528 6560
rect 12208 6495 12528 6496
rect 23472 6560 23792 6561
rect 23472 6496 23480 6560
rect 23544 6496 23560 6560
rect 23624 6496 23640 6560
rect 23704 6496 23720 6560
rect 23784 6496 23792 6560
rect 23472 6495 23792 6496
rect 35200 6068 36000 6308
rect 6576 6016 6896 6017
rect 6576 5952 6584 6016
rect 6648 5952 6664 6016
rect 6728 5952 6744 6016
rect 6808 5952 6824 6016
rect 6888 5952 6896 6016
rect 6576 5951 6896 5952
rect 17840 6016 18160 6017
rect 17840 5952 17848 6016
rect 17912 5952 17928 6016
rect 17992 5952 18008 6016
rect 18072 5952 18088 6016
rect 18152 5952 18160 6016
rect 17840 5951 18160 5952
rect 29104 6016 29424 6017
rect 29104 5952 29112 6016
rect 29176 5952 29192 6016
rect 29256 5952 29272 6016
rect 29336 5952 29352 6016
rect 29416 5952 29424 6016
rect 29104 5951 29424 5952
rect 0 5538 800 5628
rect 1853 5538 1919 5541
rect 0 5536 1919 5538
rect 0 5480 1858 5536
rect 1914 5480 1919 5536
rect 0 5478 1919 5480
rect 0 5388 800 5478
rect 1853 5475 1919 5478
rect 12208 5472 12528 5473
rect 12208 5408 12216 5472
rect 12280 5408 12296 5472
rect 12360 5408 12376 5472
rect 12440 5408 12456 5472
rect 12520 5408 12528 5472
rect 12208 5407 12528 5408
rect 23472 5472 23792 5473
rect 23472 5408 23480 5472
rect 23544 5408 23560 5472
rect 23624 5408 23640 5472
rect 23704 5408 23720 5472
rect 23784 5408 23792 5472
rect 23472 5407 23792 5408
rect 35200 5388 36000 5628
rect 0 4858 800 4948
rect 6576 4928 6896 4929
rect 6576 4864 6584 4928
rect 6648 4864 6664 4928
rect 6728 4864 6744 4928
rect 6808 4864 6824 4928
rect 6888 4864 6896 4928
rect 6576 4863 6896 4864
rect 17840 4928 18160 4929
rect 17840 4864 17848 4928
rect 17912 4864 17928 4928
rect 17992 4864 18008 4928
rect 18072 4864 18088 4928
rect 18152 4864 18160 4928
rect 17840 4863 18160 4864
rect 29104 4928 29424 4929
rect 29104 4864 29112 4928
rect 29176 4864 29192 4928
rect 29256 4864 29272 4928
rect 29336 4864 29352 4928
rect 29416 4864 29424 4928
rect 29104 4863 29424 4864
rect 3049 4858 3115 4861
rect 0 4856 3115 4858
rect 0 4800 3054 4856
rect 3110 4800 3115 4856
rect 0 4798 3115 4800
rect 0 4708 800 4798
rect 3049 4795 3115 4798
rect 34145 4858 34211 4861
rect 35200 4858 36000 4948
rect 34145 4856 36000 4858
rect 34145 4800 34150 4856
rect 34206 4800 36000 4856
rect 34145 4798 36000 4800
rect 34145 4795 34211 4798
rect 35200 4708 36000 4798
rect 12208 4384 12528 4385
rect 12208 4320 12216 4384
rect 12280 4320 12296 4384
rect 12360 4320 12376 4384
rect 12440 4320 12456 4384
rect 12520 4320 12528 4384
rect 12208 4319 12528 4320
rect 23472 4384 23792 4385
rect 23472 4320 23480 4384
rect 23544 4320 23560 4384
rect 23624 4320 23640 4384
rect 23704 4320 23720 4384
rect 23784 4320 23792 4384
rect 23472 4319 23792 4320
rect 0 4178 800 4268
rect 2957 4178 3023 4181
rect 0 4176 3023 4178
rect 0 4120 2962 4176
rect 3018 4120 3023 4176
rect 0 4118 3023 4120
rect 0 4028 800 4118
rect 2957 4115 3023 4118
rect 34145 4178 34211 4181
rect 35200 4178 36000 4268
rect 34145 4176 36000 4178
rect 34145 4120 34150 4176
rect 34206 4120 36000 4176
rect 34145 4118 36000 4120
rect 34145 4115 34211 4118
rect 35200 4028 36000 4118
rect 6576 3840 6896 3841
rect 6576 3776 6584 3840
rect 6648 3776 6664 3840
rect 6728 3776 6744 3840
rect 6808 3776 6824 3840
rect 6888 3776 6896 3840
rect 6576 3775 6896 3776
rect 17840 3840 18160 3841
rect 17840 3776 17848 3840
rect 17912 3776 17928 3840
rect 17992 3776 18008 3840
rect 18072 3776 18088 3840
rect 18152 3776 18160 3840
rect 17840 3775 18160 3776
rect 29104 3840 29424 3841
rect 29104 3776 29112 3840
rect 29176 3776 29192 3840
rect 29256 3776 29272 3840
rect 29336 3776 29352 3840
rect 29416 3776 29424 3840
rect 29104 3775 29424 3776
rect 0 3498 800 3588
rect 3233 3498 3299 3501
rect 0 3496 3299 3498
rect 0 3440 3238 3496
rect 3294 3440 3299 3496
rect 0 3438 3299 3440
rect 0 3348 800 3438
rect 3233 3435 3299 3438
rect 33041 3498 33107 3501
rect 35200 3498 36000 3588
rect 33041 3496 36000 3498
rect 33041 3440 33046 3496
rect 33102 3440 36000 3496
rect 33041 3438 36000 3440
rect 33041 3435 33107 3438
rect 35200 3348 36000 3438
rect 12208 3296 12528 3297
rect 12208 3232 12216 3296
rect 12280 3232 12296 3296
rect 12360 3232 12376 3296
rect 12440 3232 12456 3296
rect 12520 3232 12528 3296
rect 12208 3231 12528 3232
rect 23472 3296 23792 3297
rect 23472 3232 23480 3296
rect 23544 3232 23560 3296
rect 23624 3232 23640 3296
rect 23704 3232 23720 3296
rect 23784 3232 23792 3296
rect 23472 3231 23792 3232
rect 0 2818 800 2908
rect 2773 2818 2839 2821
rect 0 2816 2839 2818
rect 0 2760 2778 2816
rect 2834 2760 2839 2816
rect 0 2758 2839 2760
rect 0 2668 800 2758
rect 2773 2755 2839 2758
rect 6576 2752 6896 2753
rect 6576 2688 6584 2752
rect 6648 2688 6664 2752
rect 6728 2688 6744 2752
rect 6808 2688 6824 2752
rect 6888 2688 6896 2752
rect 6576 2687 6896 2688
rect 17840 2752 18160 2753
rect 17840 2688 17848 2752
rect 17912 2688 17928 2752
rect 17992 2688 18008 2752
rect 18072 2688 18088 2752
rect 18152 2688 18160 2752
rect 17840 2687 18160 2688
rect 29104 2752 29424 2753
rect 29104 2688 29112 2752
rect 29176 2688 29192 2752
rect 29256 2688 29272 2752
rect 29336 2688 29352 2752
rect 29416 2688 29424 2752
rect 29104 2687 29424 2688
rect 35200 2668 36000 2908
rect 0 2138 800 2228
rect 12208 2208 12528 2209
rect 12208 2144 12216 2208
rect 12280 2144 12296 2208
rect 12360 2144 12376 2208
rect 12440 2144 12456 2208
rect 12520 2144 12528 2208
rect 12208 2143 12528 2144
rect 23472 2208 23792 2209
rect 23472 2144 23480 2208
rect 23544 2144 23560 2208
rect 23624 2144 23640 2208
rect 23704 2144 23720 2208
rect 23784 2144 23792 2208
rect 23472 2143 23792 2144
rect 2865 2138 2931 2141
rect 0 2136 2931 2138
rect 0 2080 2870 2136
rect 2926 2080 2931 2136
rect 0 2078 2931 2080
rect 0 1988 800 2078
rect 2865 2075 2931 2078
rect 32029 2138 32095 2141
rect 35200 2138 36000 2228
rect 32029 2136 36000 2138
rect 32029 2080 32034 2136
rect 32090 2080 36000 2136
rect 32029 2078 36000 2080
rect 32029 2075 32095 2078
rect 35200 1988 36000 2078
rect 0 1458 800 1548
rect 3417 1458 3483 1461
rect 0 1456 3483 1458
rect 0 1400 3422 1456
rect 3478 1400 3483 1456
rect 0 1398 3483 1400
rect 0 1308 800 1398
rect 3417 1395 3483 1398
rect 0 628 800 868
rect 34421 778 34487 781
rect 35200 778 36000 868
rect 34421 776 36000 778
rect 34421 720 34426 776
rect 34482 720 36000 776
rect 34421 718 36000 720
rect 34421 715 34487 718
rect 35200 628 36000 718
rect 32581 98 32647 101
rect 35200 98 36000 188
rect 32581 96 36000 98
rect 32581 40 32586 96
rect 32642 40 36000 96
rect 32581 38 36000 40
rect 32581 35 32647 38
rect 35200 -52 36000 38
<< via3 >>
rect 14596 40836 14660 40900
rect 18460 40428 18524 40492
rect 12020 39748 12084 39812
rect 6584 39740 6648 39744
rect 6584 39684 6588 39740
rect 6588 39684 6644 39740
rect 6644 39684 6648 39740
rect 6584 39680 6648 39684
rect 6664 39740 6728 39744
rect 6664 39684 6668 39740
rect 6668 39684 6724 39740
rect 6724 39684 6728 39740
rect 6664 39680 6728 39684
rect 6744 39740 6808 39744
rect 6744 39684 6748 39740
rect 6748 39684 6804 39740
rect 6804 39684 6808 39740
rect 6744 39680 6808 39684
rect 6824 39740 6888 39744
rect 6824 39684 6828 39740
rect 6828 39684 6884 39740
rect 6884 39684 6888 39740
rect 6824 39680 6888 39684
rect 17848 39740 17912 39744
rect 17848 39684 17852 39740
rect 17852 39684 17908 39740
rect 17908 39684 17912 39740
rect 17848 39680 17912 39684
rect 17928 39740 17992 39744
rect 17928 39684 17932 39740
rect 17932 39684 17988 39740
rect 17988 39684 17992 39740
rect 17928 39680 17992 39684
rect 18008 39740 18072 39744
rect 18008 39684 18012 39740
rect 18012 39684 18068 39740
rect 18068 39684 18072 39740
rect 18008 39680 18072 39684
rect 18088 39740 18152 39744
rect 18088 39684 18092 39740
rect 18092 39684 18148 39740
rect 18148 39684 18152 39740
rect 18088 39680 18152 39684
rect 29112 39740 29176 39744
rect 29112 39684 29116 39740
rect 29116 39684 29172 39740
rect 29172 39684 29176 39740
rect 29112 39680 29176 39684
rect 29192 39740 29256 39744
rect 29192 39684 29196 39740
rect 29196 39684 29252 39740
rect 29252 39684 29256 39740
rect 29192 39680 29256 39684
rect 29272 39740 29336 39744
rect 29272 39684 29276 39740
rect 29276 39684 29332 39740
rect 29332 39684 29336 39740
rect 29272 39680 29336 39684
rect 29352 39740 29416 39744
rect 29352 39684 29356 39740
rect 29356 39684 29412 39740
rect 29412 39684 29416 39740
rect 29352 39680 29416 39684
rect 12216 39196 12280 39200
rect 12216 39140 12220 39196
rect 12220 39140 12276 39196
rect 12276 39140 12280 39196
rect 12216 39136 12280 39140
rect 12296 39196 12360 39200
rect 12296 39140 12300 39196
rect 12300 39140 12356 39196
rect 12356 39140 12360 39196
rect 12296 39136 12360 39140
rect 12376 39196 12440 39200
rect 12376 39140 12380 39196
rect 12380 39140 12436 39196
rect 12436 39140 12440 39196
rect 12376 39136 12440 39140
rect 12456 39196 12520 39200
rect 12456 39140 12460 39196
rect 12460 39140 12516 39196
rect 12516 39140 12520 39196
rect 12456 39136 12520 39140
rect 18460 39068 18524 39132
rect 23480 39196 23544 39200
rect 23480 39140 23484 39196
rect 23484 39140 23540 39196
rect 23540 39140 23544 39196
rect 23480 39136 23544 39140
rect 23560 39196 23624 39200
rect 23560 39140 23564 39196
rect 23564 39140 23620 39196
rect 23620 39140 23624 39196
rect 23560 39136 23624 39140
rect 23640 39196 23704 39200
rect 23640 39140 23644 39196
rect 23644 39140 23700 39196
rect 23700 39140 23704 39196
rect 23640 39136 23704 39140
rect 23720 39196 23784 39200
rect 23720 39140 23724 39196
rect 23724 39140 23780 39196
rect 23780 39140 23784 39196
rect 23720 39136 23784 39140
rect 12756 38796 12820 38860
rect 6584 38652 6648 38656
rect 6584 38596 6588 38652
rect 6588 38596 6644 38652
rect 6644 38596 6648 38652
rect 6584 38592 6648 38596
rect 6664 38652 6728 38656
rect 6664 38596 6668 38652
rect 6668 38596 6724 38652
rect 6724 38596 6728 38652
rect 6664 38592 6728 38596
rect 6744 38652 6808 38656
rect 6744 38596 6748 38652
rect 6748 38596 6804 38652
rect 6804 38596 6808 38652
rect 6744 38592 6808 38596
rect 6824 38652 6888 38656
rect 6824 38596 6828 38652
rect 6828 38596 6884 38652
rect 6884 38596 6888 38652
rect 6824 38592 6888 38596
rect 12020 38524 12084 38588
rect 17848 38652 17912 38656
rect 17848 38596 17852 38652
rect 17852 38596 17908 38652
rect 17908 38596 17912 38652
rect 17848 38592 17912 38596
rect 17928 38652 17992 38656
rect 17928 38596 17932 38652
rect 17932 38596 17988 38652
rect 17988 38596 17992 38652
rect 17928 38592 17992 38596
rect 18008 38652 18072 38656
rect 18008 38596 18012 38652
rect 18012 38596 18068 38652
rect 18068 38596 18072 38652
rect 18008 38592 18072 38596
rect 18088 38652 18152 38656
rect 18088 38596 18092 38652
rect 18092 38596 18148 38652
rect 18148 38596 18152 38652
rect 18088 38592 18152 38596
rect 29112 38652 29176 38656
rect 29112 38596 29116 38652
rect 29116 38596 29172 38652
rect 29172 38596 29176 38652
rect 29112 38592 29176 38596
rect 29192 38652 29256 38656
rect 29192 38596 29196 38652
rect 29196 38596 29252 38652
rect 29252 38596 29256 38652
rect 29192 38592 29256 38596
rect 29272 38652 29336 38656
rect 29272 38596 29276 38652
rect 29276 38596 29332 38652
rect 29332 38596 29336 38652
rect 29272 38592 29336 38596
rect 29352 38652 29416 38656
rect 29352 38596 29356 38652
rect 29356 38596 29412 38652
rect 29412 38596 29416 38652
rect 29352 38592 29416 38596
rect 12216 38108 12280 38112
rect 12216 38052 12220 38108
rect 12220 38052 12276 38108
rect 12276 38052 12280 38108
rect 12216 38048 12280 38052
rect 12296 38108 12360 38112
rect 12296 38052 12300 38108
rect 12300 38052 12356 38108
rect 12356 38052 12360 38108
rect 12296 38048 12360 38052
rect 12376 38108 12440 38112
rect 12376 38052 12380 38108
rect 12380 38052 12436 38108
rect 12436 38052 12440 38108
rect 12376 38048 12440 38052
rect 12456 38108 12520 38112
rect 12456 38052 12460 38108
rect 12460 38052 12516 38108
rect 12516 38052 12520 38108
rect 12456 38048 12520 38052
rect 23480 38108 23544 38112
rect 23480 38052 23484 38108
rect 23484 38052 23540 38108
rect 23540 38052 23544 38108
rect 23480 38048 23544 38052
rect 23560 38108 23624 38112
rect 23560 38052 23564 38108
rect 23564 38052 23620 38108
rect 23620 38052 23624 38108
rect 23560 38048 23624 38052
rect 23640 38108 23704 38112
rect 23640 38052 23644 38108
rect 23644 38052 23700 38108
rect 23700 38052 23704 38108
rect 23640 38048 23704 38052
rect 23720 38108 23784 38112
rect 23720 38052 23724 38108
rect 23724 38052 23780 38108
rect 23780 38052 23784 38108
rect 23720 38048 23784 38052
rect 6584 37564 6648 37568
rect 6584 37508 6588 37564
rect 6588 37508 6644 37564
rect 6644 37508 6648 37564
rect 6584 37504 6648 37508
rect 6664 37564 6728 37568
rect 6664 37508 6668 37564
rect 6668 37508 6724 37564
rect 6724 37508 6728 37564
rect 6664 37504 6728 37508
rect 6744 37564 6808 37568
rect 6744 37508 6748 37564
rect 6748 37508 6804 37564
rect 6804 37508 6808 37564
rect 6744 37504 6808 37508
rect 6824 37564 6888 37568
rect 6824 37508 6828 37564
rect 6828 37508 6884 37564
rect 6884 37508 6888 37564
rect 6824 37504 6888 37508
rect 17848 37564 17912 37568
rect 17848 37508 17852 37564
rect 17852 37508 17908 37564
rect 17908 37508 17912 37564
rect 17848 37504 17912 37508
rect 17928 37564 17992 37568
rect 17928 37508 17932 37564
rect 17932 37508 17988 37564
rect 17988 37508 17992 37564
rect 17928 37504 17992 37508
rect 18008 37564 18072 37568
rect 18008 37508 18012 37564
rect 18012 37508 18068 37564
rect 18068 37508 18072 37564
rect 18008 37504 18072 37508
rect 18088 37564 18152 37568
rect 18088 37508 18092 37564
rect 18092 37508 18148 37564
rect 18148 37508 18152 37564
rect 18088 37504 18152 37508
rect 29112 37564 29176 37568
rect 29112 37508 29116 37564
rect 29116 37508 29172 37564
rect 29172 37508 29176 37564
rect 29112 37504 29176 37508
rect 29192 37564 29256 37568
rect 29192 37508 29196 37564
rect 29196 37508 29252 37564
rect 29252 37508 29256 37564
rect 29192 37504 29256 37508
rect 29272 37564 29336 37568
rect 29272 37508 29276 37564
rect 29276 37508 29332 37564
rect 29332 37508 29336 37564
rect 29272 37504 29336 37508
rect 29352 37564 29416 37568
rect 29352 37508 29356 37564
rect 29356 37508 29412 37564
rect 29412 37508 29416 37564
rect 29352 37504 29416 37508
rect 17540 37496 17604 37500
rect 17540 37440 17590 37496
rect 17590 37440 17604 37496
rect 17540 37436 17604 37440
rect 12216 37020 12280 37024
rect 12216 36964 12220 37020
rect 12220 36964 12276 37020
rect 12276 36964 12280 37020
rect 12216 36960 12280 36964
rect 12296 37020 12360 37024
rect 12296 36964 12300 37020
rect 12300 36964 12356 37020
rect 12356 36964 12360 37020
rect 12296 36960 12360 36964
rect 12376 37020 12440 37024
rect 12376 36964 12380 37020
rect 12380 36964 12436 37020
rect 12436 36964 12440 37020
rect 12376 36960 12440 36964
rect 12456 37020 12520 37024
rect 12456 36964 12460 37020
rect 12460 36964 12516 37020
rect 12516 36964 12520 37020
rect 12456 36960 12520 36964
rect 23480 37020 23544 37024
rect 23480 36964 23484 37020
rect 23484 36964 23540 37020
rect 23540 36964 23544 37020
rect 23480 36960 23544 36964
rect 23560 37020 23624 37024
rect 23560 36964 23564 37020
rect 23564 36964 23620 37020
rect 23620 36964 23624 37020
rect 23560 36960 23624 36964
rect 23640 37020 23704 37024
rect 23640 36964 23644 37020
rect 23644 36964 23700 37020
rect 23700 36964 23704 37020
rect 23640 36960 23704 36964
rect 23720 37020 23784 37024
rect 23720 36964 23724 37020
rect 23724 36964 23780 37020
rect 23780 36964 23784 37020
rect 23720 36960 23784 36964
rect 6584 36476 6648 36480
rect 6584 36420 6588 36476
rect 6588 36420 6644 36476
rect 6644 36420 6648 36476
rect 6584 36416 6648 36420
rect 6664 36476 6728 36480
rect 6664 36420 6668 36476
rect 6668 36420 6724 36476
rect 6724 36420 6728 36476
rect 6664 36416 6728 36420
rect 6744 36476 6808 36480
rect 6744 36420 6748 36476
rect 6748 36420 6804 36476
rect 6804 36420 6808 36476
rect 6744 36416 6808 36420
rect 6824 36476 6888 36480
rect 6824 36420 6828 36476
rect 6828 36420 6884 36476
rect 6884 36420 6888 36476
rect 6824 36416 6888 36420
rect 17848 36476 17912 36480
rect 17848 36420 17852 36476
rect 17852 36420 17908 36476
rect 17908 36420 17912 36476
rect 17848 36416 17912 36420
rect 17928 36476 17992 36480
rect 17928 36420 17932 36476
rect 17932 36420 17988 36476
rect 17988 36420 17992 36476
rect 17928 36416 17992 36420
rect 18008 36476 18072 36480
rect 18008 36420 18012 36476
rect 18012 36420 18068 36476
rect 18068 36420 18072 36476
rect 18008 36416 18072 36420
rect 18088 36476 18152 36480
rect 18088 36420 18092 36476
rect 18092 36420 18148 36476
rect 18148 36420 18152 36476
rect 18088 36416 18152 36420
rect 29112 36476 29176 36480
rect 29112 36420 29116 36476
rect 29116 36420 29172 36476
rect 29172 36420 29176 36476
rect 29112 36416 29176 36420
rect 29192 36476 29256 36480
rect 29192 36420 29196 36476
rect 29196 36420 29252 36476
rect 29252 36420 29256 36476
rect 29192 36416 29256 36420
rect 29272 36476 29336 36480
rect 29272 36420 29276 36476
rect 29276 36420 29332 36476
rect 29332 36420 29336 36476
rect 29272 36416 29336 36420
rect 29352 36476 29416 36480
rect 29352 36420 29356 36476
rect 29356 36420 29412 36476
rect 29412 36420 29416 36476
rect 29352 36416 29416 36420
rect 12216 35932 12280 35936
rect 12216 35876 12220 35932
rect 12220 35876 12276 35932
rect 12276 35876 12280 35932
rect 12216 35872 12280 35876
rect 12296 35932 12360 35936
rect 12296 35876 12300 35932
rect 12300 35876 12356 35932
rect 12356 35876 12360 35932
rect 12296 35872 12360 35876
rect 12376 35932 12440 35936
rect 12376 35876 12380 35932
rect 12380 35876 12436 35932
rect 12436 35876 12440 35932
rect 12376 35872 12440 35876
rect 12456 35932 12520 35936
rect 12456 35876 12460 35932
rect 12460 35876 12516 35932
rect 12516 35876 12520 35932
rect 12456 35872 12520 35876
rect 23480 35932 23544 35936
rect 23480 35876 23484 35932
rect 23484 35876 23540 35932
rect 23540 35876 23544 35932
rect 23480 35872 23544 35876
rect 23560 35932 23624 35936
rect 23560 35876 23564 35932
rect 23564 35876 23620 35932
rect 23620 35876 23624 35932
rect 23560 35872 23624 35876
rect 23640 35932 23704 35936
rect 23640 35876 23644 35932
rect 23644 35876 23700 35932
rect 23700 35876 23704 35932
rect 23640 35872 23704 35876
rect 23720 35932 23784 35936
rect 23720 35876 23724 35932
rect 23724 35876 23780 35932
rect 23780 35876 23784 35932
rect 23720 35872 23784 35876
rect 17356 35532 17420 35596
rect 6584 35388 6648 35392
rect 6584 35332 6588 35388
rect 6588 35332 6644 35388
rect 6644 35332 6648 35388
rect 6584 35328 6648 35332
rect 6664 35388 6728 35392
rect 6664 35332 6668 35388
rect 6668 35332 6724 35388
rect 6724 35332 6728 35388
rect 6664 35328 6728 35332
rect 6744 35388 6808 35392
rect 6744 35332 6748 35388
rect 6748 35332 6804 35388
rect 6804 35332 6808 35388
rect 6744 35328 6808 35332
rect 6824 35388 6888 35392
rect 6824 35332 6828 35388
rect 6828 35332 6884 35388
rect 6884 35332 6888 35388
rect 6824 35328 6888 35332
rect 17848 35388 17912 35392
rect 17848 35332 17852 35388
rect 17852 35332 17908 35388
rect 17908 35332 17912 35388
rect 17848 35328 17912 35332
rect 17928 35388 17992 35392
rect 17928 35332 17932 35388
rect 17932 35332 17988 35388
rect 17988 35332 17992 35388
rect 17928 35328 17992 35332
rect 18008 35388 18072 35392
rect 18008 35332 18012 35388
rect 18012 35332 18068 35388
rect 18068 35332 18072 35388
rect 18008 35328 18072 35332
rect 18088 35388 18152 35392
rect 18088 35332 18092 35388
rect 18092 35332 18148 35388
rect 18148 35332 18152 35388
rect 18088 35328 18152 35332
rect 29112 35388 29176 35392
rect 29112 35332 29116 35388
rect 29116 35332 29172 35388
rect 29172 35332 29176 35388
rect 29112 35328 29176 35332
rect 29192 35388 29256 35392
rect 29192 35332 29196 35388
rect 29196 35332 29252 35388
rect 29252 35332 29256 35388
rect 29192 35328 29256 35332
rect 29272 35388 29336 35392
rect 29272 35332 29276 35388
rect 29276 35332 29332 35388
rect 29332 35332 29336 35388
rect 29272 35328 29336 35332
rect 29352 35388 29416 35392
rect 29352 35332 29356 35388
rect 29356 35332 29412 35388
rect 29412 35332 29416 35388
rect 29352 35328 29416 35332
rect 17356 35260 17420 35324
rect 31524 35184 31588 35188
rect 31524 35128 31574 35184
rect 31574 35128 31588 35184
rect 31524 35124 31588 35128
rect 14228 34988 14292 35052
rect 15332 34988 15396 35052
rect 12216 34844 12280 34848
rect 12216 34788 12220 34844
rect 12220 34788 12276 34844
rect 12276 34788 12280 34844
rect 12216 34784 12280 34788
rect 12296 34844 12360 34848
rect 12296 34788 12300 34844
rect 12300 34788 12356 34844
rect 12356 34788 12360 34844
rect 12296 34784 12360 34788
rect 12376 34844 12440 34848
rect 12376 34788 12380 34844
rect 12380 34788 12436 34844
rect 12436 34788 12440 34844
rect 12376 34784 12440 34788
rect 12456 34844 12520 34848
rect 12456 34788 12460 34844
rect 12460 34788 12516 34844
rect 12516 34788 12520 34844
rect 12456 34784 12520 34788
rect 23480 34844 23544 34848
rect 23480 34788 23484 34844
rect 23484 34788 23540 34844
rect 23540 34788 23544 34844
rect 23480 34784 23544 34788
rect 23560 34844 23624 34848
rect 23560 34788 23564 34844
rect 23564 34788 23620 34844
rect 23620 34788 23624 34844
rect 23560 34784 23624 34788
rect 23640 34844 23704 34848
rect 23640 34788 23644 34844
rect 23644 34788 23700 34844
rect 23700 34788 23704 34844
rect 23640 34784 23704 34788
rect 23720 34844 23784 34848
rect 23720 34788 23724 34844
rect 23724 34788 23780 34844
rect 23780 34788 23784 34844
rect 23720 34784 23784 34788
rect 12756 34776 12820 34780
rect 12756 34720 12770 34776
rect 12770 34720 12820 34776
rect 12756 34716 12820 34720
rect 14596 34580 14660 34644
rect 6584 34300 6648 34304
rect 6584 34244 6588 34300
rect 6588 34244 6644 34300
rect 6644 34244 6648 34300
rect 6584 34240 6648 34244
rect 6664 34300 6728 34304
rect 6664 34244 6668 34300
rect 6668 34244 6724 34300
rect 6724 34244 6728 34300
rect 6664 34240 6728 34244
rect 6744 34300 6808 34304
rect 6744 34244 6748 34300
rect 6748 34244 6804 34300
rect 6804 34244 6808 34300
rect 6744 34240 6808 34244
rect 6824 34300 6888 34304
rect 6824 34244 6828 34300
rect 6828 34244 6884 34300
rect 6884 34244 6888 34300
rect 6824 34240 6888 34244
rect 17848 34300 17912 34304
rect 17848 34244 17852 34300
rect 17852 34244 17908 34300
rect 17908 34244 17912 34300
rect 17848 34240 17912 34244
rect 17928 34300 17992 34304
rect 17928 34244 17932 34300
rect 17932 34244 17988 34300
rect 17988 34244 17992 34300
rect 17928 34240 17992 34244
rect 18008 34300 18072 34304
rect 18008 34244 18012 34300
rect 18012 34244 18068 34300
rect 18068 34244 18072 34300
rect 18008 34240 18072 34244
rect 18088 34300 18152 34304
rect 18088 34244 18092 34300
rect 18092 34244 18148 34300
rect 18148 34244 18152 34300
rect 18088 34240 18152 34244
rect 29112 34300 29176 34304
rect 29112 34244 29116 34300
rect 29116 34244 29172 34300
rect 29172 34244 29176 34300
rect 29112 34240 29176 34244
rect 29192 34300 29256 34304
rect 29192 34244 29196 34300
rect 29196 34244 29252 34300
rect 29252 34244 29256 34300
rect 29192 34240 29256 34244
rect 29272 34300 29336 34304
rect 29272 34244 29276 34300
rect 29276 34244 29332 34300
rect 29332 34244 29336 34300
rect 29272 34240 29336 34244
rect 29352 34300 29416 34304
rect 29352 34244 29356 34300
rect 29356 34244 29412 34300
rect 29412 34244 29416 34300
rect 29352 34240 29416 34244
rect 18460 34172 18524 34236
rect 14228 34036 14292 34100
rect 14596 34096 14660 34100
rect 14596 34040 14610 34096
rect 14610 34040 14660 34096
rect 14596 34036 14660 34040
rect 15884 33900 15948 33964
rect 20852 33764 20916 33828
rect 12216 33756 12280 33760
rect 12216 33700 12220 33756
rect 12220 33700 12276 33756
rect 12276 33700 12280 33756
rect 12216 33696 12280 33700
rect 12296 33756 12360 33760
rect 12296 33700 12300 33756
rect 12300 33700 12356 33756
rect 12356 33700 12360 33756
rect 12296 33696 12360 33700
rect 12376 33756 12440 33760
rect 12376 33700 12380 33756
rect 12380 33700 12436 33756
rect 12436 33700 12440 33756
rect 12376 33696 12440 33700
rect 12456 33756 12520 33760
rect 12456 33700 12460 33756
rect 12460 33700 12516 33756
rect 12516 33700 12520 33756
rect 12456 33696 12520 33700
rect 23480 33756 23544 33760
rect 23480 33700 23484 33756
rect 23484 33700 23540 33756
rect 23540 33700 23544 33756
rect 23480 33696 23544 33700
rect 23560 33756 23624 33760
rect 23560 33700 23564 33756
rect 23564 33700 23620 33756
rect 23620 33700 23624 33756
rect 23560 33696 23624 33700
rect 23640 33756 23704 33760
rect 23640 33700 23644 33756
rect 23644 33700 23700 33756
rect 23700 33700 23704 33756
rect 23640 33696 23704 33700
rect 23720 33756 23784 33760
rect 23720 33700 23724 33756
rect 23724 33700 23780 33756
rect 23780 33700 23784 33756
rect 23720 33696 23784 33700
rect 18460 33628 18524 33692
rect 15884 33492 15948 33556
rect 18276 33356 18340 33420
rect 18460 33356 18524 33420
rect 18276 33220 18340 33284
rect 31524 33416 31588 33420
rect 31524 33360 31574 33416
rect 31574 33360 31588 33416
rect 31524 33356 31588 33360
rect 6584 33212 6648 33216
rect 6584 33156 6588 33212
rect 6588 33156 6644 33212
rect 6644 33156 6648 33212
rect 6584 33152 6648 33156
rect 6664 33212 6728 33216
rect 6664 33156 6668 33212
rect 6668 33156 6724 33212
rect 6724 33156 6728 33212
rect 6664 33152 6728 33156
rect 6744 33212 6808 33216
rect 6744 33156 6748 33212
rect 6748 33156 6804 33212
rect 6804 33156 6808 33212
rect 6744 33152 6808 33156
rect 6824 33212 6888 33216
rect 6824 33156 6828 33212
rect 6828 33156 6884 33212
rect 6884 33156 6888 33212
rect 6824 33152 6888 33156
rect 17848 33212 17912 33216
rect 17848 33156 17852 33212
rect 17852 33156 17908 33212
rect 17908 33156 17912 33212
rect 17848 33152 17912 33156
rect 17928 33212 17992 33216
rect 17928 33156 17932 33212
rect 17932 33156 17988 33212
rect 17988 33156 17992 33212
rect 17928 33152 17992 33156
rect 18008 33212 18072 33216
rect 18008 33156 18012 33212
rect 18012 33156 18068 33212
rect 18068 33156 18072 33212
rect 18008 33152 18072 33156
rect 18088 33212 18152 33216
rect 18088 33156 18092 33212
rect 18092 33156 18148 33212
rect 18148 33156 18152 33212
rect 18088 33152 18152 33156
rect 29112 33212 29176 33216
rect 29112 33156 29116 33212
rect 29116 33156 29172 33212
rect 29172 33156 29176 33212
rect 29112 33152 29176 33156
rect 29192 33212 29256 33216
rect 29192 33156 29196 33212
rect 29196 33156 29252 33212
rect 29252 33156 29256 33212
rect 29192 33152 29256 33156
rect 29272 33212 29336 33216
rect 29272 33156 29276 33212
rect 29276 33156 29332 33212
rect 29332 33156 29336 33212
rect 29272 33152 29336 33156
rect 29352 33212 29416 33216
rect 29352 33156 29356 33212
rect 29356 33156 29412 33212
rect 29412 33156 29416 33212
rect 29352 33152 29416 33156
rect 16068 32948 16132 33012
rect 16436 33084 16500 33148
rect 12216 32668 12280 32672
rect 12216 32612 12220 32668
rect 12220 32612 12276 32668
rect 12276 32612 12280 32668
rect 12216 32608 12280 32612
rect 12296 32668 12360 32672
rect 12296 32612 12300 32668
rect 12300 32612 12356 32668
rect 12356 32612 12360 32668
rect 12296 32608 12360 32612
rect 12376 32668 12440 32672
rect 12376 32612 12380 32668
rect 12380 32612 12436 32668
rect 12436 32612 12440 32668
rect 12376 32608 12440 32612
rect 12456 32668 12520 32672
rect 12456 32612 12460 32668
rect 12460 32612 12516 32668
rect 12516 32612 12520 32668
rect 12456 32608 12520 32612
rect 17540 32676 17604 32740
rect 18276 32676 18340 32740
rect 23480 32668 23544 32672
rect 23480 32612 23484 32668
rect 23484 32612 23540 32668
rect 23540 32612 23544 32668
rect 23480 32608 23544 32612
rect 23560 32668 23624 32672
rect 23560 32612 23564 32668
rect 23564 32612 23620 32668
rect 23620 32612 23624 32668
rect 23560 32608 23624 32612
rect 23640 32668 23704 32672
rect 23640 32612 23644 32668
rect 23644 32612 23700 32668
rect 23700 32612 23704 32668
rect 23640 32608 23704 32612
rect 23720 32668 23784 32672
rect 23720 32612 23724 32668
rect 23724 32612 23780 32668
rect 23780 32612 23784 32668
rect 23720 32608 23784 32612
rect 18460 32404 18524 32468
rect 18644 32404 18708 32468
rect 14780 32132 14844 32196
rect 17356 32132 17420 32196
rect 18276 32192 18340 32196
rect 18276 32136 18290 32192
rect 18290 32136 18340 32192
rect 18276 32132 18340 32136
rect 18460 32132 18524 32196
rect 30420 32192 30484 32196
rect 30420 32136 30470 32192
rect 30470 32136 30484 32192
rect 30420 32132 30484 32136
rect 30788 32192 30852 32196
rect 30788 32136 30838 32192
rect 30838 32136 30852 32192
rect 30788 32132 30852 32136
rect 6584 32124 6648 32128
rect 6584 32068 6588 32124
rect 6588 32068 6644 32124
rect 6644 32068 6648 32124
rect 6584 32064 6648 32068
rect 6664 32124 6728 32128
rect 6664 32068 6668 32124
rect 6668 32068 6724 32124
rect 6724 32068 6728 32124
rect 6664 32064 6728 32068
rect 6744 32124 6808 32128
rect 6744 32068 6748 32124
rect 6748 32068 6804 32124
rect 6804 32068 6808 32124
rect 6744 32064 6808 32068
rect 6824 32124 6888 32128
rect 6824 32068 6828 32124
rect 6828 32068 6884 32124
rect 6884 32068 6888 32124
rect 6824 32064 6888 32068
rect 17848 32124 17912 32128
rect 17848 32068 17852 32124
rect 17852 32068 17908 32124
rect 17908 32068 17912 32124
rect 17848 32064 17912 32068
rect 17928 32124 17992 32128
rect 17928 32068 17932 32124
rect 17932 32068 17988 32124
rect 17988 32068 17992 32124
rect 17928 32064 17992 32068
rect 18008 32124 18072 32128
rect 18008 32068 18012 32124
rect 18012 32068 18068 32124
rect 18068 32068 18072 32124
rect 18008 32064 18072 32068
rect 18088 32124 18152 32128
rect 18088 32068 18092 32124
rect 18092 32068 18148 32124
rect 18148 32068 18152 32124
rect 18088 32064 18152 32068
rect 29112 32124 29176 32128
rect 29112 32068 29116 32124
rect 29116 32068 29172 32124
rect 29172 32068 29176 32124
rect 29112 32064 29176 32068
rect 29192 32124 29256 32128
rect 29192 32068 29196 32124
rect 29196 32068 29252 32124
rect 29252 32068 29256 32124
rect 29192 32064 29256 32068
rect 29272 32124 29336 32128
rect 29272 32068 29276 32124
rect 29276 32068 29332 32124
rect 29332 32068 29336 32124
rect 29272 32064 29336 32068
rect 29352 32124 29416 32128
rect 29352 32068 29356 32124
rect 29356 32068 29412 32124
rect 29412 32068 29416 32124
rect 29352 32064 29416 32068
rect 18828 31996 18892 32060
rect 16252 31724 16316 31788
rect 16436 31724 16500 31788
rect 12216 31580 12280 31584
rect 12216 31524 12220 31580
rect 12220 31524 12276 31580
rect 12276 31524 12280 31580
rect 12216 31520 12280 31524
rect 12296 31580 12360 31584
rect 12296 31524 12300 31580
rect 12300 31524 12356 31580
rect 12356 31524 12360 31580
rect 12296 31520 12360 31524
rect 12376 31580 12440 31584
rect 12376 31524 12380 31580
rect 12380 31524 12436 31580
rect 12436 31524 12440 31580
rect 12376 31520 12440 31524
rect 12456 31580 12520 31584
rect 12456 31524 12460 31580
rect 12460 31524 12516 31580
rect 12516 31524 12520 31580
rect 12456 31520 12520 31524
rect 23480 31580 23544 31584
rect 23480 31524 23484 31580
rect 23484 31524 23540 31580
rect 23540 31524 23544 31580
rect 23480 31520 23544 31524
rect 23560 31580 23624 31584
rect 23560 31524 23564 31580
rect 23564 31524 23620 31580
rect 23620 31524 23624 31580
rect 23560 31520 23624 31524
rect 23640 31580 23704 31584
rect 23640 31524 23644 31580
rect 23644 31524 23700 31580
rect 23700 31524 23704 31580
rect 23640 31520 23704 31524
rect 23720 31580 23784 31584
rect 23720 31524 23724 31580
rect 23724 31524 23780 31580
rect 23780 31524 23784 31580
rect 23720 31520 23784 31524
rect 17540 31044 17604 31108
rect 6584 31036 6648 31040
rect 6584 30980 6588 31036
rect 6588 30980 6644 31036
rect 6644 30980 6648 31036
rect 6584 30976 6648 30980
rect 6664 31036 6728 31040
rect 6664 30980 6668 31036
rect 6668 30980 6724 31036
rect 6724 30980 6728 31036
rect 6664 30976 6728 30980
rect 6744 31036 6808 31040
rect 6744 30980 6748 31036
rect 6748 30980 6804 31036
rect 6804 30980 6808 31036
rect 6744 30976 6808 30980
rect 6824 31036 6888 31040
rect 6824 30980 6828 31036
rect 6828 30980 6884 31036
rect 6884 30980 6888 31036
rect 6824 30976 6888 30980
rect 17848 31036 17912 31040
rect 17848 30980 17852 31036
rect 17852 30980 17908 31036
rect 17908 30980 17912 31036
rect 17848 30976 17912 30980
rect 17928 31036 17992 31040
rect 17928 30980 17932 31036
rect 17932 30980 17988 31036
rect 17988 30980 17992 31036
rect 17928 30976 17992 30980
rect 18008 31036 18072 31040
rect 18008 30980 18012 31036
rect 18012 30980 18068 31036
rect 18068 30980 18072 31036
rect 18008 30976 18072 30980
rect 18088 31036 18152 31040
rect 18088 30980 18092 31036
rect 18092 30980 18148 31036
rect 18148 30980 18152 31036
rect 18088 30976 18152 30980
rect 18460 30908 18524 30972
rect 18644 30908 18708 30972
rect 21772 31044 21836 31108
rect 23060 31044 23124 31108
rect 27660 31044 27724 31108
rect 29112 31036 29176 31040
rect 29112 30980 29116 31036
rect 29116 30980 29172 31036
rect 29172 30980 29176 31036
rect 29112 30976 29176 30980
rect 29192 31036 29256 31040
rect 29192 30980 29196 31036
rect 29196 30980 29252 31036
rect 29252 30980 29256 31036
rect 29192 30976 29256 30980
rect 29272 31036 29336 31040
rect 29272 30980 29276 31036
rect 29276 30980 29332 31036
rect 29332 30980 29336 31036
rect 29272 30976 29336 30980
rect 29352 31036 29416 31040
rect 29352 30980 29356 31036
rect 29356 30980 29412 31036
rect 29412 30980 29416 31036
rect 29352 30976 29416 30980
rect 21220 30772 21284 30836
rect 21220 30636 21284 30700
rect 12216 30492 12280 30496
rect 12216 30436 12220 30492
rect 12220 30436 12276 30492
rect 12276 30436 12280 30492
rect 12216 30432 12280 30436
rect 12296 30492 12360 30496
rect 12296 30436 12300 30492
rect 12300 30436 12356 30492
rect 12356 30436 12360 30492
rect 12296 30432 12360 30436
rect 12376 30492 12440 30496
rect 12376 30436 12380 30492
rect 12380 30436 12436 30492
rect 12436 30436 12440 30492
rect 12376 30432 12440 30436
rect 12456 30492 12520 30496
rect 12456 30436 12460 30492
rect 12460 30436 12516 30492
rect 12516 30436 12520 30492
rect 12456 30432 12520 30436
rect 18828 30364 18892 30428
rect 23060 30500 23124 30564
rect 28580 30636 28644 30700
rect 30420 30500 30484 30564
rect 23480 30492 23544 30496
rect 23480 30436 23484 30492
rect 23484 30436 23540 30492
rect 23540 30436 23544 30492
rect 23480 30432 23544 30436
rect 23560 30492 23624 30496
rect 23560 30436 23564 30492
rect 23564 30436 23620 30492
rect 23620 30436 23624 30492
rect 23560 30432 23624 30436
rect 23640 30492 23704 30496
rect 23640 30436 23644 30492
rect 23644 30436 23700 30492
rect 23700 30436 23704 30492
rect 23640 30432 23704 30436
rect 23720 30492 23784 30496
rect 23720 30436 23724 30492
rect 23724 30436 23780 30492
rect 23780 30436 23784 30492
rect 23720 30432 23784 30436
rect 18460 29956 18524 30020
rect 22692 29956 22756 30020
rect 6584 29948 6648 29952
rect 6584 29892 6588 29948
rect 6588 29892 6644 29948
rect 6644 29892 6648 29948
rect 6584 29888 6648 29892
rect 6664 29948 6728 29952
rect 6664 29892 6668 29948
rect 6668 29892 6724 29948
rect 6724 29892 6728 29948
rect 6664 29888 6728 29892
rect 6744 29948 6808 29952
rect 6744 29892 6748 29948
rect 6748 29892 6804 29948
rect 6804 29892 6808 29948
rect 6744 29888 6808 29892
rect 6824 29948 6888 29952
rect 6824 29892 6828 29948
rect 6828 29892 6884 29948
rect 6884 29892 6888 29948
rect 6824 29888 6888 29892
rect 17848 29948 17912 29952
rect 17848 29892 17852 29948
rect 17852 29892 17908 29948
rect 17908 29892 17912 29948
rect 17848 29888 17912 29892
rect 17928 29948 17992 29952
rect 17928 29892 17932 29948
rect 17932 29892 17988 29948
rect 17988 29892 17992 29948
rect 17928 29888 17992 29892
rect 18008 29948 18072 29952
rect 18008 29892 18012 29948
rect 18012 29892 18068 29948
rect 18068 29892 18072 29948
rect 18008 29888 18072 29892
rect 18088 29948 18152 29952
rect 18088 29892 18092 29948
rect 18092 29892 18148 29948
rect 18148 29892 18152 29948
rect 18088 29888 18152 29892
rect 17540 29820 17604 29884
rect 18276 29880 18340 29884
rect 18276 29824 18290 29880
rect 18290 29824 18340 29880
rect 18276 29820 18340 29824
rect 23244 29820 23308 29884
rect 29112 29948 29176 29952
rect 29112 29892 29116 29948
rect 29116 29892 29172 29948
rect 29172 29892 29176 29948
rect 29112 29888 29176 29892
rect 29192 29948 29256 29952
rect 29192 29892 29196 29948
rect 29196 29892 29252 29948
rect 29252 29892 29256 29948
rect 29192 29888 29256 29892
rect 29272 29948 29336 29952
rect 29272 29892 29276 29948
rect 29276 29892 29332 29948
rect 29332 29892 29336 29948
rect 29272 29888 29336 29892
rect 29352 29948 29416 29952
rect 29352 29892 29356 29948
rect 29356 29892 29412 29948
rect 29412 29892 29416 29948
rect 29352 29888 29416 29892
rect 28580 29880 28644 29884
rect 28580 29824 28594 29880
rect 28594 29824 28644 29880
rect 28580 29820 28644 29824
rect 30788 29880 30852 29884
rect 30788 29824 30838 29880
rect 30838 29824 30852 29880
rect 30788 29820 30852 29824
rect 23244 29412 23308 29476
rect 12216 29404 12280 29408
rect 12216 29348 12220 29404
rect 12220 29348 12276 29404
rect 12276 29348 12280 29404
rect 12216 29344 12280 29348
rect 12296 29404 12360 29408
rect 12296 29348 12300 29404
rect 12300 29348 12356 29404
rect 12356 29348 12360 29404
rect 12296 29344 12360 29348
rect 12376 29404 12440 29408
rect 12376 29348 12380 29404
rect 12380 29348 12436 29404
rect 12436 29348 12440 29404
rect 12376 29344 12440 29348
rect 12456 29404 12520 29408
rect 12456 29348 12460 29404
rect 12460 29348 12516 29404
rect 12516 29348 12520 29404
rect 12456 29344 12520 29348
rect 23480 29404 23544 29408
rect 23480 29348 23484 29404
rect 23484 29348 23540 29404
rect 23540 29348 23544 29404
rect 23480 29344 23544 29348
rect 23560 29404 23624 29408
rect 23560 29348 23564 29404
rect 23564 29348 23620 29404
rect 23620 29348 23624 29404
rect 23560 29344 23624 29348
rect 23640 29404 23704 29408
rect 23640 29348 23644 29404
rect 23644 29348 23700 29404
rect 23700 29348 23704 29404
rect 23640 29344 23704 29348
rect 23720 29404 23784 29408
rect 23720 29348 23724 29404
rect 23724 29348 23780 29404
rect 23780 29348 23784 29404
rect 23720 29344 23784 29348
rect 20852 29064 20916 29068
rect 20852 29008 20902 29064
rect 20902 29008 20916 29064
rect 20852 29004 20916 29008
rect 6584 28860 6648 28864
rect 6584 28804 6588 28860
rect 6588 28804 6644 28860
rect 6644 28804 6648 28860
rect 6584 28800 6648 28804
rect 6664 28860 6728 28864
rect 6664 28804 6668 28860
rect 6668 28804 6724 28860
rect 6724 28804 6728 28860
rect 6664 28800 6728 28804
rect 6744 28860 6808 28864
rect 6744 28804 6748 28860
rect 6748 28804 6804 28860
rect 6804 28804 6808 28860
rect 6744 28800 6808 28804
rect 6824 28860 6888 28864
rect 6824 28804 6828 28860
rect 6828 28804 6884 28860
rect 6884 28804 6888 28860
rect 6824 28800 6888 28804
rect 17848 28860 17912 28864
rect 17848 28804 17852 28860
rect 17852 28804 17908 28860
rect 17908 28804 17912 28860
rect 17848 28800 17912 28804
rect 17928 28860 17992 28864
rect 17928 28804 17932 28860
rect 17932 28804 17988 28860
rect 17988 28804 17992 28860
rect 17928 28800 17992 28804
rect 18008 28860 18072 28864
rect 18008 28804 18012 28860
rect 18012 28804 18068 28860
rect 18068 28804 18072 28860
rect 18008 28800 18072 28804
rect 18088 28860 18152 28864
rect 18088 28804 18092 28860
rect 18092 28804 18148 28860
rect 18148 28804 18152 28860
rect 18088 28800 18152 28804
rect 29868 28868 29932 28932
rect 29112 28860 29176 28864
rect 29112 28804 29116 28860
rect 29116 28804 29172 28860
rect 29172 28804 29176 28860
rect 29112 28800 29176 28804
rect 29192 28860 29256 28864
rect 29192 28804 29196 28860
rect 29196 28804 29252 28860
rect 29252 28804 29256 28860
rect 29192 28800 29256 28804
rect 29272 28860 29336 28864
rect 29272 28804 29276 28860
rect 29276 28804 29332 28860
rect 29332 28804 29336 28860
rect 29272 28800 29336 28804
rect 29352 28860 29416 28864
rect 29352 28804 29356 28860
rect 29356 28804 29412 28860
rect 29412 28804 29416 28860
rect 29352 28800 29416 28804
rect 16804 28596 16868 28660
rect 14228 28384 14292 28388
rect 14228 28328 14278 28384
rect 14278 28328 14292 28384
rect 14228 28324 14292 28328
rect 12216 28316 12280 28320
rect 12216 28260 12220 28316
rect 12220 28260 12276 28316
rect 12276 28260 12280 28316
rect 12216 28256 12280 28260
rect 12296 28316 12360 28320
rect 12296 28260 12300 28316
rect 12300 28260 12356 28316
rect 12356 28260 12360 28316
rect 12296 28256 12360 28260
rect 12376 28316 12440 28320
rect 12376 28260 12380 28316
rect 12380 28260 12436 28316
rect 12436 28260 12440 28316
rect 12376 28256 12440 28260
rect 12456 28316 12520 28320
rect 12456 28260 12460 28316
rect 12460 28260 12516 28316
rect 12516 28260 12520 28316
rect 12456 28256 12520 28260
rect 23480 28316 23544 28320
rect 23480 28260 23484 28316
rect 23484 28260 23540 28316
rect 23540 28260 23544 28316
rect 23480 28256 23544 28260
rect 23560 28316 23624 28320
rect 23560 28260 23564 28316
rect 23564 28260 23620 28316
rect 23620 28260 23624 28316
rect 23560 28256 23624 28260
rect 23640 28316 23704 28320
rect 23640 28260 23644 28316
rect 23644 28260 23700 28316
rect 23700 28260 23704 28316
rect 23640 28256 23704 28260
rect 23720 28316 23784 28320
rect 23720 28260 23724 28316
rect 23724 28260 23780 28316
rect 23780 28260 23784 28316
rect 23720 28256 23784 28260
rect 30052 28188 30116 28252
rect 15332 27916 15396 27980
rect 6584 27772 6648 27776
rect 6584 27716 6588 27772
rect 6588 27716 6644 27772
rect 6644 27716 6648 27772
rect 6584 27712 6648 27716
rect 6664 27772 6728 27776
rect 6664 27716 6668 27772
rect 6668 27716 6724 27772
rect 6724 27716 6728 27772
rect 6664 27712 6728 27716
rect 6744 27772 6808 27776
rect 6744 27716 6748 27772
rect 6748 27716 6804 27772
rect 6804 27716 6808 27772
rect 6744 27712 6808 27716
rect 6824 27772 6888 27776
rect 6824 27716 6828 27772
rect 6828 27716 6884 27772
rect 6884 27716 6888 27772
rect 6824 27712 6888 27716
rect 17848 27772 17912 27776
rect 17848 27716 17852 27772
rect 17852 27716 17908 27772
rect 17908 27716 17912 27772
rect 17848 27712 17912 27716
rect 17928 27772 17992 27776
rect 17928 27716 17932 27772
rect 17932 27716 17988 27772
rect 17988 27716 17992 27772
rect 17928 27712 17992 27716
rect 18008 27772 18072 27776
rect 18008 27716 18012 27772
rect 18012 27716 18068 27772
rect 18068 27716 18072 27772
rect 18008 27712 18072 27716
rect 18088 27772 18152 27776
rect 18088 27716 18092 27772
rect 18092 27716 18148 27772
rect 18148 27716 18152 27772
rect 18088 27712 18152 27716
rect 29112 27772 29176 27776
rect 29112 27716 29116 27772
rect 29116 27716 29172 27772
rect 29172 27716 29176 27772
rect 29112 27712 29176 27716
rect 29192 27772 29256 27776
rect 29192 27716 29196 27772
rect 29196 27716 29252 27772
rect 29252 27716 29256 27772
rect 29192 27712 29256 27716
rect 29272 27772 29336 27776
rect 29272 27716 29276 27772
rect 29276 27716 29332 27772
rect 29332 27716 29336 27772
rect 29272 27712 29336 27716
rect 29352 27772 29416 27776
rect 29352 27716 29356 27772
rect 29356 27716 29412 27772
rect 29412 27716 29416 27772
rect 29352 27712 29416 27716
rect 16068 27508 16132 27572
rect 12216 27228 12280 27232
rect 12216 27172 12220 27228
rect 12220 27172 12276 27228
rect 12276 27172 12280 27228
rect 12216 27168 12280 27172
rect 12296 27228 12360 27232
rect 12296 27172 12300 27228
rect 12300 27172 12356 27228
rect 12356 27172 12360 27228
rect 12296 27168 12360 27172
rect 12376 27228 12440 27232
rect 12376 27172 12380 27228
rect 12380 27172 12436 27228
rect 12436 27172 12440 27228
rect 12376 27168 12440 27172
rect 12456 27228 12520 27232
rect 12456 27172 12460 27228
rect 12460 27172 12516 27228
rect 12516 27172 12520 27228
rect 12456 27168 12520 27172
rect 16620 27236 16684 27300
rect 30420 27236 30484 27300
rect 23480 27228 23544 27232
rect 23480 27172 23484 27228
rect 23484 27172 23540 27228
rect 23540 27172 23544 27228
rect 23480 27168 23544 27172
rect 23560 27228 23624 27232
rect 23560 27172 23564 27228
rect 23564 27172 23620 27228
rect 23620 27172 23624 27228
rect 23560 27168 23624 27172
rect 23640 27228 23704 27232
rect 23640 27172 23644 27228
rect 23644 27172 23700 27228
rect 23700 27172 23704 27228
rect 23640 27168 23704 27172
rect 23720 27228 23784 27232
rect 23720 27172 23724 27228
rect 23724 27172 23780 27228
rect 23780 27172 23784 27228
rect 23720 27168 23784 27172
rect 30788 27160 30852 27164
rect 30788 27104 30838 27160
rect 30838 27104 30852 27160
rect 30788 27100 30852 27104
rect 29500 26888 29564 26892
rect 29500 26832 29550 26888
rect 29550 26832 29564 26888
rect 29500 26828 29564 26832
rect 6584 26684 6648 26688
rect 6584 26628 6588 26684
rect 6588 26628 6644 26684
rect 6644 26628 6648 26684
rect 6584 26624 6648 26628
rect 6664 26684 6728 26688
rect 6664 26628 6668 26684
rect 6668 26628 6724 26684
rect 6724 26628 6728 26684
rect 6664 26624 6728 26628
rect 6744 26684 6808 26688
rect 6744 26628 6748 26684
rect 6748 26628 6804 26684
rect 6804 26628 6808 26684
rect 6744 26624 6808 26628
rect 6824 26684 6888 26688
rect 6824 26628 6828 26684
rect 6828 26628 6884 26684
rect 6884 26628 6888 26684
rect 6824 26624 6888 26628
rect 17848 26684 17912 26688
rect 17848 26628 17852 26684
rect 17852 26628 17908 26684
rect 17908 26628 17912 26684
rect 17848 26624 17912 26628
rect 17928 26684 17992 26688
rect 17928 26628 17932 26684
rect 17932 26628 17988 26684
rect 17988 26628 17992 26684
rect 17928 26624 17992 26628
rect 18008 26684 18072 26688
rect 18008 26628 18012 26684
rect 18012 26628 18068 26684
rect 18068 26628 18072 26684
rect 18008 26624 18072 26628
rect 18088 26684 18152 26688
rect 18088 26628 18092 26684
rect 18092 26628 18148 26684
rect 18148 26628 18152 26684
rect 18088 26624 18152 26628
rect 29112 26684 29176 26688
rect 29112 26628 29116 26684
rect 29116 26628 29172 26684
rect 29172 26628 29176 26684
rect 29112 26624 29176 26628
rect 29192 26684 29256 26688
rect 29192 26628 29196 26684
rect 29196 26628 29252 26684
rect 29252 26628 29256 26684
rect 29192 26624 29256 26628
rect 29272 26684 29336 26688
rect 29272 26628 29276 26684
rect 29276 26628 29332 26684
rect 29332 26628 29336 26684
rect 29272 26624 29336 26628
rect 29352 26684 29416 26688
rect 29352 26628 29356 26684
rect 29356 26628 29412 26684
rect 29412 26628 29416 26684
rect 29352 26624 29416 26628
rect 12216 26140 12280 26144
rect 12216 26084 12220 26140
rect 12220 26084 12276 26140
rect 12276 26084 12280 26140
rect 12216 26080 12280 26084
rect 12296 26140 12360 26144
rect 12296 26084 12300 26140
rect 12300 26084 12356 26140
rect 12356 26084 12360 26140
rect 12296 26080 12360 26084
rect 12376 26140 12440 26144
rect 12376 26084 12380 26140
rect 12380 26084 12436 26140
rect 12436 26084 12440 26140
rect 12376 26080 12440 26084
rect 12456 26140 12520 26144
rect 12456 26084 12460 26140
rect 12460 26084 12516 26140
rect 12516 26084 12520 26140
rect 12456 26080 12520 26084
rect 23480 26140 23544 26144
rect 23480 26084 23484 26140
rect 23484 26084 23540 26140
rect 23540 26084 23544 26140
rect 23480 26080 23544 26084
rect 23560 26140 23624 26144
rect 23560 26084 23564 26140
rect 23564 26084 23620 26140
rect 23620 26084 23624 26140
rect 23560 26080 23624 26084
rect 23640 26140 23704 26144
rect 23640 26084 23644 26140
rect 23644 26084 23700 26140
rect 23700 26084 23704 26140
rect 23640 26080 23704 26084
rect 23720 26140 23784 26144
rect 23720 26084 23724 26140
rect 23724 26084 23780 26140
rect 23780 26084 23784 26140
rect 23720 26080 23784 26084
rect 31708 25876 31772 25940
rect 6584 25596 6648 25600
rect 6584 25540 6588 25596
rect 6588 25540 6644 25596
rect 6644 25540 6648 25596
rect 6584 25536 6648 25540
rect 6664 25596 6728 25600
rect 6664 25540 6668 25596
rect 6668 25540 6724 25596
rect 6724 25540 6728 25596
rect 6664 25536 6728 25540
rect 6744 25596 6808 25600
rect 6744 25540 6748 25596
rect 6748 25540 6804 25596
rect 6804 25540 6808 25596
rect 6744 25536 6808 25540
rect 6824 25596 6888 25600
rect 6824 25540 6828 25596
rect 6828 25540 6884 25596
rect 6884 25540 6888 25596
rect 6824 25536 6888 25540
rect 17848 25596 17912 25600
rect 17848 25540 17852 25596
rect 17852 25540 17908 25596
rect 17908 25540 17912 25596
rect 17848 25536 17912 25540
rect 17928 25596 17992 25600
rect 17928 25540 17932 25596
rect 17932 25540 17988 25596
rect 17988 25540 17992 25596
rect 17928 25536 17992 25540
rect 18008 25596 18072 25600
rect 18008 25540 18012 25596
rect 18012 25540 18068 25596
rect 18068 25540 18072 25596
rect 18008 25536 18072 25540
rect 18088 25596 18152 25600
rect 18088 25540 18092 25596
rect 18092 25540 18148 25596
rect 18148 25540 18152 25596
rect 18088 25536 18152 25540
rect 29112 25596 29176 25600
rect 29112 25540 29116 25596
rect 29116 25540 29172 25596
rect 29172 25540 29176 25596
rect 29112 25536 29176 25540
rect 29192 25596 29256 25600
rect 29192 25540 29196 25596
rect 29196 25540 29252 25596
rect 29252 25540 29256 25596
rect 29192 25536 29256 25540
rect 29272 25596 29336 25600
rect 29272 25540 29276 25596
rect 29276 25540 29332 25596
rect 29332 25540 29336 25596
rect 29272 25536 29336 25540
rect 29352 25596 29416 25600
rect 29352 25540 29356 25596
rect 29356 25540 29412 25596
rect 29412 25540 29416 25596
rect 29352 25536 29416 25540
rect 12216 25052 12280 25056
rect 12216 24996 12220 25052
rect 12220 24996 12276 25052
rect 12276 24996 12280 25052
rect 12216 24992 12280 24996
rect 12296 25052 12360 25056
rect 12296 24996 12300 25052
rect 12300 24996 12356 25052
rect 12356 24996 12360 25052
rect 12296 24992 12360 24996
rect 12376 25052 12440 25056
rect 12376 24996 12380 25052
rect 12380 24996 12436 25052
rect 12436 24996 12440 25052
rect 12376 24992 12440 24996
rect 12456 25052 12520 25056
rect 12456 24996 12460 25052
rect 12460 24996 12516 25052
rect 12516 24996 12520 25052
rect 12456 24992 12520 24996
rect 23480 25052 23544 25056
rect 23480 24996 23484 25052
rect 23484 24996 23540 25052
rect 23540 24996 23544 25052
rect 23480 24992 23544 24996
rect 23560 25052 23624 25056
rect 23560 24996 23564 25052
rect 23564 24996 23620 25052
rect 23620 24996 23624 25052
rect 23560 24992 23624 24996
rect 23640 25052 23704 25056
rect 23640 24996 23644 25052
rect 23644 24996 23700 25052
rect 23700 24996 23704 25052
rect 23640 24992 23704 24996
rect 23720 25052 23784 25056
rect 23720 24996 23724 25052
rect 23724 24996 23780 25052
rect 23780 24996 23784 25052
rect 23720 24992 23784 24996
rect 27660 24788 27724 24852
rect 29684 24576 29748 24580
rect 29684 24520 29734 24576
rect 29734 24520 29748 24576
rect 29684 24516 29748 24520
rect 6584 24508 6648 24512
rect 6584 24452 6588 24508
rect 6588 24452 6644 24508
rect 6644 24452 6648 24508
rect 6584 24448 6648 24452
rect 6664 24508 6728 24512
rect 6664 24452 6668 24508
rect 6668 24452 6724 24508
rect 6724 24452 6728 24508
rect 6664 24448 6728 24452
rect 6744 24508 6808 24512
rect 6744 24452 6748 24508
rect 6748 24452 6804 24508
rect 6804 24452 6808 24508
rect 6744 24448 6808 24452
rect 6824 24508 6888 24512
rect 6824 24452 6828 24508
rect 6828 24452 6884 24508
rect 6884 24452 6888 24508
rect 6824 24448 6888 24452
rect 17848 24508 17912 24512
rect 17848 24452 17852 24508
rect 17852 24452 17908 24508
rect 17908 24452 17912 24508
rect 17848 24448 17912 24452
rect 17928 24508 17992 24512
rect 17928 24452 17932 24508
rect 17932 24452 17988 24508
rect 17988 24452 17992 24508
rect 17928 24448 17992 24452
rect 18008 24508 18072 24512
rect 18008 24452 18012 24508
rect 18012 24452 18068 24508
rect 18068 24452 18072 24508
rect 18008 24448 18072 24452
rect 18088 24508 18152 24512
rect 18088 24452 18092 24508
rect 18092 24452 18148 24508
rect 18148 24452 18152 24508
rect 18088 24448 18152 24452
rect 29112 24508 29176 24512
rect 29112 24452 29116 24508
rect 29116 24452 29172 24508
rect 29172 24452 29176 24508
rect 29112 24448 29176 24452
rect 29192 24508 29256 24512
rect 29192 24452 29196 24508
rect 29196 24452 29252 24508
rect 29252 24452 29256 24508
rect 29192 24448 29256 24452
rect 29272 24508 29336 24512
rect 29272 24452 29276 24508
rect 29276 24452 29332 24508
rect 29332 24452 29336 24508
rect 29272 24448 29336 24452
rect 29352 24508 29416 24512
rect 29352 24452 29356 24508
rect 29356 24452 29412 24508
rect 29412 24452 29416 24508
rect 29352 24448 29416 24452
rect 12216 23964 12280 23968
rect 12216 23908 12220 23964
rect 12220 23908 12276 23964
rect 12276 23908 12280 23964
rect 12216 23904 12280 23908
rect 12296 23964 12360 23968
rect 12296 23908 12300 23964
rect 12300 23908 12356 23964
rect 12356 23908 12360 23964
rect 12296 23904 12360 23908
rect 12376 23964 12440 23968
rect 12376 23908 12380 23964
rect 12380 23908 12436 23964
rect 12436 23908 12440 23964
rect 12376 23904 12440 23908
rect 12456 23964 12520 23968
rect 12456 23908 12460 23964
rect 12460 23908 12516 23964
rect 12516 23908 12520 23964
rect 12456 23904 12520 23908
rect 23480 23964 23544 23968
rect 23480 23908 23484 23964
rect 23484 23908 23540 23964
rect 23540 23908 23544 23964
rect 23480 23904 23544 23908
rect 23560 23964 23624 23968
rect 23560 23908 23564 23964
rect 23564 23908 23620 23964
rect 23620 23908 23624 23964
rect 23560 23904 23624 23908
rect 23640 23964 23704 23968
rect 23640 23908 23644 23964
rect 23644 23908 23700 23964
rect 23700 23908 23704 23964
rect 23640 23904 23704 23908
rect 23720 23964 23784 23968
rect 23720 23908 23724 23964
rect 23724 23908 23780 23964
rect 23780 23908 23784 23964
rect 23720 23904 23784 23908
rect 32628 23836 32692 23900
rect 6584 23420 6648 23424
rect 6584 23364 6588 23420
rect 6588 23364 6644 23420
rect 6644 23364 6648 23420
rect 6584 23360 6648 23364
rect 6664 23420 6728 23424
rect 6664 23364 6668 23420
rect 6668 23364 6724 23420
rect 6724 23364 6728 23420
rect 6664 23360 6728 23364
rect 6744 23420 6808 23424
rect 6744 23364 6748 23420
rect 6748 23364 6804 23420
rect 6804 23364 6808 23420
rect 6744 23360 6808 23364
rect 6824 23420 6888 23424
rect 6824 23364 6828 23420
rect 6828 23364 6884 23420
rect 6884 23364 6888 23420
rect 6824 23360 6888 23364
rect 17848 23420 17912 23424
rect 17848 23364 17852 23420
rect 17852 23364 17908 23420
rect 17908 23364 17912 23420
rect 17848 23360 17912 23364
rect 17928 23420 17992 23424
rect 17928 23364 17932 23420
rect 17932 23364 17988 23420
rect 17988 23364 17992 23420
rect 17928 23360 17992 23364
rect 18008 23420 18072 23424
rect 18008 23364 18012 23420
rect 18012 23364 18068 23420
rect 18068 23364 18072 23420
rect 18008 23360 18072 23364
rect 18088 23420 18152 23424
rect 18088 23364 18092 23420
rect 18092 23364 18148 23420
rect 18148 23364 18152 23420
rect 18088 23360 18152 23364
rect 29112 23420 29176 23424
rect 29112 23364 29116 23420
rect 29116 23364 29172 23420
rect 29172 23364 29176 23420
rect 29112 23360 29176 23364
rect 29192 23420 29256 23424
rect 29192 23364 29196 23420
rect 29196 23364 29252 23420
rect 29252 23364 29256 23420
rect 29192 23360 29256 23364
rect 29272 23420 29336 23424
rect 29272 23364 29276 23420
rect 29276 23364 29332 23420
rect 29332 23364 29336 23420
rect 29272 23360 29336 23364
rect 29352 23420 29416 23424
rect 29352 23364 29356 23420
rect 29356 23364 29412 23420
rect 29412 23364 29416 23420
rect 29352 23360 29416 23364
rect 32812 22884 32876 22948
rect 12216 22876 12280 22880
rect 12216 22820 12220 22876
rect 12220 22820 12276 22876
rect 12276 22820 12280 22876
rect 12216 22816 12280 22820
rect 12296 22876 12360 22880
rect 12296 22820 12300 22876
rect 12300 22820 12356 22876
rect 12356 22820 12360 22876
rect 12296 22816 12360 22820
rect 12376 22876 12440 22880
rect 12376 22820 12380 22876
rect 12380 22820 12436 22876
rect 12436 22820 12440 22876
rect 12376 22816 12440 22820
rect 12456 22876 12520 22880
rect 12456 22820 12460 22876
rect 12460 22820 12516 22876
rect 12516 22820 12520 22876
rect 12456 22816 12520 22820
rect 23480 22876 23544 22880
rect 23480 22820 23484 22876
rect 23484 22820 23540 22876
rect 23540 22820 23544 22876
rect 23480 22816 23544 22820
rect 23560 22876 23624 22880
rect 23560 22820 23564 22876
rect 23564 22820 23620 22876
rect 23620 22820 23624 22876
rect 23560 22816 23624 22820
rect 23640 22876 23704 22880
rect 23640 22820 23644 22876
rect 23644 22820 23700 22876
rect 23700 22820 23704 22876
rect 23640 22816 23704 22820
rect 23720 22876 23784 22880
rect 23720 22820 23724 22876
rect 23724 22820 23780 22876
rect 23780 22820 23784 22876
rect 23720 22816 23784 22820
rect 29868 22748 29932 22812
rect 30788 22612 30852 22676
rect 30236 22340 30300 22404
rect 31892 22536 31956 22540
rect 31892 22480 31906 22536
rect 31906 22480 31956 22536
rect 31892 22476 31956 22480
rect 31708 22400 31772 22404
rect 31708 22344 31758 22400
rect 31758 22344 31772 22400
rect 31708 22340 31772 22344
rect 6584 22332 6648 22336
rect 6584 22276 6588 22332
rect 6588 22276 6644 22332
rect 6644 22276 6648 22332
rect 6584 22272 6648 22276
rect 6664 22332 6728 22336
rect 6664 22276 6668 22332
rect 6668 22276 6724 22332
rect 6724 22276 6728 22332
rect 6664 22272 6728 22276
rect 6744 22332 6808 22336
rect 6744 22276 6748 22332
rect 6748 22276 6804 22332
rect 6804 22276 6808 22332
rect 6744 22272 6808 22276
rect 6824 22332 6888 22336
rect 6824 22276 6828 22332
rect 6828 22276 6884 22332
rect 6884 22276 6888 22332
rect 6824 22272 6888 22276
rect 17848 22332 17912 22336
rect 17848 22276 17852 22332
rect 17852 22276 17908 22332
rect 17908 22276 17912 22332
rect 17848 22272 17912 22276
rect 17928 22332 17992 22336
rect 17928 22276 17932 22332
rect 17932 22276 17988 22332
rect 17988 22276 17992 22332
rect 17928 22272 17992 22276
rect 18008 22332 18072 22336
rect 18008 22276 18012 22332
rect 18012 22276 18068 22332
rect 18068 22276 18072 22332
rect 18008 22272 18072 22276
rect 18088 22332 18152 22336
rect 18088 22276 18092 22332
rect 18092 22276 18148 22332
rect 18148 22276 18152 22332
rect 18088 22272 18152 22276
rect 29112 22332 29176 22336
rect 29112 22276 29116 22332
rect 29116 22276 29172 22332
rect 29172 22276 29176 22332
rect 29112 22272 29176 22276
rect 29192 22332 29256 22336
rect 29192 22276 29196 22332
rect 29196 22276 29252 22332
rect 29252 22276 29256 22332
rect 29192 22272 29256 22276
rect 29272 22332 29336 22336
rect 29272 22276 29276 22332
rect 29276 22276 29332 22332
rect 29332 22276 29336 22332
rect 29272 22272 29336 22276
rect 29352 22332 29416 22336
rect 29352 22276 29356 22332
rect 29356 22276 29412 22332
rect 29412 22276 29416 22332
rect 29352 22272 29416 22276
rect 25268 22068 25332 22132
rect 32628 22068 32692 22132
rect 30236 21992 30300 21996
rect 30236 21936 30286 21992
rect 30286 21936 30300 21992
rect 30236 21932 30300 21936
rect 32812 21796 32876 21860
rect 12216 21788 12280 21792
rect 12216 21732 12220 21788
rect 12220 21732 12276 21788
rect 12276 21732 12280 21788
rect 12216 21728 12280 21732
rect 12296 21788 12360 21792
rect 12296 21732 12300 21788
rect 12300 21732 12356 21788
rect 12356 21732 12360 21788
rect 12296 21728 12360 21732
rect 12376 21788 12440 21792
rect 12376 21732 12380 21788
rect 12380 21732 12436 21788
rect 12436 21732 12440 21788
rect 12376 21728 12440 21732
rect 12456 21788 12520 21792
rect 12456 21732 12460 21788
rect 12460 21732 12516 21788
rect 12516 21732 12520 21788
rect 12456 21728 12520 21732
rect 23480 21788 23544 21792
rect 23480 21732 23484 21788
rect 23484 21732 23540 21788
rect 23540 21732 23544 21788
rect 23480 21728 23544 21732
rect 23560 21788 23624 21792
rect 23560 21732 23564 21788
rect 23564 21732 23620 21788
rect 23620 21732 23624 21788
rect 23560 21728 23624 21732
rect 23640 21788 23704 21792
rect 23640 21732 23644 21788
rect 23644 21732 23700 21788
rect 23700 21732 23704 21788
rect 23640 21728 23704 21732
rect 23720 21788 23784 21792
rect 23720 21732 23724 21788
rect 23724 21732 23780 21788
rect 23780 21732 23784 21788
rect 23720 21728 23784 21732
rect 30420 21312 30484 21316
rect 30420 21256 30470 21312
rect 30470 21256 30484 21312
rect 30420 21252 30484 21256
rect 6584 21244 6648 21248
rect 6584 21188 6588 21244
rect 6588 21188 6644 21244
rect 6644 21188 6648 21244
rect 6584 21184 6648 21188
rect 6664 21244 6728 21248
rect 6664 21188 6668 21244
rect 6668 21188 6724 21244
rect 6724 21188 6728 21244
rect 6664 21184 6728 21188
rect 6744 21244 6808 21248
rect 6744 21188 6748 21244
rect 6748 21188 6804 21244
rect 6804 21188 6808 21244
rect 6744 21184 6808 21188
rect 6824 21244 6888 21248
rect 6824 21188 6828 21244
rect 6828 21188 6884 21244
rect 6884 21188 6888 21244
rect 6824 21184 6888 21188
rect 17848 21244 17912 21248
rect 17848 21188 17852 21244
rect 17852 21188 17908 21244
rect 17908 21188 17912 21244
rect 17848 21184 17912 21188
rect 17928 21244 17992 21248
rect 17928 21188 17932 21244
rect 17932 21188 17988 21244
rect 17988 21188 17992 21244
rect 17928 21184 17992 21188
rect 18008 21244 18072 21248
rect 18008 21188 18012 21244
rect 18012 21188 18068 21244
rect 18068 21188 18072 21244
rect 18008 21184 18072 21188
rect 18088 21244 18152 21248
rect 18088 21188 18092 21244
rect 18092 21188 18148 21244
rect 18148 21188 18152 21244
rect 18088 21184 18152 21188
rect 29112 21244 29176 21248
rect 29112 21188 29116 21244
rect 29116 21188 29172 21244
rect 29172 21188 29176 21244
rect 29112 21184 29176 21188
rect 29192 21244 29256 21248
rect 29192 21188 29196 21244
rect 29196 21188 29252 21244
rect 29252 21188 29256 21244
rect 29192 21184 29256 21188
rect 29272 21244 29336 21248
rect 29272 21188 29276 21244
rect 29276 21188 29332 21244
rect 29332 21188 29336 21244
rect 29272 21184 29336 21188
rect 29352 21244 29416 21248
rect 29352 21188 29356 21244
rect 29356 21188 29412 21244
rect 29412 21188 29416 21244
rect 29352 21184 29416 21188
rect 25268 21176 25332 21180
rect 25268 21120 25318 21176
rect 25318 21120 25332 21176
rect 25268 21116 25332 21120
rect 12216 20700 12280 20704
rect 12216 20644 12220 20700
rect 12220 20644 12276 20700
rect 12276 20644 12280 20700
rect 12216 20640 12280 20644
rect 12296 20700 12360 20704
rect 12296 20644 12300 20700
rect 12300 20644 12356 20700
rect 12356 20644 12360 20700
rect 12296 20640 12360 20644
rect 12376 20700 12440 20704
rect 12376 20644 12380 20700
rect 12380 20644 12436 20700
rect 12436 20644 12440 20700
rect 12376 20640 12440 20644
rect 12456 20700 12520 20704
rect 12456 20644 12460 20700
rect 12460 20644 12516 20700
rect 12516 20644 12520 20700
rect 12456 20640 12520 20644
rect 23480 20700 23544 20704
rect 23480 20644 23484 20700
rect 23484 20644 23540 20700
rect 23540 20644 23544 20700
rect 23480 20640 23544 20644
rect 23560 20700 23624 20704
rect 23560 20644 23564 20700
rect 23564 20644 23620 20700
rect 23620 20644 23624 20700
rect 23560 20640 23624 20644
rect 23640 20700 23704 20704
rect 23640 20644 23644 20700
rect 23644 20644 23700 20700
rect 23700 20644 23704 20700
rect 23640 20640 23704 20644
rect 23720 20700 23784 20704
rect 23720 20644 23724 20700
rect 23724 20644 23780 20700
rect 23780 20644 23784 20700
rect 23720 20640 23784 20644
rect 31892 20496 31956 20500
rect 31892 20440 31906 20496
rect 31906 20440 31956 20496
rect 31892 20436 31956 20440
rect 6584 20156 6648 20160
rect 6584 20100 6588 20156
rect 6588 20100 6644 20156
rect 6644 20100 6648 20156
rect 6584 20096 6648 20100
rect 6664 20156 6728 20160
rect 6664 20100 6668 20156
rect 6668 20100 6724 20156
rect 6724 20100 6728 20156
rect 6664 20096 6728 20100
rect 6744 20156 6808 20160
rect 6744 20100 6748 20156
rect 6748 20100 6804 20156
rect 6804 20100 6808 20156
rect 6744 20096 6808 20100
rect 6824 20156 6888 20160
rect 6824 20100 6828 20156
rect 6828 20100 6884 20156
rect 6884 20100 6888 20156
rect 6824 20096 6888 20100
rect 17848 20156 17912 20160
rect 17848 20100 17852 20156
rect 17852 20100 17908 20156
rect 17908 20100 17912 20156
rect 17848 20096 17912 20100
rect 17928 20156 17992 20160
rect 17928 20100 17932 20156
rect 17932 20100 17988 20156
rect 17988 20100 17992 20156
rect 17928 20096 17992 20100
rect 18008 20156 18072 20160
rect 18008 20100 18012 20156
rect 18012 20100 18068 20156
rect 18068 20100 18072 20156
rect 18008 20096 18072 20100
rect 18088 20156 18152 20160
rect 18088 20100 18092 20156
rect 18092 20100 18148 20156
rect 18148 20100 18152 20156
rect 18088 20096 18152 20100
rect 29112 20156 29176 20160
rect 29112 20100 29116 20156
rect 29116 20100 29172 20156
rect 29172 20100 29176 20156
rect 29112 20096 29176 20100
rect 29192 20156 29256 20160
rect 29192 20100 29196 20156
rect 29196 20100 29252 20156
rect 29252 20100 29256 20156
rect 29192 20096 29256 20100
rect 29272 20156 29336 20160
rect 29272 20100 29276 20156
rect 29276 20100 29332 20156
rect 29332 20100 29336 20156
rect 29272 20096 29336 20100
rect 29352 20156 29416 20160
rect 29352 20100 29356 20156
rect 29356 20100 29412 20156
rect 29412 20100 29416 20156
rect 29352 20096 29416 20100
rect 29684 19620 29748 19684
rect 12216 19612 12280 19616
rect 12216 19556 12220 19612
rect 12220 19556 12276 19612
rect 12276 19556 12280 19612
rect 12216 19552 12280 19556
rect 12296 19612 12360 19616
rect 12296 19556 12300 19612
rect 12300 19556 12356 19612
rect 12356 19556 12360 19612
rect 12296 19552 12360 19556
rect 12376 19612 12440 19616
rect 12376 19556 12380 19612
rect 12380 19556 12436 19612
rect 12436 19556 12440 19612
rect 12376 19552 12440 19556
rect 12456 19612 12520 19616
rect 12456 19556 12460 19612
rect 12460 19556 12516 19612
rect 12516 19556 12520 19612
rect 12456 19552 12520 19556
rect 23480 19612 23544 19616
rect 23480 19556 23484 19612
rect 23484 19556 23540 19612
rect 23540 19556 23544 19612
rect 23480 19552 23544 19556
rect 23560 19612 23624 19616
rect 23560 19556 23564 19612
rect 23564 19556 23620 19612
rect 23620 19556 23624 19612
rect 23560 19552 23624 19556
rect 23640 19612 23704 19616
rect 23640 19556 23644 19612
rect 23644 19556 23700 19612
rect 23700 19556 23704 19612
rect 23640 19552 23704 19556
rect 23720 19612 23784 19616
rect 23720 19556 23724 19612
rect 23724 19556 23780 19612
rect 23780 19556 23784 19612
rect 23720 19552 23784 19556
rect 29500 19408 29564 19412
rect 29500 19352 29550 19408
rect 29550 19352 29564 19408
rect 29500 19348 29564 19352
rect 30420 19348 30484 19412
rect 6584 19068 6648 19072
rect 6584 19012 6588 19068
rect 6588 19012 6644 19068
rect 6644 19012 6648 19068
rect 6584 19008 6648 19012
rect 6664 19068 6728 19072
rect 6664 19012 6668 19068
rect 6668 19012 6724 19068
rect 6724 19012 6728 19068
rect 6664 19008 6728 19012
rect 6744 19068 6808 19072
rect 6744 19012 6748 19068
rect 6748 19012 6804 19068
rect 6804 19012 6808 19068
rect 6744 19008 6808 19012
rect 6824 19068 6888 19072
rect 6824 19012 6828 19068
rect 6828 19012 6884 19068
rect 6884 19012 6888 19068
rect 6824 19008 6888 19012
rect 17848 19068 17912 19072
rect 17848 19012 17852 19068
rect 17852 19012 17908 19068
rect 17908 19012 17912 19068
rect 17848 19008 17912 19012
rect 17928 19068 17992 19072
rect 17928 19012 17932 19068
rect 17932 19012 17988 19068
rect 17988 19012 17992 19068
rect 17928 19008 17992 19012
rect 18008 19068 18072 19072
rect 18008 19012 18012 19068
rect 18012 19012 18068 19068
rect 18068 19012 18072 19068
rect 18008 19008 18072 19012
rect 18088 19068 18152 19072
rect 18088 19012 18092 19068
rect 18092 19012 18148 19068
rect 18148 19012 18152 19068
rect 18088 19008 18152 19012
rect 29112 19068 29176 19072
rect 29112 19012 29116 19068
rect 29116 19012 29172 19068
rect 29172 19012 29176 19068
rect 29112 19008 29176 19012
rect 29192 19068 29256 19072
rect 29192 19012 29196 19068
rect 29196 19012 29252 19068
rect 29252 19012 29256 19068
rect 29192 19008 29256 19012
rect 29272 19068 29336 19072
rect 29272 19012 29276 19068
rect 29276 19012 29332 19068
rect 29332 19012 29336 19068
rect 29272 19008 29336 19012
rect 29352 19068 29416 19072
rect 29352 19012 29356 19068
rect 29356 19012 29412 19068
rect 29412 19012 29416 19068
rect 29352 19008 29416 19012
rect 30052 18592 30116 18596
rect 30052 18536 30102 18592
rect 30102 18536 30116 18592
rect 30052 18532 30116 18536
rect 12216 18524 12280 18528
rect 12216 18468 12220 18524
rect 12220 18468 12276 18524
rect 12276 18468 12280 18524
rect 12216 18464 12280 18468
rect 12296 18524 12360 18528
rect 12296 18468 12300 18524
rect 12300 18468 12356 18524
rect 12356 18468 12360 18524
rect 12296 18464 12360 18468
rect 12376 18524 12440 18528
rect 12376 18468 12380 18524
rect 12380 18468 12436 18524
rect 12436 18468 12440 18524
rect 12376 18464 12440 18468
rect 12456 18524 12520 18528
rect 12456 18468 12460 18524
rect 12460 18468 12516 18524
rect 12516 18468 12520 18524
rect 12456 18464 12520 18468
rect 23480 18524 23544 18528
rect 23480 18468 23484 18524
rect 23484 18468 23540 18524
rect 23540 18468 23544 18524
rect 23480 18464 23544 18468
rect 23560 18524 23624 18528
rect 23560 18468 23564 18524
rect 23564 18468 23620 18524
rect 23620 18468 23624 18524
rect 23560 18464 23624 18468
rect 23640 18524 23704 18528
rect 23640 18468 23644 18524
rect 23644 18468 23700 18524
rect 23700 18468 23704 18524
rect 23640 18464 23704 18468
rect 23720 18524 23784 18528
rect 23720 18468 23724 18524
rect 23724 18468 23780 18524
rect 23780 18468 23784 18524
rect 23720 18464 23784 18468
rect 6584 17980 6648 17984
rect 6584 17924 6588 17980
rect 6588 17924 6644 17980
rect 6644 17924 6648 17980
rect 6584 17920 6648 17924
rect 6664 17980 6728 17984
rect 6664 17924 6668 17980
rect 6668 17924 6724 17980
rect 6724 17924 6728 17980
rect 6664 17920 6728 17924
rect 6744 17980 6808 17984
rect 6744 17924 6748 17980
rect 6748 17924 6804 17980
rect 6804 17924 6808 17980
rect 6744 17920 6808 17924
rect 6824 17980 6888 17984
rect 6824 17924 6828 17980
rect 6828 17924 6884 17980
rect 6884 17924 6888 17980
rect 6824 17920 6888 17924
rect 17848 17980 17912 17984
rect 17848 17924 17852 17980
rect 17852 17924 17908 17980
rect 17908 17924 17912 17980
rect 17848 17920 17912 17924
rect 17928 17980 17992 17984
rect 17928 17924 17932 17980
rect 17932 17924 17988 17980
rect 17988 17924 17992 17980
rect 17928 17920 17992 17924
rect 18008 17980 18072 17984
rect 18008 17924 18012 17980
rect 18012 17924 18068 17980
rect 18068 17924 18072 17980
rect 18008 17920 18072 17924
rect 18088 17980 18152 17984
rect 18088 17924 18092 17980
rect 18092 17924 18148 17980
rect 18148 17924 18152 17980
rect 18088 17920 18152 17924
rect 29112 17980 29176 17984
rect 29112 17924 29116 17980
rect 29116 17924 29172 17980
rect 29172 17924 29176 17980
rect 29112 17920 29176 17924
rect 29192 17980 29256 17984
rect 29192 17924 29196 17980
rect 29196 17924 29252 17980
rect 29252 17924 29256 17980
rect 29192 17920 29256 17924
rect 29272 17980 29336 17984
rect 29272 17924 29276 17980
rect 29276 17924 29332 17980
rect 29332 17924 29336 17980
rect 29272 17920 29336 17924
rect 29352 17980 29416 17984
rect 29352 17924 29356 17980
rect 29356 17924 29412 17980
rect 29412 17924 29416 17980
rect 29352 17920 29416 17924
rect 12216 17436 12280 17440
rect 12216 17380 12220 17436
rect 12220 17380 12276 17436
rect 12276 17380 12280 17436
rect 12216 17376 12280 17380
rect 12296 17436 12360 17440
rect 12296 17380 12300 17436
rect 12300 17380 12356 17436
rect 12356 17380 12360 17436
rect 12296 17376 12360 17380
rect 12376 17436 12440 17440
rect 12376 17380 12380 17436
rect 12380 17380 12436 17436
rect 12436 17380 12440 17436
rect 12376 17376 12440 17380
rect 12456 17436 12520 17440
rect 12456 17380 12460 17436
rect 12460 17380 12516 17436
rect 12516 17380 12520 17436
rect 12456 17376 12520 17380
rect 23480 17436 23544 17440
rect 23480 17380 23484 17436
rect 23484 17380 23540 17436
rect 23540 17380 23544 17436
rect 23480 17376 23544 17380
rect 23560 17436 23624 17440
rect 23560 17380 23564 17436
rect 23564 17380 23620 17436
rect 23620 17380 23624 17436
rect 23560 17376 23624 17380
rect 23640 17436 23704 17440
rect 23640 17380 23644 17436
rect 23644 17380 23700 17436
rect 23700 17380 23704 17436
rect 23640 17376 23704 17380
rect 23720 17436 23784 17440
rect 23720 17380 23724 17436
rect 23724 17380 23780 17436
rect 23780 17380 23784 17436
rect 23720 17376 23784 17380
rect 6584 16892 6648 16896
rect 6584 16836 6588 16892
rect 6588 16836 6644 16892
rect 6644 16836 6648 16892
rect 6584 16832 6648 16836
rect 6664 16892 6728 16896
rect 6664 16836 6668 16892
rect 6668 16836 6724 16892
rect 6724 16836 6728 16892
rect 6664 16832 6728 16836
rect 6744 16892 6808 16896
rect 6744 16836 6748 16892
rect 6748 16836 6804 16892
rect 6804 16836 6808 16892
rect 6744 16832 6808 16836
rect 6824 16892 6888 16896
rect 6824 16836 6828 16892
rect 6828 16836 6884 16892
rect 6884 16836 6888 16892
rect 6824 16832 6888 16836
rect 17848 16892 17912 16896
rect 17848 16836 17852 16892
rect 17852 16836 17908 16892
rect 17908 16836 17912 16892
rect 17848 16832 17912 16836
rect 17928 16892 17992 16896
rect 17928 16836 17932 16892
rect 17932 16836 17988 16892
rect 17988 16836 17992 16892
rect 17928 16832 17992 16836
rect 18008 16892 18072 16896
rect 18008 16836 18012 16892
rect 18012 16836 18068 16892
rect 18068 16836 18072 16892
rect 18008 16832 18072 16836
rect 18088 16892 18152 16896
rect 18088 16836 18092 16892
rect 18092 16836 18148 16892
rect 18148 16836 18152 16892
rect 18088 16832 18152 16836
rect 29112 16892 29176 16896
rect 29112 16836 29116 16892
rect 29116 16836 29172 16892
rect 29172 16836 29176 16892
rect 29112 16832 29176 16836
rect 29192 16892 29256 16896
rect 29192 16836 29196 16892
rect 29196 16836 29252 16892
rect 29252 16836 29256 16892
rect 29192 16832 29256 16836
rect 29272 16892 29336 16896
rect 29272 16836 29276 16892
rect 29276 16836 29332 16892
rect 29332 16836 29336 16892
rect 29272 16832 29336 16836
rect 29352 16892 29416 16896
rect 29352 16836 29356 16892
rect 29356 16836 29412 16892
rect 29412 16836 29416 16892
rect 29352 16832 29416 16836
rect 12216 16348 12280 16352
rect 12216 16292 12220 16348
rect 12220 16292 12276 16348
rect 12276 16292 12280 16348
rect 12216 16288 12280 16292
rect 12296 16348 12360 16352
rect 12296 16292 12300 16348
rect 12300 16292 12356 16348
rect 12356 16292 12360 16348
rect 12296 16288 12360 16292
rect 12376 16348 12440 16352
rect 12376 16292 12380 16348
rect 12380 16292 12436 16348
rect 12436 16292 12440 16348
rect 12376 16288 12440 16292
rect 12456 16348 12520 16352
rect 12456 16292 12460 16348
rect 12460 16292 12516 16348
rect 12516 16292 12520 16348
rect 12456 16288 12520 16292
rect 23480 16348 23544 16352
rect 23480 16292 23484 16348
rect 23484 16292 23540 16348
rect 23540 16292 23544 16348
rect 23480 16288 23544 16292
rect 23560 16348 23624 16352
rect 23560 16292 23564 16348
rect 23564 16292 23620 16348
rect 23620 16292 23624 16348
rect 23560 16288 23624 16292
rect 23640 16348 23704 16352
rect 23640 16292 23644 16348
rect 23644 16292 23700 16348
rect 23700 16292 23704 16348
rect 23640 16288 23704 16292
rect 23720 16348 23784 16352
rect 23720 16292 23724 16348
rect 23724 16292 23780 16348
rect 23780 16292 23784 16348
rect 23720 16288 23784 16292
rect 6584 15804 6648 15808
rect 6584 15748 6588 15804
rect 6588 15748 6644 15804
rect 6644 15748 6648 15804
rect 6584 15744 6648 15748
rect 6664 15804 6728 15808
rect 6664 15748 6668 15804
rect 6668 15748 6724 15804
rect 6724 15748 6728 15804
rect 6664 15744 6728 15748
rect 6744 15804 6808 15808
rect 6744 15748 6748 15804
rect 6748 15748 6804 15804
rect 6804 15748 6808 15804
rect 6744 15744 6808 15748
rect 6824 15804 6888 15808
rect 6824 15748 6828 15804
rect 6828 15748 6884 15804
rect 6884 15748 6888 15804
rect 6824 15744 6888 15748
rect 17848 15804 17912 15808
rect 17848 15748 17852 15804
rect 17852 15748 17908 15804
rect 17908 15748 17912 15804
rect 17848 15744 17912 15748
rect 17928 15804 17992 15808
rect 17928 15748 17932 15804
rect 17932 15748 17988 15804
rect 17988 15748 17992 15804
rect 17928 15744 17992 15748
rect 18008 15804 18072 15808
rect 18008 15748 18012 15804
rect 18012 15748 18068 15804
rect 18068 15748 18072 15804
rect 18008 15744 18072 15748
rect 18088 15804 18152 15808
rect 18088 15748 18092 15804
rect 18092 15748 18148 15804
rect 18148 15748 18152 15804
rect 18088 15744 18152 15748
rect 29112 15804 29176 15808
rect 29112 15748 29116 15804
rect 29116 15748 29172 15804
rect 29172 15748 29176 15804
rect 29112 15744 29176 15748
rect 29192 15804 29256 15808
rect 29192 15748 29196 15804
rect 29196 15748 29252 15804
rect 29252 15748 29256 15804
rect 29192 15744 29256 15748
rect 29272 15804 29336 15808
rect 29272 15748 29276 15804
rect 29276 15748 29332 15804
rect 29332 15748 29336 15804
rect 29272 15744 29336 15748
rect 29352 15804 29416 15808
rect 29352 15748 29356 15804
rect 29356 15748 29412 15804
rect 29412 15748 29416 15804
rect 29352 15744 29416 15748
rect 12216 15260 12280 15264
rect 12216 15204 12220 15260
rect 12220 15204 12276 15260
rect 12276 15204 12280 15260
rect 12216 15200 12280 15204
rect 12296 15260 12360 15264
rect 12296 15204 12300 15260
rect 12300 15204 12356 15260
rect 12356 15204 12360 15260
rect 12296 15200 12360 15204
rect 12376 15260 12440 15264
rect 12376 15204 12380 15260
rect 12380 15204 12436 15260
rect 12436 15204 12440 15260
rect 12376 15200 12440 15204
rect 12456 15260 12520 15264
rect 12456 15204 12460 15260
rect 12460 15204 12516 15260
rect 12516 15204 12520 15260
rect 12456 15200 12520 15204
rect 23480 15260 23544 15264
rect 23480 15204 23484 15260
rect 23484 15204 23540 15260
rect 23540 15204 23544 15260
rect 23480 15200 23544 15204
rect 23560 15260 23624 15264
rect 23560 15204 23564 15260
rect 23564 15204 23620 15260
rect 23620 15204 23624 15260
rect 23560 15200 23624 15204
rect 23640 15260 23704 15264
rect 23640 15204 23644 15260
rect 23644 15204 23700 15260
rect 23700 15204 23704 15260
rect 23640 15200 23704 15204
rect 23720 15260 23784 15264
rect 23720 15204 23724 15260
rect 23724 15204 23780 15260
rect 23780 15204 23784 15260
rect 23720 15200 23784 15204
rect 6584 14716 6648 14720
rect 6584 14660 6588 14716
rect 6588 14660 6644 14716
rect 6644 14660 6648 14716
rect 6584 14656 6648 14660
rect 6664 14716 6728 14720
rect 6664 14660 6668 14716
rect 6668 14660 6724 14716
rect 6724 14660 6728 14716
rect 6664 14656 6728 14660
rect 6744 14716 6808 14720
rect 6744 14660 6748 14716
rect 6748 14660 6804 14716
rect 6804 14660 6808 14716
rect 6744 14656 6808 14660
rect 6824 14716 6888 14720
rect 6824 14660 6828 14716
rect 6828 14660 6884 14716
rect 6884 14660 6888 14716
rect 6824 14656 6888 14660
rect 17848 14716 17912 14720
rect 17848 14660 17852 14716
rect 17852 14660 17908 14716
rect 17908 14660 17912 14716
rect 17848 14656 17912 14660
rect 17928 14716 17992 14720
rect 17928 14660 17932 14716
rect 17932 14660 17988 14716
rect 17988 14660 17992 14716
rect 17928 14656 17992 14660
rect 18008 14716 18072 14720
rect 18008 14660 18012 14716
rect 18012 14660 18068 14716
rect 18068 14660 18072 14716
rect 18008 14656 18072 14660
rect 18088 14716 18152 14720
rect 18088 14660 18092 14716
rect 18092 14660 18148 14716
rect 18148 14660 18152 14716
rect 18088 14656 18152 14660
rect 29112 14716 29176 14720
rect 29112 14660 29116 14716
rect 29116 14660 29172 14716
rect 29172 14660 29176 14716
rect 29112 14656 29176 14660
rect 29192 14716 29256 14720
rect 29192 14660 29196 14716
rect 29196 14660 29252 14716
rect 29252 14660 29256 14716
rect 29192 14656 29256 14660
rect 29272 14716 29336 14720
rect 29272 14660 29276 14716
rect 29276 14660 29332 14716
rect 29332 14660 29336 14716
rect 29272 14656 29336 14660
rect 29352 14716 29416 14720
rect 29352 14660 29356 14716
rect 29356 14660 29412 14716
rect 29412 14660 29416 14716
rect 29352 14656 29416 14660
rect 12216 14172 12280 14176
rect 12216 14116 12220 14172
rect 12220 14116 12276 14172
rect 12276 14116 12280 14172
rect 12216 14112 12280 14116
rect 12296 14172 12360 14176
rect 12296 14116 12300 14172
rect 12300 14116 12356 14172
rect 12356 14116 12360 14172
rect 12296 14112 12360 14116
rect 12376 14172 12440 14176
rect 12376 14116 12380 14172
rect 12380 14116 12436 14172
rect 12436 14116 12440 14172
rect 12376 14112 12440 14116
rect 12456 14172 12520 14176
rect 12456 14116 12460 14172
rect 12460 14116 12516 14172
rect 12516 14116 12520 14172
rect 12456 14112 12520 14116
rect 23480 14172 23544 14176
rect 23480 14116 23484 14172
rect 23484 14116 23540 14172
rect 23540 14116 23544 14172
rect 23480 14112 23544 14116
rect 23560 14172 23624 14176
rect 23560 14116 23564 14172
rect 23564 14116 23620 14172
rect 23620 14116 23624 14172
rect 23560 14112 23624 14116
rect 23640 14172 23704 14176
rect 23640 14116 23644 14172
rect 23644 14116 23700 14172
rect 23700 14116 23704 14172
rect 23640 14112 23704 14116
rect 23720 14172 23784 14176
rect 23720 14116 23724 14172
rect 23724 14116 23780 14172
rect 23780 14116 23784 14172
rect 23720 14112 23784 14116
rect 6584 13628 6648 13632
rect 6584 13572 6588 13628
rect 6588 13572 6644 13628
rect 6644 13572 6648 13628
rect 6584 13568 6648 13572
rect 6664 13628 6728 13632
rect 6664 13572 6668 13628
rect 6668 13572 6724 13628
rect 6724 13572 6728 13628
rect 6664 13568 6728 13572
rect 6744 13628 6808 13632
rect 6744 13572 6748 13628
rect 6748 13572 6804 13628
rect 6804 13572 6808 13628
rect 6744 13568 6808 13572
rect 6824 13628 6888 13632
rect 6824 13572 6828 13628
rect 6828 13572 6884 13628
rect 6884 13572 6888 13628
rect 6824 13568 6888 13572
rect 17848 13628 17912 13632
rect 17848 13572 17852 13628
rect 17852 13572 17908 13628
rect 17908 13572 17912 13628
rect 17848 13568 17912 13572
rect 17928 13628 17992 13632
rect 17928 13572 17932 13628
rect 17932 13572 17988 13628
rect 17988 13572 17992 13628
rect 17928 13568 17992 13572
rect 18008 13628 18072 13632
rect 18008 13572 18012 13628
rect 18012 13572 18068 13628
rect 18068 13572 18072 13628
rect 18008 13568 18072 13572
rect 18088 13628 18152 13632
rect 18088 13572 18092 13628
rect 18092 13572 18148 13628
rect 18148 13572 18152 13628
rect 18088 13568 18152 13572
rect 29112 13628 29176 13632
rect 29112 13572 29116 13628
rect 29116 13572 29172 13628
rect 29172 13572 29176 13628
rect 29112 13568 29176 13572
rect 29192 13628 29256 13632
rect 29192 13572 29196 13628
rect 29196 13572 29252 13628
rect 29252 13572 29256 13628
rect 29192 13568 29256 13572
rect 29272 13628 29336 13632
rect 29272 13572 29276 13628
rect 29276 13572 29332 13628
rect 29332 13572 29336 13628
rect 29272 13568 29336 13572
rect 29352 13628 29416 13632
rect 29352 13572 29356 13628
rect 29356 13572 29412 13628
rect 29412 13572 29416 13628
rect 29352 13568 29416 13572
rect 12216 13084 12280 13088
rect 12216 13028 12220 13084
rect 12220 13028 12276 13084
rect 12276 13028 12280 13084
rect 12216 13024 12280 13028
rect 12296 13084 12360 13088
rect 12296 13028 12300 13084
rect 12300 13028 12356 13084
rect 12356 13028 12360 13084
rect 12296 13024 12360 13028
rect 12376 13084 12440 13088
rect 12376 13028 12380 13084
rect 12380 13028 12436 13084
rect 12436 13028 12440 13084
rect 12376 13024 12440 13028
rect 12456 13084 12520 13088
rect 12456 13028 12460 13084
rect 12460 13028 12516 13084
rect 12516 13028 12520 13084
rect 12456 13024 12520 13028
rect 23480 13084 23544 13088
rect 23480 13028 23484 13084
rect 23484 13028 23540 13084
rect 23540 13028 23544 13084
rect 23480 13024 23544 13028
rect 23560 13084 23624 13088
rect 23560 13028 23564 13084
rect 23564 13028 23620 13084
rect 23620 13028 23624 13084
rect 23560 13024 23624 13028
rect 23640 13084 23704 13088
rect 23640 13028 23644 13084
rect 23644 13028 23700 13084
rect 23700 13028 23704 13084
rect 23640 13024 23704 13028
rect 23720 13084 23784 13088
rect 23720 13028 23724 13084
rect 23724 13028 23780 13084
rect 23780 13028 23784 13084
rect 23720 13024 23784 13028
rect 6584 12540 6648 12544
rect 6584 12484 6588 12540
rect 6588 12484 6644 12540
rect 6644 12484 6648 12540
rect 6584 12480 6648 12484
rect 6664 12540 6728 12544
rect 6664 12484 6668 12540
rect 6668 12484 6724 12540
rect 6724 12484 6728 12540
rect 6664 12480 6728 12484
rect 6744 12540 6808 12544
rect 6744 12484 6748 12540
rect 6748 12484 6804 12540
rect 6804 12484 6808 12540
rect 6744 12480 6808 12484
rect 6824 12540 6888 12544
rect 6824 12484 6828 12540
rect 6828 12484 6884 12540
rect 6884 12484 6888 12540
rect 6824 12480 6888 12484
rect 17848 12540 17912 12544
rect 17848 12484 17852 12540
rect 17852 12484 17908 12540
rect 17908 12484 17912 12540
rect 17848 12480 17912 12484
rect 17928 12540 17992 12544
rect 17928 12484 17932 12540
rect 17932 12484 17988 12540
rect 17988 12484 17992 12540
rect 17928 12480 17992 12484
rect 18008 12540 18072 12544
rect 18008 12484 18012 12540
rect 18012 12484 18068 12540
rect 18068 12484 18072 12540
rect 18008 12480 18072 12484
rect 18088 12540 18152 12544
rect 18088 12484 18092 12540
rect 18092 12484 18148 12540
rect 18148 12484 18152 12540
rect 18088 12480 18152 12484
rect 29112 12540 29176 12544
rect 29112 12484 29116 12540
rect 29116 12484 29172 12540
rect 29172 12484 29176 12540
rect 29112 12480 29176 12484
rect 29192 12540 29256 12544
rect 29192 12484 29196 12540
rect 29196 12484 29252 12540
rect 29252 12484 29256 12540
rect 29192 12480 29256 12484
rect 29272 12540 29336 12544
rect 29272 12484 29276 12540
rect 29276 12484 29332 12540
rect 29332 12484 29336 12540
rect 29272 12480 29336 12484
rect 29352 12540 29416 12544
rect 29352 12484 29356 12540
rect 29356 12484 29412 12540
rect 29412 12484 29416 12540
rect 29352 12480 29416 12484
rect 12216 11996 12280 12000
rect 12216 11940 12220 11996
rect 12220 11940 12276 11996
rect 12276 11940 12280 11996
rect 12216 11936 12280 11940
rect 12296 11996 12360 12000
rect 12296 11940 12300 11996
rect 12300 11940 12356 11996
rect 12356 11940 12360 11996
rect 12296 11936 12360 11940
rect 12376 11996 12440 12000
rect 12376 11940 12380 11996
rect 12380 11940 12436 11996
rect 12436 11940 12440 11996
rect 12376 11936 12440 11940
rect 12456 11996 12520 12000
rect 12456 11940 12460 11996
rect 12460 11940 12516 11996
rect 12516 11940 12520 11996
rect 12456 11936 12520 11940
rect 23480 11996 23544 12000
rect 23480 11940 23484 11996
rect 23484 11940 23540 11996
rect 23540 11940 23544 11996
rect 23480 11936 23544 11940
rect 23560 11996 23624 12000
rect 23560 11940 23564 11996
rect 23564 11940 23620 11996
rect 23620 11940 23624 11996
rect 23560 11936 23624 11940
rect 23640 11996 23704 12000
rect 23640 11940 23644 11996
rect 23644 11940 23700 11996
rect 23700 11940 23704 11996
rect 23640 11936 23704 11940
rect 23720 11996 23784 12000
rect 23720 11940 23724 11996
rect 23724 11940 23780 11996
rect 23780 11940 23784 11996
rect 23720 11936 23784 11940
rect 6584 11452 6648 11456
rect 6584 11396 6588 11452
rect 6588 11396 6644 11452
rect 6644 11396 6648 11452
rect 6584 11392 6648 11396
rect 6664 11452 6728 11456
rect 6664 11396 6668 11452
rect 6668 11396 6724 11452
rect 6724 11396 6728 11452
rect 6664 11392 6728 11396
rect 6744 11452 6808 11456
rect 6744 11396 6748 11452
rect 6748 11396 6804 11452
rect 6804 11396 6808 11452
rect 6744 11392 6808 11396
rect 6824 11452 6888 11456
rect 6824 11396 6828 11452
rect 6828 11396 6884 11452
rect 6884 11396 6888 11452
rect 6824 11392 6888 11396
rect 17848 11452 17912 11456
rect 17848 11396 17852 11452
rect 17852 11396 17908 11452
rect 17908 11396 17912 11452
rect 17848 11392 17912 11396
rect 17928 11452 17992 11456
rect 17928 11396 17932 11452
rect 17932 11396 17988 11452
rect 17988 11396 17992 11452
rect 17928 11392 17992 11396
rect 18008 11452 18072 11456
rect 18008 11396 18012 11452
rect 18012 11396 18068 11452
rect 18068 11396 18072 11452
rect 18008 11392 18072 11396
rect 18088 11452 18152 11456
rect 18088 11396 18092 11452
rect 18092 11396 18148 11452
rect 18148 11396 18152 11452
rect 18088 11392 18152 11396
rect 29112 11452 29176 11456
rect 29112 11396 29116 11452
rect 29116 11396 29172 11452
rect 29172 11396 29176 11452
rect 29112 11392 29176 11396
rect 29192 11452 29256 11456
rect 29192 11396 29196 11452
rect 29196 11396 29252 11452
rect 29252 11396 29256 11452
rect 29192 11392 29256 11396
rect 29272 11452 29336 11456
rect 29272 11396 29276 11452
rect 29276 11396 29332 11452
rect 29332 11396 29336 11452
rect 29272 11392 29336 11396
rect 29352 11452 29416 11456
rect 29352 11396 29356 11452
rect 29356 11396 29412 11452
rect 29412 11396 29416 11452
rect 29352 11392 29416 11396
rect 12216 10908 12280 10912
rect 12216 10852 12220 10908
rect 12220 10852 12276 10908
rect 12276 10852 12280 10908
rect 12216 10848 12280 10852
rect 12296 10908 12360 10912
rect 12296 10852 12300 10908
rect 12300 10852 12356 10908
rect 12356 10852 12360 10908
rect 12296 10848 12360 10852
rect 12376 10908 12440 10912
rect 12376 10852 12380 10908
rect 12380 10852 12436 10908
rect 12436 10852 12440 10908
rect 12376 10848 12440 10852
rect 12456 10908 12520 10912
rect 12456 10852 12460 10908
rect 12460 10852 12516 10908
rect 12516 10852 12520 10908
rect 12456 10848 12520 10852
rect 23480 10908 23544 10912
rect 23480 10852 23484 10908
rect 23484 10852 23540 10908
rect 23540 10852 23544 10908
rect 23480 10848 23544 10852
rect 23560 10908 23624 10912
rect 23560 10852 23564 10908
rect 23564 10852 23620 10908
rect 23620 10852 23624 10908
rect 23560 10848 23624 10852
rect 23640 10908 23704 10912
rect 23640 10852 23644 10908
rect 23644 10852 23700 10908
rect 23700 10852 23704 10908
rect 23640 10848 23704 10852
rect 23720 10908 23784 10912
rect 23720 10852 23724 10908
rect 23724 10852 23780 10908
rect 23780 10852 23784 10908
rect 23720 10848 23784 10852
rect 6584 10364 6648 10368
rect 6584 10308 6588 10364
rect 6588 10308 6644 10364
rect 6644 10308 6648 10364
rect 6584 10304 6648 10308
rect 6664 10364 6728 10368
rect 6664 10308 6668 10364
rect 6668 10308 6724 10364
rect 6724 10308 6728 10364
rect 6664 10304 6728 10308
rect 6744 10364 6808 10368
rect 6744 10308 6748 10364
rect 6748 10308 6804 10364
rect 6804 10308 6808 10364
rect 6744 10304 6808 10308
rect 6824 10364 6888 10368
rect 6824 10308 6828 10364
rect 6828 10308 6884 10364
rect 6884 10308 6888 10364
rect 6824 10304 6888 10308
rect 17848 10364 17912 10368
rect 17848 10308 17852 10364
rect 17852 10308 17908 10364
rect 17908 10308 17912 10364
rect 17848 10304 17912 10308
rect 17928 10364 17992 10368
rect 17928 10308 17932 10364
rect 17932 10308 17988 10364
rect 17988 10308 17992 10364
rect 17928 10304 17992 10308
rect 18008 10364 18072 10368
rect 18008 10308 18012 10364
rect 18012 10308 18068 10364
rect 18068 10308 18072 10364
rect 18008 10304 18072 10308
rect 18088 10364 18152 10368
rect 18088 10308 18092 10364
rect 18092 10308 18148 10364
rect 18148 10308 18152 10364
rect 18088 10304 18152 10308
rect 29112 10364 29176 10368
rect 29112 10308 29116 10364
rect 29116 10308 29172 10364
rect 29172 10308 29176 10364
rect 29112 10304 29176 10308
rect 29192 10364 29256 10368
rect 29192 10308 29196 10364
rect 29196 10308 29252 10364
rect 29252 10308 29256 10364
rect 29192 10304 29256 10308
rect 29272 10364 29336 10368
rect 29272 10308 29276 10364
rect 29276 10308 29332 10364
rect 29332 10308 29336 10364
rect 29272 10304 29336 10308
rect 29352 10364 29416 10368
rect 29352 10308 29356 10364
rect 29356 10308 29412 10364
rect 29412 10308 29416 10364
rect 29352 10304 29416 10308
rect 12216 9820 12280 9824
rect 12216 9764 12220 9820
rect 12220 9764 12276 9820
rect 12276 9764 12280 9820
rect 12216 9760 12280 9764
rect 12296 9820 12360 9824
rect 12296 9764 12300 9820
rect 12300 9764 12356 9820
rect 12356 9764 12360 9820
rect 12296 9760 12360 9764
rect 12376 9820 12440 9824
rect 12376 9764 12380 9820
rect 12380 9764 12436 9820
rect 12436 9764 12440 9820
rect 12376 9760 12440 9764
rect 12456 9820 12520 9824
rect 12456 9764 12460 9820
rect 12460 9764 12516 9820
rect 12516 9764 12520 9820
rect 12456 9760 12520 9764
rect 23480 9820 23544 9824
rect 23480 9764 23484 9820
rect 23484 9764 23540 9820
rect 23540 9764 23544 9820
rect 23480 9760 23544 9764
rect 23560 9820 23624 9824
rect 23560 9764 23564 9820
rect 23564 9764 23620 9820
rect 23620 9764 23624 9820
rect 23560 9760 23624 9764
rect 23640 9820 23704 9824
rect 23640 9764 23644 9820
rect 23644 9764 23700 9820
rect 23700 9764 23704 9820
rect 23640 9760 23704 9764
rect 23720 9820 23784 9824
rect 23720 9764 23724 9820
rect 23724 9764 23780 9820
rect 23780 9764 23784 9820
rect 23720 9760 23784 9764
rect 6584 9276 6648 9280
rect 6584 9220 6588 9276
rect 6588 9220 6644 9276
rect 6644 9220 6648 9276
rect 6584 9216 6648 9220
rect 6664 9276 6728 9280
rect 6664 9220 6668 9276
rect 6668 9220 6724 9276
rect 6724 9220 6728 9276
rect 6664 9216 6728 9220
rect 6744 9276 6808 9280
rect 6744 9220 6748 9276
rect 6748 9220 6804 9276
rect 6804 9220 6808 9276
rect 6744 9216 6808 9220
rect 6824 9276 6888 9280
rect 6824 9220 6828 9276
rect 6828 9220 6884 9276
rect 6884 9220 6888 9276
rect 6824 9216 6888 9220
rect 17848 9276 17912 9280
rect 17848 9220 17852 9276
rect 17852 9220 17908 9276
rect 17908 9220 17912 9276
rect 17848 9216 17912 9220
rect 17928 9276 17992 9280
rect 17928 9220 17932 9276
rect 17932 9220 17988 9276
rect 17988 9220 17992 9276
rect 17928 9216 17992 9220
rect 18008 9276 18072 9280
rect 18008 9220 18012 9276
rect 18012 9220 18068 9276
rect 18068 9220 18072 9276
rect 18008 9216 18072 9220
rect 18088 9276 18152 9280
rect 18088 9220 18092 9276
rect 18092 9220 18148 9276
rect 18148 9220 18152 9276
rect 18088 9216 18152 9220
rect 29112 9276 29176 9280
rect 29112 9220 29116 9276
rect 29116 9220 29172 9276
rect 29172 9220 29176 9276
rect 29112 9216 29176 9220
rect 29192 9276 29256 9280
rect 29192 9220 29196 9276
rect 29196 9220 29252 9276
rect 29252 9220 29256 9276
rect 29192 9216 29256 9220
rect 29272 9276 29336 9280
rect 29272 9220 29276 9276
rect 29276 9220 29332 9276
rect 29332 9220 29336 9276
rect 29272 9216 29336 9220
rect 29352 9276 29416 9280
rect 29352 9220 29356 9276
rect 29356 9220 29412 9276
rect 29412 9220 29416 9276
rect 29352 9216 29416 9220
rect 12216 8732 12280 8736
rect 12216 8676 12220 8732
rect 12220 8676 12276 8732
rect 12276 8676 12280 8732
rect 12216 8672 12280 8676
rect 12296 8732 12360 8736
rect 12296 8676 12300 8732
rect 12300 8676 12356 8732
rect 12356 8676 12360 8732
rect 12296 8672 12360 8676
rect 12376 8732 12440 8736
rect 12376 8676 12380 8732
rect 12380 8676 12436 8732
rect 12436 8676 12440 8732
rect 12376 8672 12440 8676
rect 12456 8732 12520 8736
rect 12456 8676 12460 8732
rect 12460 8676 12516 8732
rect 12516 8676 12520 8732
rect 12456 8672 12520 8676
rect 23480 8732 23544 8736
rect 23480 8676 23484 8732
rect 23484 8676 23540 8732
rect 23540 8676 23544 8732
rect 23480 8672 23544 8676
rect 23560 8732 23624 8736
rect 23560 8676 23564 8732
rect 23564 8676 23620 8732
rect 23620 8676 23624 8732
rect 23560 8672 23624 8676
rect 23640 8732 23704 8736
rect 23640 8676 23644 8732
rect 23644 8676 23700 8732
rect 23700 8676 23704 8732
rect 23640 8672 23704 8676
rect 23720 8732 23784 8736
rect 23720 8676 23724 8732
rect 23724 8676 23780 8732
rect 23780 8676 23784 8732
rect 23720 8672 23784 8676
rect 6584 8188 6648 8192
rect 6584 8132 6588 8188
rect 6588 8132 6644 8188
rect 6644 8132 6648 8188
rect 6584 8128 6648 8132
rect 6664 8188 6728 8192
rect 6664 8132 6668 8188
rect 6668 8132 6724 8188
rect 6724 8132 6728 8188
rect 6664 8128 6728 8132
rect 6744 8188 6808 8192
rect 6744 8132 6748 8188
rect 6748 8132 6804 8188
rect 6804 8132 6808 8188
rect 6744 8128 6808 8132
rect 6824 8188 6888 8192
rect 6824 8132 6828 8188
rect 6828 8132 6884 8188
rect 6884 8132 6888 8188
rect 6824 8128 6888 8132
rect 17848 8188 17912 8192
rect 17848 8132 17852 8188
rect 17852 8132 17908 8188
rect 17908 8132 17912 8188
rect 17848 8128 17912 8132
rect 17928 8188 17992 8192
rect 17928 8132 17932 8188
rect 17932 8132 17988 8188
rect 17988 8132 17992 8188
rect 17928 8128 17992 8132
rect 18008 8188 18072 8192
rect 18008 8132 18012 8188
rect 18012 8132 18068 8188
rect 18068 8132 18072 8188
rect 18008 8128 18072 8132
rect 18088 8188 18152 8192
rect 18088 8132 18092 8188
rect 18092 8132 18148 8188
rect 18148 8132 18152 8188
rect 18088 8128 18152 8132
rect 29112 8188 29176 8192
rect 29112 8132 29116 8188
rect 29116 8132 29172 8188
rect 29172 8132 29176 8188
rect 29112 8128 29176 8132
rect 29192 8188 29256 8192
rect 29192 8132 29196 8188
rect 29196 8132 29252 8188
rect 29252 8132 29256 8188
rect 29192 8128 29256 8132
rect 29272 8188 29336 8192
rect 29272 8132 29276 8188
rect 29276 8132 29332 8188
rect 29332 8132 29336 8188
rect 29272 8128 29336 8132
rect 29352 8188 29416 8192
rect 29352 8132 29356 8188
rect 29356 8132 29412 8188
rect 29412 8132 29416 8188
rect 29352 8128 29416 8132
rect 12216 7644 12280 7648
rect 12216 7588 12220 7644
rect 12220 7588 12276 7644
rect 12276 7588 12280 7644
rect 12216 7584 12280 7588
rect 12296 7644 12360 7648
rect 12296 7588 12300 7644
rect 12300 7588 12356 7644
rect 12356 7588 12360 7644
rect 12296 7584 12360 7588
rect 12376 7644 12440 7648
rect 12376 7588 12380 7644
rect 12380 7588 12436 7644
rect 12436 7588 12440 7644
rect 12376 7584 12440 7588
rect 12456 7644 12520 7648
rect 12456 7588 12460 7644
rect 12460 7588 12516 7644
rect 12516 7588 12520 7644
rect 12456 7584 12520 7588
rect 23480 7644 23544 7648
rect 23480 7588 23484 7644
rect 23484 7588 23540 7644
rect 23540 7588 23544 7644
rect 23480 7584 23544 7588
rect 23560 7644 23624 7648
rect 23560 7588 23564 7644
rect 23564 7588 23620 7644
rect 23620 7588 23624 7644
rect 23560 7584 23624 7588
rect 23640 7644 23704 7648
rect 23640 7588 23644 7644
rect 23644 7588 23700 7644
rect 23700 7588 23704 7644
rect 23640 7584 23704 7588
rect 23720 7644 23784 7648
rect 23720 7588 23724 7644
rect 23724 7588 23780 7644
rect 23780 7588 23784 7644
rect 23720 7584 23784 7588
rect 6584 7100 6648 7104
rect 6584 7044 6588 7100
rect 6588 7044 6644 7100
rect 6644 7044 6648 7100
rect 6584 7040 6648 7044
rect 6664 7100 6728 7104
rect 6664 7044 6668 7100
rect 6668 7044 6724 7100
rect 6724 7044 6728 7100
rect 6664 7040 6728 7044
rect 6744 7100 6808 7104
rect 6744 7044 6748 7100
rect 6748 7044 6804 7100
rect 6804 7044 6808 7100
rect 6744 7040 6808 7044
rect 6824 7100 6888 7104
rect 6824 7044 6828 7100
rect 6828 7044 6884 7100
rect 6884 7044 6888 7100
rect 6824 7040 6888 7044
rect 17848 7100 17912 7104
rect 17848 7044 17852 7100
rect 17852 7044 17908 7100
rect 17908 7044 17912 7100
rect 17848 7040 17912 7044
rect 17928 7100 17992 7104
rect 17928 7044 17932 7100
rect 17932 7044 17988 7100
rect 17988 7044 17992 7100
rect 17928 7040 17992 7044
rect 18008 7100 18072 7104
rect 18008 7044 18012 7100
rect 18012 7044 18068 7100
rect 18068 7044 18072 7100
rect 18008 7040 18072 7044
rect 18088 7100 18152 7104
rect 18088 7044 18092 7100
rect 18092 7044 18148 7100
rect 18148 7044 18152 7100
rect 18088 7040 18152 7044
rect 29112 7100 29176 7104
rect 29112 7044 29116 7100
rect 29116 7044 29172 7100
rect 29172 7044 29176 7100
rect 29112 7040 29176 7044
rect 29192 7100 29256 7104
rect 29192 7044 29196 7100
rect 29196 7044 29252 7100
rect 29252 7044 29256 7100
rect 29192 7040 29256 7044
rect 29272 7100 29336 7104
rect 29272 7044 29276 7100
rect 29276 7044 29332 7100
rect 29332 7044 29336 7100
rect 29272 7040 29336 7044
rect 29352 7100 29416 7104
rect 29352 7044 29356 7100
rect 29356 7044 29412 7100
rect 29412 7044 29416 7100
rect 29352 7040 29416 7044
rect 12216 6556 12280 6560
rect 12216 6500 12220 6556
rect 12220 6500 12276 6556
rect 12276 6500 12280 6556
rect 12216 6496 12280 6500
rect 12296 6556 12360 6560
rect 12296 6500 12300 6556
rect 12300 6500 12356 6556
rect 12356 6500 12360 6556
rect 12296 6496 12360 6500
rect 12376 6556 12440 6560
rect 12376 6500 12380 6556
rect 12380 6500 12436 6556
rect 12436 6500 12440 6556
rect 12376 6496 12440 6500
rect 12456 6556 12520 6560
rect 12456 6500 12460 6556
rect 12460 6500 12516 6556
rect 12516 6500 12520 6556
rect 12456 6496 12520 6500
rect 23480 6556 23544 6560
rect 23480 6500 23484 6556
rect 23484 6500 23540 6556
rect 23540 6500 23544 6556
rect 23480 6496 23544 6500
rect 23560 6556 23624 6560
rect 23560 6500 23564 6556
rect 23564 6500 23620 6556
rect 23620 6500 23624 6556
rect 23560 6496 23624 6500
rect 23640 6556 23704 6560
rect 23640 6500 23644 6556
rect 23644 6500 23700 6556
rect 23700 6500 23704 6556
rect 23640 6496 23704 6500
rect 23720 6556 23784 6560
rect 23720 6500 23724 6556
rect 23724 6500 23780 6556
rect 23780 6500 23784 6556
rect 23720 6496 23784 6500
rect 6584 6012 6648 6016
rect 6584 5956 6588 6012
rect 6588 5956 6644 6012
rect 6644 5956 6648 6012
rect 6584 5952 6648 5956
rect 6664 6012 6728 6016
rect 6664 5956 6668 6012
rect 6668 5956 6724 6012
rect 6724 5956 6728 6012
rect 6664 5952 6728 5956
rect 6744 6012 6808 6016
rect 6744 5956 6748 6012
rect 6748 5956 6804 6012
rect 6804 5956 6808 6012
rect 6744 5952 6808 5956
rect 6824 6012 6888 6016
rect 6824 5956 6828 6012
rect 6828 5956 6884 6012
rect 6884 5956 6888 6012
rect 6824 5952 6888 5956
rect 17848 6012 17912 6016
rect 17848 5956 17852 6012
rect 17852 5956 17908 6012
rect 17908 5956 17912 6012
rect 17848 5952 17912 5956
rect 17928 6012 17992 6016
rect 17928 5956 17932 6012
rect 17932 5956 17988 6012
rect 17988 5956 17992 6012
rect 17928 5952 17992 5956
rect 18008 6012 18072 6016
rect 18008 5956 18012 6012
rect 18012 5956 18068 6012
rect 18068 5956 18072 6012
rect 18008 5952 18072 5956
rect 18088 6012 18152 6016
rect 18088 5956 18092 6012
rect 18092 5956 18148 6012
rect 18148 5956 18152 6012
rect 18088 5952 18152 5956
rect 29112 6012 29176 6016
rect 29112 5956 29116 6012
rect 29116 5956 29172 6012
rect 29172 5956 29176 6012
rect 29112 5952 29176 5956
rect 29192 6012 29256 6016
rect 29192 5956 29196 6012
rect 29196 5956 29252 6012
rect 29252 5956 29256 6012
rect 29192 5952 29256 5956
rect 29272 6012 29336 6016
rect 29272 5956 29276 6012
rect 29276 5956 29332 6012
rect 29332 5956 29336 6012
rect 29272 5952 29336 5956
rect 29352 6012 29416 6016
rect 29352 5956 29356 6012
rect 29356 5956 29412 6012
rect 29412 5956 29416 6012
rect 29352 5952 29416 5956
rect 12216 5468 12280 5472
rect 12216 5412 12220 5468
rect 12220 5412 12276 5468
rect 12276 5412 12280 5468
rect 12216 5408 12280 5412
rect 12296 5468 12360 5472
rect 12296 5412 12300 5468
rect 12300 5412 12356 5468
rect 12356 5412 12360 5468
rect 12296 5408 12360 5412
rect 12376 5468 12440 5472
rect 12376 5412 12380 5468
rect 12380 5412 12436 5468
rect 12436 5412 12440 5468
rect 12376 5408 12440 5412
rect 12456 5468 12520 5472
rect 12456 5412 12460 5468
rect 12460 5412 12516 5468
rect 12516 5412 12520 5468
rect 12456 5408 12520 5412
rect 23480 5468 23544 5472
rect 23480 5412 23484 5468
rect 23484 5412 23540 5468
rect 23540 5412 23544 5468
rect 23480 5408 23544 5412
rect 23560 5468 23624 5472
rect 23560 5412 23564 5468
rect 23564 5412 23620 5468
rect 23620 5412 23624 5468
rect 23560 5408 23624 5412
rect 23640 5468 23704 5472
rect 23640 5412 23644 5468
rect 23644 5412 23700 5468
rect 23700 5412 23704 5468
rect 23640 5408 23704 5412
rect 23720 5468 23784 5472
rect 23720 5412 23724 5468
rect 23724 5412 23780 5468
rect 23780 5412 23784 5468
rect 23720 5408 23784 5412
rect 6584 4924 6648 4928
rect 6584 4868 6588 4924
rect 6588 4868 6644 4924
rect 6644 4868 6648 4924
rect 6584 4864 6648 4868
rect 6664 4924 6728 4928
rect 6664 4868 6668 4924
rect 6668 4868 6724 4924
rect 6724 4868 6728 4924
rect 6664 4864 6728 4868
rect 6744 4924 6808 4928
rect 6744 4868 6748 4924
rect 6748 4868 6804 4924
rect 6804 4868 6808 4924
rect 6744 4864 6808 4868
rect 6824 4924 6888 4928
rect 6824 4868 6828 4924
rect 6828 4868 6884 4924
rect 6884 4868 6888 4924
rect 6824 4864 6888 4868
rect 17848 4924 17912 4928
rect 17848 4868 17852 4924
rect 17852 4868 17908 4924
rect 17908 4868 17912 4924
rect 17848 4864 17912 4868
rect 17928 4924 17992 4928
rect 17928 4868 17932 4924
rect 17932 4868 17988 4924
rect 17988 4868 17992 4924
rect 17928 4864 17992 4868
rect 18008 4924 18072 4928
rect 18008 4868 18012 4924
rect 18012 4868 18068 4924
rect 18068 4868 18072 4924
rect 18008 4864 18072 4868
rect 18088 4924 18152 4928
rect 18088 4868 18092 4924
rect 18092 4868 18148 4924
rect 18148 4868 18152 4924
rect 18088 4864 18152 4868
rect 29112 4924 29176 4928
rect 29112 4868 29116 4924
rect 29116 4868 29172 4924
rect 29172 4868 29176 4924
rect 29112 4864 29176 4868
rect 29192 4924 29256 4928
rect 29192 4868 29196 4924
rect 29196 4868 29252 4924
rect 29252 4868 29256 4924
rect 29192 4864 29256 4868
rect 29272 4924 29336 4928
rect 29272 4868 29276 4924
rect 29276 4868 29332 4924
rect 29332 4868 29336 4924
rect 29272 4864 29336 4868
rect 29352 4924 29416 4928
rect 29352 4868 29356 4924
rect 29356 4868 29412 4924
rect 29412 4868 29416 4924
rect 29352 4864 29416 4868
rect 12216 4380 12280 4384
rect 12216 4324 12220 4380
rect 12220 4324 12276 4380
rect 12276 4324 12280 4380
rect 12216 4320 12280 4324
rect 12296 4380 12360 4384
rect 12296 4324 12300 4380
rect 12300 4324 12356 4380
rect 12356 4324 12360 4380
rect 12296 4320 12360 4324
rect 12376 4380 12440 4384
rect 12376 4324 12380 4380
rect 12380 4324 12436 4380
rect 12436 4324 12440 4380
rect 12376 4320 12440 4324
rect 12456 4380 12520 4384
rect 12456 4324 12460 4380
rect 12460 4324 12516 4380
rect 12516 4324 12520 4380
rect 12456 4320 12520 4324
rect 23480 4380 23544 4384
rect 23480 4324 23484 4380
rect 23484 4324 23540 4380
rect 23540 4324 23544 4380
rect 23480 4320 23544 4324
rect 23560 4380 23624 4384
rect 23560 4324 23564 4380
rect 23564 4324 23620 4380
rect 23620 4324 23624 4380
rect 23560 4320 23624 4324
rect 23640 4380 23704 4384
rect 23640 4324 23644 4380
rect 23644 4324 23700 4380
rect 23700 4324 23704 4380
rect 23640 4320 23704 4324
rect 23720 4380 23784 4384
rect 23720 4324 23724 4380
rect 23724 4324 23780 4380
rect 23780 4324 23784 4380
rect 23720 4320 23784 4324
rect 6584 3836 6648 3840
rect 6584 3780 6588 3836
rect 6588 3780 6644 3836
rect 6644 3780 6648 3836
rect 6584 3776 6648 3780
rect 6664 3836 6728 3840
rect 6664 3780 6668 3836
rect 6668 3780 6724 3836
rect 6724 3780 6728 3836
rect 6664 3776 6728 3780
rect 6744 3836 6808 3840
rect 6744 3780 6748 3836
rect 6748 3780 6804 3836
rect 6804 3780 6808 3836
rect 6744 3776 6808 3780
rect 6824 3836 6888 3840
rect 6824 3780 6828 3836
rect 6828 3780 6884 3836
rect 6884 3780 6888 3836
rect 6824 3776 6888 3780
rect 17848 3836 17912 3840
rect 17848 3780 17852 3836
rect 17852 3780 17908 3836
rect 17908 3780 17912 3836
rect 17848 3776 17912 3780
rect 17928 3836 17992 3840
rect 17928 3780 17932 3836
rect 17932 3780 17988 3836
rect 17988 3780 17992 3836
rect 17928 3776 17992 3780
rect 18008 3836 18072 3840
rect 18008 3780 18012 3836
rect 18012 3780 18068 3836
rect 18068 3780 18072 3836
rect 18008 3776 18072 3780
rect 18088 3836 18152 3840
rect 18088 3780 18092 3836
rect 18092 3780 18148 3836
rect 18148 3780 18152 3836
rect 18088 3776 18152 3780
rect 29112 3836 29176 3840
rect 29112 3780 29116 3836
rect 29116 3780 29172 3836
rect 29172 3780 29176 3836
rect 29112 3776 29176 3780
rect 29192 3836 29256 3840
rect 29192 3780 29196 3836
rect 29196 3780 29252 3836
rect 29252 3780 29256 3836
rect 29192 3776 29256 3780
rect 29272 3836 29336 3840
rect 29272 3780 29276 3836
rect 29276 3780 29332 3836
rect 29332 3780 29336 3836
rect 29272 3776 29336 3780
rect 29352 3836 29416 3840
rect 29352 3780 29356 3836
rect 29356 3780 29412 3836
rect 29412 3780 29416 3836
rect 29352 3776 29416 3780
rect 12216 3292 12280 3296
rect 12216 3236 12220 3292
rect 12220 3236 12276 3292
rect 12276 3236 12280 3292
rect 12216 3232 12280 3236
rect 12296 3292 12360 3296
rect 12296 3236 12300 3292
rect 12300 3236 12356 3292
rect 12356 3236 12360 3292
rect 12296 3232 12360 3236
rect 12376 3292 12440 3296
rect 12376 3236 12380 3292
rect 12380 3236 12436 3292
rect 12436 3236 12440 3292
rect 12376 3232 12440 3236
rect 12456 3292 12520 3296
rect 12456 3236 12460 3292
rect 12460 3236 12516 3292
rect 12516 3236 12520 3292
rect 12456 3232 12520 3236
rect 23480 3292 23544 3296
rect 23480 3236 23484 3292
rect 23484 3236 23540 3292
rect 23540 3236 23544 3292
rect 23480 3232 23544 3236
rect 23560 3292 23624 3296
rect 23560 3236 23564 3292
rect 23564 3236 23620 3292
rect 23620 3236 23624 3292
rect 23560 3232 23624 3236
rect 23640 3292 23704 3296
rect 23640 3236 23644 3292
rect 23644 3236 23700 3292
rect 23700 3236 23704 3292
rect 23640 3232 23704 3236
rect 23720 3292 23784 3296
rect 23720 3236 23724 3292
rect 23724 3236 23780 3292
rect 23780 3236 23784 3292
rect 23720 3232 23784 3236
rect 6584 2748 6648 2752
rect 6584 2692 6588 2748
rect 6588 2692 6644 2748
rect 6644 2692 6648 2748
rect 6584 2688 6648 2692
rect 6664 2748 6728 2752
rect 6664 2692 6668 2748
rect 6668 2692 6724 2748
rect 6724 2692 6728 2748
rect 6664 2688 6728 2692
rect 6744 2748 6808 2752
rect 6744 2692 6748 2748
rect 6748 2692 6804 2748
rect 6804 2692 6808 2748
rect 6744 2688 6808 2692
rect 6824 2748 6888 2752
rect 6824 2692 6828 2748
rect 6828 2692 6884 2748
rect 6884 2692 6888 2748
rect 6824 2688 6888 2692
rect 17848 2748 17912 2752
rect 17848 2692 17852 2748
rect 17852 2692 17908 2748
rect 17908 2692 17912 2748
rect 17848 2688 17912 2692
rect 17928 2748 17992 2752
rect 17928 2692 17932 2748
rect 17932 2692 17988 2748
rect 17988 2692 17992 2748
rect 17928 2688 17992 2692
rect 18008 2748 18072 2752
rect 18008 2692 18012 2748
rect 18012 2692 18068 2748
rect 18068 2692 18072 2748
rect 18008 2688 18072 2692
rect 18088 2748 18152 2752
rect 18088 2692 18092 2748
rect 18092 2692 18148 2748
rect 18148 2692 18152 2748
rect 18088 2688 18152 2692
rect 29112 2748 29176 2752
rect 29112 2692 29116 2748
rect 29116 2692 29172 2748
rect 29172 2692 29176 2748
rect 29112 2688 29176 2692
rect 29192 2748 29256 2752
rect 29192 2692 29196 2748
rect 29196 2692 29252 2748
rect 29252 2692 29256 2748
rect 29192 2688 29256 2692
rect 29272 2748 29336 2752
rect 29272 2692 29276 2748
rect 29276 2692 29332 2748
rect 29332 2692 29336 2748
rect 29272 2688 29336 2692
rect 29352 2748 29416 2752
rect 29352 2692 29356 2748
rect 29356 2692 29412 2748
rect 29412 2692 29416 2748
rect 29352 2688 29416 2692
rect 12216 2204 12280 2208
rect 12216 2148 12220 2204
rect 12220 2148 12276 2204
rect 12276 2148 12280 2204
rect 12216 2144 12280 2148
rect 12296 2204 12360 2208
rect 12296 2148 12300 2204
rect 12300 2148 12356 2204
rect 12356 2148 12360 2204
rect 12296 2144 12360 2148
rect 12376 2204 12440 2208
rect 12376 2148 12380 2204
rect 12380 2148 12436 2204
rect 12436 2148 12440 2204
rect 12376 2144 12440 2148
rect 12456 2204 12520 2208
rect 12456 2148 12460 2204
rect 12460 2148 12516 2204
rect 12516 2148 12520 2204
rect 12456 2144 12520 2148
rect 23480 2204 23544 2208
rect 23480 2148 23484 2204
rect 23484 2148 23540 2204
rect 23540 2148 23544 2204
rect 23480 2144 23544 2148
rect 23560 2204 23624 2208
rect 23560 2148 23564 2204
rect 23564 2148 23620 2204
rect 23620 2148 23624 2204
rect 23560 2144 23624 2148
rect 23640 2204 23704 2208
rect 23640 2148 23644 2204
rect 23644 2148 23700 2204
rect 23700 2148 23704 2204
rect 23640 2144 23704 2148
rect 23720 2204 23784 2208
rect 23720 2148 23724 2204
rect 23724 2148 23780 2204
rect 23780 2148 23784 2204
rect 23720 2144 23784 2148
<< metal4 >>
rect 14595 40900 14661 40901
rect 14595 40836 14596 40900
rect 14660 40836 14661 40900
rect 14595 40835 14661 40836
rect 12019 39812 12085 39813
rect 6576 39744 6896 39760
rect 12019 39748 12020 39812
rect 12084 39748 12085 39812
rect 12019 39747 12085 39748
rect 6576 39680 6584 39744
rect 6648 39680 6664 39744
rect 6728 39680 6744 39744
rect 6808 39680 6824 39744
rect 6888 39680 6896 39744
rect 6576 38656 6896 39680
rect 6576 38592 6584 38656
rect 6648 38592 6664 38656
rect 6728 38592 6744 38656
rect 6808 38592 6824 38656
rect 6888 38592 6896 38656
rect 6576 37568 6896 38592
rect 12022 38589 12082 39747
rect 12208 39200 12528 39760
rect 12208 39136 12216 39200
rect 12280 39136 12296 39200
rect 12360 39136 12376 39200
rect 12440 39136 12456 39200
rect 12520 39136 12528 39200
rect 12019 38588 12085 38589
rect 12019 38524 12020 38588
rect 12084 38524 12085 38588
rect 12019 38523 12085 38524
rect 6576 37504 6584 37568
rect 6648 37504 6664 37568
rect 6728 37504 6744 37568
rect 6808 37504 6824 37568
rect 6888 37504 6896 37568
rect 6576 36480 6896 37504
rect 6576 36416 6584 36480
rect 6648 36416 6664 36480
rect 6728 36416 6744 36480
rect 6808 36416 6824 36480
rect 6888 36416 6896 36480
rect 6576 35392 6896 36416
rect 6576 35328 6584 35392
rect 6648 35328 6664 35392
rect 6728 35328 6744 35392
rect 6808 35328 6824 35392
rect 6888 35328 6896 35392
rect 6576 34304 6896 35328
rect 6576 34240 6584 34304
rect 6648 34240 6664 34304
rect 6728 34240 6744 34304
rect 6808 34240 6824 34304
rect 6888 34240 6896 34304
rect 6576 33216 6896 34240
rect 6576 33152 6584 33216
rect 6648 33152 6664 33216
rect 6728 33152 6744 33216
rect 6808 33152 6824 33216
rect 6888 33152 6896 33216
rect 6576 32128 6896 33152
rect 6576 32064 6584 32128
rect 6648 32064 6664 32128
rect 6728 32064 6744 32128
rect 6808 32064 6824 32128
rect 6888 32064 6896 32128
rect 6576 31040 6896 32064
rect 6576 30976 6584 31040
rect 6648 30976 6664 31040
rect 6728 30976 6744 31040
rect 6808 30976 6824 31040
rect 6888 30976 6896 31040
rect 6576 29952 6896 30976
rect 6576 29888 6584 29952
rect 6648 29888 6664 29952
rect 6728 29888 6744 29952
rect 6808 29888 6824 29952
rect 6888 29888 6896 29952
rect 6576 28864 6896 29888
rect 6576 28800 6584 28864
rect 6648 28800 6664 28864
rect 6728 28800 6744 28864
rect 6808 28800 6824 28864
rect 6888 28800 6896 28864
rect 6576 27776 6896 28800
rect 6576 27712 6584 27776
rect 6648 27712 6664 27776
rect 6728 27712 6744 27776
rect 6808 27712 6824 27776
rect 6888 27712 6896 27776
rect 6576 26688 6896 27712
rect 6576 26624 6584 26688
rect 6648 26624 6664 26688
rect 6728 26624 6744 26688
rect 6808 26624 6824 26688
rect 6888 26624 6896 26688
rect 6576 25600 6896 26624
rect 6576 25536 6584 25600
rect 6648 25536 6664 25600
rect 6728 25536 6744 25600
rect 6808 25536 6824 25600
rect 6888 25536 6896 25600
rect 6576 24512 6896 25536
rect 6576 24448 6584 24512
rect 6648 24448 6664 24512
rect 6728 24448 6744 24512
rect 6808 24448 6824 24512
rect 6888 24448 6896 24512
rect 6576 23424 6896 24448
rect 6576 23360 6584 23424
rect 6648 23360 6664 23424
rect 6728 23360 6744 23424
rect 6808 23360 6824 23424
rect 6888 23360 6896 23424
rect 6576 22336 6896 23360
rect 6576 22272 6584 22336
rect 6648 22272 6664 22336
rect 6728 22272 6744 22336
rect 6808 22272 6824 22336
rect 6888 22272 6896 22336
rect 6576 21248 6896 22272
rect 6576 21184 6584 21248
rect 6648 21184 6664 21248
rect 6728 21184 6744 21248
rect 6808 21184 6824 21248
rect 6888 21184 6896 21248
rect 6576 20160 6896 21184
rect 6576 20096 6584 20160
rect 6648 20096 6664 20160
rect 6728 20096 6744 20160
rect 6808 20096 6824 20160
rect 6888 20096 6896 20160
rect 6576 19072 6896 20096
rect 6576 19008 6584 19072
rect 6648 19008 6664 19072
rect 6728 19008 6744 19072
rect 6808 19008 6824 19072
rect 6888 19008 6896 19072
rect 6576 17984 6896 19008
rect 6576 17920 6584 17984
rect 6648 17920 6664 17984
rect 6728 17920 6744 17984
rect 6808 17920 6824 17984
rect 6888 17920 6896 17984
rect 6576 16896 6896 17920
rect 6576 16832 6584 16896
rect 6648 16832 6664 16896
rect 6728 16832 6744 16896
rect 6808 16832 6824 16896
rect 6888 16832 6896 16896
rect 6576 15808 6896 16832
rect 6576 15744 6584 15808
rect 6648 15744 6664 15808
rect 6728 15744 6744 15808
rect 6808 15744 6824 15808
rect 6888 15744 6896 15808
rect 6576 14720 6896 15744
rect 6576 14656 6584 14720
rect 6648 14656 6664 14720
rect 6728 14656 6744 14720
rect 6808 14656 6824 14720
rect 6888 14656 6896 14720
rect 6576 13632 6896 14656
rect 6576 13568 6584 13632
rect 6648 13568 6664 13632
rect 6728 13568 6744 13632
rect 6808 13568 6824 13632
rect 6888 13568 6896 13632
rect 6576 12544 6896 13568
rect 6576 12480 6584 12544
rect 6648 12480 6664 12544
rect 6728 12480 6744 12544
rect 6808 12480 6824 12544
rect 6888 12480 6896 12544
rect 6576 11456 6896 12480
rect 6576 11392 6584 11456
rect 6648 11392 6664 11456
rect 6728 11392 6744 11456
rect 6808 11392 6824 11456
rect 6888 11392 6896 11456
rect 6576 10368 6896 11392
rect 6576 10304 6584 10368
rect 6648 10304 6664 10368
rect 6728 10304 6744 10368
rect 6808 10304 6824 10368
rect 6888 10304 6896 10368
rect 6576 9280 6896 10304
rect 6576 9216 6584 9280
rect 6648 9216 6664 9280
rect 6728 9216 6744 9280
rect 6808 9216 6824 9280
rect 6888 9216 6896 9280
rect 6576 8192 6896 9216
rect 6576 8128 6584 8192
rect 6648 8128 6664 8192
rect 6728 8128 6744 8192
rect 6808 8128 6824 8192
rect 6888 8128 6896 8192
rect 6576 7104 6896 8128
rect 6576 7040 6584 7104
rect 6648 7040 6664 7104
rect 6728 7040 6744 7104
rect 6808 7040 6824 7104
rect 6888 7040 6896 7104
rect 6576 6016 6896 7040
rect 6576 5952 6584 6016
rect 6648 5952 6664 6016
rect 6728 5952 6744 6016
rect 6808 5952 6824 6016
rect 6888 5952 6896 6016
rect 6576 4928 6896 5952
rect 6576 4864 6584 4928
rect 6648 4864 6664 4928
rect 6728 4864 6744 4928
rect 6808 4864 6824 4928
rect 6888 4864 6896 4928
rect 6576 3840 6896 4864
rect 6576 3776 6584 3840
rect 6648 3776 6664 3840
rect 6728 3776 6744 3840
rect 6808 3776 6824 3840
rect 6888 3776 6896 3840
rect 6576 2752 6896 3776
rect 6576 2688 6584 2752
rect 6648 2688 6664 2752
rect 6728 2688 6744 2752
rect 6808 2688 6824 2752
rect 6888 2688 6896 2752
rect 6576 2128 6896 2688
rect 12208 38112 12528 39136
rect 12755 38860 12821 38861
rect 12755 38796 12756 38860
rect 12820 38796 12821 38860
rect 12755 38795 12821 38796
rect 12208 38048 12216 38112
rect 12280 38048 12296 38112
rect 12360 38048 12376 38112
rect 12440 38048 12456 38112
rect 12520 38048 12528 38112
rect 12208 37024 12528 38048
rect 12208 36960 12216 37024
rect 12280 36960 12296 37024
rect 12360 36960 12376 37024
rect 12440 36960 12456 37024
rect 12520 36960 12528 37024
rect 12208 35936 12528 36960
rect 12208 35872 12216 35936
rect 12280 35872 12296 35936
rect 12360 35872 12376 35936
rect 12440 35872 12456 35936
rect 12520 35872 12528 35936
rect 12208 34848 12528 35872
rect 12208 34784 12216 34848
rect 12280 34784 12296 34848
rect 12360 34784 12376 34848
rect 12440 34784 12456 34848
rect 12520 34784 12528 34848
rect 12208 33760 12528 34784
rect 12758 34781 12818 38795
rect 14227 35052 14293 35053
rect 14227 34988 14228 35052
rect 14292 34988 14293 35052
rect 14227 34987 14293 34988
rect 12755 34780 12821 34781
rect 12755 34716 12756 34780
rect 12820 34716 12821 34780
rect 12755 34715 12821 34716
rect 14230 34101 14290 34987
rect 14598 34645 14658 40835
rect 18459 40492 18525 40493
rect 18459 40428 18460 40492
rect 18524 40428 18525 40492
rect 18459 40427 18525 40428
rect 17840 39744 18160 39760
rect 17840 39680 17848 39744
rect 17912 39680 17928 39744
rect 17992 39680 18008 39744
rect 18072 39680 18088 39744
rect 18152 39680 18160 39744
rect 17840 38656 18160 39680
rect 18462 39133 18522 40427
rect 23472 39200 23792 39760
rect 23472 39136 23480 39200
rect 23544 39136 23560 39200
rect 23624 39136 23640 39200
rect 23704 39136 23720 39200
rect 23784 39136 23792 39200
rect 18459 39132 18525 39133
rect 18459 39068 18460 39132
rect 18524 39068 18525 39132
rect 18459 39067 18525 39068
rect 17840 38592 17848 38656
rect 17912 38592 17928 38656
rect 17992 38592 18008 38656
rect 18072 38592 18088 38656
rect 18152 38592 18160 38656
rect 17840 37568 18160 38592
rect 17840 37504 17848 37568
rect 17912 37504 17928 37568
rect 17992 37504 18008 37568
rect 18072 37504 18088 37568
rect 18152 37504 18160 37568
rect 17539 37500 17605 37501
rect 17539 37436 17540 37500
rect 17604 37436 17605 37500
rect 17539 37435 17605 37436
rect 17355 35596 17421 35597
rect 17355 35532 17356 35596
rect 17420 35532 17421 35596
rect 17355 35531 17421 35532
rect 17358 35325 17418 35531
rect 17355 35324 17421 35325
rect 17355 35260 17356 35324
rect 17420 35260 17421 35324
rect 17355 35259 17421 35260
rect 15331 35052 15397 35053
rect 15331 34988 15332 35052
rect 15396 34988 15397 35052
rect 15331 34987 15397 34988
rect 14595 34644 14661 34645
rect 14595 34580 14596 34644
rect 14660 34580 14661 34644
rect 14595 34579 14661 34580
rect 14227 34100 14293 34101
rect 14227 34036 14228 34100
rect 14292 34036 14293 34100
rect 14227 34035 14293 34036
rect 14595 34100 14661 34101
rect 14595 34036 14596 34100
rect 14660 34036 14661 34100
rect 14595 34035 14661 34036
rect 12208 33696 12216 33760
rect 12280 33696 12296 33760
rect 12360 33696 12376 33760
rect 12440 33696 12456 33760
rect 12520 33696 12528 33760
rect 12208 32672 12528 33696
rect 12208 32608 12216 32672
rect 12280 32608 12296 32672
rect 12360 32608 12376 32672
rect 12440 32608 12456 32672
rect 12520 32608 12528 32672
rect 12208 31584 12528 32608
rect 12208 31520 12216 31584
rect 12280 31520 12296 31584
rect 12360 31520 12376 31584
rect 12440 31520 12456 31584
rect 12520 31520 12528 31584
rect 12208 30496 12528 31520
rect 12208 30432 12216 30496
rect 12280 30432 12296 30496
rect 12360 30432 12376 30496
rect 12440 30432 12456 30496
rect 12520 30432 12528 30496
rect 12208 29408 12528 30432
rect 12208 29344 12216 29408
rect 12280 29344 12296 29408
rect 12360 29344 12376 29408
rect 12440 29344 12456 29408
rect 12520 29344 12528 29408
rect 12208 28320 12528 29344
rect 14230 28389 14290 34035
rect 14598 33690 14658 34035
rect 15334 33826 15394 34987
rect 17542 34098 17602 37435
rect 16438 34038 17602 34098
rect 17840 36480 18160 37504
rect 17840 36416 17848 36480
rect 17912 36416 17928 36480
rect 17992 36416 18008 36480
rect 18072 36416 18088 36480
rect 18152 36416 18160 36480
rect 17840 35392 18160 36416
rect 17840 35328 17848 35392
rect 17912 35328 17928 35392
rect 17992 35328 18008 35392
rect 18072 35328 18088 35392
rect 18152 35328 18160 35392
rect 17840 34304 18160 35328
rect 17840 34240 17848 34304
rect 17912 34240 17928 34304
rect 17992 34240 18008 34304
rect 18072 34240 18088 34304
rect 18152 34240 18160 34304
rect 15883 33964 15949 33965
rect 15883 33900 15884 33964
rect 15948 33962 15949 33964
rect 16438 33962 16498 34038
rect 15948 33902 16498 33962
rect 15948 33900 15949 33902
rect 15883 33899 15949 33900
rect 15334 33766 16498 33826
rect 14598 33630 15946 33690
rect 15886 33557 15946 33630
rect 15883 33556 15949 33557
rect 15883 33492 15884 33556
rect 15948 33492 15949 33556
rect 15883 33491 15949 33492
rect 16438 33149 16498 33766
rect 17840 33216 18160 34240
rect 23472 38112 23792 39136
rect 23472 38048 23480 38112
rect 23544 38048 23560 38112
rect 23624 38048 23640 38112
rect 23704 38048 23720 38112
rect 23784 38048 23792 38112
rect 23472 37024 23792 38048
rect 23472 36960 23480 37024
rect 23544 36960 23560 37024
rect 23624 36960 23640 37024
rect 23704 36960 23720 37024
rect 23784 36960 23792 37024
rect 23472 35936 23792 36960
rect 23472 35872 23480 35936
rect 23544 35872 23560 35936
rect 23624 35872 23640 35936
rect 23704 35872 23720 35936
rect 23784 35872 23792 35936
rect 23472 34848 23792 35872
rect 23472 34784 23480 34848
rect 23544 34784 23560 34848
rect 23624 34784 23640 34848
rect 23704 34784 23720 34848
rect 23784 34784 23792 34848
rect 18459 34236 18525 34237
rect 18459 34234 18460 34236
rect 18278 34174 18460 34234
rect 18278 33421 18338 34174
rect 18459 34172 18460 34174
rect 18524 34172 18525 34236
rect 18459 34171 18525 34172
rect 20851 33828 20917 33829
rect 20851 33764 20852 33828
rect 20916 33764 20917 33828
rect 20851 33763 20917 33764
rect 18459 33692 18525 33693
rect 18459 33628 18460 33692
rect 18524 33628 18525 33692
rect 18459 33627 18525 33628
rect 18462 33421 18522 33627
rect 18275 33420 18341 33421
rect 18275 33356 18276 33420
rect 18340 33356 18341 33420
rect 18275 33355 18341 33356
rect 18459 33420 18525 33421
rect 18459 33356 18460 33420
rect 18524 33356 18525 33420
rect 18459 33355 18525 33356
rect 18275 33284 18341 33285
rect 18275 33220 18276 33284
rect 18340 33220 18341 33284
rect 18275 33219 18341 33220
rect 17840 33152 17848 33216
rect 17912 33152 17928 33216
rect 17992 33152 18008 33216
rect 18072 33152 18088 33216
rect 18152 33152 18160 33216
rect 16435 33148 16501 33149
rect 16435 33084 16436 33148
rect 16500 33084 16501 33148
rect 16435 33083 16501 33084
rect 16067 33012 16133 33013
rect 16067 32948 16068 33012
rect 16132 33010 16133 33012
rect 16132 32950 17602 33010
rect 16132 32948 16133 32950
rect 16067 32947 16133 32948
rect 17542 32741 17602 32950
rect 17539 32740 17605 32741
rect 17539 32676 17540 32740
rect 17604 32676 17605 32740
rect 17539 32675 17605 32676
rect 14779 32196 14845 32197
rect 14779 32132 14780 32196
rect 14844 32194 14845 32196
rect 17355 32196 17421 32197
rect 14844 32134 16498 32194
rect 14844 32132 14845 32134
rect 14779 32131 14845 32132
rect 16438 31789 16498 32134
rect 17355 32132 17356 32196
rect 17420 32132 17421 32196
rect 17355 32131 17421 32132
rect 16251 31788 16317 31789
rect 16251 31724 16252 31788
rect 16316 31724 16317 31788
rect 16251 31723 16317 31724
rect 16435 31788 16501 31789
rect 16435 31724 16436 31788
rect 16500 31724 16501 31788
rect 16435 31723 16501 31724
rect 16254 31650 16314 31723
rect 17358 31650 17418 32131
rect 16254 31590 17418 31650
rect 17840 32128 18160 33152
rect 18278 32741 18338 33219
rect 18275 32740 18341 32741
rect 18275 32676 18276 32740
rect 18340 32676 18341 32740
rect 18275 32675 18341 32676
rect 18459 32468 18525 32469
rect 18459 32404 18460 32468
rect 18524 32404 18525 32468
rect 18459 32403 18525 32404
rect 18643 32468 18709 32469
rect 18643 32404 18644 32468
rect 18708 32404 18709 32468
rect 18643 32403 18709 32404
rect 18462 32197 18522 32403
rect 18275 32196 18341 32197
rect 18275 32132 18276 32196
rect 18340 32194 18341 32196
rect 18459 32196 18525 32197
rect 18340 32132 18384 32194
rect 18275 32131 18384 32132
rect 18459 32132 18460 32196
rect 18524 32132 18525 32196
rect 18459 32131 18525 32132
rect 17840 32064 17848 32128
rect 17912 32064 17928 32128
rect 17992 32064 18008 32128
rect 18072 32064 18088 32128
rect 18152 32064 18160 32128
rect 17539 31108 17605 31109
rect 17539 31044 17540 31108
rect 17604 31044 17605 31108
rect 17539 31043 17605 31044
rect 17542 29885 17602 31043
rect 17840 31040 18160 32064
rect 18324 32058 18384 32131
rect 18646 32058 18706 32403
rect 18324 31998 18706 32058
rect 18827 32060 18893 32061
rect 18827 31996 18828 32060
rect 18892 31996 18893 32060
rect 18827 31995 18893 31996
rect 17840 30976 17848 31040
rect 17912 30976 17928 31040
rect 17992 30976 18008 31040
rect 18072 30976 18088 31040
rect 18152 30976 18160 31040
rect 17840 29952 18160 30976
rect 18459 30972 18525 30973
rect 18459 30908 18460 30972
rect 18524 30908 18525 30972
rect 18459 30907 18525 30908
rect 18643 30972 18709 30973
rect 18643 30908 18644 30972
rect 18708 30908 18709 30972
rect 18643 30907 18709 30908
rect 18462 30021 18522 30907
rect 18459 30020 18525 30021
rect 18459 29956 18460 30020
rect 18524 29956 18525 30020
rect 18459 29955 18525 29956
rect 17840 29888 17848 29952
rect 17912 29888 17928 29952
rect 17992 29888 18008 29952
rect 18072 29888 18088 29952
rect 18152 29888 18160 29952
rect 17539 29884 17605 29885
rect 17539 29820 17540 29884
rect 17604 29820 17605 29884
rect 17539 29819 17605 29820
rect 17840 28864 18160 29888
rect 18275 29884 18341 29885
rect 18275 29820 18276 29884
rect 18340 29882 18341 29884
rect 18646 29882 18706 30907
rect 18830 30429 18890 31995
rect 18827 30428 18893 30429
rect 18827 30364 18828 30428
rect 18892 30364 18893 30428
rect 18827 30363 18893 30364
rect 18340 29822 18706 29882
rect 18340 29820 18341 29822
rect 18275 29819 18341 29820
rect 20854 29069 20914 33763
rect 23472 33760 23792 34784
rect 23472 33696 23480 33760
rect 23544 33696 23560 33760
rect 23624 33696 23640 33760
rect 23704 33696 23720 33760
rect 23784 33696 23792 33760
rect 23472 32672 23792 33696
rect 23472 32608 23480 32672
rect 23544 32608 23560 32672
rect 23624 32608 23640 32672
rect 23704 32608 23720 32672
rect 23784 32608 23792 32672
rect 23472 31584 23792 32608
rect 23472 31520 23480 31584
rect 23544 31520 23560 31584
rect 23624 31520 23640 31584
rect 23704 31520 23720 31584
rect 23784 31520 23792 31584
rect 21771 31108 21837 31109
rect 21771 31044 21772 31108
rect 21836 31044 21837 31108
rect 21771 31043 21837 31044
rect 23059 31108 23125 31109
rect 23059 31044 23060 31108
rect 23124 31044 23125 31108
rect 23059 31043 23125 31044
rect 21219 30836 21285 30837
rect 21219 30772 21220 30836
rect 21284 30834 21285 30836
rect 21774 30834 21834 31043
rect 21284 30774 21834 30834
rect 21284 30772 21285 30774
rect 21219 30771 21285 30772
rect 21219 30700 21285 30701
rect 21219 30636 21220 30700
rect 21284 30636 21285 30700
rect 21219 30635 21285 30636
rect 21222 30290 21282 30635
rect 23062 30565 23122 31043
rect 23059 30564 23125 30565
rect 23059 30500 23060 30564
rect 23124 30500 23125 30564
rect 23059 30499 23125 30500
rect 23472 30496 23792 31520
rect 29104 39744 29424 39760
rect 29104 39680 29112 39744
rect 29176 39680 29192 39744
rect 29256 39680 29272 39744
rect 29336 39680 29352 39744
rect 29416 39680 29424 39744
rect 29104 38656 29424 39680
rect 29104 38592 29112 38656
rect 29176 38592 29192 38656
rect 29256 38592 29272 38656
rect 29336 38592 29352 38656
rect 29416 38592 29424 38656
rect 29104 37568 29424 38592
rect 29104 37504 29112 37568
rect 29176 37504 29192 37568
rect 29256 37504 29272 37568
rect 29336 37504 29352 37568
rect 29416 37504 29424 37568
rect 29104 36480 29424 37504
rect 29104 36416 29112 36480
rect 29176 36416 29192 36480
rect 29256 36416 29272 36480
rect 29336 36416 29352 36480
rect 29416 36416 29424 36480
rect 29104 35392 29424 36416
rect 29104 35328 29112 35392
rect 29176 35328 29192 35392
rect 29256 35328 29272 35392
rect 29336 35328 29352 35392
rect 29416 35328 29424 35392
rect 29104 34304 29424 35328
rect 31523 35188 31589 35189
rect 31523 35124 31524 35188
rect 31588 35124 31589 35188
rect 31523 35123 31589 35124
rect 29104 34240 29112 34304
rect 29176 34240 29192 34304
rect 29256 34240 29272 34304
rect 29336 34240 29352 34304
rect 29416 34240 29424 34304
rect 29104 33216 29424 34240
rect 31526 33421 31586 35123
rect 31523 33420 31589 33421
rect 31523 33356 31524 33420
rect 31588 33356 31589 33420
rect 31523 33355 31589 33356
rect 29104 33152 29112 33216
rect 29176 33152 29192 33216
rect 29256 33152 29272 33216
rect 29336 33152 29352 33216
rect 29416 33152 29424 33216
rect 29104 32128 29424 33152
rect 30419 32196 30485 32197
rect 30419 32132 30420 32196
rect 30484 32132 30485 32196
rect 30419 32131 30485 32132
rect 30787 32196 30853 32197
rect 30787 32132 30788 32196
rect 30852 32132 30853 32196
rect 30787 32131 30853 32132
rect 29104 32064 29112 32128
rect 29176 32064 29192 32128
rect 29256 32064 29272 32128
rect 29336 32064 29352 32128
rect 29416 32064 29424 32128
rect 27659 31108 27725 31109
rect 27659 31044 27660 31108
rect 27724 31044 27725 31108
rect 27659 31043 27725 31044
rect 23472 30432 23480 30496
rect 23544 30432 23560 30496
rect 23624 30432 23640 30496
rect 23704 30432 23720 30496
rect 23784 30432 23792 30496
rect 21222 30230 22754 30290
rect 22694 30021 22754 30230
rect 22691 30020 22757 30021
rect 22691 29956 22692 30020
rect 22756 29956 22757 30020
rect 22691 29955 22757 29956
rect 23243 29884 23309 29885
rect 23243 29820 23244 29884
rect 23308 29820 23309 29884
rect 23243 29819 23309 29820
rect 23246 29477 23306 29819
rect 23243 29476 23309 29477
rect 23243 29412 23244 29476
rect 23308 29412 23309 29476
rect 23243 29411 23309 29412
rect 23472 29408 23792 30432
rect 23472 29344 23480 29408
rect 23544 29344 23560 29408
rect 23624 29344 23640 29408
rect 23704 29344 23720 29408
rect 23784 29344 23792 29408
rect 20851 29068 20917 29069
rect 20851 29004 20852 29068
rect 20916 29004 20917 29068
rect 20851 29003 20917 29004
rect 17840 28800 17848 28864
rect 17912 28800 17928 28864
rect 17992 28800 18008 28864
rect 18072 28800 18088 28864
rect 18152 28800 18160 28864
rect 16803 28660 16869 28661
rect 16803 28596 16804 28660
rect 16868 28596 16869 28660
rect 16803 28595 16869 28596
rect 14227 28388 14293 28389
rect 14227 28324 14228 28388
rect 14292 28324 14293 28388
rect 16806 28386 16866 28595
rect 14227 28323 14293 28324
rect 15334 28326 16866 28386
rect 12208 28256 12216 28320
rect 12280 28256 12296 28320
rect 12360 28256 12376 28320
rect 12440 28256 12456 28320
rect 12520 28256 12528 28320
rect 12208 27232 12528 28256
rect 15334 27981 15394 28326
rect 15331 27980 15397 27981
rect 15331 27916 15332 27980
rect 15396 27916 15397 27980
rect 15331 27915 15397 27916
rect 17840 27776 18160 28800
rect 17840 27712 17848 27776
rect 17912 27712 17928 27776
rect 17992 27712 18008 27776
rect 18072 27712 18088 27776
rect 18152 27712 18160 27776
rect 16067 27572 16133 27573
rect 16067 27508 16068 27572
rect 16132 27570 16133 27572
rect 16132 27510 16682 27570
rect 16132 27508 16133 27510
rect 16067 27507 16133 27508
rect 16622 27301 16682 27510
rect 16619 27300 16685 27301
rect 16619 27236 16620 27300
rect 16684 27236 16685 27300
rect 16619 27235 16685 27236
rect 12208 27168 12216 27232
rect 12280 27168 12296 27232
rect 12360 27168 12376 27232
rect 12440 27168 12456 27232
rect 12520 27168 12528 27232
rect 12208 26144 12528 27168
rect 12208 26080 12216 26144
rect 12280 26080 12296 26144
rect 12360 26080 12376 26144
rect 12440 26080 12456 26144
rect 12520 26080 12528 26144
rect 12208 25056 12528 26080
rect 12208 24992 12216 25056
rect 12280 24992 12296 25056
rect 12360 24992 12376 25056
rect 12440 24992 12456 25056
rect 12520 24992 12528 25056
rect 12208 23968 12528 24992
rect 12208 23904 12216 23968
rect 12280 23904 12296 23968
rect 12360 23904 12376 23968
rect 12440 23904 12456 23968
rect 12520 23904 12528 23968
rect 12208 22880 12528 23904
rect 12208 22816 12216 22880
rect 12280 22816 12296 22880
rect 12360 22816 12376 22880
rect 12440 22816 12456 22880
rect 12520 22816 12528 22880
rect 12208 21792 12528 22816
rect 12208 21728 12216 21792
rect 12280 21728 12296 21792
rect 12360 21728 12376 21792
rect 12440 21728 12456 21792
rect 12520 21728 12528 21792
rect 12208 20704 12528 21728
rect 12208 20640 12216 20704
rect 12280 20640 12296 20704
rect 12360 20640 12376 20704
rect 12440 20640 12456 20704
rect 12520 20640 12528 20704
rect 12208 19616 12528 20640
rect 12208 19552 12216 19616
rect 12280 19552 12296 19616
rect 12360 19552 12376 19616
rect 12440 19552 12456 19616
rect 12520 19552 12528 19616
rect 12208 18528 12528 19552
rect 12208 18464 12216 18528
rect 12280 18464 12296 18528
rect 12360 18464 12376 18528
rect 12440 18464 12456 18528
rect 12520 18464 12528 18528
rect 12208 17440 12528 18464
rect 12208 17376 12216 17440
rect 12280 17376 12296 17440
rect 12360 17376 12376 17440
rect 12440 17376 12456 17440
rect 12520 17376 12528 17440
rect 12208 16352 12528 17376
rect 12208 16288 12216 16352
rect 12280 16288 12296 16352
rect 12360 16288 12376 16352
rect 12440 16288 12456 16352
rect 12520 16288 12528 16352
rect 12208 15264 12528 16288
rect 12208 15200 12216 15264
rect 12280 15200 12296 15264
rect 12360 15200 12376 15264
rect 12440 15200 12456 15264
rect 12520 15200 12528 15264
rect 12208 14176 12528 15200
rect 12208 14112 12216 14176
rect 12280 14112 12296 14176
rect 12360 14112 12376 14176
rect 12440 14112 12456 14176
rect 12520 14112 12528 14176
rect 12208 13088 12528 14112
rect 12208 13024 12216 13088
rect 12280 13024 12296 13088
rect 12360 13024 12376 13088
rect 12440 13024 12456 13088
rect 12520 13024 12528 13088
rect 12208 12000 12528 13024
rect 12208 11936 12216 12000
rect 12280 11936 12296 12000
rect 12360 11936 12376 12000
rect 12440 11936 12456 12000
rect 12520 11936 12528 12000
rect 12208 10912 12528 11936
rect 12208 10848 12216 10912
rect 12280 10848 12296 10912
rect 12360 10848 12376 10912
rect 12440 10848 12456 10912
rect 12520 10848 12528 10912
rect 12208 9824 12528 10848
rect 12208 9760 12216 9824
rect 12280 9760 12296 9824
rect 12360 9760 12376 9824
rect 12440 9760 12456 9824
rect 12520 9760 12528 9824
rect 12208 8736 12528 9760
rect 12208 8672 12216 8736
rect 12280 8672 12296 8736
rect 12360 8672 12376 8736
rect 12440 8672 12456 8736
rect 12520 8672 12528 8736
rect 12208 7648 12528 8672
rect 12208 7584 12216 7648
rect 12280 7584 12296 7648
rect 12360 7584 12376 7648
rect 12440 7584 12456 7648
rect 12520 7584 12528 7648
rect 12208 6560 12528 7584
rect 12208 6496 12216 6560
rect 12280 6496 12296 6560
rect 12360 6496 12376 6560
rect 12440 6496 12456 6560
rect 12520 6496 12528 6560
rect 12208 5472 12528 6496
rect 12208 5408 12216 5472
rect 12280 5408 12296 5472
rect 12360 5408 12376 5472
rect 12440 5408 12456 5472
rect 12520 5408 12528 5472
rect 12208 4384 12528 5408
rect 12208 4320 12216 4384
rect 12280 4320 12296 4384
rect 12360 4320 12376 4384
rect 12440 4320 12456 4384
rect 12520 4320 12528 4384
rect 12208 3296 12528 4320
rect 12208 3232 12216 3296
rect 12280 3232 12296 3296
rect 12360 3232 12376 3296
rect 12440 3232 12456 3296
rect 12520 3232 12528 3296
rect 12208 2208 12528 3232
rect 12208 2144 12216 2208
rect 12280 2144 12296 2208
rect 12360 2144 12376 2208
rect 12440 2144 12456 2208
rect 12520 2144 12528 2208
rect 12208 2128 12528 2144
rect 17840 26688 18160 27712
rect 17840 26624 17848 26688
rect 17912 26624 17928 26688
rect 17992 26624 18008 26688
rect 18072 26624 18088 26688
rect 18152 26624 18160 26688
rect 17840 25600 18160 26624
rect 17840 25536 17848 25600
rect 17912 25536 17928 25600
rect 17992 25536 18008 25600
rect 18072 25536 18088 25600
rect 18152 25536 18160 25600
rect 17840 24512 18160 25536
rect 17840 24448 17848 24512
rect 17912 24448 17928 24512
rect 17992 24448 18008 24512
rect 18072 24448 18088 24512
rect 18152 24448 18160 24512
rect 17840 23424 18160 24448
rect 17840 23360 17848 23424
rect 17912 23360 17928 23424
rect 17992 23360 18008 23424
rect 18072 23360 18088 23424
rect 18152 23360 18160 23424
rect 17840 22336 18160 23360
rect 17840 22272 17848 22336
rect 17912 22272 17928 22336
rect 17992 22272 18008 22336
rect 18072 22272 18088 22336
rect 18152 22272 18160 22336
rect 17840 21248 18160 22272
rect 17840 21184 17848 21248
rect 17912 21184 17928 21248
rect 17992 21184 18008 21248
rect 18072 21184 18088 21248
rect 18152 21184 18160 21248
rect 17840 20160 18160 21184
rect 17840 20096 17848 20160
rect 17912 20096 17928 20160
rect 17992 20096 18008 20160
rect 18072 20096 18088 20160
rect 18152 20096 18160 20160
rect 17840 19072 18160 20096
rect 17840 19008 17848 19072
rect 17912 19008 17928 19072
rect 17992 19008 18008 19072
rect 18072 19008 18088 19072
rect 18152 19008 18160 19072
rect 17840 17984 18160 19008
rect 17840 17920 17848 17984
rect 17912 17920 17928 17984
rect 17992 17920 18008 17984
rect 18072 17920 18088 17984
rect 18152 17920 18160 17984
rect 17840 16896 18160 17920
rect 17840 16832 17848 16896
rect 17912 16832 17928 16896
rect 17992 16832 18008 16896
rect 18072 16832 18088 16896
rect 18152 16832 18160 16896
rect 17840 15808 18160 16832
rect 17840 15744 17848 15808
rect 17912 15744 17928 15808
rect 17992 15744 18008 15808
rect 18072 15744 18088 15808
rect 18152 15744 18160 15808
rect 17840 14720 18160 15744
rect 17840 14656 17848 14720
rect 17912 14656 17928 14720
rect 17992 14656 18008 14720
rect 18072 14656 18088 14720
rect 18152 14656 18160 14720
rect 17840 13632 18160 14656
rect 17840 13568 17848 13632
rect 17912 13568 17928 13632
rect 17992 13568 18008 13632
rect 18072 13568 18088 13632
rect 18152 13568 18160 13632
rect 17840 12544 18160 13568
rect 17840 12480 17848 12544
rect 17912 12480 17928 12544
rect 17992 12480 18008 12544
rect 18072 12480 18088 12544
rect 18152 12480 18160 12544
rect 17840 11456 18160 12480
rect 17840 11392 17848 11456
rect 17912 11392 17928 11456
rect 17992 11392 18008 11456
rect 18072 11392 18088 11456
rect 18152 11392 18160 11456
rect 17840 10368 18160 11392
rect 17840 10304 17848 10368
rect 17912 10304 17928 10368
rect 17992 10304 18008 10368
rect 18072 10304 18088 10368
rect 18152 10304 18160 10368
rect 17840 9280 18160 10304
rect 17840 9216 17848 9280
rect 17912 9216 17928 9280
rect 17992 9216 18008 9280
rect 18072 9216 18088 9280
rect 18152 9216 18160 9280
rect 17840 8192 18160 9216
rect 17840 8128 17848 8192
rect 17912 8128 17928 8192
rect 17992 8128 18008 8192
rect 18072 8128 18088 8192
rect 18152 8128 18160 8192
rect 17840 7104 18160 8128
rect 17840 7040 17848 7104
rect 17912 7040 17928 7104
rect 17992 7040 18008 7104
rect 18072 7040 18088 7104
rect 18152 7040 18160 7104
rect 17840 6016 18160 7040
rect 17840 5952 17848 6016
rect 17912 5952 17928 6016
rect 17992 5952 18008 6016
rect 18072 5952 18088 6016
rect 18152 5952 18160 6016
rect 17840 4928 18160 5952
rect 17840 4864 17848 4928
rect 17912 4864 17928 4928
rect 17992 4864 18008 4928
rect 18072 4864 18088 4928
rect 18152 4864 18160 4928
rect 17840 3840 18160 4864
rect 17840 3776 17848 3840
rect 17912 3776 17928 3840
rect 17992 3776 18008 3840
rect 18072 3776 18088 3840
rect 18152 3776 18160 3840
rect 17840 2752 18160 3776
rect 17840 2688 17848 2752
rect 17912 2688 17928 2752
rect 17992 2688 18008 2752
rect 18072 2688 18088 2752
rect 18152 2688 18160 2752
rect 17840 2128 18160 2688
rect 23472 28320 23792 29344
rect 23472 28256 23480 28320
rect 23544 28256 23560 28320
rect 23624 28256 23640 28320
rect 23704 28256 23720 28320
rect 23784 28256 23792 28320
rect 23472 27232 23792 28256
rect 23472 27168 23480 27232
rect 23544 27168 23560 27232
rect 23624 27168 23640 27232
rect 23704 27168 23720 27232
rect 23784 27168 23792 27232
rect 23472 26144 23792 27168
rect 23472 26080 23480 26144
rect 23544 26080 23560 26144
rect 23624 26080 23640 26144
rect 23704 26080 23720 26144
rect 23784 26080 23792 26144
rect 23472 25056 23792 26080
rect 23472 24992 23480 25056
rect 23544 24992 23560 25056
rect 23624 24992 23640 25056
rect 23704 24992 23720 25056
rect 23784 24992 23792 25056
rect 23472 23968 23792 24992
rect 27662 24853 27722 31043
rect 29104 31040 29424 32064
rect 29104 30976 29112 31040
rect 29176 30976 29192 31040
rect 29256 30976 29272 31040
rect 29336 30976 29352 31040
rect 29416 30976 29424 31040
rect 28579 30700 28645 30701
rect 28579 30636 28580 30700
rect 28644 30636 28645 30700
rect 28579 30635 28645 30636
rect 28582 29885 28642 30635
rect 29104 29952 29424 30976
rect 30422 30565 30482 32131
rect 30419 30564 30485 30565
rect 30419 30500 30420 30564
rect 30484 30500 30485 30564
rect 30419 30499 30485 30500
rect 29104 29888 29112 29952
rect 29176 29888 29192 29952
rect 29256 29888 29272 29952
rect 29336 29888 29352 29952
rect 29416 29888 29424 29952
rect 28579 29884 28645 29885
rect 28579 29820 28580 29884
rect 28644 29820 28645 29884
rect 28579 29819 28645 29820
rect 29104 28864 29424 29888
rect 30790 29885 30850 32131
rect 30787 29884 30853 29885
rect 30787 29820 30788 29884
rect 30852 29820 30853 29884
rect 30787 29819 30853 29820
rect 29867 28932 29933 28933
rect 29867 28868 29868 28932
rect 29932 28868 29933 28932
rect 29867 28867 29933 28868
rect 29104 28800 29112 28864
rect 29176 28800 29192 28864
rect 29256 28800 29272 28864
rect 29336 28800 29352 28864
rect 29416 28800 29424 28864
rect 29104 27776 29424 28800
rect 29104 27712 29112 27776
rect 29176 27712 29192 27776
rect 29256 27712 29272 27776
rect 29336 27712 29352 27776
rect 29416 27712 29424 27776
rect 29104 26688 29424 27712
rect 29499 26892 29565 26893
rect 29499 26828 29500 26892
rect 29564 26828 29565 26892
rect 29499 26827 29565 26828
rect 29104 26624 29112 26688
rect 29176 26624 29192 26688
rect 29256 26624 29272 26688
rect 29336 26624 29352 26688
rect 29416 26624 29424 26688
rect 29104 25600 29424 26624
rect 29104 25536 29112 25600
rect 29176 25536 29192 25600
rect 29256 25536 29272 25600
rect 29336 25536 29352 25600
rect 29416 25536 29424 25600
rect 27659 24852 27725 24853
rect 27659 24788 27660 24852
rect 27724 24788 27725 24852
rect 27659 24787 27725 24788
rect 23472 23904 23480 23968
rect 23544 23904 23560 23968
rect 23624 23904 23640 23968
rect 23704 23904 23720 23968
rect 23784 23904 23792 23968
rect 23472 22880 23792 23904
rect 23472 22816 23480 22880
rect 23544 22816 23560 22880
rect 23624 22816 23640 22880
rect 23704 22816 23720 22880
rect 23784 22816 23792 22880
rect 23472 21792 23792 22816
rect 29104 24512 29424 25536
rect 29104 24448 29112 24512
rect 29176 24448 29192 24512
rect 29256 24448 29272 24512
rect 29336 24448 29352 24512
rect 29416 24448 29424 24512
rect 29104 23424 29424 24448
rect 29104 23360 29112 23424
rect 29176 23360 29192 23424
rect 29256 23360 29272 23424
rect 29336 23360 29352 23424
rect 29416 23360 29424 23424
rect 29104 22336 29424 23360
rect 29104 22272 29112 22336
rect 29176 22272 29192 22336
rect 29256 22272 29272 22336
rect 29336 22272 29352 22336
rect 29416 22272 29424 22336
rect 25267 22132 25333 22133
rect 25267 22068 25268 22132
rect 25332 22068 25333 22132
rect 25267 22067 25333 22068
rect 23472 21728 23480 21792
rect 23544 21728 23560 21792
rect 23624 21728 23640 21792
rect 23704 21728 23720 21792
rect 23784 21728 23792 21792
rect 23472 20704 23792 21728
rect 25270 21181 25330 22067
rect 29104 21248 29424 22272
rect 29104 21184 29112 21248
rect 29176 21184 29192 21248
rect 29256 21184 29272 21248
rect 29336 21184 29352 21248
rect 29416 21184 29424 21248
rect 25267 21180 25333 21181
rect 25267 21116 25268 21180
rect 25332 21116 25333 21180
rect 25267 21115 25333 21116
rect 23472 20640 23480 20704
rect 23544 20640 23560 20704
rect 23624 20640 23640 20704
rect 23704 20640 23720 20704
rect 23784 20640 23792 20704
rect 23472 19616 23792 20640
rect 23472 19552 23480 19616
rect 23544 19552 23560 19616
rect 23624 19552 23640 19616
rect 23704 19552 23720 19616
rect 23784 19552 23792 19616
rect 23472 18528 23792 19552
rect 23472 18464 23480 18528
rect 23544 18464 23560 18528
rect 23624 18464 23640 18528
rect 23704 18464 23720 18528
rect 23784 18464 23792 18528
rect 23472 17440 23792 18464
rect 23472 17376 23480 17440
rect 23544 17376 23560 17440
rect 23624 17376 23640 17440
rect 23704 17376 23720 17440
rect 23784 17376 23792 17440
rect 23472 16352 23792 17376
rect 23472 16288 23480 16352
rect 23544 16288 23560 16352
rect 23624 16288 23640 16352
rect 23704 16288 23720 16352
rect 23784 16288 23792 16352
rect 23472 15264 23792 16288
rect 23472 15200 23480 15264
rect 23544 15200 23560 15264
rect 23624 15200 23640 15264
rect 23704 15200 23720 15264
rect 23784 15200 23792 15264
rect 23472 14176 23792 15200
rect 23472 14112 23480 14176
rect 23544 14112 23560 14176
rect 23624 14112 23640 14176
rect 23704 14112 23720 14176
rect 23784 14112 23792 14176
rect 23472 13088 23792 14112
rect 23472 13024 23480 13088
rect 23544 13024 23560 13088
rect 23624 13024 23640 13088
rect 23704 13024 23720 13088
rect 23784 13024 23792 13088
rect 23472 12000 23792 13024
rect 23472 11936 23480 12000
rect 23544 11936 23560 12000
rect 23624 11936 23640 12000
rect 23704 11936 23720 12000
rect 23784 11936 23792 12000
rect 23472 10912 23792 11936
rect 23472 10848 23480 10912
rect 23544 10848 23560 10912
rect 23624 10848 23640 10912
rect 23704 10848 23720 10912
rect 23784 10848 23792 10912
rect 23472 9824 23792 10848
rect 23472 9760 23480 9824
rect 23544 9760 23560 9824
rect 23624 9760 23640 9824
rect 23704 9760 23720 9824
rect 23784 9760 23792 9824
rect 23472 8736 23792 9760
rect 23472 8672 23480 8736
rect 23544 8672 23560 8736
rect 23624 8672 23640 8736
rect 23704 8672 23720 8736
rect 23784 8672 23792 8736
rect 23472 7648 23792 8672
rect 23472 7584 23480 7648
rect 23544 7584 23560 7648
rect 23624 7584 23640 7648
rect 23704 7584 23720 7648
rect 23784 7584 23792 7648
rect 23472 6560 23792 7584
rect 23472 6496 23480 6560
rect 23544 6496 23560 6560
rect 23624 6496 23640 6560
rect 23704 6496 23720 6560
rect 23784 6496 23792 6560
rect 23472 5472 23792 6496
rect 23472 5408 23480 5472
rect 23544 5408 23560 5472
rect 23624 5408 23640 5472
rect 23704 5408 23720 5472
rect 23784 5408 23792 5472
rect 23472 4384 23792 5408
rect 23472 4320 23480 4384
rect 23544 4320 23560 4384
rect 23624 4320 23640 4384
rect 23704 4320 23720 4384
rect 23784 4320 23792 4384
rect 23472 3296 23792 4320
rect 23472 3232 23480 3296
rect 23544 3232 23560 3296
rect 23624 3232 23640 3296
rect 23704 3232 23720 3296
rect 23784 3232 23792 3296
rect 23472 2208 23792 3232
rect 23472 2144 23480 2208
rect 23544 2144 23560 2208
rect 23624 2144 23640 2208
rect 23704 2144 23720 2208
rect 23784 2144 23792 2208
rect 23472 2128 23792 2144
rect 29104 20160 29424 21184
rect 29104 20096 29112 20160
rect 29176 20096 29192 20160
rect 29256 20096 29272 20160
rect 29336 20096 29352 20160
rect 29416 20096 29424 20160
rect 29104 19072 29424 20096
rect 29502 19413 29562 26827
rect 29683 24580 29749 24581
rect 29683 24516 29684 24580
rect 29748 24516 29749 24580
rect 29683 24515 29749 24516
rect 29686 19685 29746 24515
rect 29870 22813 29930 28867
rect 30051 28252 30117 28253
rect 30051 28188 30052 28252
rect 30116 28188 30117 28252
rect 30051 28187 30117 28188
rect 29867 22812 29933 22813
rect 29867 22748 29868 22812
rect 29932 22748 29933 22812
rect 29867 22747 29933 22748
rect 29683 19684 29749 19685
rect 29683 19620 29684 19684
rect 29748 19620 29749 19684
rect 29683 19619 29749 19620
rect 29499 19412 29565 19413
rect 29499 19348 29500 19412
rect 29564 19348 29565 19412
rect 29499 19347 29565 19348
rect 29104 19008 29112 19072
rect 29176 19008 29192 19072
rect 29256 19008 29272 19072
rect 29336 19008 29352 19072
rect 29416 19008 29424 19072
rect 29104 17984 29424 19008
rect 30054 18597 30114 28187
rect 30419 27300 30485 27301
rect 30419 27236 30420 27300
rect 30484 27236 30485 27300
rect 30419 27235 30485 27236
rect 30235 22404 30301 22405
rect 30235 22340 30236 22404
rect 30300 22340 30301 22404
rect 30235 22339 30301 22340
rect 30238 21997 30298 22339
rect 30235 21996 30301 21997
rect 30235 21932 30236 21996
rect 30300 21932 30301 21996
rect 30235 21931 30301 21932
rect 30422 21317 30482 27235
rect 30787 27164 30853 27165
rect 30787 27100 30788 27164
rect 30852 27100 30853 27164
rect 30787 27099 30853 27100
rect 30790 22677 30850 27099
rect 31707 25940 31773 25941
rect 31707 25876 31708 25940
rect 31772 25876 31773 25940
rect 31707 25875 31773 25876
rect 30787 22676 30853 22677
rect 30787 22612 30788 22676
rect 30852 22612 30853 22676
rect 30787 22611 30853 22612
rect 31710 22405 31770 25875
rect 32627 23900 32693 23901
rect 32627 23836 32628 23900
rect 32692 23836 32693 23900
rect 32627 23835 32693 23836
rect 31891 22540 31957 22541
rect 31891 22476 31892 22540
rect 31956 22476 31957 22540
rect 31891 22475 31957 22476
rect 31707 22404 31773 22405
rect 31707 22340 31708 22404
rect 31772 22340 31773 22404
rect 31707 22339 31773 22340
rect 30419 21316 30485 21317
rect 30419 21252 30420 21316
rect 30484 21252 30485 21316
rect 30419 21251 30485 21252
rect 30422 19413 30482 21251
rect 31894 20501 31954 22475
rect 32630 22133 32690 23835
rect 32811 22948 32877 22949
rect 32811 22884 32812 22948
rect 32876 22884 32877 22948
rect 32811 22883 32877 22884
rect 32627 22132 32693 22133
rect 32627 22068 32628 22132
rect 32692 22068 32693 22132
rect 32627 22067 32693 22068
rect 32814 21861 32874 22883
rect 32811 21860 32877 21861
rect 32811 21796 32812 21860
rect 32876 21796 32877 21860
rect 32811 21795 32877 21796
rect 31891 20500 31957 20501
rect 31891 20436 31892 20500
rect 31956 20436 31957 20500
rect 31891 20435 31957 20436
rect 30419 19412 30485 19413
rect 30419 19348 30420 19412
rect 30484 19348 30485 19412
rect 30419 19347 30485 19348
rect 30051 18596 30117 18597
rect 30051 18532 30052 18596
rect 30116 18532 30117 18596
rect 30051 18531 30117 18532
rect 29104 17920 29112 17984
rect 29176 17920 29192 17984
rect 29256 17920 29272 17984
rect 29336 17920 29352 17984
rect 29416 17920 29424 17984
rect 29104 16896 29424 17920
rect 29104 16832 29112 16896
rect 29176 16832 29192 16896
rect 29256 16832 29272 16896
rect 29336 16832 29352 16896
rect 29416 16832 29424 16896
rect 29104 15808 29424 16832
rect 29104 15744 29112 15808
rect 29176 15744 29192 15808
rect 29256 15744 29272 15808
rect 29336 15744 29352 15808
rect 29416 15744 29424 15808
rect 29104 14720 29424 15744
rect 29104 14656 29112 14720
rect 29176 14656 29192 14720
rect 29256 14656 29272 14720
rect 29336 14656 29352 14720
rect 29416 14656 29424 14720
rect 29104 13632 29424 14656
rect 29104 13568 29112 13632
rect 29176 13568 29192 13632
rect 29256 13568 29272 13632
rect 29336 13568 29352 13632
rect 29416 13568 29424 13632
rect 29104 12544 29424 13568
rect 29104 12480 29112 12544
rect 29176 12480 29192 12544
rect 29256 12480 29272 12544
rect 29336 12480 29352 12544
rect 29416 12480 29424 12544
rect 29104 11456 29424 12480
rect 29104 11392 29112 11456
rect 29176 11392 29192 11456
rect 29256 11392 29272 11456
rect 29336 11392 29352 11456
rect 29416 11392 29424 11456
rect 29104 10368 29424 11392
rect 29104 10304 29112 10368
rect 29176 10304 29192 10368
rect 29256 10304 29272 10368
rect 29336 10304 29352 10368
rect 29416 10304 29424 10368
rect 29104 9280 29424 10304
rect 29104 9216 29112 9280
rect 29176 9216 29192 9280
rect 29256 9216 29272 9280
rect 29336 9216 29352 9280
rect 29416 9216 29424 9280
rect 29104 8192 29424 9216
rect 29104 8128 29112 8192
rect 29176 8128 29192 8192
rect 29256 8128 29272 8192
rect 29336 8128 29352 8192
rect 29416 8128 29424 8192
rect 29104 7104 29424 8128
rect 29104 7040 29112 7104
rect 29176 7040 29192 7104
rect 29256 7040 29272 7104
rect 29336 7040 29352 7104
rect 29416 7040 29424 7104
rect 29104 6016 29424 7040
rect 29104 5952 29112 6016
rect 29176 5952 29192 6016
rect 29256 5952 29272 6016
rect 29336 5952 29352 6016
rect 29416 5952 29424 6016
rect 29104 4928 29424 5952
rect 29104 4864 29112 4928
rect 29176 4864 29192 4928
rect 29256 4864 29272 4928
rect 29336 4864 29352 4928
rect 29416 4864 29424 4928
rect 29104 3840 29424 4864
rect 29104 3776 29112 3840
rect 29176 3776 29192 3840
rect 29256 3776 29272 3840
rect 29336 3776 29352 3840
rect 29416 3776 29424 3840
rect 29104 2752 29424 3776
rect 29104 2688 29112 2752
rect 29176 2688 29192 2752
rect 29256 2688 29272 2752
rect 29336 2688 29352 2752
rect 29416 2688 29424 2752
rect 29104 2128 29424 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 12604 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1644511149
transform -1 0 12972 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1644511149
transform 1 0 23736 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1644511149
transform -1 0 13892 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1644511149
transform -1 0 31004 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51
timestamp 1644511149
transform 1 0 5796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55
timestamp 1644511149
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8280 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_108
timestamp 1644511149
transform 1 0 11040 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_113 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_125
timestamp 1644511149
transform 1 0 12604 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_134
timestamp 1644511149
transform 1 0 13432 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_144
timestamp 1644511149
transform 1 0 14352 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_156 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15456 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_162
timestamp 1644511149
transform 1 0 16008 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_174 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17112 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_182
timestamp 1644511149
transform 1 0 17848 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_189
timestamp 1644511149
transform 1 0 18492 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1644511149
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_220
timestamp 1644511149
transform 1 0 21344 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_228
timestamp 1644511149
transform 1 0 22080 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_240
timestamp 1644511149
transform 1 0 23184 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_253
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_265
timestamp 1644511149
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1644511149
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_281
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_293
timestamp 1644511149
transform 1 0 28060 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_304
timestamp 1644511149
transform 1 0 29072 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1644511149
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_332
timestamp 1644511149
transform 1 0 31648 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1644511149
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_360
timestamp 1644511149
transform 1 0 34224 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_3
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_9
timestamp 1644511149
transform 1 0 1932 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_34
timestamp 1644511149
transform 1 0 4232 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_41
timestamp 1644511149
transform 1 0 4876 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1644511149
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_78
timestamp 1644511149
transform 1 0 8280 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_86
timestamp 1644511149
transform 1 0 9016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_108
timestamp 1644511149
transform 1 0 11040 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_113
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_117
timestamp 1644511149
transform 1 0 11868 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_139
timestamp 1644511149
transform 1 0 13892 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_164
timestamp 1644511149
transform 1 0 16192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_192
timestamp 1644511149
transform 1 0 18768 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_198
timestamp 1644511149
transform 1 0 19320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_220
timestamp 1644511149
transform 1 0 21344 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_228
timestamp 1644511149
transform 1 0 22080 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_243
timestamp 1644511149
transform 1 0 23460 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_268
timestamp 1644511149
transform 1 0 25760 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_281
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_292
timestamp 1644511149
transform 1 0 27968 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_299
timestamp 1644511149
transform 1 0 28612 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_306
timestamp 1644511149
transform 1 0 29256 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_331
timestamp 1644511149
transform 1 0 31556 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1644511149
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_337
timestamp 1644511149
transform 1 0 32108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_360
timestamp 1644511149
transform 1 0 34224 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_24
timestamp 1644511149
transform 1 0 3312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_32
timestamp 1644511149
transform 1 0 4048 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_57
timestamp 1644511149
transform 1 0 6348 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_64
timestamp 1644511149
transform 1 0 6992 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_72
timestamp 1644511149
transform 1 0 7728 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1644511149
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1644511149
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_88
timestamp 1644511149
transform 1 0 9200 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_113
timestamp 1644511149
transform 1 0 11500 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_120
timestamp 1644511149
transform 1 0 12144 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_128
timestamp 1644511149
transform 1 0 12880 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_132
timestamp 1644511149
transform 1 0 13248 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_146
timestamp 1644511149
transform 1 0 14536 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_154
timestamp 1644511149
transform 1 0 15272 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_177
timestamp 1644511149
transform 1 0 17388 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_184
timestamp 1644511149
transform 1 0 18032 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_202
timestamp 1644511149
transform 1 0 19688 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_206
timestamp 1644511149
transform 1 0 20056 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_210
timestamp 1644511149
transform 1 0 20424 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_235
timestamp 1644511149
transform 1 0 22724 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_247
timestamp 1644511149
transform 1 0 23828 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1644511149
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_256
timestamp 1644511149
transform 1 0 24656 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_268
timestamp 1644511149
transform 1 0 25760 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_280
timestamp 1644511149
transform 1 0 26864 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_286
timestamp 1644511149
transform 1 0 27416 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_290
timestamp 1644511149
transform 1 0 27784 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_297
timestamp 1644511149
transform 1 0 28428 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_304
timestamp 1644511149
transform 1 0 29072 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_315
timestamp 1644511149
transform 1 0 30084 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_340
timestamp 1644511149
transform 1 0 32384 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_358
timestamp 1644511149
transform 1 0 34040 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_28
timestamp 1644511149
transform 1 0 3680 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_35
timestamp 1644511149
transform 1 0 4324 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_42
timestamp 1644511149
transform 1 0 4968 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_49
timestamp 1644511149
transform 1 0 5612 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1644511149
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_60
timestamp 1644511149
transform 1 0 6624 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_67
timestamp 1644511149
transform 1 0 7268 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_71
timestamp 1644511149
transform 1 0 7636 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_93
timestamp 1644511149
transform 1 0 9660 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_3_102
timestamp 1644511149
transform 1 0 10488 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1644511149
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_113
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_125
timestamp 1644511149
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_137
timestamp 1644511149
transform 1 0 13708 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_143
timestamp 1644511149
transform 1 0 14260 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_147
timestamp 1644511149
transform 1 0 14628 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_155
timestamp 1644511149
transform 1 0 15364 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_160
timestamp 1644511149
transform 1 0 15824 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_169
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_181
timestamp 1644511149
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_193
timestamp 1644511149
transform 1 0 18860 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_199
timestamp 1644511149
transform 1 0 19412 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_203
timestamp 1644511149
transform 1 0 19780 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_213
timestamp 1644511149
transform 1 0 20700 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_220
timestamp 1644511149
transform 1 0 21344 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_225
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_237
timestamp 1644511149
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_249
timestamp 1644511149
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_261
timestamp 1644511149
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1644511149
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1644511149
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_281
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_293
timestamp 1644511149
transform 1 0 28060 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_300
timestamp 1644511149
transform 1 0 28704 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_307
timestamp 1644511149
transform 1 0 29348 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_332
timestamp 1644511149
transform 1 0 31648 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_358
timestamp 1644511149
transform 1 0 34040 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_7
timestamp 1644511149
transform 1 0 1748 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_11
timestamp 1644511149
transform 1 0 2116 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_4_20
timestamp 1644511149
transform 1 0 2944 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_32
timestamp 1644511149
transform 1 0 4048 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_39
timestamp 1644511149
transform 1 0 4692 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_43
timestamp 1644511149
transform 1 0 5060 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_65
timestamp 1644511149
transform 1 0 7084 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_76
timestamp 1644511149
transform 1 0 8096 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_85
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_96
timestamp 1644511149
transform 1 0 9936 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_103
timestamp 1644511149
transform 1 0 10580 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_115
timestamp 1644511149
transform 1 0 11684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_127
timestamp 1644511149
transform 1 0 12788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1644511149
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_153
timestamp 1644511149
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_165
timestamp 1644511149
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_177
timestamp 1644511149
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1644511149
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1644511149
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_197
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_209
timestamp 1644511149
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_221
timestamp 1644511149
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_233
timestamp 1644511149
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1644511149
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1644511149
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_253
timestamp 1644511149
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_265
timestamp 1644511149
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_277
timestamp 1644511149
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_289
timestamp 1644511149
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1644511149
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1644511149
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_309
timestamp 1644511149
transform 1 0 29532 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_333
timestamp 1644511149
transform 1 0 31740 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_360
timestamp 1644511149
transform 1 0 34224 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_10
timestamp 1644511149
transform 1 0 2024 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_37
timestamp 1644511149
transform 1 0 4508 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_44
timestamp 1644511149
transform 1 0 5152 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1644511149
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1644511149
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_60
timestamp 1644511149
transform 1 0 6624 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_72
timestamp 1644511149
transform 1 0 7728 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_84
timestamp 1644511149
transform 1 0 8832 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_96
timestamp 1644511149
transform 1 0 9936 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_108
timestamp 1644511149
transform 1 0 11040 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_113
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_125
timestamp 1644511149
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_137
timestamp 1644511149
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_149
timestamp 1644511149
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1644511149
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1644511149
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_169
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_181
timestamp 1644511149
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_193
timestamp 1644511149
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_205
timestamp 1644511149
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1644511149
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1644511149
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_225
timestamp 1644511149
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_237
timestamp 1644511149
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_249
timestamp 1644511149
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_261
timestamp 1644511149
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1644511149
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1644511149
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_281
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_293
timestamp 1644511149
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_305
timestamp 1644511149
transform 1 0 29164 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_311
timestamp 1644511149
transform 1 0 29716 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_318
timestamp 1644511149
transform 1 0 30360 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_325
timestamp 1644511149
transform 1 0 31004 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_332
timestamp 1644511149
transform 1 0 31648 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_337
timestamp 1644511149
transform 1 0 32108 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_360
timestamp 1644511149
transform 1 0 34224 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp 1644511149
transform 1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_50
timestamp 1644511149
transform 1 0 5704 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_57
timestamp 1644511149
transform 1 0 6348 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_69
timestamp 1644511149
transform 1 0 7452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_81
timestamp 1644511149
transform 1 0 8556 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_97
timestamp 1644511149
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_109
timestamp 1644511149
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_121
timestamp 1644511149
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1644511149
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1644511149
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_153
timestamp 1644511149
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_165
timestamp 1644511149
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_177
timestamp 1644511149
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1644511149
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1644511149
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_197
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_209
timestamp 1644511149
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_221
timestamp 1644511149
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_233
timestamp 1644511149
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1644511149
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1644511149
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_253
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_265
timestamp 1644511149
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_277
timestamp 1644511149
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_289
timestamp 1644511149
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1644511149
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1644511149
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_309
timestamp 1644511149
transform 1 0 29532 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_317
timestamp 1644511149
transform 1 0 30268 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_321
timestamp 1644511149
transform 1 0 30636 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_328
timestamp 1644511149
transform 1 0 31280 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_353
timestamp 1644511149
transform 1 0 33580 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_360
timestamp 1644511149
transform 1 0 34224 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_6
timestamp 1644511149
transform 1 0 1656 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_31
timestamp 1644511149
transform 1 0 3956 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_38
timestamp 1644511149
transform 1 0 4600 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_45
timestamp 1644511149
transform 1 0 5244 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_53
timestamp 1644511149
transform 1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1644511149
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_81
timestamp 1644511149
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1644511149
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1644511149
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1644511149
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_113
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_125
timestamp 1644511149
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_137
timestamp 1644511149
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_149
timestamp 1644511149
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1644511149
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1644511149
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_169
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_181
timestamp 1644511149
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_193
timestamp 1644511149
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_205
timestamp 1644511149
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1644511149
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1644511149
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_225
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_237
timestamp 1644511149
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_249
timestamp 1644511149
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_261
timestamp 1644511149
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1644511149
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1644511149
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_293
timestamp 1644511149
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_305
timestamp 1644511149
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_317
timestamp 1644511149
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_332
timestamp 1644511149
transform 1 0 31648 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_337
timestamp 1644511149
transform 1 0 32108 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_342
timestamp 1644511149
transform 1 0 32568 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_349
timestamp 1644511149
transform 1 0 33212 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_356
timestamp 1644511149
transform 1 0 33856 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_12
timestamp 1644511149
transform 1 0 2208 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_19
timestamp 1644511149
transform 1 0 2852 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1644511149
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1644511149
transform 1 0 4048 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1644511149
transform 1 0 5152 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_56
timestamp 1644511149
transform 1 0 6256 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_68
timestamp 1644511149
transform 1 0 7360 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_80
timestamp 1644511149
transform 1 0 8464 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_97
timestamp 1644511149
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_109
timestamp 1644511149
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_121
timestamp 1644511149
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1644511149
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1644511149
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_153
timestamp 1644511149
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_165
timestamp 1644511149
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_177
timestamp 1644511149
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1644511149
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1644511149
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_197
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_209
timestamp 1644511149
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_221
timestamp 1644511149
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_233
timestamp 1644511149
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1644511149
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1644511149
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_253
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_265
timestamp 1644511149
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_277
timestamp 1644511149
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_289
timestamp 1644511149
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1644511149
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1644511149
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_309
timestamp 1644511149
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_321
timestamp 1644511149
transform 1 0 30636 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_329
timestamp 1644511149
transform 1 0 31372 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_335
timestamp 1644511149
transform 1 0 31924 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_360
timestamp 1644511149
transform 1 0 34224 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_26
timestamp 1644511149
transform 1 0 3496 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_33
timestamp 1644511149
transform 1 0 4140 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_45
timestamp 1644511149
transform 1 0 5244 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_53
timestamp 1644511149
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_69
timestamp 1644511149
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_81
timestamp 1644511149
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_93
timestamp 1644511149
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1644511149
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1644511149
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_113
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_125
timestamp 1644511149
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_137
timestamp 1644511149
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_149
timestamp 1644511149
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1644511149
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1644511149
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_181
timestamp 1644511149
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_193
timestamp 1644511149
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_205
timestamp 1644511149
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1644511149
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1644511149
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_225
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_237
timestamp 1644511149
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_249
timestamp 1644511149
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_261
timestamp 1644511149
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1644511149
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1644511149
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_281
timestamp 1644511149
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_293
timestamp 1644511149
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_305
timestamp 1644511149
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_317
timestamp 1644511149
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1644511149
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1644511149
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_337
timestamp 1644511149
transform 1 0 32108 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_345
timestamp 1644511149
transform 1 0 32844 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_351
timestamp 1644511149
transform 1 0 33396 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_358
timestamp 1644511149
transform 1 0 34040 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_10_3
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_12
timestamp 1644511149
transform 1 0 2208 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_19
timestamp 1644511149
transform 1 0 2852 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1644511149
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1644511149
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_53
timestamp 1644511149
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_65
timestamp 1644511149
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1644511149
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1644511149
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_97
timestamp 1644511149
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_109
timestamp 1644511149
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_121
timestamp 1644511149
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1644511149
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1644511149
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_153
timestamp 1644511149
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_165
timestamp 1644511149
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_177
timestamp 1644511149
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1644511149
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1644511149
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_197
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_209
timestamp 1644511149
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_221
timestamp 1644511149
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_233
timestamp 1644511149
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1644511149
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1644511149
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_253
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_265
timestamp 1644511149
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_277
timestamp 1644511149
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_289
timestamp 1644511149
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1644511149
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1644511149
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_309
timestamp 1644511149
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_321
timestamp 1644511149
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_333
timestamp 1644511149
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_345
timestamp 1644511149
transform 1 0 32844 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_353
timestamp 1644511149
transform 1 0 33580 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_358
timestamp 1644511149
transform 1 0 34040 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_7
timestamp 1644511149
transform 1 0 1748 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_11
timestamp 1644511149
transform 1 0 2116 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_18
timestamp 1644511149
transform 1 0 2760 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_30
timestamp 1644511149
transform 1 0 3864 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_42
timestamp 1644511149
transform 1 0 4968 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1644511149
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_69
timestamp 1644511149
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_81
timestamp 1644511149
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_93
timestamp 1644511149
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1644511149
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1644511149
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_113
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_125
timestamp 1644511149
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_137
timestamp 1644511149
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_149
timestamp 1644511149
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1644511149
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1644511149
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_169
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_181
timestamp 1644511149
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_193
timestamp 1644511149
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_205
timestamp 1644511149
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1644511149
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1644511149
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_225
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_237
timestamp 1644511149
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_249
timestamp 1644511149
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_261
timestamp 1644511149
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1644511149
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1644511149
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_281
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_293
timestamp 1644511149
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_305
timestamp 1644511149
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_317
timestamp 1644511149
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1644511149
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1644511149
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_337
timestamp 1644511149
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_349
timestamp 1644511149
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_361
timestamp 1644511149
transform 1 0 34316 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_24
timestamp 1644511149
transform 1 0 3312 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_41
timestamp 1644511149
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_53
timestamp 1644511149
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_65
timestamp 1644511149
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1644511149
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1644511149
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_85
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_97
timestamp 1644511149
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_109
timestamp 1644511149
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_121
timestamp 1644511149
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1644511149
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1644511149
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_153
timestamp 1644511149
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_165
timestamp 1644511149
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_177
timestamp 1644511149
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1644511149
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1644511149
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_197
timestamp 1644511149
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_209
timestamp 1644511149
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_221
timestamp 1644511149
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_233
timestamp 1644511149
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1644511149
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1644511149
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_253
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_265
timestamp 1644511149
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_277
timestamp 1644511149
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_289
timestamp 1644511149
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1644511149
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1644511149
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_309
timestamp 1644511149
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_321
timestamp 1644511149
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_333
timestamp 1644511149
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_345
timestamp 1644511149
transform 1 0 32844 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_353
timestamp 1644511149
transform 1 0 33580 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_358
timestamp 1644511149
transform 1 0 34040 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_25
timestamp 1644511149
transform 1 0 3404 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_37
timestamp 1644511149
transform 1 0 4508 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_49
timestamp 1644511149
transform 1 0 5612 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1644511149
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_69
timestamp 1644511149
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_81
timestamp 1644511149
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_93
timestamp 1644511149
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1644511149
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1644511149
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_113
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_125
timestamp 1644511149
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_137
timestamp 1644511149
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_149
timestamp 1644511149
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1644511149
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1644511149
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_169
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_181
timestamp 1644511149
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_193
timestamp 1644511149
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_205
timestamp 1644511149
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1644511149
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1644511149
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_225
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_237
timestamp 1644511149
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_249
timestamp 1644511149
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_261
timestamp 1644511149
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1644511149
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1644511149
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_281
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_293
timestamp 1644511149
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_305
timestamp 1644511149
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_317
timestamp 1644511149
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1644511149
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1644511149
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_337
timestamp 1644511149
transform 1 0 32108 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_360
timestamp 1644511149
transform 1 0 34224 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_3
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_10
timestamp 1644511149
transform 1 0 2024 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_17
timestamp 1644511149
transform 1 0 2668 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_25
timestamp 1644511149
transform 1 0 3404 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_53
timestamp 1644511149
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_65
timestamp 1644511149
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1644511149
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1644511149
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_97
timestamp 1644511149
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_109
timestamp 1644511149
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_121
timestamp 1644511149
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1644511149
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1644511149
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_153
timestamp 1644511149
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_165
timestamp 1644511149
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_177
timestamp 1644511149
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1644511149
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1644511149
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_197
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_209
timestamp 1644511149
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_221
timestamp 1644511149
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_233
timestamp 1644511149
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1644511149
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1644511149
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_253
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_265
timestamp 1644511149
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_277
timestamp 1644511149
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_289
timestamp 1644511149
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1644511149
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1644511149
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_309
timestamp 1644511149
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_321
timestamp 1644511149
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_333
timestamp 1644511149
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_345
timestamp 1644511149
transform 1 0 32844 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_352
timestamp 1644511149
transform 1 0 33488 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_360
timestamp 1644511149
transform 1 0 34224 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_3
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_7
timestamp 1644511149
transform 1 0 1748 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_11
timestamp 1644511149
transform 1 0 2116 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_18
timestamp 1644511149
transform 1 0 2760 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_30
timestamp 1644511149
transform 1 0 3864 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_42
timestamp 1644511149
transform 1 0 4968 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 1644511149
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1644511149
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_81
timestamp 1644511149
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_93
timestamp 1644511149
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1644511149
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1644511149
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_113
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_125
timestamp 1644511149
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_137
timestamp 1644511149
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_149
timestamp 1644511149
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1644511149
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1644511149
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_169
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_181
timestamp 1644511149
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_193
timestamp 1644511149
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_205
timestamp 1644511149
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1644511149
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1644511149
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_225
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_237
timestamp 1644511149
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_249
timestamp 1644511149
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_261
timestamp 1644511149
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1644511149
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1644511149
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_281
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_293
timestamp 1644511149
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_305
timestamp 1644511149
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_317
timestamp 1644511149
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1644511149
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1644511149
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_337
timestamp 1644511149
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_349
timestamp 1644511149
transform 1 0 33212 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_15_358
timestamp 1644511149
transform 1 0 34040 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_24
timestamp 1644511149
transform 1 0 3312 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1644511149
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_53
timestamp 1644511149
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_65
timestamp 1644511149
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1644511149
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1644511149
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_85
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_97
timestamp 1644511149
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_109
timestamp 1644511149
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_121
timestamp 1644511149
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1644511149
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1644511149
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_141
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_153
timestamp 1644511149
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_165
timestamp 1644511149
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_177
timestamp 1644511149
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1644511149
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1644511149
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_197
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_209
timestamp 1644511149
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_221
timestamp 1644511149
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_233
timestamp 1644511149
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1644511149
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1644511149
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_253
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_265
timestamp 1644511149
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_277
timestamp 1644511149
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_289
timestamp 1644511149
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1644511149
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1644511149
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_309
timestamp 1644511149
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_321
timestamp 1644511149
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_333
timestamp 1644511149
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_345
timestamp 1644511149
transform 1 0 32844 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_356
timestamp 1644511149
transform 1 0 33856 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_26
timestamp 1644511149
transform 1 0 3496 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_38
timestamp 1644511149
transform 1 0 4600 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_50
timestamp 1644511149
transform 1 0 5704 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_69
timestamp 1644511149
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_81
timestamp 1644511149
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_93
timestamp 1644511149
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1644511149
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1644511149
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_113
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_125
timestamp 1644511149
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_137
timestamp 1644511149
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_149
timestamp 1644511149
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1644511149
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1644511149
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_169
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_181
timestamp 1644511149
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_193
timestamp 1644511149
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_205
timestamp 1644511149
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1644511149
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1644511149
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_225
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_237
timestamp 1644511149
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_249
timestamp 1644511149
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_261
timestamp 1644511149
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1644511149
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1644511149
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_281
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_293
timestamp 1644511149
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_305
timestamp 1644511149
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_317
timestamp 1644511149
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1644511149
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1644511149
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_337
timestamp 1644511149
transform 1 0 32108 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_360
timestamp 1644511149
transform 1 0 34224 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_3
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_18_12
timestamp 1644511149
transform 1 0 2208 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_24
timestamp 1644511149
transform 1 0 3312 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1644511149
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_53
timestamp 1644511149
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_65
timestamp 1644511149
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1644511149
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1644511149
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_85
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_97
timestamp 1644511149
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_109
timestamp 1644511149
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_121
timestamp 1644511149
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1644511149
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1644511149
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_153
timestamp 1644511149
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_165
timestamp 1644511149
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_177
timestamp 1644511149
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1644511149
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1644511149
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_197
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_209
timestamp 1644511149
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_221
timestamp 1644511149
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_233
timestamp 1644511149
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1644511149
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1644511149
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_253
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_265
timestamp 1644511149
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_277
timestamp 1644511149
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_289
timestamp 1644511149
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1644511149
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1644511149
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_309
timestamp 1644511149
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_321
timestamp 1644511149
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_333
timestamp 1644511149
transform 1 0 31740 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_360
timestamp 1644511149
transform 1 0 34224 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_3
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_9
timestamp 1644511149
transform 1 0 1932 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_21
timestamp 1644511149
transform 1 0 3036 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_33
timestamp 1644511149
transform 1 0 4140 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_45
timestamp 1644511149
transform 1 0 5244 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_53
timestamp 1644511149
transform 1 0 5980 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 1644511149
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_81
timestamp 1644511149
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_93
timestamp 1644511149
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1644511149
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1644511149
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_113
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_125
timestamp 1644511149
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_137
timestamp 1644511149
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_149
timestamp 1644511149
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1644511149
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1644511149
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_169
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_181
timestamp 1644511149
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_193
timestamp 1644511149
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_205
timestamp 1644511149
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1644511149
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1644511149
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_225
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_237
timestamp 1644511149
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_249
timestamp 1644511149
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_261
timestamp 1644511149
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1644511149
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1644511149
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_281
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_293
timestamp 1644511149
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_305
timestamp 1644511149
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_317
timestamp 1644511149
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1644511149
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1644511149
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_337
timestamp 1644511149
transform 1 0 32108 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_360
timestamp 1644511149
transform 1 0 34224 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_24
timestamp 1644511149
transform 1 0 3312 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1644511149
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 1644511149
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1644511149
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1644511149
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1644511149
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_97
timestamp 1644511149
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_109
timestamp 1644511149
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_121
timestamp 1644511149
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1644511149
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1644511149
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_153
timestamp 1644511149
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_165
timestamp 1644511149
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_177
timestamp 1644511149
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1644511149
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1644511149
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_197
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_209
timestamp 1644511149
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_221
timestamp 1644511149
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_233
timestamp 1644511149
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1644511149
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1644511149
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_253
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_265
timestamp 1644511149
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_277
timestamp 1644511149
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_289
timestamp 1644511149
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1644511149
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1644511149
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_309
timestamp 1644511149
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_321
timestamp 1644511149
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_333
timestamp 1644511149
transform 1 0 31740 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_342
timestamp 1644511149
transform 1 0 32568 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_349
timestamp 1644511149
transform 1 0 33212 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_356
timestamp 1644511149
transform 1 0 33856 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_3
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_10
timestamp 1644511149
transform 1 0 2024 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_19
timestamp 1644511149
transform 1 0 2852 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_26
timestamp 1644511149
transform 1 0 3496 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_38
timestamp 1644511149
transform 1 0 4600 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_50
timestamp 1644511149
transform 1 0 5704 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_81
timestamp 1644511149
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_93
timestamp 1644511149
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1644511149
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1644511149
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_113
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_125
timestamp 1644511149
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_137
timestamp 1644511149
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_149
timestamp 1644511149
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1644511149
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1644511149
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_169
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_181
timestamp 1644511149
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_193
timestamp 1644511149
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_205
timestamp 1644511149
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1644511149
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1644511149
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_225
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_237
timestamp 1644511149
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_249
timestamp 1644511149
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_261
timestamp 1644511149
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1644511149
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1644511149
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_281
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_293
timestamp 1644511149
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_305
timestamp 1644511149
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_317
timestamp 1644511149
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_332
timestamp 1644511149
transform 1 0 31648 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_337
timestamp 1644511149
transform 1 0 32108 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_360
timestamp 1644511149
transform 1 0 34224 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_24
timestamp 1644511149
transform 1 0 3312 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1644511149
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_53
timestamp 1644511149
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_65
timestamp 1644511149
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1644511149
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1644511149
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_85
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_97
timestamp 1644511149
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_109
timestamp 1644511149
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_121
timestamp 1644511149
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1644511149
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1644511149
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_141
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_153
timestamp 1644511149
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_165
timestamp 1644511149
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_177
timestamp 1644511149
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1644511149
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1644511149
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_197
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_209
timestamp 1644511149
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_221
timestamp 1644511149
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_233
timestamp 1644511149
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1644511149
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1644511149
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_253
timestamp 1644511149
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_265
timestamp 1644511149
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_277
timestamp 1644511149
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_289
timestamp 1644511149
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1644511149
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1644511149
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_309
timestamp 1644511149
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_321
timestamp 1644511149
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_333
timestamp 1644511149
transform 1 0 31740 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_360
timestamp 1644511149
transform 1 0 34224 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_12
timestamp 1644511149
transform 1 0 2208 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_19
timestamp 1644511149
transform 1 0 2852 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_31
timestamp 1644511149
transform 1 0 3956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_43
timestamp 1644511149
transform 1 0 5060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1644511149
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1644511149
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_81
timestamp 1644511149
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_93
timestamp 1644511149
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1644511149
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1644511149
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_113
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_125
timestamp 1644511149
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_137
timestamp 1644511149
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_149
timestamp 1644511149
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1644511149
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1644511149
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_169
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_181
timestamp 1644511149
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_193
timestamp 1644511149
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_205
timestamp 1644511149
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1644511149
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1644511149
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_225
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_237
timestamp 1644511149
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_249
timestamp 1644511149
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_261
timestamp 1644511149
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1644511149
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1644511149
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_281
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_293
timestamp 1644511149
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_305
timestamp 1644511149
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_317
timestamp 1644511149
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1644511149
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1644511149
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_337
timestamp 1644511149
transform 1 0 32108 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_343
timestamp 1644511149
transform 1 0 32660 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_350
timestamp 1644511149
transform 1 0 33304 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_357
timestamp 1644511149
transform 1 0 33948 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_363
timestamp 1644511149
transform 1 0 34500 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_24
timestamp 1644511149
transform 1 0 3312 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1644511149
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_53
timestamp 1644511149
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_65
timestamp 1644511149
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1644511149
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1644511149
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_85
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_97
timestamp 1644511149
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_109
timestamp 1644511149
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_121
timestamp 1644511149
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1644511149
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1644511149
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_153
timestamp 1644511149
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_165
timestamp 1644511149
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_177
timestamp 1644511149
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1644511149
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1644511149
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_197
timestamp 1644511149
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_209
timestamp 1644511149
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_221
timestamp 1644511149
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_233
timestamp 1644511149
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1644511149
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1644511149
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_253
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_265
timestamp 1644511149
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_277
timestamp 1644511149
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_289
timestamp 1644511149
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1644511149
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1644511149
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_309
timestamp 1644511149
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_321
timestamp 1644511149
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_333
timestamp 1644511149
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_345
timestamp 1644511149
transform 1 0 32844 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_349
timestamp 1644511149
transform 1 0 33212 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_356
timestamp 1644511149
transform 1 0 33856 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_3
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_9
timestamp 1644511149
transform 1 0 1932 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_21
timestamp 1644511149
transform 1 0 3036 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_33
timestamp 1644511149
transform 1 0 4140 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_45
timestamp 1644511149
transform 1 0 5244 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_53
timestamp 1644511149
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_69
timestamp 1644511149
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_81
timestamp 1644511149
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_93
timestamp 1644511149
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1644511149
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1644511149
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_113
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_125
timestamp 1644511149
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_137
timestamp 1644511149
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_149
timestamp 1644511149
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1644511149
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1644511149
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_169
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_181
timestamp 1644511149
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_193
timestamp 1644511149
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_205
timestamp 1644511149
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1644511149
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1644511149
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_225
timestamp 1644511149
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_237
timestamp 1644511149
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_249
timestamp 1644511149
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_261
timestamp 1644511149
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1644511149
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1644511149
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_281
timestamp 1644511149
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_293
timestamp 1644511149
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_305
timestamp 1644511149
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_317
timestamp 1644511149
transform 1 0 30268 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_321
timestamp 1644511149
transform 1 0 30636 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_325
timestamp 1644511149
transform 1 0 31004 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_332
timestamp 1644511149
transform 1 0 31648 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_337
timestamp 1644511149
transform 1 0 32108 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_360
timestamp 1644511149
transform 1 0 34224 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_3
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_10
timestamp 1644511149
transform 1 0 2024 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_17
timestamp 1644511149
transform 1 0 2668 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_25
timestamp 1644511149
transform 1 0 3404 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1644511149
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_53
timestamp 1644511149
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_65
timestamp 1644511149
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1644511149
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1644511149
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_85
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_97
timestamp 1644511149
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_109
timestamp 1644511149
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_121
timestamp 1644511149
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1644511149
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1644511149
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_153
timestamp 1644511149
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_165
timestamp 1644511149
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_177
timestamp 1644511149
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1644511149
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1644511149
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_197
timestamp 1644511149
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_209
timestamp 1644511149
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_221
timestamp 1644511149
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_233
timestamp 1644511149
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1644511149
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1644511149
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_253
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_265
timestamp 1644511149
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_277
timestamp 1644511149
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_289
timestamp 1644511149
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1644511149
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1644511149
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_309
timestamp 1644511149
transform 1 0 29532 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_315
timestamp 1644511149
transform 1 0 30084 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_319
timestamp 1644511149
transform 1 0 30452 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_326
timestamp 1644511149
transform 1 0 31096 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_333
timestamp 1644511149
transform 1 0 31740 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_340
timestamp 1644511149
transform 1 0 32384 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_346
timestamp 1644511149
transform 1 0 32936 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_350
timestamp 1644511149
transform 1 0 33304 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1644511149
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1644511149
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_3
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_25
timestamp 1644511149
transform 1 0 3404 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_37
timestamp 1644511149
transform 1 0 4508 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_49
timestamp 1644511149
transform 1 0 5612 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1644511149
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_69
timestamp 1644511149
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_81
timestamp 1644511149
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_93
timestamp 1644511149
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1644511149
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1644511149
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_113
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_125
timestamp 1644511149
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_137
timestamp 1644511149
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_149
timestamp 1644511149
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1644511149
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1644511149
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_169
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_181
timestamp 1644511149
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_193
timestamp 1644511149
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_205
timestamp 1644511149
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1644511149
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1644511149
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_225
timestamp 1644511149
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_237
timestamp 1644511149
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_249
timestamp 1644511149
transform 1 0 24012 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_255
timestamp 1644511149
transform 1 0 24564 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_260
timestamp 1644511149
transform 1 0 25024 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_267
timestamp 1644511149
transform 1 0 25668 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1644511149
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_281
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_289
timestamp 1644511149
transform 1 0 27692 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_293
timestamp 1644511149
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_305
timestamp 1644511149
transform 1 0 29164 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_311
timestamp 1644511149
transform 1 0 29716 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_318
timestamp 1644511149
transform 1 0 30360 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_325
timestamp 1644511149
transform 1 0 31004 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_332
timestamp 1644511149
transform 1 0 31648 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_337
timestamp 1644511149
transform 1 0 32108 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_360
timestamp 1644511149
transform 1 0 34224 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_3
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_10
timestamp 1644511149
transform 1 0 2024 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_22
timestamp 1644511149
transform 1 0 3128 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_41
timestamp 1644511149
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_53
timestamp 1644511149
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_65
timestamp 1644511149
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1644511149
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1644511149
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_85
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_97
timestamp 1644511149
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_109
timestamp 1644511149
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_121
timestamp 1644511149
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1644511149
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1644511149
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_141
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_153
timestamp 1644511149
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_165
timestamp 1644511149
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_177
timestamp 1644511149
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1644511149
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1644511149
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_197
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_209
timestamp 1644511149
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_221
timestamp 1644511149
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_233
timestamp 1644511149
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1644511149
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1644511149
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_253
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_263
timestamp 1644511149
transform 1 0 25300 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_271
timestamp 1644511149
transform 1 0 26036 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_278
timestamp 1644511149
transform 1 0 26680 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_284
timestamp 1644511149
transform 1 0 27232 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_289
timestamp 1644511149
transform 1 0 27692 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_297
timestamp 1644511149
transform 1 0 28428 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1644511149
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1644511149
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_309
timestamp 1644511149
transform 1 0 29532 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_316
timestamp 1644511149
transform 1 0 30176 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_323
timestamp 1644511149
transform 1 0 30820 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_330
timestamp 1644511149
transform 1 0 31464 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_338
timestamp 1644511149
transform 1 0 32200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_360
timestamp 1644511149
transform 1 0 34224 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_3
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_25
timestamp 1644511149
transform 1 0 3404 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_37
timestamp 1644511149
transform 1 0 4508 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_49
timestamp 1644511149
transform 1 0 5612 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1644511149
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_69
timestamp 1644511149
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_81
timestamp 1644511149
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_93
timestamp 1644511149
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1644511149
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1644511149
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_113
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_125
timestamp 1644511149
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_137
timestamp 1644511149
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_149
timestamp 1644511149
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1644511149
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1644511149
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_169
timestamp 1644511149
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_181
timestamp 1644511149
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_193
timestamp 1644511149
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_205
timestamp 1644511149
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1644511149
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1644511149
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_225
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_29_234
timestamp 1644511149
transform 1 0 22632 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_249
timestamp 1644511149
transform 1 0 24012 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_256
timestamp 1644511149
transform 1 0 24656 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_276
timestamp 1644511149
transform 1 0 26496 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_297
timestamp 1644511149
transform 1 0 28428 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_305
timestamp 1644511149
transform 1 0 29164 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_312
timestamp 1644511149
transform 1 0 29808 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_319
timestamp 1644511149
transform 1 0 30452 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_327
timestamp 1644511149
transform 1 0 31188 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_332
timestamp 1644511149
transform 1 0 31648 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_337
timestamp 1644511149
transform 1 0 32108 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_344
timestamp 1644511149
transform 1 0 32752 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_352
timestamp 1644511149
transform 1 0 33488 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_356
timestamp 1644511149
transform 1 0 33856 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_3
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_7
timestamp 1644511149
transform 1 0 1748 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_13
timestamp 1644511149
transform 1 0 2300 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_17
timestamp 1644511149
transform 1 0 2668 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_25
timestamp 1644511149
transform 1 0 3404 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1644511149
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_53
timestamp 1644511149
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_65
timestamp 1644511149
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1644511149
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1644511149
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_97
timestamp 1644511149
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_109
timestamp 1644511149
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_121
timestamp 1644511149
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1644511149
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1644511149
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_141
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_153
timestamp 1644511149
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_165
timestamp 1644511149
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_177
timestamp 1644511149
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1644511149
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1644511149
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_197
timestamp 1644511149
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_209
timestamp 1644511149
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_221
timestamp 1644511149
transform 1 0 21436 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_227
timestamp 1644511149
transform 1 0 21988 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_236
timestamp 1644511149
transform 1 0 22816 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_247
timestamp 1644511149
transform 1 0 23828 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1644511149
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_253
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_258
timestamp 1644511149
transform 1 0 24840 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_278
timestamp 1644511149
transform 1 0 26680 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_284
timestamp 1644511149
transform 1 0 27232 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1644511149
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1644511149
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_325
timestamp 1644511149
transform 1 0 31004 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_332
timestamp 1644511149
transform 1 0 31648 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_338
timestamp 1644511149
transform 1 0 32200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_360
timestamp 1644511149
transform 1 0 34224 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_28
timestamp 1644511149
transform 1 0 3680 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_40
timestamp 1644511149
transform 1 0 4784 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_52
timestamp 1644511149
transform 1 0 5888 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_69
timestamp 1644511149
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_81
timestamp 1644511149
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_93
timestamp 1644511149
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1644511149
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1644511149
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_113
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_125
timestamp 1644511149
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_137
timestamp 1644511149
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_149
timestamp 1644511149
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1644511149
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1644511149
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_169
timestamp 1644511149
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_181
timestamp 1644511149
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_193
timestamp 1644511149
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_205
timestamp 1644511149
transform 1 0 19964 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_211
timestamp 1644511149
transform 1 0 20516 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_215
timestamp 1644511149
transform 1 0 20884 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1644511149
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_225
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_235
timestamp 1644511149
transform 1 0 22724 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_246
timestamp 1644511149
transform 1 0 23736 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_255
timestamp 1644511149
transform 1 0 24564 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_269
timestamp 1644511149
transform 1 0 25852 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_276
timestamp 1644511149
transform 1 0 26496 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_281
timestamp 1644511149
transform 1 0 26956 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_288
timestamp 1644511149
transform 1 0 27600 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_297
timestamp 1644511149
transform 1 0 28428 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_305
timestamp 1644511149
transform 1 0 29164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_322
timestamp 1644511149
transform 1 0 30728 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1644511149
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1644511149
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_340
timestamp 1644511149
transform 1 0 32384 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_351
timestamp 1644511149
transform 1 0 33396 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_355
timestamp 1644511149
transform 1 0 33764 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_359
timestamp 1644511149
transform 1 0 34132 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_363
timestamp 1644511149
transform 1 0 34500 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_3
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_10
timestamp 1644511149
transform 1 0 2024 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_22
timestamp 1644511149
transform 1 0 3128 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_41
timestamp 1644511149
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_53
timestamp 1644511149
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_65
timestamp 1644511149
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1644511149
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1644511149
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_85
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_97
timestamp 1644511149
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_109
timestamp 1644511149
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_121
timestamp 1644511149
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1644511149
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1644511149
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_141
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_153
timestamp 1644511149
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_165
timestamp 1644511149
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_177
timestamp 1644511149
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1644511149
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1644511149
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_197
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_209
timestamp 1644511149
transform 1 0 20332 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_213
timestamp 1644511149
transform 1 0 20700 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_223
timestamp 1644511149
transform 1 0 21620 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_234
timestamp 1644511149
transform 1 0 22632 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_247
timestamp 1644511149
transform 1 0 23828 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1644511149
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_260
timestamp 1644511149
transform 1 0 25024 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_268
timestamp 1644511149
transform 1 0 25760 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_275
timestamp 1644511149
transform 1 0 26404 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_286
timestamp 1644511149
transform 1 0 27416 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_296
timestamp 1644511149
transform 1 0 28336 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_304
timestamp 1644511149
transform 1 0 29072 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_315
timestamp 1644511149
transform 1 0 30084 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_323
timestamp 1644511149
transform 1 0 30820 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_330
timestamp 1644511149
transform 1 0 31464 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_338
timestamp 1644511149
transform 1 0 32200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_360
timestamp 1644511149
transform 1 0 34224 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1644511149
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1644511149
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1644511149
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1644511149
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1644511149
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_57
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_69
timestamp 1644511149
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_81
timestamp 1644511149
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_93
timestamp 1644511149
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1644511149
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1644511149
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_113
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_125
timestamp 1644511149
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_137
timestamp 1644511149
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_149
timestamp 1644511149
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1644511149
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1644511149
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_169
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_181
timestamp 1644511149
transform 1 0 17756 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_190
timestamp 1644511149
transform 1 0 18584 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_202
timestamp 1644511149
transform 1 0 19688 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_213
timestamp 1644511149
transform 1 0 20700 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_220
timestamp 1644511149
transform 1 0 21344 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_229
timestamp 1644511149
transform 1 0 22172 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_240
timestamp 1644511149
transform 1 0 23184 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_252
timestamp 1644511149
transform 1 0 24288 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_266
timestamp 1644511149
transform 1 0 25576 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_276
timestamp 1644511149
transform 1 0 26496 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_290
timestamp 1644511149
transform 1 0 27784 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_302
timestamp 1644511149
transform 1 0 28888 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_311
timestamp 1644511149
transform 1 0 29716 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_319
timestamp 1644511149
transform 1 0 30452 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_327
timestamp 1644511149
transform 1 0 31188 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1644511149
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_337
timestamp 1644511149
transform 1 0 32108 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_360
timestamp 1644511149
transform 1 0 34224 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1644511149
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1644511149
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_41
timestamp 1644511149
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_53
timestamp 1644511149
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_65
timestamp 1644511149
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1644511149
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1644511149
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_85
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_97
timestamp 1644511149
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_109
timestamp 1644511149
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_121
timestamp 1644511149
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1644511149
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1644511149
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_141
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_153
timestamp 1644511149
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_165
timestamp 1644511149
transform 1 0 16284 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_176
timestamp 1644511149
transform 1 0 17296 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_183
timestamp 1644511149
transform 1 0 17940 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_192
timestamp 1644511149
transform 1 0 18768 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_197
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_206
timestamp 1644511149
transform 1 0 20056 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_213
timestamp 1644511149
transform 1 0 20700 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_233
timestamp 1644511149
transform 1 0 22540 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1644511149
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1644511149
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_253
timestamp 1644511149
transform 1 0 24380 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_260
timestamp 1644511149
transform 1 0 25024 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_280
timestamp 1644511149
transform 1 0 26864 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_291
timestamp 1644511149
transform 1 0 27876 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1644511149
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1644511149
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_325
timestamp 1644511149
transform 1 0 31004 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_333
timestamp 1644511149
transform 1 0 31740 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_340
timestamp 1644511149
transform 1 0 32384 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_348
timestamp 1644511149
transform 1 0 33120 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_352
timestamp 1644511149
transform 1 0 33488 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_359
timestamp 1644511149
transform 1 0 34132 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1644511149
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1644511149
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1644511149
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1644511149
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1644511149
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1644511149
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1644511149
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_57
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_69
timestamp 1644511149
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_81
timestamp 1644511149
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_93
timestamp 1644511149
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1644511149
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1644511149
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_113
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_125
timestamp 1644511149
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_137
timestamp 1644511149
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_149
timestamp 1644511149
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1644511149
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1644511149
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_169
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_180
timestamp 1644511149
transform 1 0 17664 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_200
timestamp 1644511149
transform 1 0 19504 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_220
timestamp 1644511149
transform 1 0 21344 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_230
timestamp 1644511149
transform 1 0 22264 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_240
timestamp 1644511149
transform 1 0 23184 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_250
timestamp 1644511149
transform 1 0 24104 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_262
timestamp 1644511149
transform 1 0 25208 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1644511149
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1644511149
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_281
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_292
timestamp 1644511149
transform 1 0 27968 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_300
timestamp 1644511149
transform 1 0 28704 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_311
timestamp 1644511149
transform 1 0 29716 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_319
timestamp 1644511149
transform 1 0 30452 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_327
timestamp 1644511149
transform 1 0 31188 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1644511149
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_341
timestamp 1644511149
transform 1 0 32476 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_349
timestamp 1644511149
transform 1 0 33212 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_353
timestamp 1644511149
transform 1 0 33580 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_360
timestamp 1644511149
transform 1 0 34224 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1644511149
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1644511149
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_41
timestamp 1644511149
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_53
timestamp 1644511149
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_65
timestamp 1644511149
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1644511149
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1644511149
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_85
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_97
timestamp 1644511149
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_109
timestamp 1644511149
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_121
timestamp 1644511149
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1644511149
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1644511149
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_141
timestamp 1644511149
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_153
timestamp 1644511149
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_165
timestamp 1644511149
transform 1 0 16284 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_182
timestamp 1644511149
transform 1 0 17848 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_191
timestamp 1644511149
transform 1 0 18676 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1644511149
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_203
timestamp 1644511149
transform 1 0 19780 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_212
timestamp 1644511149
transform 1 0 20608 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_220
timestamp 1644511149
transform 1 0 21344 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_231
timestamp 1644511149
transform 1 0 22356 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1644511149
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1644511149
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_260
timestamp 1644511149
transform 1 0 25024 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_267
timestamp 1644511149
transform 1 0 25668 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_287
timestamp 1644511149
transform 1 0 27508 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_298
timestamp 1644511149
transform 1 0 28520 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_306
timestamp 1644511149
transform 1 0 29256 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_314
timestamp 1644511149
transform 1 0 29992 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_322
timestamp 1644511149
transform 1 0 30728 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_330
timestamp 1644511149
transform 1 0 31464 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_338
timestamp 1644511149
transform 1 0 32200 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_346
timestamp 1644511149
transform 1 0 32936 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_352
timestamp 1644511149
transform 1 0 33488 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_356
timestamp 1644511149
transform 1 0 33856 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1644511149
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1644511149
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1644511149
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1644511149
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1644511149
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_57
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_69
timestamp 1644511149
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_81
timestamp 1644511149
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_93
timestamp 1644511149
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1644511149
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1644511149
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_113
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_125
timestamp 1644511149
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_137
timestamp 1644511149
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_149
timestamp 1644511149
transform 1 0 14812 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_155
timestamp 1644511149
transform 1 0 15364 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_164
timestamp 1644511149
transform 1 0 16192 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_185
timestamp 1644511149
transform 1 0 18124 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_193
timestamp 1644511149
transform 1 0 18860 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_202
timestamp 1644511149
transform 1 0 19688 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_210
timestamp 1644511149
transform 1 0 20424 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_220
timestamp 1644511149
transform 1 0 21344 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_225
timestamp 1644511149
transform 1 0 21804 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_245
timestamp 1644511149
transform 1 0 23644 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_252
timestamp 1644511149
transform 1 0 24288 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_264
timestamp 1644511149
transform 1 0 25392 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_275
timestamp 1644511149
transform 1 0 26404 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1644511149
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_37_281
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_294
timestamp 1644511149
transform 1 0 28152 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_301
timestamp 1644511149
transform 1 0 28796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_321
timestamp 1644511149
transform 1 0 30636 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1644511149
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1644511149
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_341
timestamp 1644511149
transform 1 0 32476 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_349
timestamp 1644511149
transform 1 0 33212 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_357
timestamp 1644511149
transform 1 0 33948 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_363
timestamp 1644511149
transform 1 0 34500 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1644511149
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1644511149
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1644511149
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_41
timestamp 1644511149
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_53
timestamp 1644511149
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_65
timestamp 1644511149
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1644511149
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1644511149
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_85
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_97
timestamp 1644511149
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_109
timestamp 1644511149
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_121
timestamp 1644511149
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1644511149
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1644511149
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_141
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_148
timestamp 1644511149
transform 1 0 14720 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_155
timestamp 1644511149
transform 1 0 15364 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_164
timestamp 1644511149
transform 1 0 16192 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_184
timestamp 1644511149
transform 1 0 18032 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_192
timestamp 1644511149
transform 1 0 18768 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_213
timestamp 1644511149
transform 1 0 20700 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_221
timestamp 1644511149
transform 1 0 21436 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_234
timestamp 1644511149
transform 1 0 22632 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_248
timestamp 1644511149
transform 1 0 23920 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_253
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_257
timestamp 1644511149
transform 1 0 24748 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_265
timestamp 1644511149
transform 1 0 25484 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_287
timestamp 1644511149
transform 1 0 27508 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_298
timestamp 1644511149
transform 1 0 28520 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_306
timestamp 1644511149
transform 1 0 29256 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_325
timestamp 1644511149
transform 1 0 31004 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_333
timestamp 1644511149
transform 1 0 31740 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_360
timestamp 1644511149
transform 1 0 34224 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1644511149
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_27
timestamp 1644511149
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_39
timestamp 1644511149
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1644511149
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1644511149
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_69
timestamp 1644511149
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_81
timestamp 1644511149
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_93
timestamp 1644511149
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1644511149
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1644511149
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_113
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_125
timestamp 1644511149
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_137
timestamp 1644511149
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_152
timestamp 1644511149
transform 1 0 15088 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_158
timestamp 1644511149
transform 1 0 15640 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_164
timestamp 1644511149
transform 1 0 16192 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_169
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_180
timestamp 1644511149
transform 1 0 17664 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_200
timestamp 1644511149
transform 1 0 19504 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_220
timestamp 1644511149
transform 1 0 21344 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_233
timestamp 1644511149
transform 1 0 22540 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_244
timestamp 1644511149
transform 1 0 23552 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_254
timestamp 1644511149
transform 1 0 24472 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_39_271
timestamp 1644511149
transform 1 0 26036 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1644511149
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_281
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_288
timestamp 1644511149
transform 1 0 27600 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_292
timestamp 1644511149
transform 1 0 27968 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_299
timestamp 1644511149
transform 1 0 28612 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_313
timestamp 1644511149
transform 1 0 29900 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_321
timestamp 1644511149
transform 1 0 30636 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_327
timestamp 1644511149
transform 1 0 31188 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1644511149
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_337
timestamp 1644511149
transform 1 0 32108 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_360
timestamp 1644511149
transform 1 0 34224 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1644511149
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1644511149
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1644511149
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_41
timestamp 1644511149
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_53
timestamp 1644511149
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_65
timestamp 1644511149
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1644511149
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1644511149
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_85
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_97
timestamp 1644511149
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_109
timestamp 1644511149
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_121
timestamp 1644511149
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1644511149
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1644511149
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_141
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_147
timestamp 1644511149
transform 1 0 14628 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_151
timestamp 1644511149
transform 1 0 14996 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_159
timestamp 1644511149
transform 1 0 15732 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_179
timestamp 1644511149
transform 1 0 17572 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1644511149
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1644511149
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_207
timestamp 1644511149
transform 1 0 20148 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_215
timestamp 1644511149
transform 1 0 20884 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_222
timestamp 1644511149
transform 1 0 21528 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_226
timestamp 1644511149
transform 1 0 21896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_233
timestamp 1644511149
transform 1 0 22540 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_237
timestamp 1644511149
transform 1 0 22908 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_244
timestamp 1644511149
transform 1 0 23552 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_253
timestamp 1644511149
transform 1 0 24380 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_272
timestamp 1644511149
transform 1 0 26128 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_281
timestamp 1644511149
transform 1 0 26956 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_287
timestamp 1644511149
transform 1 0 27508 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_304
timestamp 1644511149
transform 1 0 29072 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_313
timestamp 1644511149
transform 1 0 29900 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_317
timestamp 1644511149
transform 1 0 30268 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_334
timestamp 1644511149
transform 1 0 31832 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_338
timestamp 1644511149
transform 1 0 32200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_360
timestamp 1644511149
transform 1 0 34224 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_3
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_7
timestamp 1644511149
transform 1 0 1748 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_11
timestamp 1644511149
transform 1 0 2116 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_15
timestamp 1644511149
transform 1 0 2484 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_19
timestamp 1644511149
transform 1 0 2852 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_31
timestamp 1644511149
transform 1 0 3956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_43
timestamp 1644511149
transform 1 0 5060 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1644511149
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_69
timestamp 1644511149
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_81
timestamp 1644511149
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_93
timestamp 1644511149
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1644511149
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1644511149
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_113
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_125
timestamp 1644511149
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_140
timestamp 1644511149
transform 1 0 13984 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_147
timestamp 1644511149
transform 1 0 14628 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_155
timestamp 1644511149
transform 1 0 15364 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_164
timestamp 1644511149
transform 1 0 16192 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_169
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_180
timestamp 1644511149
transform 1 0 17664 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_200
timestamp 1644511149
transform 1 0 19504 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_208
timestamp 1644511149
transform 1 0 20240 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_220
timestamp 1644511149
transform 1 0 21344 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_230
timestamp 1644511149
transform 1 0 22264 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_239
timestamp 1644511149
transform 1 0 23092 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_41_255
timestamp 1644511149
transform 1 0 24564 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_269
timestamp 1644511149
transform 1 0 25852 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_276
timestamp 1644511149
transform 1 0 26496 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_281
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_286
timestamp 1644511149
transform 1 0 27416 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_295
timestamp 1644511149
transform 1 0 28244 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_303
timestamp 1644511149
transform 1 0 28980 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_312
timestamp 1644511149
transform 1 0 29808 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_332
timestamp 1644511149
transform 1 0 31648 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_353
timestamp 1644511149
transform 1 0 33580 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_360
timestamp 1644511149
transform 1 0 34224 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_24
timestamp 1644511149
transform 1 0 3312 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_41
timestamp 1644511149
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_53
timestamp 1644511149
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_65
timestamp 1644511149
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1644511149
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1644511149
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_85
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_97
timestamp 1644511149
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_109
timestamp 1644511149
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_121
timestamp 1644511149
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1644511149
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1644511149
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_42_141
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_147
timestamp 1644511149
transform 1 0 14628 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_155
timestamp 1644511149
transform 1 0 15364 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_175
timestamp 1644511149
transform 1 0 17204 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_183
timestamp 1644511149
transform 1 0 17940 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_192
timestamp 1644511149
transform 1 0 18768 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_197
timestamp 1644511149
transform 1 0 19228 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_201
timestamp 1644511149
transform 1 0 19596 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_207
timestamp 1644511149
transform 1 0 20148 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_213
timestamp 1644511149
transform 1 0 20700 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_230
timestamp 1644511149
transform 1 0 22264 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_239
timestamp 1644511149
transform 1 0 23092 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_248
timestamp 1644511149
transform 1 0 23920 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_258
timestamp 1644511149
transform 1 0 24840 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_262
timestamp 1644511149
transform 1 0 25208 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_267
timestamp 1644511149
transform 1 0 25668 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_276
timestamp 1644511149
transform 1 0 26496 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_286
timestamp 1644511149
transform 1 0 27416 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_294
timestamp 1644511149
transform 1 0 28152 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_298
timestamp 1644511149
transform 1 0 28520 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_304
timestamp 1644511149
transform 1 0 29072 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_325
timestamp 1644511149
transform 1 0 31004 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_335
timestamp 1644511149
transform 1 0 31924 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_360
timestamp 1644511149
transform 1 0 34224 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1644511149
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1644511149
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_39
timestamp 1644511149
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1644511149
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1644511149
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_57
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_69
timestamp 1644511149
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_81
timestamp 1644511149
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_93
timestamp 1644511149
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1644511149
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1644511149
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_113
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_125
timestamp 1644511149
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_137
timestamp 1644511149
transform 1 0 13708 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_141
timestamp 1644511149
transform 1 0 14076 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_148
timestamp 1644511149
transform 1 0 14720 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_156
timestamp 1644511149
transform 1 0 15456 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_164
timestamp 1644511149
transform 1 0 16192 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_169
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_173
timestamp 1644511149
transform 1 0 17020 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_190
timestamp 1644511149
transform 1 0 18584 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_198
timestamp 1644511149
transform 1 0 19320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_215
timestamp 1644511149
transform 1 0 20884 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1644511149
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_43_225
timestamp 1644511149
transform 1 0 21804 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_242
timestamp 1644511149
transform 1 0 23368 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_262
timestamp 1644511149
transform 1 0 25208 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_272
timestamp 1644511149
transform 1 0 26128 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_43_287
timestamp 1644511149
transform 1 0 27508 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_295
timestamp 1644511149
transform 1 0 28244 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_312
timestamp 1644511149
transform 1 0 29808 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_321
timestamp 1644511149
transform 1 0 30636 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_325
timestamp 1644511149
transform 1 0 31004 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_332
timestamp 1644511149
transform 1 0 31648 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_337
timestamp 1644511149
transform 1 0 32108 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_360
timestamp 1644511149
transform 1 0 34224 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1644511149
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1644511149
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_41
timestamp 1644511149
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_53
timestamp 1644511149
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_65
timestamp 1644511149
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1644511149
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1644511149
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_85
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_97
timestamp 1644511149
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_109
timestamp 1644511149
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_121
timestamp 1644511149
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1644511149
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1644511149
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_141
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_146
timestamp 1644511149
transform 1 0 14536 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_153
timestamp 1644511149
transform 1 0 15180 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_173
timestamp 1644511149
transform 1 0 17020 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_183
timestamp 1644511149
transform 1 0 17940 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_192
timestamp 1644511149
transform 1 0 18768 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_213
timestamp 1644511149
transform 1 0 20700 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_223
timestamp 1644511149
transform 1 0 21620 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_237
timestamp 1644511149
transform 1 0 22908 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_246
timestamp 1644511149
transform 1 0 23736 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_253
timestamp 1644511149
transform 1 0 24380 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_257
timestamp 1644511149
transform 1 0 24748 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_274
timestamp 1644511149
transform 1 0 26312 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_294
timestamp 1644511149
transform 1 0 28152 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_298
timestamp 1644511149
transform 1 0 28520 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_304
timestamp 1644511149
transform 1 0 29072 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_309
timestamp 1644511149
transform 1 0 29532 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_320
timestamp 1644511149
transform 1 0 30544 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_330
timestamp 1644511149
transform 1 0 31464 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_338
timestamp 1644511149
transform 1 0 32200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_355
timestamp 1644511149
transform 1 0 33764 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1644511149
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1644511149
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1644511149
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_27
timestamp 1644511149
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_39
timestamp 1644511149
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1644511149
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1644511149
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_69
timestamp 1644511149
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_81
timestamp 1644511149
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_93
timestamp 1644511149
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1644511149
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1644511149
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_113
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_125
timestamp 1644511149
transform 1 0 12604 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_136
timestamp 1644511149
transform 1 0 13616 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_143
timestamp 1644511149
transform 1 0 14260 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_150
timestamp 1644511149
transform 1 0 14904 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_157
timestamp 1644511149
transform 1 0 15548 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_164
timestamp 1644511149
transform 1 0 16192 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_173
timestamp 1644511149
transform 1 0 17020 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_184
timestamp 1644511149
transform 1 0 18032 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_190
timestamp 1644511149
transform 1 0 18584 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_199
timestamp 1644511149
transform 1 0 19412 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_203
timestamp 1644511149
transform 1 0 19780 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_220
timestamp 1644511149
transform 1 0 21344 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_225
timestamp 1644511149
transform 1 0 21804 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_235
timestamp 1644511149
transform 1 0 22724 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_243
timestamp 1644511149
transform 1 0 23460 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_263
timestamp 1644511149
transform 1 0 25300 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_272
timestamp 1644511149
transform 1 0 26128 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_297
timestamp 1644511149
transform 1 0 28428 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_307
timestamp 1644511149
transform 1 0 29348 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_321
timestamp 1644511149
transform 1 0 30636 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_332
timestamp 1644511149
transform 1 0 31648 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_340
timestamp 1644511149
transform 1 0 32384 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_353
timestamp 1644511149
transform 1 0 33580 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_360
timestamp 1644511149
transform 1 0 34224 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1644511149
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1644511149
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_41
timestamp 1644511149
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_53
timestamp 1644511149
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_65
timestamp 1644511149
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1644511149
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1644511149
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_85
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_97
timestamp 1644511149
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_109
timestamp 1644511149
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_121
timestamp 1644511149
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_136
timestamp 1644511149
transform 1 0 13616 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_141
timestamp 1644511149
transform 1 0 14076 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_150
timestamp 1644511149
transform 1 0 14904 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_157
timestamp 1644511149
transform 1 0 15548 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_161
timestamp 1644511149
transform 1 0 15916 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_165
timestamp 1644511149
transform 1 0 16284 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_174
timestamp 1644511149
transform 1 0 17112 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_183
timestamp 1644511149
transform 1 0 17940 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_192
timestamp 1644511149
transform 1 0 18768 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_203
timestamp 1644511149
transform 1 0 19780 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_211
timestamp 1644511149
transform 1 0 20516 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_220
timestamp 1644511149
transform 1 0 21344 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_234
timestamp 1644511149
transform 1 0 22632 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_242
timestamp 1644511149
transform 1 0 23368 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_248
timestamp 1644511149
transform 1 0 23920 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_260
timestamp 1644511149
transform 1 0 25024 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_268
timestamp 1644511149
transform 1 0 25760 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_277
timestamp 1644511149
transform 1 0 26588 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_285
timestamp 1644511149
transform 1 0 27324 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_293
timestamp 1644511149
transform 1 0 28060 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_297
timestamp 1644511149
transform 1 0 28428 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_304
timestamp 1644511149
transform 1 0 29072 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_319
timestamp 1644511149
transform 1 0 30452 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_327
timestamp 1644511149
transform 1 0 31188 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_340
timestamp 1644511149
transform 1 0 32384 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_360
timestamp 1644511149
transform 1 0 34224 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1644511149
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1644511149
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1644511149
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_39
timestamp 1644511149
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1644511149
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1644511149
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_69
timestamp 1644511149
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_81
timestamp 1644511149
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_93
timestamp 1644511149
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1644511149
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1644511149
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_113
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_125
timestamp 1644511149
transform 1 0 12604 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_131
timestamp 1644511149
transform 1 0 13156 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_135
timestamp 1644511149
transform 1 0 13524 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_142
timestamp 1644511149
transform 1 0 14168 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_149
timestamp 1644511149
transform 1 0 14812 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_156
timestamp 1644511149
transform 1 0 15456 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_164
timestamp 1644511149
transform 1 0 16192 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_47_169
timestamp 1644511149
transform 1 0 16652 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_47_177
timestamp 1644511149
transform 1 0 17388 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_183
timestamp 1644511149
transform 1 0 17940 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_200
timestamp 1644511149
transform 1 0 19504 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_220
timestamp 1644511149
transform 1 0 21344 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_225
timestamp 1644511149
transform 1 0 21804 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_231
timestamp 1644511149
transform 1 0 22356 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_243
timestamp 1644511149
transform 1 0 23460 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_253
timestamp 1644511149
transform 1 0 24380 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_266
timestamp 1644511149
transform 1 0 25576 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_275
timestamp 1644511149
transform 1 0 26404 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1644511149
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_288
timestamp 1644511149
transform 1 0 27600 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_294
timestamp 1644511149
transform 1 0 28152 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_311
timestamp 1644511149
transform 1 0 29716 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_322
timestamp 1644511149
transform 1 0 30728 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_332
timestamp 1644511149
transform 1 0 31648 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_337
timestamp 1644511149
transform 1 0 32108 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_360
timestamp 1644511149
transform 1 0 34224 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1644511149
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1644511149
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1644511149
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1644511149
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_53
timestamp 1644511149
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_65
timestamp 1644511149
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1644511149
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1644511149
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_85
timestamp 1644511149
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_97
timestamp 1644511149
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_109
timestamp 1644511149
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_121
timestamp 1644511149
transform 1 0 12236 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_125
timestamp 1644511149
transform 1 0 12604 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_129
timestamp 1644511149
transform 1 0 12972 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_136
timestamp 1644511149
transform 1 0 13616 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_141
timestamp 1644511149
transform 1 0 14076 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_150
timestamp 1644511149
transform 1 0 14904 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_157
timestamp 1644511149
transform 1 0 15548 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_181
timestamp 1644511149
transform 1 0 17756 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_192
timestamp 1644511149
transform 1 0 18768 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_213
timestamp 1644511149
transform 1 0 20700 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_223
timestamp 1644511149
transform 1 0 21620 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_231
timestamp 1644511149
transform 1 0 22356 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_248
timestamp 1644511149
transform 1 0 23920 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_253
timestamp 1644511149
transform 1 0 24380 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_277
timestamp 1644511149
transform 1 0 26588 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_293
timestamp 1644511149
transform 1 0 28060 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_297
timestamp 1644511149
transform 1 0 28428 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_304
timestamp 1644511149
transform 1 0 29072 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_309
timestamp 1644511149
transform 1 0 29532 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_331
timestamp 1644511149
transform 1 0 31556 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_343
timestamp 1644511149
transform 1 0 32660 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1644511149
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1644511149
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1644511149
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_15
timestamp 1644511149
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_27
timestamp 1644511149
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_39
timestamp 1644511149
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1644511149
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1644511149
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_69
timestamp 1644511149
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_81
timestamp 1644511149
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_93
timestamp 1644511149
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1644511149
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1644511149
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_113
timestamp 1644511149
transform 1 0 11500 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_117
timestamp 1644511149
transform 1 0 11868 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_121
timestamp 1644511149
transform 1 0 12236 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_125
timestamp 1644511149
transform 1 0 12604 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_135
timestamp 1644511149
transform 1 0 13524 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_142
timestamp 1644511149
transform 1 0 14168 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_149
timestamp 1644511149
transform 1 0 14812 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_156
timestamp 1644511149
transform 1 0 15456 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_164
timestamp 1644511149
transform 1 0 16192 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_49_169
timestamp 1644511149
transform 1 0 16652 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_188
timestamp 1644511149
transform 1 0 18400 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_197
timestamp 1644511149
transform 1 0 19228 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_206
timestamp 1644511149
transform 1 0 20056 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_214
timestamp 1644511149
transform 1 0 20792 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_220
timestamp 1644511149
transform 1 0 21344 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_230
timestamp 1644511149
transform 1 0 22264 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_234
timestamp 1644511149
transform 1 0 22632 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_243
timestamp 1644511149
transform 1 0 23460 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_249
timestamp 1644511149
transform 1 0 24012 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_266
timestamp 1644511149
transform 1 0 25576 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_276
timestamp 1644511149
transform 1 0 26496 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_297
timestamp 1644511149
transform 1 0 28428 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_317
timestamp 1644511149
transform 1 0 30268 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_332
timestamp 1644511149
transform 1 0 31648 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_341
timestamp 1644511149
transform 1 0 32476 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_353
timestamp 1644511149
transform 1 0 33580 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_360
timestamp 1644511149
transform 1 0 34224 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_3
timestamp 1644511149
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_15
timestamp 1644511149
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1644511149
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_29
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_41
timestamp 1644511149
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_53
timestamp 1644511149
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_65
timestamp 1644511149
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1644511149
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1644511149
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_85
timestamp 1644511149
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_97
timestamp 1644511149
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_109
timestamp 1644511149
transform 1 0 11132 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_117
timestamp 1644511149
transform 1 0 11868 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_122
timestamp 1644511149
transform 1 0 12328 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_129
timestamp 1644511149
transform 1 0 12972 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_136
timestamp 1644511149
transform 1 0 13616 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_144
timestamp 1644511149
transform 1 0 14352 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_151
timestamp 1644511149
transform 1 0 14996 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_158
timestamp 1644511149
transform 1 0 15640 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_178
timestamp 1644511149
transform 1 0 17480 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_187
timestamp 1644511149
transform 1 0 18308 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1644511149
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_50_197
timestamp 1644511149
transform 1 0 19228 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_216
timestamp 1644511149
transform 1 0 20976 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_228
timestamp 1644511149
transform 1 0 22080 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_238
timestamp 1644511149
transform 1 0 23000 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_247
timestamp 1644511149
transform 1 0 23828 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1644511149
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_258
timestamp 1644511149
transform 1 0 24840 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_262
timestamp 1644511149
transform 1 0 25208 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_268
timestamp 1644511149
transform 1 0 25760 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_279
timestamp 1644511149
transform 1 0 26772 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_290
timestamp 1644511149
transform 1 0 27784 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_304
timestamp 1644511149
transform 1 0 29072 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_316
timestamp 1644511149
transform 1 0 30176 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_324
timestamp 1644511149
transform 1 0 30912 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_333
timestamp 1644511149
transform 1 0 31740 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_340
timestamp 1644511149
transform 1 0 32384 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_360
timestamp 1644511149
transform 1 0 34224 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1644511149
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_15
timestamp 1644511149
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_27
timestamp 1644511149
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_39
timestamp 1644511149
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1644511149
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1644511149
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_69
timestamp 1644511149
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_81
timestamp 1644511149
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_93
timestamp 1644511149
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1644511149
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1644511149
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_113
timestamp 1644511149
transform 1 0 11500 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_120
timestamp 1644511149
transform 1 0 12144 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_127
timestamp 1644511149
transform 1 0 12788 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_134
timestamp 1644511149
transform 1 0 13432 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_141
timestamp 1644511149
transform 1 0 14076 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_148
timestamp 1644511149
transform 1 0 14720 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_156
timestamp 1644511149
transform 1 0 15456 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_164
timestamp 1644511149
transform 1 0 16192 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_51_169
timestamp 1644511149
transform 1 0 16652 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_176
timestamp 1644511149
transform 1 0 17296 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_196
timestamp 1644511149
transform 1 0 19136 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_216
timestamp 1644511149
transform 1 0 20976 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_233
timestamp 1644511149
transform 1 0 22540 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_244
timestamp 1644511149
transform 1 0 23552 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_251
timestamp 1644511149
transform 1 0 24196 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_262
timestamp 1644511149
transform 1 0 25208 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_270
timestamp 1644511149
transform 1 0 25944 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_276
timestamp 1644511149
transform 1 0 26496 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_281
timestamp 1644511149
transform 1 0 26956 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_288
timestamp 1644511149
transform 1 0 27600 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_308
timestamp 1644511149
transform 1 0 29440 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_312
timestamp 1644511149
transform 1 0 29808 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_321
timestamp 1644511149
transform 1 0 30636 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_325
timestamp 1644511149
transform 1 0 31004 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_332
timestamp 1644511149
transform 1 0 31648 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_337
timestamp 1644511149
transform 1 0 32108 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_346
timestamp 1644511149
transform 1 0 32936 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_356
timestamp 1644511149
transform 1 0 33856 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_3
timestamp 1644511149
transform 1 0 1380 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_10
timestamp 1644511149
transform 1 0 2024 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_22
timestamp 1644511149
transform 1 0 3128 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_52_29
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_41
timestamp 1644511149
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_53
timestamp 1644511149
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_65
timestamp 1644511149
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1644511149
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1644511149
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_85
timestamp 1644511149
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_97
timestamp 1644511149
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_109
timestamp 1644511149
transform 1 0 11132 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_115
timestamp 1644511149
transform 1 0 11684 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_122
timestamp 1644511149
transform 1 0 12328 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_129
timestamp 1644511149
transform 1 0 12972 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_136
timestamp 1644511149
transform 1 0 13616 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_141
timestamp 1644511149
transform 1 0 14076 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_151
timestamp 1644511149
transform 1 0 14996 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_159
timestamp 1644511149
transform 1 0 15732 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_168
timestamp 1644511149
transform 1 0 16560 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_192
timestamp 1644511149
transform 1 0 18768 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_202
timestamp 1644511149
transform 1 0 19688 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_206
timestamp 1644511149
transform 1 0 20056 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_211
timestamp 1644511149
transform 1 0 20516 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_223
timestamp 1644511149
transform 1 0 21620 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_234
timestamp 1644511149
transform 1 0 22632 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1644511149
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1644511149
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_253
timestamp 1644511149
transform 1 0 24380 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_262
timestamp 1644511149
transform 1 0 25208 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_272
timestamp 1644511149
transform 1 0 26128 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_292
timestamp 1644511149
transform 1 0 27968 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_296
timestamp 1644511149
transform 1 0 28336 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_304
timestamp 1644511149
transform 1 0 29072 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_309
timestamp 1644511149
transform 1 0 29532 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_331
timestamp 1644511149
transform 1 0 31556 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_342
timestamp 1644511149
transform 1 0 32568 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_352
timestamp 1644511149
transform 1 0 33488 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_360
timestamp 1644511149
transform 1 0 34224 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_3
timestamp 1644511149
transform 1 0 1380 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_25
timestamp 1644511149
transform 1 0 3404 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_37
timestamp 1644511149
transform 1 0 4508 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_49
timestamp 1644511149
transform 1 0 5612 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1644511149
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_57
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_69
timestamp 1644511149
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_81
timestamp 1644511149
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_93
timestamp 1644511149
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1644511149
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1644511149
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_113
timestamp 1644511149
transform 1 0 11500 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_122
timestamp 1644511149
transform 1 0 12328 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_126
timestamp 1644511149
transform 1 0 12696 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_130
timestamp 1644511149
transform 1 0 13064 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_137
timestamp 1644511149
transform 1 0 13708 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_144
timestamp 1644511149
transform 1 0 14352 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_164
timestamp 1644511149
transform 1 0 16192 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_173
timestamp 1644511149
transform 1 0 17020 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_182
timestamp 1644511149
transform 1 0 17848 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_192
timestamp 1644511149
transform 1 0 18768 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_204
timestamp 1644511149
transform 1 0 19872 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_212
timestamp 1644511149
transform 1 0 20608 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_220
timestamp 1644511149
transform 1 0 21344 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_232
timestamp 1644511149
transform 1 0 22448 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_239
timestamp 1644511149
transform 1 0 23092 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_250
timestamp 1644511149
transform 1 0 24104 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_262
timestamp 1644511149
transform 1 0 25208 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1644511149
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1644511149
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_281
timestamp 1644511149
transform 1 0 26956 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_53_308
timestamp 1644511149
transform 1 0 29440 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_323
timestamp 1644511149
transform 1 0 30820 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_332
timestamp 1644511149
transform 1 0 31648 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_337
timestamp 1644511149
transform 1 0 32108 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_360
timestamp 1644511149
transform 1 0 34224 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_3
timestamp 1644511149
transform 1 0 1380 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_7
timestamp 1644511149
transform 1 0 1748 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_19
timestamp 1644511149
transform 1 0 2852 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1644511149
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_29
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_41
timestamp 1644511149
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_53
timestamp 1644511149
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_65
timestamp 1644511149
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1644511149
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1644511149
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_85
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_97
timestamp 1644511149
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_109
timestamp 1644511149
transform 1 0 11132 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_116
timestamp 1644511149
transform 1 0 11776 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_123
timestamp 1644511149
transform 1 0 12420 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_130
timestamp 1644511149
transform 1 0 13064 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_138
timestamp 1644511149
transform 1 0 13800 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_141
timestamp 1644511149
transform 1 0 14076 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_145
timestamp 1644511149
transform 1 0 14444 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_150
timestamp 1644511149
transform 1 0 14904 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_170
timestamp 1644511149
transform 1 0 16744 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_181
timestamp 1644511149
transform 1 0 17756 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_185
timestamp 1644511149
transform 1 0 18124 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_192
timestamp 1644511149
transform 1 0 18768 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_54_197
timestamp 1644511149
transform 1 0 19228 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_54_204
timestamp 1644511149
transform 1 0 19872 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_210
timestamp 1644511149
transform 1 0 20424 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_217
timestamp 1644511149
transform 1 0 21068 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_225
timestamp 1644511149
transform 1 0 21804 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_234
timestamp 1644511149
transform 1 0 22632 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_248
timestamp 1644511149
transform 1 0 23920 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_261
timestamp 1644511149
transform 1 0 25116 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_271
timestamp 1644511149
transform 1 0 26036 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_283
timestamp 1644511149
transform 1 0 27140 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_294
timestamp 1644511149
transform 1 0 28152 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_304
timestamp 1644511149
transform 1 0 29072 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_309
timestamp 1644511149
transform 1 0 29532 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_54_322
timestamp 1644511149
transform 1 0 30728 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_335
timestamp 1644511149
transform 1 0 31924 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_360
timestamp 1644511149
transform 1 0 34224 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_3
timestamp 1644511149
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_15
timestamp 1644511149
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_27
timestamp 1644511149
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_39
timestamp 1644511149
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1644511149
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1644511149
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_69
timestamp 1644511149
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_81
timestamp 1644511149
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_93
timestamp 1644511149
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1644511149
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1644511149
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_55_113
timestamp 1644511149
transform 1 0 11500 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_117
timestamp 1644511149
transform 1 0 11868 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_124
timestamp 1644511149
transform 1 0 12512 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_131
timestamp 1644511149
transform 1 0 13156 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_138
timestamp 1644511149
transform 1 0 13800 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_145
timestamp 1644511149
transform 1 0 14444 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_154
timestamp 1644511149
transform 1 0 15272 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_164
timestamp 1644511149
transform 1 0 16192 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_173
timestamp 1644511149
transform 1 0 17020 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_185
timestamp 1644511149
transform 1 0 18124 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_205
timestamp 1644511149
transform 1 0 19964 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_211
timestamp 1644511149
transform 1 0 20516 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_220
timestamp 1644511149
transform 1 0 21344 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_232
timestamp 1644511149
transform 1 0 22448 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_239
timestamp 1644511149
transform 1 0 23092 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_259
timestamp 1644511149
transform 1 0 24932 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_267
timestamp 1644511149
transform 1 0 25668 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_276
timestamp 1644511149
transform 1 0 26496 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_281
timestamp 1644511149
transform 1 0 26956 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_291
timestamp 1644511149
transform 1 0 27876 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_302
timestamp 1644511149
transform 1 0 28888 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_313
timestamp 1644511149
transform 1 0 29900 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_321
timestamp 1644511149
transform 1 0 30636 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_332
timestamp 1644511149
transform 1 0 31648 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_337
timestamp 1644511149
transform 1 0 32108 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_360
timestamp 1644511149
transform 1 0 34224 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_3
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_15
timestamp 1644511149
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1644511149
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_29
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_41
timestamp 1644511149
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_53
timestamp 1644511149
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_65
timestamp 1644511149
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1644511149
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1644511149
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_85
timestamp 1644511149
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_97
timestamp 1644511149
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_109
timestamp 1644511149
transform 1 0 11132 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_117
timestamp 1644511149
transform 1 0 11868 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_122
timestamp 1644511149
transform 1 0 12328 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_129
timestamp 1644511149
transform 1 0 12972 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_136
timestamp 1644511149
transform 1 0 13616 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_141
timestamp 1644511149
transform 1 0 14076 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_148
timestamp 1644511149
transform 1 0 14720 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_168
timestamp 1644511149
transform 1 0 16560 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_192
timestamp 1644511149
transform 1 0 18768 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_213
timestamp 1644511149
transform 1 0 20700 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_219
timestamp 1644511149
transform 1 0 21252 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_229
timestamp 1644511149
transform 1 0 22172 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_239
timestamp 1644511149
transform 1 0 23092 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_248
timestamp 1644511149
transform 1 0 23920 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_253
timestamp 1644511149
transform 1 0 24380 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_258
timestamp 1644511149
transform 1 0 24840 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_267
timestamp 1644511149
transform 1 0 25668 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_276
timestamp 1644511149
transform 1 0 26496 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_290
timestamp 1644511149
transform 1 0 27784 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_303
timestamp 1644511149
transform 1 0 28980 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1644511149
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_312
timestamp 1644511149
transform 1 0 29808 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_323
timestamp 1644511149
transform 1 0 30820 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_329
timestamp 1644511149
transform 1 0 31372 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_339
timestamp 1644511149
transform 1 0 32292 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_359
timestamp 1644511149
transform 1 0 34132 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1644511149
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_3
timestamp 1644511149
transform 1 0 1380 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_7
timestamp 1644511149
transform 1 0 1748 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_11
timestamp 1644511149
transform 1 0 2116 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_18
timestamp 1644511149
transform 1 0 2760 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_30
timestamp 1644511149
transform 1 0 3864 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_42
timestamp 1644511149
transform 1 0 4968 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_54
timestamp 1644511149
transform 1 0 6072 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1644511149
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_81
timestamp 1644511149
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_93
timestamp 1644511149
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1644511149
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1644511149
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_113
timestamp 1644511149
transform 1 0 11500 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_122
timestamp 1644511149
transform 1 0 12328 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_129
timestamp 1644511149
transform 1 0 12972 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_136
timestamp 1644511149
transform 1 0 13616 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_140
timestamp 1644511149
transform 1 0 13984 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_144
timestamp 1644511149
transform 1 0 14352 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_164
timestamp 1644511149
transform 1 0 16192 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_174
timestamp 1644511149
transform 1 0 17112 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_180
timestamp 1644511149
transform 1 0 17664 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_186
timestamp 1644511149
transform 1 0 18216 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_195
timestamp 1644511149
transform 1 0 19044 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_201
timestamp 1644511149
transform 1 0 19596 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_207
timestamp 1644511149
transform 1 0 20148 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1644511149
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1644511149
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_232
timestamp 1644511149
transform 1 0 22448 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_241
timestamp 1644511149
transform 1 0 23276 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_245
timestamp 1644511149
transform 1 0 23644 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_248
timestamp 1644511149
transform 1 0 23920 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_266
timestamp 1644511149
transform 1 0 25576 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_270
timestamp 1644511149
transform 1 0 25944 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_276
timestamp 1644511149
transform 1 0 26496 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_281
timestamp 1644511149
transform 1 0 26956 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_285
timestamp 1644511149
transform 1 0 27324 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_294
timestamp 1644511149
transform 1 0 28152 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_305
timestamp 1644511149
transform 1 0 29164 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_309
timestamp 1644511149
transform 1 0 29532 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_318
timestamp 1644511149
transform 1 0 30360 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_332
timestamp 1644511149
transform 1 0 31648 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_337
timestamp 1644511149
transform 1 0 32108 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_360
timestamp 1644511149
transform 1 0 34224 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_24
timestamp 1644511149
transform 1 0 3312 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1644511149
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_41
timestamp 1644511149
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_53
timestamp 1644511149
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_65
timestamp 1644511149
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1644511149
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1644511149
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_85
timestamp 1644511149
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_97
timestamp 1644511149
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_109
timestamp 1644511149
transform 1 0 11132 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_117
timestamp 1644511149
transform 1 0 11868 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_122
timestamp 1644511149
transform 1 0 12328 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_129
timestamp 1644511149
transform 1 0 12972 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_136
timestamp 1644511149
transform 1 0 13616 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_144
timestamp 1644511149
transform 1 0 14352 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_151
timestamp 1644511149
transform 1 0 14996 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_158
timestamp 1644511149
transform 1 0 15640 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_165
timestamp 1644511149
transform 1 0 16284 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_185
timestamp 1644511149
transform 1 0 18124 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_192
timestamp 1644511149
transform 1 0 18768 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_213
timestamp 1644511149
transform 1 0 20700 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_221
timestamp 1644511149
transform 1 0 21436 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_229
timestamp 1644511149
transform 1 0 22172 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_237
timestamp 1644511149
transform 1 0 22908 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1644511149
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1644511149
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_58_253
timestamp 1644511149
transform 1 0 24380 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_259
timestamp 1644511149
transform 1 0 24932 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_279
timestamp 1644511149
transform 1 0 26772 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_299
timestamp 1644511149
transform 1 0 28612 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1644511149
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_318
timestamp 1644511149
transform 1 0 30360 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_330
timestamp 1644511149
transform 1 0 31464 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_338
timestamp 1644511149
transform 1 0 32200 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_360
timestamp 1644511149
transform 1 0 34224 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_3
timestamp 1644511149
transform 1 0 1380 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_8
timestamp 1644511149
transform 1 0 1840 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_15
timestamp 1644511149
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_27
timestamp 1644511149
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_39
timestamp 1644511149
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1644511149
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1644511149
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_69
timestamp 1644511149
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_81
timestamp 1644511149
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_93
timestamp 1644511149
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1644511149
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1644511149
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_113
timestamp 1644511149
transform 1 0 11500 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_122
timestamp 1644511149
transform 1 0 12328 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_129
timestamp 1644511149
transform 1 0 12972 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_136
timestamp 1644511149
transform 1 0 13616 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_143
timestamp 1644511149
transform 1 0 14260 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_150
timestamp 1644511149
transform 1 0 14904 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_157
timestamp 1644511149
transform 1 0 15548 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_164
timestamp 1644511149
transform 1 0 16192 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_174
timestamp 1644511149
transform 1 0 17112 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_184
timestamp 1644511149
transform 1 0 18032 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_193
timestamp 1644511149
transform 1 0 18860 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1644511149
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1644511149
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_59_225
timestamp 1644511149
transform 1 0 21804 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_244
timestamp 1644511149
transform 1 0 23552 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_264
timestamp 1644511149
transform 1 0 25392 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1644511149
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1644511149
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_285
timestamp 1644511149
transform 1 0 27324 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_295
timestamp 1644511149
transform 1 0 28244 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_305
timestamp 1644511149
transform 1 0 29164 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_309
timestamp 1644511149
transform 1 0 29532 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_326
timestamp 1644511149
transform 1 0 31096 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_334
timestamp 1644511149
transform 1 0 31832 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_345
timestamp 1644511149
transform 1 0 32844 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_355
timestamp 1644511149
transform 1 0 33764 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_363
timestamp 1644511149
transform 1 0 34500 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_24
timestamp 1644511149
transform 1 0 3312 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_29
timestamp 1644511149
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_41
timestamp 1644511149
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_53
timestamp 1644511149
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_65
timestamp 1644511149
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1644511149
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1644511149
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_85
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_97
timestamp 1644511149
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_109
timestamp 1644511149
transform 1 0 11132 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_120
timestamp 1644511149
transform 1 0 12144 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_127
timestamp 1644511149
transform 1 0 12788 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_134
timestamp 1644511149
transform 1 0 13432 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_60_141
timestamp 1644511149
transform 1 0 14076 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_146
timestamp 1644511149
transform 1 0 14536 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_153
timestamp 1644511149
transform 1 0 15180 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_173
timestamp 1644511149
transform 1 0 17020 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_184
timestamp 1644511149
transform 1 0 18032 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_192
timestamp 1644511149
transform 1 0 18768 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_205
timestamp 1644511149
transform 1 0 19964 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_214
timestamp 1644511149
transform 1 0 20792 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_238
timestamp 1644511149
transform 1 0 23000 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_248
timestamp 1644511149
transform 1 0 23920 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_261
timestamp 1644511149
transform 1 0 25116 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_283
timestamp 1644511149
transform 1 0 27140 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_295
timestamp 1644511149
transform 1 0 28244 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_304
timestamp 1644511149
transform 1 0 29072 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_315
timestamp 1644511149
transform 1 0 30084 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_335
timestamp 1644511149
transform 1 0 31924 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_360
timestamp 1644511149
transform 1 0 34224 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_7
timestamp 1644511149
transform 1 0 1748 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_14
timestamp 1644511149
transform 1 0 2392 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_20
timestamp 1644511149
transform 1 0 2944 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_25
timestamp 1644511149
transform 1 0 3404 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_32
timestamp 1644511149
transform 1 0 4048 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_39
timestamp 1644511149
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1644511149
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1644511149
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_57
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_69
timestamp 1644511149
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_81
timestamp 1644511149
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_93
timestamp 1644511149
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1644511149
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1644511149
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_113
timestamp 1644511149
transform 1 0 11500 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_120
timestamp 1644511149
transform 1 0 12144 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_127
timestamp 1644511149
transform 1 0 12788 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_134
timestamp 1644511149
transform 1 0 13432 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_141
timestamp 1644511149
transform 1 0 14076 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_148
timestamp 1644511149
transform 1 0 14720 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_155
timestamp 1644511149
transform 1 0 15364 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_164
timestamp 1644511149
transform 1 0 16192 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_185
timestamp 1644511149
transform 1 0 18124 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_194
timestamp 1644511149
transform 1 0 18952 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_205
timestamp 1644511149
transform 1 0 19964 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_214
timestamp 1644511149
transform 1 0 20792 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_222
timestamp 1644511149
transform 1 0 21528 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_241
timestamp 1644511149
transform 1 0 23276 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_248
timestamp 1644511149
transform 1 0 23920 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_268
timestamp 1644511149
transform 1 0 25760 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_276
timestamp 1644511149
transform 1 0 26496 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_61_281
timestamp 1644511149
transform 1 0 26956 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_300
timestamp 1644511149
transform 1 0 28704 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_320
timestamp 1644511149
transform 1 0 30544 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_326
timestamp 1644511149
transform 1 0 31096 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_332
timestamp 1644511149
transform 1 0 31648 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_342
timestamp 1644511149
transform 1 0 32568 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_360
timestamp 1644511149
transform 1 0 34224 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_24
timestamp 1644511149
transform 1 0 3312 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_38
timestamp 1644511149
transform 1 0 4600 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_45
timestamp 1644511149
transform 1 0 5244 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_57
timestamp 1644511149
transform 1 0 6348 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_69
timestamp 1644511149
transform 1 0 7452 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_81
timestamp 1644511149
transform 1 0 8556 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_85
timestamp 1644511149
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_97
timestamp 1644511149
transform 1 0 10028 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_108
timestamp 1644511149
transform 1 0 11040 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_115
timestamp 1644511149
transform 1 0 11684 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_122
timestamp 1644511149
transform 1 0 12328 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_129
timestamp 1644511149
transform 1 0 12972 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_136
timestamp 1644511149
transform 1 0 13616 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_141
timestamp 1644511149
transform 1 0 14076 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_151
timestamp 1644511149
transform 1 0 14996 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_159
timestamp 1644511149
transform 1 0 15732 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_163
timestamp 1644511149
transform 1 0 16100 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_172
timestamp 1644511149
transform 1 0 16928 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_192
timestamp 1644511149
transform 1 0 18768 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_62_197
timestamp 1644511149
transform 1 0 19228 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_216
timestamp 1644511149
transform 1 0 20976 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_236
timestamp 1644511149
transform 1 0 22816 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1644511149
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1644511149
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_269
timestamp 1644511149
transform 1 0 25852 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_280
timestamp 1644511149
transform 1 0 26864 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_286
timestamp 1644511149
transform 1 0 27416 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_294
timestamp 1644511149
transform 1 0 28152 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_304
timestamp 1644511149
transform 1 0 29072 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_318
timestamp 1644511149
transform 1 0 30360 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_331
timestamp 1644511149
transform 1 0 31556 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_360
timestamp 1644511149
transform 1 0 34224 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_3
timestamp 1644511149
transform 1 0 1380 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_7
timestamp 1644511149
transform 1 0 1748 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_32
timestamp 1644511149
transform 1 0 4048 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_45
timestamp 1644511149
transform 1 0 5244 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_52
timestamp 1644511149
transform 1 0 5888 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_57
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_69
timestamp 1644511149
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_81
timestamp 1644511149
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_93
timestamp 1644511149
transform 1 0 9660 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_97
timestamp 1644511149
transform 1 0 10028 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_101
timestamp 1644511149
transform 1 0 10396 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_108
timestamp 1644511149
transform 1 0 11040 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_113
timestamp 1644511149
transform 1 0 11500 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_117
timestamp 1644511149
transform 1 0 11868 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_124
timestamp 1644511149
transform 1 0 12512 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_131
timestamp 1644511149
transform 1 0 13156 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_138
timestamp 1644511149
transform 1 0 13800 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_154
timestamp 1644511149
transform 1 0 15272 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_160
timestamp 1644511149
transform 1 0 15824 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_164
timestamp 1644511149
transform 1 0 16192 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_185
timestamp 1644511149
transform 1 0 18124 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_205
timestamp 1644511149
transform 1 0 19964 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_214
timestamp 1644511149
transform 1 0 20792 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_222
timestamp 1644511149
transform 1 0 21528 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_228
timestamp 1644511149
transform 1 0 22080 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_238
timestamp 1644511149
transform 1 0 23000 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_247
timestamp 1644511149
transform 1 0 23828 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_256
timestamp 1644511149
transform 1 0 24656 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_264
timestamp 1644511149
transform 1 0 25392 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_272
timestamp 1644511149
transform 1 0 26128 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_281
timestamp 1644511149
transform 1 0 26956 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_299
timestamp 1644511149
transform 1 0 28612 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_312
timestamp 1644511149
transform 1 0 29808 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_325
timestamp 1644511149
transform 1 0 31004 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_332
timestamp 1644511149
transform 1 0 31648 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_337
timestamp 1644511149
transform 1 0 32108 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_360
timestamp 1644511149
transform 1 0 34224 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_3
timestamp 1644511149
transform 1 0 1380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_8
timestamp 1644511149
transform 1 0 1840 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_24
timestamp 1644511149
transform 1 0 3312 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_41
timestamp 1644511149
transform 1 0 4876 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_54
timestamp 1644511149
transform 1 0 6072 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_66
timestamp 1644511149
transform 1 0 7176 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_70
timestamp 1644511149
transform 1 0 7544 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1644511149
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1644511149
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_85
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_89
timestamp 1644511149
transform 1 0 9292 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_93
timestamp 1644511149
transform 1 0 9660 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_100
timestamp 1644511149
transform 1 0 10304 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_107
timestamp 1644511149
transform 1 0 10948 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_114
timestamp 1644511149
transform 1 0 11592 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_121
timestamp 1644511149
transform 1 0 12236 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_128
timestamp 1644511149
transform 1 0 12880 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_136
timestamp 1644511149
transform 1 0 13616 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_141
timestamp 1644511149
transform 1 0 14076 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_154
timestamp 1644511149
transform 1 0 15272 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_167
timestamp 1644511149
transform 1 0 16468 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_176
timestamp 1644511149
transform 1 0 17296 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_183
timestamp 1644511149
transform 1 0 17940 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_192
timestamp 1644511149
transform 1 0 18768 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_197
timestamp 1644511149
transform 1 0 19228 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_204
timestamp 1644511149
transform 1 0 19872 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_213
timestamp 1644511149
transform 1 0 20700 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_222
timestamp 1644511149
transform 1 0 21528 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_230
timestamp 1644511149
transform 1 0 22264 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_247
timestamp 1644511149
transform 1 0 23828 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1644511149
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_253
timestamp 1644511149
transform 1 0 24380 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_273
timestamp 1644511149
transform 1 0 26220 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_293
timestamp 1644511149
transform 1 0 28060 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_297
timestamp 1644511149
transform 1 0 28428 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_304
timestamp 1644511149
transform 1 0 29072 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_309
timestamp 1644511149
transform 1 0 29532 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_324
timestamp 1644511149
transform 1 0 30912 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_333
timestamp 1644511149
transform 1 0 31740 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_358
timestamp 1644511149
transform 1 0 34040 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_65_3
timestamp 1644511149
transform 1 0 1380 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_7
timestamp 1644511149
transform 1 0 1748 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_11
timestamp 1644511149
transform 1 0 2116 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_15
timestamp 1644511149
transform 1 0 2484 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_37
timestamp 1644511149
transform 1 0 4508 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_65_48
timestamp 1644511149
transform 1 0 5520 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_57
timestamp 1644511149
transform 1 0 6348 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_62
timestamp 1644511149
transform 1 0 6808 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_87
timestamp 1644511149
transform 1 0 9108 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_94
timestamp 1644511149
transform 1 0 9752 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_101
timestamp 1644511149
transform 1 0 10396 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_108
timestamp 1644511149
transform 1 0 11040 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_113
timestamp 1644511149
transform 1 0 11500 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_117
timestamp 1644511149
transform 1 0 11868 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_124
timestamp 1644511149
transform 1 0 12512 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_131
timestamp 1644511149
transform 1 0 13156 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_138
timestamp 1644511149
transform 1 0 13800 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_151
timestamp 1644511149
transform 1 0 14996 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_159
timestamp 1644511149
transform 1 0 15732 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_164
timestamp 1644511149
transform 1 0 16192 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_185
timestamp 1644511149
transform 1 0 18124 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_205
timestamp 1644511149
transform 1 0 19964 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_214
timestamp 1644511149
transform 1 0 20792 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_222
timestamp 1644511149
transform 1 0 21528 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_241
timestamp 1644511149
transform 1 0 23276 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_252
timestamp 1644511149
transform 1 0 24288 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_261
timestamp 1644511149
transform 1 0 25116 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_270
timestamp 1644511149
transform 1 0 25944 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_278
timestamp 1644511149
transform 1 0 26680 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_65_286
timestamp 1644511149
transform 1 0 27416 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_294
timestamp 1644511149
transform 1 0 28152 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_307
timestamp 1644511149
transform 1 0 29348 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_332
timestamp 1644511149
transform 1 0 31648 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_337
timestamp 1644511149
transform 1 0 32108 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_360
timestamp 1644511149
transform 1 0 34224 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_24
timestamp 1644511149
transform 1 0 3312 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_29
timestamp 1644511149
transform 1 0 3772 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_33
timestamp 1644511149
transform 1 0 4140 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_55
timestamp 1644511149
transform 1 0 6164 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_80
timestamp 1644511149
transform 1 0 8464 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_106
timestamp 1644511149
transform 1 0 10856 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_66_115
timestamp 1644511149
transform 1 0 11684 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_122
timestamp 1644511149
transform 1 0 12328 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_129
timestamp 1644511149
transform 1 0 12972 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_136
timestamp 1644511149
transform 1 0 13616 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_66_141
timestamp 1644511149
transform 1 0 14076 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_66_147
timestamp 1644511149
transform 1 0 14628 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_155
timestamp 1644511149
transform 1 0 15364 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_177
timestamp 1644511149
transform 1 0 17388 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_186
timestamp 1644511149
transform 1 0 18216 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_194
timestamp 1644511149
transform 1 0 18952 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_66_200
timestamp 1644511149
transform 1 0 19504 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_66_227
timestamp 1644511149
transform 1 0 21988 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_247
timestamp 1644511149
transform 1 0 23828 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1644511149
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_257
timestamp 1644511149
transform 1 0 24748 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_282
timestamp 1644511149
transform 1 0 27048 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_291
timestamp 1644511149
transform 1 0 27876 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_304
timestamp 1644511149
transform 1 0 29072 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_330
timestamp 1644511149
transform 1 0 31464 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_338
timestamp 1644511149
transform 1 0 32200 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_360
timestamp 1644511149
transform 1 0 34224 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_3
timestamp 1644511149
transform 1 0 1380 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_25
timestamp 1644511149
transform 1 0 3404 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_50
timestamp 1644511149
transform 1 0 5704 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_67_57
timestamp 1644511149
transform 1 0 6348 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_62
timestamp 1644511149
transform 1 0 6808 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_66
timestamp 1644511149
transform 1 0 7176 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_70
timestamp 1644511149
transform 1 0 7544 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_77
timestamp 1644511149
transform 1 0 8188 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_102
timestamp 1644511149
transform 1 0 10488 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_110
timestamp 1644511149
transform 1 0 11224 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_67_113
timestamp 1644511149
transform 1 0 11500 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_117
timestamp 1644511149
transform 1 0 11868 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_124
timestamp 1644511149
transform 1 0 12512 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_131
timestamp 1644511149
transform 1 0 13156 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_138
timestamp 1644511149
transform 1 0 13800 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_163
timestamp 1644511149
transform 1 0 16100 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1644511149
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_174
timestamp 1644511149
transform 1 0 17112 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_199
timestamp 1644511149
transform 1 0 19412 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_203
timestamp 1644511149
transform 1 0 19780 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_220
timestamp 1644511149
transform 1 0 21344 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_225
timestamp 1644511149
transform 1 0 21804 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_250
timestamp 1644511149
transform 1 0 24104 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_275
timestamp 1644511149
transform 1 0 26404 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_279
timestamp 1644511149
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_285
timestamp 1644511149
transform 1 0 27324 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_310
timestamp 1644511149
transform 1 0 29624 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_319
timestamp 1644511149
transform 1 0 30452 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_327
timestamp 1644511149
transform 1 0 31188 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1644511149
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_337
timestamp 1644511149
transform 1 0 32108 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_360
timestamp 1644511149
transform 1 0 34224 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_13
timestamp 1644511149
transform 1 0 2300 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_68_24
timestamp 1644511149
transform 1 0 3312 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_32
timestamp 1644511149
transform 1 0 4048 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_39
timestamp 1644511149
transform 1 0 4692 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_46
timestamp 1644511149
transform 1 0 5336 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_54
timestamp 1644511149
transform 1 0 6072 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_68_60
timestamp 1644511149
transform 1 0 6624 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_68_69
timestamp 1644511149
transform 1 0 7452 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_68_80
timestamp 1644511149
transform 1 0 8464 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_88
timestamp 1644511149
transform 1 0 9200 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_96
timestamp 1644511149
transform 1 0 9936 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_101
timestamp 1644511149
transform 1 0 10396 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_108
timestamp 1644511149
transform 1 0 11040 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_113
timestamp 1644511149
transform 1 0 11500 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_68_122
timestamp 1644511149
transform 1 0 12328 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_129
timestamp 1644511149
transform 1 0 12972 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_136
timestamp 1644511149
transform 1 0 13616 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_141
timestamp 1644511149
transform 1 0 14076 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_148
timestamp 1644511149
transform 1 0 14720 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_155
timestamp 1644511149
transform 1 0 15364 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_164
timestamp 1644511149
transform 1 0 16192 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_190
timestamp 1644511149
transform 1 0 18584 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_68_197
timestamp 1644511149
transform 1 0 19228 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_220
timestamp 1644511149
transform 1 0 21344 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_230
timestamp 1644511149
transform 1 0 22264 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_237
timestamp 1644511149
transform 1 0 22908 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_68_248
timestamp 1644511149
transform 1 0 23920 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_253
timestamp 1644511149
transform 1 0 24380 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_259
timestamp 1644511149
transform 1 0 24932 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_267
timestamp 1644511149
transform 1 0 25668 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_276
timestamp 1644511149
transform 1 0 26496 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_302
timestamp 1644511149
transform 1 0 28888 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_68_309
timestamp 1644511149
transform 1 0 29532 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_317
timestamp 1644511149
transform 1 0 30268 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_324
timestamp 1644511149
transform 1 0 30912 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_332
timestamp 1644511149
transform 1 0 31648 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_337
timestamp 1644511149
transform 1 0 32108 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_360
timestamp 1644511149
transform 1 0 34224 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 34868 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 34868 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 34868 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 34868 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 34868 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 34868 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 34868 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 34868 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 34868 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 34868 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 34868 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 34868 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 34868 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 34868 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 34868 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 34868 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 34868 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 34868 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 34868 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 34868 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 34868 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 34868 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 34868 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 34868 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 34868 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 34868 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 34868 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 34868 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 34868 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 34868 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 34868 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 34868 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 34868 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 34868 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 34868 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 34868 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 34868 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 34868 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 34868 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 34868 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 34868 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 34868 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 34868 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 34868 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 34868 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 34868 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 34868 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 34868 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 34868 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 34868 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 34868 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 34868 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 34868 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 34868 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 34868 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 34868 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 34868 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 34868 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 34868 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 34868 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 34868 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 34868 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 34868 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 34868 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 34868 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1644511149
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1644511149
transform -1 0 34868 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1644511149
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1644511149
transform -1 0 34868 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1644511149
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1644511149
transform -1 0 34868 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1644511149
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1644511149
transform -1 0 34868 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1644511149
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1644511149
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1644511149
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1644511149
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1644511149
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1644511149
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1644511149
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1644511149
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1644511149
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1644511149
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1644511149
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1644511149
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1644511149
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1644511149
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1644511149
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1644511149
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1644511149
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1644511149
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1644511149
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1644511149
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1644511149
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1644511149
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1644511149
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1644511149
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1644511149
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1644511149
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1644511149
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1644511149
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1644511149
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1644511149
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1644511149
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1644511149
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1644511149
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1644511149
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1644511149
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1644511149
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1644511149
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1644511149
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1644511149
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1644511149
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1644511149
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1644511149
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1644511149
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1644511149
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1644511149
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1644511149
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1644511149
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1644511149
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1644511149
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1644511149
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1644511149
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1644511149
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1644511149
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1644511149
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1644511149
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1644511149
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1644511149
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1644511149
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1644511149
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1644511149
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1644511149
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1644511149
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1644511149
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1644511149
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1644511149
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1644511149
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1644511149
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1644511149
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1644511149
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1644511149
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1644511149
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1644511149
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1644511149
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1644511149
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1644511149
transform 1 0 6256 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1644511149
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1644511149
transform 1 0 11408 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1644511149
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1644511149
transform 1 0 16560 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1644511149
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1644511149
transform 1 0 21712 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1644511149
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1644511149
transform 1 0 26864 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1644511149
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1644511149
transform 1 0 32016 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _0708_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26128 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _0709_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29532 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _0710_
timestamp 1644511149
transform 1 0 29532 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0711_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5612 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0712_
timestamp 1644511149
transform 1 0 1932 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0713_
timestamp 1644511149
transform 1 0 15732 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0714_
timestamp 1644511149
transform 1 0 1932 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0715_
timestamp 1644511149
transform 1 0 28980 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0716_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32936 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0717_
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0718_
timestamp 1644511149
transform 1 0 33580 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0719_
timestamp 1644511149
transform 1 0 1840 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0720_
timestamp 1644511149
transform 1 0 1840 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0721_
timestamp 1644511149
transform 1 0 31372 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0722_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 13248 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  _0723_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14168 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0724_
timestamp 1644511149
transform 1 0 19228 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0725_
timestamp 1644511149
transform 1 0 16836 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0726_
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0727_
timestamp 1644511149
transform 1 0 33580 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0728_
timestamp 1644511149
transform 1 0 33580 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0729_
timestamp 1644511149
transform 1 0 15640 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0730_
timestamp 1644511149
transform 1 0 23644 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0731_
timestamp 1644511149
transform 1 0 33948 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0732_
timestamp 1644511149
transform 1 0 1564 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0733_
timestamp 1644511149
transform 1 0 33580 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0734_
timestamp 1644511149
transform 1 0 1840 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0735_
timestamp 1644511149
transform 1 0 14168 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0736_
timestamp 1644511149
transform 1 0 29532 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0737_
timestamp 1644511149
transform 1 0 22632 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0738_
timestamp 1644511149
transform 1 0 10212 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0739_
timestamp 1644511149
transform 1 0 33672 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0740_
timestamp 1644511149
transform 1 0 33580 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0741_
timestamp 1644511149
transform 1 0 14168 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0742_
timestamp 1644511149
transform 1 0 4600 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0743_
timestamp 1644511149
transform 1 0 30636 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0744_
timestamp 1644511149
transform 1 0 33948 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0745_
timestamp 1644511149
transform 1 0 23644 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0746_
timestamp 1644511149
transform 1 0 1472 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0747_
timestamp 1644511149
transform 1 0 14168 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0748_
timestamp 1644511149
transform 1 0 4692 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0749_
timestamp 1644511149
transform 1 0 33580 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0750_
timestamp 1644511149
transform 1 0 2484 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0751_
timestamp 1644511149
transform 1 0 33948 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0752_
timestamp 1644511149
transform 1 0 14352 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0753_
timestamp 1644511149
transform 1 0 29900 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  _0754_
timestamp 1644511149
transform 1 0 28980 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0755_
timestamp 1644511149
transform 1 0 21804 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0756_
timestamp 1644511149
transform 1 0 1932 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0757_
timestamp 1644511149
transform 1 0 14260 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0758_
timestamp 1644511149
transform 1 0 1932 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0759_
timestamp 1644511149
transform 1 0 33948 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0760_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28520 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0761_
timestamp 1644511149
transform 1 0 33304 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0762_
timestamp 1644511149
transform 1 0 22816 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0763_
timestamp 1644511149
transform 1 0 22816 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0764_
timestamp 1644511149
transform 1 0 32108 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0765_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 33580 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  _0766_
timestamp 1644511149
transform 1 0 28244 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0767_
timestamp 1644511149
transform 1 0 29440 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0768_
timestamp 1644511149
transform 1 0 1748 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0769_
timestamp 1644511149
transform 1 0 1748 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0770_
timestamp 1644511149
transform 1 0 17664 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0771_
timestamp 1644511149
transform 1 0 1748 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  _0772_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29900 0 1 36992
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _0773_
timestamp 1644511149
transform 1 0 23184 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0774_
timestamp 1644511149
transform 1 0 33212 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0775_
timestamp 1644511149
transform 1 0 21804 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0776_
timestamp 1644511149
transform 1 0 17020 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0777_
timestamp 1644511149
transform 1 0 20332 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  _0778_
timestamp 1644511149
transform 1 0 28244 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0779_
timestamp 1644511149
transform 1 0 15916 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0780_
timestamp 1644511149
transform 1 0 33212 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0781_
timestamp 1644511149
transform 1 0 2116 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0782_
timestamp 1644511149
transform 1 0 32108 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0783_
timestamp 1644511149
transform 1 0 1840 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0784_
timestamp 1644511149
transform 1 0 3036 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  _0785_
timestamp 1644511149
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0786_
timestamp 1644511149
transform 1 0 23920 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0787_
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0788_
timestamp 1644511149
transform 1 0 7912 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0789_
timestamp 1644511149
transform 1 0 32936 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0790_
timestamp 1644511149
transform 1 0 15916 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0791_
timestamp 1644511149
transform 1 0 3772 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0792_
timestamp 1644511149
transform 1 0 28336 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0793_
timestamp 1644511149
transform 1 0 18492 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0794_
timestamp 1644511149
transform 1 0 19412 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0795_
timestamp 1644511149
transform 1 0 28796 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0796_
timestamp 1644511149
transform 1 0 2576 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0797_
timestamp 1644511149
transform 1 0 4416 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0798_
timestamp 1644511149
transform 1 0 33028 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0799_
timestamp 1644511149
transform 1 0 6532 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0800_
timestamp 1644511149
transform 1 0 33672 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0801_
timestamp 1644511149
transform 1 0 33028 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0802_
timestamp 1644511149
transform 1 0 2668 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0803_
timestamp 1644511149
transform 1 0 2208 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0804_
timestamp 1644511149
transform 1 0 33948 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0805_
timestamp 1644511149
transform 1 0 7268 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0806_
timestamp 1644511149
transform 1 0 2576 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0807_
timestamp 1644511149
transform 1 0 31372 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0808_
timestamp 1644511149
transform 1 0 7912 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0809_
timestamp 1644511149
transform 1 0 5244 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0810_
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0811_
timestamp 1644511149
transform 1 0 15088 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0812_
timestamp 1644511149
transform 1 0 7268 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0813_
timestamp 1644511149
transform 1 0 33120 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0814_
timestamp 1644511149
transform 1 0 3036 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0815_
timestamp 1644511149
transform 1 0 29532 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0816_
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0817_
timestamp 1644511149
transform 1 0 14444 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0818_
timestamp 1644511149
transform 1 0 13524 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0819_
timestamp 1644511149
transform 1 0 3772 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0820_
timestamp 1644511149
transform 1 0 26220 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0821_
timestamp 1644511149
transform 1 0 30176 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0822_
timestamp 1644511149
transform 1 0 28796 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0823_
timestamp 1644511149
transform 1 0 27692 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0824_
timestamp 1644511149
transform 1 0 2392 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0825_
timestamp 1644511149
transform 1 0 15824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0826_
timestamp 1644511149
transform 1 0 29072 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0827_
timestamp 1644511149
transform 1 0 30728 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0828_
timestamp 1644511149
transform 1 0 16008 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0829_
timestamp 1644511149
transform 1 0 5244 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0830_
timestamp 1644511149
transform 1 0 1748 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0831_
timestamp 1644511149
transform 1 0 1748 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0832_
timestamp 1644511149
transform 1 0 1748 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0833_
timestamp 1644511149
transform 1 0 29532 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0834_
timestamp 1644511149
transform 1 0 15364 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0835_
timestamp 1644511149
transform 1 0 1656 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0836_
timestamp 1644511149
transform 1 0 4048 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0837_
timestamp 1644511149
transform 1 0 13156 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0838_
timestamp 1644511149
transform 1 0 4416 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0839_
timestamp 1644511149
transform 1 0 30728 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0840_
timestamp 1644511149
transform 1 0 21804 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0841_
timestamp 1644511149
transform 1 0 15088 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0842_
timestamp 1644511149
transform 1 0 28520 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0843_
timestamp 1644511149
transform 1 0 25300 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0844_
timestamp 1644511149
transform 1 0 24472 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _0845_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27784 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0846_
timestamp 1644511149
transform 1 0 26128 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0847_
timestamp 1644511149
transform 1 0 26220 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0848_
timestamp 1644511149
transform 1 0 31188 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0849_
timestamp 1644511149
transform 1 0 31096 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0850_
timestamp 1644511149
transform 1 0 25392 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0851_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27232 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0852_
timestamp 1644511149
transform 1 0 24012 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0853_
timestamp 1644511149
transform 1 0 20424 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0854_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23000 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__o22a_1  _0855_
timestamp 1644511149
transform 1 0 27876 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0856_
timestamp 1644511149
transform 1 0 26404 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0857_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32108 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0858_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27048 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0859_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27876 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0860_
timestamp 1644511149
transform 1 0 27232 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _0861_
timestamp 1644511149
transform 1 0 27324 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0862_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27048 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0863_
timestamp 1644511149
transform 1 0 28336 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0864_
timestamp 1644511149
transform 1 0 26772 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0865_
timestamp 1644511149
transform 1 0 28244 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _0866_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26956 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0867_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28152 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0868_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27784 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0869_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 33856 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0870_
timestamp 1644511149
transform 1 0 15180 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0871_
timestamp 1644511149
transform 1 0 14444 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0872_
timestamp 1644511149
transform 1 0 14720 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0873_
timestamp 1644511149
transform 1 0 14168 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0874_
timestamp 1644511149
transform 1 0 13800 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0875_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23460 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0876_
timestamp 1644511149
transform 1 0 15272 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0877_
timestamp 1644511149
transform 1 0 21712 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _0878_
timestamp 1644511149
transform 1 0 15916 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0879_
timestamp 1644511149
transform 1 0 16008 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0880_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20700 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0881_
timestamp 1644511149
transform 1 0 21896 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0882_
timestamp 1644511149
transform 1 0 22724 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0883_
timestamp 1644511149
transform 1 0 24380 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0884_
timestamp 1644511149
transform 1 0 24748 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0885_
timestamp 1644511149
transform 1 0 25852 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _0886_
timestamp 1644511149
transform 1 0 26956 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0887_
timestamp 1644511149
transform 1 0 32108 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0888_
timestamp 1644511149
transform 1 0 27784 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a221oi_2  _0889_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26956 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0890_
timestamp 1644511149
transform 1 0 33856 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0891_
timestamp 1644511149
transform 1 0 32476 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0892_
timestamp 1644511149
transform 1 0 13524 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0893_
timestamp 1644511149
transform 1 0 31372 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0894_
timestamp 1644511149
transform 1 0 31096 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0895_
timestamp 1644511149
transform 1 0 14076 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0896_
timestamp 1644511149
transform 1 0 15180 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0897_
timestamp 1644511149
transform 1 0 14628 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0898_
timestamp 1644511149
transform 1 0 30084 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0899_
timestamp 1644511149
transform 1 0 29532 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__o22a_1  _0900_
timestamp 1644511149
transform 1 0 29532 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0901_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30912 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0902_
timestamp 1644511149
transform 1 0 29900 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0903_
timestamp 1644511149
transform 1 0 31004 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0904_
timestamp 1644511149
transform 1 0 31556 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0905_
timestamp 1644511149
transform 1 0 31924 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _0906_
timestamp 1644511149
transform 1 0 32752 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0907_
timestamp 1644511149
transform 1 0 27048 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a211oi_2  _0908_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 33028 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0909_
timestamp 1644511149
transform 1 0 28612 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0910_
timestamp 1644511149
transform 1 0 28980 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _0911_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28520 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0912_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29532 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0913_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28060 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0914_
timestamp 1644511149
transform 1 0 30360 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0915_
timestamp 1644511149
transform 1 0 29532 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0916_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 31004 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0917_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29256 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0918_
timestamp 1644511149
transform 1 0 27692 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0919_
timestamp 1644511149
transform 1 0 30084 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0920_
timestamp 1644511149
transform 1 0 29532 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0921_
timestamp 1644511149
transform 1 0 28704 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0922_
timestamp 1644511149
transform 1 0 29532 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0923_
timestamp 1644511149
transform 1 0 30452 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0924_
timestamp 1644511149
transform 1 0 29256 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0925_
timestamp 1644511149
transform 1 0 30084 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0926_
timestamp 1644511149
transform 1 0 27968 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0927_
timestamp 1644511149
transform 1 0 28796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0928_
timestamp 1644511149
transform 1 0 27784 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0929_
timestamp 1644511149
transform 1 0 27324 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0930_
timestamp 1644511149
transform 1 0 27048 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0931_
timestamp 1644511149
transform 1 0 21988 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _0932_
timestamp 1644511149
transform 1 0 14444 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0933_
timestamp 1644511149
transform 1 0 26956 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0934_
timestamp 1644511149
transform 1 0 23092 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0935_
timestamp 1644511149
transform 1 0 21068 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0936_
timestamp 1644511149
transform 1 0 21988 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0937_
timestamp 1644511149
transform 1 0 23276 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0938_
timestamp 1644511149
transform 1 0 20976 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0939_
timestamp 1644511149
transform 1 0 23460 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0940_
timestamp 1644511149
transform 1 0 30820 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0941_
timestamp 1644511149
transform 1 0 15272 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0942_
timestamp 1644511149
transform 1 0 24380 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0943_
timestamp 1644511149
transform 1 0 20976 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0944_
timestamp 1644511149
transform 1 0 14904 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0945_
timestamp 1644511149
transform 1 0 32108 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0946_
timestamp 1644511149
transform 1 0 25668 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0947_
timestamp 1644511149
transform 1 0 15272 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0948_
timestamp 1644511149
transform 1 0 25576 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0949_
timestamp 1644511149
transform 1 0 26036 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0950_
timestamp 1644511149
transform 1 0 20424 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0951_
timestamp 1644511149
transform 1 0 21068 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0952_
timestamp 1644511149
transform 1 0 31372 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0953_
timestamp 1644511149
transform 1 0 14628 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0954_
timestamp 1644511149
transform 1 0 33856 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0955_
timestamp 1644511149
transform 1 0 26956 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0956_
timestamp 1644511149
transform 1 0 29624 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _0957_
timestamp 1644511149
transform 1 0 30176 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0958_
timestamp 1644511149
transform 1 0 31096 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0959_
timestamp 1644511149
transform 1 0 28796 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0960_
timestamp 1644511149
transform 1 0 32108 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0961_
timestamp 1644511149
transform 1 0 30176 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0962_
timestamp 1644511149
transform 1 0 30820 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0963_
timestamp 1644511149
transform 1 0 30728 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0964_
timestamp 1644511149
transform 1 0 31832 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0965_
timestamp 1644511149
transform 1 0 31372 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0966_
timestamp 1644511149
transform 1 0 29348 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0967_
timestamp 1644511149
transform 1 0 31188 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0968_
timestamp 1644511149
transform 1 0 31372 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0969_
timestamp 1644511149
transform 1 0 28612 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0970_
timestamp 1644511149
transform 1 0 32108 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0971_
timestamp 1644511149
transform 1 0 31096 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0972_
timestamp 1644511149
transform 1 0 28612 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0973_
timestamp 1644511149
transform 1 0 32844 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0974_
timestamp 1644511149
transform 1 0 31372 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0975_
timestamp 1644511149
transform 1 0 25300 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0976_
timestamp 1644511149
transform 1 0 33304 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0977_
timestamp 1644511149
transform 1 0 23644 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0978_
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0979_
timestamp 1644511149
transform 1 0 14720 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0980_
timestamp 1644511149
transform 1 0 20792 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0981_
timestamp 1644511149
transform 1 0 20976 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0982_
timestamp 1644511149
transform 1 0 22632 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0983_
timestamp 1644511149
transform 1 0 21068 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0984_
timestamp 1644511149
transform 1 0 21712 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0985_
timestamp 1644511149
transform 1 0 20424 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0986_
timestamp 1644511149
transform 1 0 25392 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0987_
timestamp 1644511149
transform 1 0 24656 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _0988_
timestamp 1644511149
transform 1 0 25300 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0989_
timestamp 1644511149
transform 1 0 20976 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0990_
timestamp 1644511149
transform 1 0 24932 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__and4b_1  _0991_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0992_
timestamp 1644511149
transform 1 0 21988 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0993_
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0994_
timestamp 1644511149
transform 1 0 21252 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0995_
timestamp 1644511149
transform 1 0 20424 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _0996_
timestamp 1644511149
transform 1 0 21804 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0997_
timestamp 1644511149
transform 1 0 19780 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0998_
timestamp 1644511149
transform 1 0 22632 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0999_
timestamp 1644511149
transform 1 0 15916 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1000_
timestamp 1644511149
transform 1 0 23000 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1001_
timestamp 1644511149
transform 1 0 17572 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1002_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22908 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1003_
timestamp 1644511149
transform 1 0 22908 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1004_
timestamp 1644511149
transform 1 0 23920 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1005_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24380 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1006_
timestamp 1644511149
transform 1 0 26496 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1007_
timestamp 1644511149
transform 1 0 24380 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1008_
timestamp 1644511149
transform 1 0 24472 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1009_
timestamp 1644511149
transform 1 0 24656 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1010_
timestamp 1644511149
transform 1 0 25392 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1011_
timestamp 1644511149
transform 1 0 25576 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1012_
timestamp 1644511149
transform 1 0 20056 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1013_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24840 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1014_
timestamp 1644511149
transform 1 0 18400 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1015_
timestamp 1644511149
transform 1 0 25208 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1016_
timestamp 1644511149
transform 1 0 23552 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1017_
timestamp 1644511149
transform 1 0 25760 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1018_
timestamp 1644511149
transform 1 0 23184 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1019_
timestamp 1644511149
transform 1 0 24104 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1020_
timestamp 1644511149
transform 1 0 20608 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1021_
timestamp 1644511149
transform 1 0 22632 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1022_
timestamp 1644511149
transform 1 0 24472 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1023_
timestamp 1644511149
transform 1 0 23092 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1024_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23552 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1025_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1026_
timestamp 1644511149
transform 1 0 24472 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1027_
timestamp 1644511149
transform 1 0 24932 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1028_
timestamp 1644511149
transform 1 0 22356 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1029_
timestamp 1644511149
transform 1 0 22356 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1030_
timestamp 1644511149
transform 1 0 21712 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1031_
timestamp 1644511149
transform 1 0 25944 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1032_
timestamp 1644511149
transform 1 0 22540 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1033_
timestamp 1644511149
transform 1 0 21988 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1034_
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1035_
timestamp 1644511149
transform 1 0 22908 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1036_
timestamp 1644511149
transform 1 0 22172 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1037_
timestamp 1644511149
transform 1 0 23184 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1038_
timestamp 1644511149
transform 1 0 23368 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1039_
timestamp 1644511149
transform 1 0 25668 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1040_
timestamp 1644511149
transform 1 0 24656 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1041_
timestamp 1644511149
transform 1 0 19688 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1042_
timestamp 1644511149
transform 1 0 15364 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1043_
timestamp 1644511149
transform 1 0 15824 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1044_
timestamp 1644511149
transform 1 0 19688 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1045_
timestamp 1644511149
transform 1 0 14260 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1046_
timestamp 1644511149
transform 1 0 20516 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1047_
timestamp 1644511149
transform 1 0 20516 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1048_
timestamp 1644511149
transform 1 0 23460 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1049_
timestamp 1644511149
transform 1 0 15916 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1050_
timestamp 1644511149
transform 1 0 21804 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1051_
timestamp 1644511149
transform 1 0 20240 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1052_
timestamp 1644511149
transform 1 0 20148 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1053_
timestamp 1644511149
transform 1 0 15824 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1054_
timestamp 1644511149
transform 1 0 21068 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1055_
timestamp 1644511149
transform 1 0 19504 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__and4b_1  _1056_
timestamp 1644511149
transform 1 0 20608 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1057_
timestamp 1644511149
transform 1 0 22540 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1058_
timestamp 1644511149
transform 1 0 26956 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1059_
timestamp 1644511149
transform 1 0 19504 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1060_
timestamp 1644511149
transform 1 0 13340 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1061_
timestamp 1644511149
transform 1 0 21344 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1062_
timestamp 1644511149
transform 1 0 12880 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1063_
timestamp 1644511149
transform 1 0 21988 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1064_
timestamp 1644511149
transform 1 0 13432 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1065_
timestamp 1644511149
transform 1 0 22724 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1066_
timestamp 1644511149
transform 1 0 21804 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1067_
timestamp 1644511149
transform 1 0 21620 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1068_
timestamp 1644511149
transform 1 0 21988 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1069_
timestamp 1644511149
transform 1 0 21804 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1070_
timestamp 1644511149
transform 1 0 14076 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1071_
timestamp 1644511149
transform 1 0 20884 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1072_
timestamp 1644511149
transform 1 0 16652 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1073_
timestamp 1644511149
transform 1 0 21804 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1074_
timestamp 1644511149
transform 1 0 14536 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1075_
timestamp 1644511149
transform 1 0 22908 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1076_
timestamp 1644511149
transform 1 0 16928 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1077_
timestamp 1644511149
transform 1 0 23368 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1078_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1079_
timestamp 1644511149
transform 1 0 21344 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1080_
timestamp 1644511149
transform 1 0 22448 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1081_
timestamp 1644511149
transform 1 0 23000 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1082_
timestamp 1644511149
transform 1 0 23460 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1083_
timestamp 1644511149
transform 1 0 24380 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1084_
timestamp 1644511149
transform 1 0 12696 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1085_
timestamp 1644511149
transform 1 0 24380 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1086_
timestamp 1644511149
transform 1 0 23184 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1087_
timestamp 1644511149
transform 1 0 24564 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1088_
timestamp 1644511149
transform 1 0 24472 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1089_
timestamp 1644511149
transform 1 0 25576 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1090_
timestamp 1644511149
transform 1 0 13892 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _1091_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1092_
timestamp 1644511149
transform 1 0 12788 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1093_
timestamp 1644511149
transform 1 0 26036 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1094_
timestamp 1644511149
transform 1 0 12788 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1095_
timestamp 1644511149
transform 1 0 25484 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1096_
timestamp 1644511149
transform 1 0 24564 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1097_
timestamp 1644511149
transform 1 0 27508 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1098_
timestamp 1644511149
transform 1 0 13156 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1099_
timestamp 1644511149
transform 1 0 26404 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1100_
timestamp 1644511149
transform 1 0 25576 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1101_
timestamp 1644511149
transform 1 0 26128 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1102_
timestamp 1644511149
transform 1 0 27140 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1103_
timestamp 1644511149
transform 1 0 14536 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _1104_
timestamp 1644511149
transform 1 0 25944 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1105_
timestamp 1644511149
transform 1 0 24472 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1106_
timestamp 1644511149
transform 1 0 14720 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1107_
timestamp 1644511149
transform 1 0 20332 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1108_
timestamp 1644511149
transform 1 0 15272 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1109_
timestamp 1644511149
transform 1 0 27232 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1110_
timestamp 1644511149
transform 1 0 27692 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1111_
timestamp 1644511149
transform 1 0 26036 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1112_
timestamp 1644511149
transform 1 0 14076 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1113_
timestamp 1644511149
transform 1 0 28520 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1114_
timestamp 1644511149
transform 1 0 26956 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1115_
timestamp 1644511149
transform 1 0 32568 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1116_
timestamp 1644511149
transform 1 0 15824 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1117_
timestamp 1644511149
transform 1 0 28520 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1118_
timestamp 1644511149
transform 1 0 30820 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__and4b_1  _1119_
timestamp 1644511149
transform 1 0 27416 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1120_
timestamp 1644511149
transform 1 0 28612 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1121_
timestamp 1644511149
transform 1 0 30728 0 -1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1122_
timestamp 1644511149
transform 1 0 31280 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1123_
timestamp 1644511149
transform 1 0 13340 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1124_
timestamp 1644511149
transform 1 0 28152 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1125_
timestamp 1644511149
transform -1 0 13524 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1126_
timestamp 1644511149
transform 1 0 28428 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1127_
timestamp 1644511149
transform 1 0 12512 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1128_
timestamp 1644511149
transform 1 0 28336 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1129_
timestamp 1644511149
transform 1 0 28244 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1130_
timestamp 1644511149
transform 1 0 28520 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1131_
timestamp 1644511149
transform 1 0 29256 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1132_
timestamp 1644511149
transform 1 0 31188 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1133_
timestamp 1644511149
transform 1 0 14076 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1134_
timestamp 1644511149
transform 1 0 29624 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1135_
timestamp 1644511149
transform 1 0 30728 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1136_
timestamp 1644511149
transform 1 0 13340 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1137_
timestamp 1644511149
transform 1 0 30084 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1138_
timestamp 1644511149
transform 1 0 25300 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1139_
timestamp 1644511149
transform -1 0 31648 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1140_
timestamp 1644511149
transform 1 0 30176 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1141_
timestamp 1644511149
transform 1 0 29900 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1142_
timestamp 1644511149
transform 1 0 27324 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1143_
timestamp 1644511149
transform 1 0 30176 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1144_
timestamp 1644511149
transform 1 0 32108 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1145_
timestamp 1644511149
transform 1 0 13340 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1146_
timestamp 1644511149
transform 1 0 31188 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1147_
timestamp 1644511149
transform 1 0 28612 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1148_
timestamp 1644511149
transform 1 0 12696 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1149_
timestamp 1644511149
transform 1 0 30912 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1150_
timestamp 1644511149
transform 1 0 32108 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1151_
timestamp 1644511149
transform 1 0 31280 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1152_
timestamp 1644511149
transform 1 0 31280 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1153_
timestamp 1644511149
transform 1 0 33212 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1154_
timestamp 1644511149
transform 1 0 14628 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1155_
timestamp 1644511149
transform 1 0 24564 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1156_
timestamp 1644511149
transform 1 0 31464 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1157_
timestamp 1644511149
transform 1 0 30544 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1158_
timestamp 1644511149
transform 1 0 25300 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1159_
timestamp 1644511149
transform 1 0 12696 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1160_
timestamp 1644511149
transform 1 0 32936 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1161_
timestamp 1644511149
transform 1 0 31924 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1162_
timestamp 1644511149
transform 1 0 32292 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1163_
timestamp 1644511149
transform 1 0 11868 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1164_
timestamp 1644511149
transform 1 0 32844 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1165_
timestamp 1644511149
transform 1 0 27048 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1166_
timestamp 1644511149
transform 1 0 31096 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1167_
timestamp 1644511149
transform 1 0 31004 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1168_
timestamp 1644511149
transform 1 0 13892 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _1169_
timestamp 1644511149
transform 1 0 28520 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1170_
timestamp 1644511149
transform 1 0 14996 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1171_
timestamp 1644511149
transform 1 0 17204 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1172_
timestamp 1644511149
transform 1 0 14352 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1173_
timestamp 1644511149
transform 1 0 18308 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1174_
timestamp 1644511149
transform 1 0 14812 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1175_
timestamp 1644511149
transform 1 0 15088 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1176_
timestamp 1644511149
transform 1 0 18216 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1177_
timestamp 1644511149
transform 1 0 18308 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1178_
timestamp 1644511149
transform 1 0 18308 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1179_
timestamp 1644511149
transform 1 0 17664 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1180_
timestamp 1644511149
transform 1 0 17204 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1181_
timestamp 1644511149
transform 1 0 17020 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1182_
timestamp 1644511149
transform 1 0 15732 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1183_
timestamp 1644511149
transform 1 0 15088 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1184_
timestamp 1644511149
transform 1 0 15732 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1185_
timestamp 1644511149
transform 1 0 14444 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1186_
timestamp 1644511149
transform 1 0 13708 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1187_
timestamp 1644511149
transform 1 0 15732 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1188_
timestamp 1644511149
transform 1 0 14352 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1189_
timestamp 1644511149
transform 1 0 26036 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1190_
timestamp 1644511149
transform 1 0 13340 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1191_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17020 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1192_
timestamp 1644511149
transform 1 0 20148 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1193_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19228 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1194_
timestamp 1644511149
transform 1 0 17940 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1195_
timestamp 1644511149
transform 1 0 19412 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1196_
timestamp 1644511149
transform 1 0 19044 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1197_
timestamp 1644511149
transform 1 0 16652 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1198_
timestamp 1644511149
transform 1 0 12052 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1199_
timestamp 1644511149
transform 1 0 16652 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1200_
timestamp 1644511149
transform 1 0 14628 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1201_
timestamp 1644511149
transform 1 0 18308 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1202_
timestamp 1644511149
transform 1 0 13800 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1203_
timestamp 1644511149
transform 1 0 17480 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1204_
timestamp 1644511149
transform 1 0 13984 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1205_
timestamp 1644511149
transform 1 0 16928 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1206_
timestamp 1644511149
transform 1 0 13248 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1207_
timestamp 1644511149
transform 1 0 16652 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1208_
timestamp 1644511149
transform 1 0 12052 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1209_
timestamp 1644511149
transform 1 0 17848 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1210_
timestamp 1644511149
transform 1 0 13340 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1211_
timestamp 1644511149
transform 1 0 18768 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1212_
timestamp 1644511149
transform 1 0 13340 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1213_
timestamp 1644511149
transform 1 0 19596 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1214_
timestamp 1644511149
transform 1 0 12696 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1215_
timestamp 1644511149
transform 1 0 18124 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1216_
timestamp 1644511149
transform 1 0 17388 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1217_
timestamp 1644511149
transform 1 0 17388 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1218_
timestamp 1644511149
transform 1 0 19228 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1219_
timestamp 1644511149
transform 1 0 18308 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1220_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18676 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1221_
timestamp 1644511149
transform 1 0 16652 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1222_
timestamp 1644511149
transform 1 0 13524 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1223_
timestamp 1644511149
transform 1 0 19228 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1224_
timestamp 1644511149
transform 1 0 12052 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1225_
timestamp 1644511149
transform 1 0 17388 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1226_
timestamp 1644511149
transform 1 0 12972 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1227_
timestamp 1644511149
transform 1 0 12236 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1228_
timestamp 1644511149
transform 1 0 17756 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1229_
timestamp 1644511149
transform 1 0 12696 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1230_
timestamp 1644511149
transform 1 0 16652 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1231_
timestamp 1644511149
transform 1 0 12052 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1232_
timestamp 1644511149
transform 1 0 14260 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1233_
timestamp 1644511149
transform 1 0 14904 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1234_
timestamp 1644511149
transform 1 0 14812 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1235_
timestamp 1644511149
transform 1 0 12144 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1236_
timestamp 1644511149
transform 1 0 16100 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1237_
timestamp 1644511149
transform 1 0 11500 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1238_
timestamp 1644511149
transform 1 0 17112 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1239_
timestamp 1644511149
transform 1 0 18584 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1240_
timestamp 1644511149
transform 1 0 18216 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1241_
timestamp 1644511149
transform 1 0 15640 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1242_
timestamp 1644511149
transform 1 0 18216 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a41o_1  _1243_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17388 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1244_
timestamp 1644511149
transform 1 0 17756 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1245_
timestamp 1644511149
transform 1 0 13340 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1246_
timestamp 1644511149
transform 1 0 14444 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1247_
timestamp 1644511149
transform 1 0 16468 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1248_
timestamp 1644511149
transform 1 0 13524 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1249_
timestamp 1644511149
transform 1 0 18492 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1250_
timestamp 1644511149
transform 1 0 13800 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1251_
timestamp 1644511149
transform 1 0 15732 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1252_
timestamp 1644511149
transform 1 0 13156 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1253_
timestamp 1644511149
transform 1 0 18400 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1254_
timestamp 1644511149
transform 1 0 14260 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1255_
timestamp 1644511149
transform 1 0 18308 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1256_
timestamp 1644511149
transform 1 0 12880 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1257_
timestamp 1644511149
transform 1 0 13340 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1258_
timestamp 1644511149
transform 1 0 20332 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1259_
timestamp 1644511149
transform 1 0 12236 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1260_
timestamp 1644511149
transform 1 0 20332 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1261_
timestamp 1644511149
transform 1 0 12696 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1262_
timestamp 1644511149
transform 1 0 19320 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1263_
timestamp 1644511149
transform 1 0 17388 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1264_
timestamp 1644511149
transform 1 0 17480 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1265_
timestamp 1644511149
transform 1 0 19320 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1266_
timestamp 1644511149
transform 1 0 20240 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1267_
timestamp 1644511149
transform 1 0 19228 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1268_
timestamp 1644511149
transform 1 0 15732 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1269_
timestamp 1644511149
transform 1 0 12880 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1270_
timestamp 1644511149
transform 1 0 20332 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1271_
timestamp 1644511149
transform 1 0 12880 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1272_
timestamp 1644511149
transform 1 0 21068 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1273_
timestamp 1644511149
transform 1 0 12696 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1274_
timestamp 1644511149
transform 1 0 21804 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1275_
timestamp 1644511149
transform 1 0 12236 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1276_
timestamp 1644511149
transform 1 0 13156 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1277_
timestamp 1644511149
transform 1 0 23368 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1278_
timestamp 1644511149
transform 1 0 12604 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1279_
timestamp 1644511149
transform 1 0 23184 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1280_
timestamp 1644511149
transform 1 0 12052 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1281_
timestamp 1644511149
transform 1 0 22816 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1282_
timestamp 1644511149
transform 1 0 13984 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1283_
timestamp 1644511149
transform 1 0 24196 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1284_
timestamp 1644511149
transform 1 0 13340 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1285_
timestamp 1644511149
transform 1 0 23000 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1286_
timestamp 1644511149
transform 1 0 23644 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1287_
timestamp 1644511149
transform 1 0 22448 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1288_
timestamp 1644511149
transform 1 0 23368 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1289_
timestamp 1644511149
transform 1 0 25760 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1290_
timestamp 1644511149
transform 1 0 24380 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1291_
timestamp 1644511149
transform 1 0 25944 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1292_
timestamp 1644511149
transform 1 0 12052 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1293_
timestamp 1644511149
transform 1 0 24656 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1294_
timestamp 1644511149
transform 1 0 11592 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1295_
timestamp 1644511149
transform 1 0 12512 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1296_
timestamp 1644511149
transform 1 0 25484 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1297_
timestamp 1644511149
transform 1 0 12512 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1298_
timestamp 1644511149
transform 1 0 26956 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1299_
timestamp 1644511149
transform 1 0 11960 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1300_
timestamp 1644511149
transform 1 0 27416 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1301_
timestamp 1644511149
transform 1 0 11316 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1302_
timestamp 1644511149
transform 1 0 29992 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1303_
timestamp 1644511149
transform 1 0 11592 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1304_
timestamp 1644511149
transform 1 0 26036 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1305_
timestamp 1644511149
transform 1 0 12696 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1306_
timestamp 1644511149
transform 1 0 26036 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1307_
timestamp 1644511149
transform 1 0 11868 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1308_
timestamp 1644511149
transform 1 0 27508 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1309_
timestamp 1644511149
transform 1 0 26220 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1310_
timestamp 1644511149
transform 1 0 25576 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1311_
timestamp 1644511149
transform 1 0 28520 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1312_
timestamp 1644511149
transform 1 0 25208 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1313_
timestamp 1644511149
transform 1 0 27508 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1314_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27600 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1315_
timestamp 1644511149
transform 1 0 29532 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1316_
timestamp 1644511149
transform 1 0 29164 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1317_
timestamp 1644511149
transform 1 0 29532 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1318_
timestamp 1644511149
transform 1 0 29256 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1319_
timestamp 1644511149
transform 1 0 29532 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1320_
timestamp 1644511149
transform 1 0 27324 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1321_
timestamp 1644511149
transform 1 0 26956 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1322_
timestamp 1644511149
transform 1 0 20792 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1323_
timestamp 1644511149
transform 1 0 19872 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1324_
timestamp 1644511149
transform 1 0 21896 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1325_
timestamp 1644511149
transform 1 0 23736 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1326_
timestamp 1644511149
transform 1 0 23828 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1327_
timestamp 1644511149
transform 1 0 24840 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1328_
timestamp 1644511149
transform 1 0 26680 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1329_
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1330_
timestamp 1644511149
transform 1 0 28336 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1331_
timestamp 1644511149
transform 1 0 28244 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1332_
timestamp 1644511149
transform 1 0 29532 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1333_
timestamp 1644511149
transform 1 0 30176 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1334_
timestamp 1644511149
transform 1 0 30360 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1335_
timestamp 1644511149
transform 1 0 32108 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1336_
timestamp 1644511149
transform 1 0 32292 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1337_
timestamp 1644511149
transform 1 0 32752 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1338_
timestamp 1644511149
transform 1 0 19872 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1339_
timestamp 1644511149
transform 1 0 24656 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1340_
timestamp 1644511149
transform 1 0 22172 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1341_
timestamp 1644511149
transform 1 0 26036 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1342_
timestamp 1644511149
transform 1 0 26036 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1343_
timestamp 1644511149
transform 1 0 25392 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1344_
timestamp 1644511149
transform 1 0 25208 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1345_
timestamp 1644511149
transform 1 0 21068 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1346_
timestamp 1644511149
transform 1 0 25024 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1347_
timestamp 1644511149
transform 1 0 19228 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1348_
timestamp 1644511149
transform 1 0 19412 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1349_
timestamp 1644511149
transform 1 0 19872 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1350_
timestamp 1644511149
transform 1 0 22448 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1351_
timestamp 1644511149
transform 1 0 19504 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1352_
timestamp 1644511149
transform 1 0 19504 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1353_
timestamp 1644511149
transform 1 0 23460 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1354_
timestamp 1644511149
transform 1 0 24104 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1355_
timestamp 1644511149
transform 1 0 26496 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1356_
timestamp 1644511149
transform 1 0 26956 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1357_
timestamp 1644511149
transform 1 0 25300 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1358_
timestamp 1644511149
transform 1 0 19596 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1359_
timestamp 1644511149
transform 1 0 28796 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1360_
timestamp 1644511149
transform 1 0 27968 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1361_
timestamp 1644511149
transform 1 0 29624 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1362_
timestamp 1644511149
transform 1 0 30084 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1363_
timestamp 1644511149
transform 1 0 30452 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1364_
timestamp 1644511149
transform 1 0 32660 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1365_
timestamp 1644511149
transform 1 0 32752 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1366_
timestamp 1644511149
transform 1 0 30084 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1367_
timestamp 1644511149
transform 1 0 18032 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1368_
timestamp 1644511149
transform 1 0 18032 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1369_
timestamp 1644511149
transform 1 0 18032 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1370_
timestamp 1644511149
transform 1 0 19872 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1371_
timestamp 1644511149
transform 1 0 16376 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1372_
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1373_
timestamp 1644511149
transform 1 0 16100 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1374_
timestamp 1644511149
transform 1 0 16560 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1375_
timestamp 1644511149
transform 1 0 27140 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1376_
timestamp 1644511149
transform 1 0 19228 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1377_
timestamp 1644511149
transform 1 0 16008 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1378_
timestamp 1644511149
transform 1 0 15548 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1379_
timestamp 1644511149
transform 1 0 15732 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1380_
timestamp 1644511149
transform 1 0 17112 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1381_
timestamp 1644511149
transform 1 0 16284 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1382_
timestamp 1644511149
transform 1 0 16928 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1383_
timestamp 1644511149
transform 1 0 19228 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1384_
timestamp 1644511149
transform 1 0 18032 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1385_
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1386_
timestamp 1644511149
transform 1 0 16652 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1387_
timestamp 1644511149
transform 1 0 17296 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1388_
timestamp 1644511149
transform 1 0 17664 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1389_
timestamp 1644511149
transform 1 0 17296 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1390_
timestamp 1644511149
transform 1 0 14720 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1391_
timestamp 1644511149
transform 1 0 15088 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1392_
timestamp 1644511149
transform 1 0 15272 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1393_
timestamp 1644511149
transform 1 0 14720 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1394_
timestamp 1644511149
transform 1 0 18492 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1395_
timestamp 1644511149
transform 1 0 16652 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1396_
timestamp 1644511149
transform 1 0 16652 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1397_
timestamp 1644511149
transform 1 0 15548 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1398_
timestamp 1644511149
transform 1 0 16652 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1399_
timestamp 1644511149
transform 1 0 17296 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1400_
timestamp 1644511149
transform 1 0 18492 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1401_
timestamp 1644511149
transform 1 0 19504 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1402_
timestamp 1644511149
transform 1 0 21344 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1403_
timestamp 1644511149
transform 1 0 19228 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1404_
timestamp 1644511149
transform 1 0 18492 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1405_
timestamp 1644511149
transform 1 0 19872 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1406_
timestamp 1644511149
transform 1 0 22356 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1407_
timestamp 1644511149
transform 1 0 21804 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1408_
timestamp 1644511149
transform 1 0 22356 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1409_
timestamp 1644511149
transform 1 0 21804 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1410_
timestamp 1644511149
transform 1 0 21528 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1411_
timestamp 1644511149
transform 1 0 22080 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1412_
timestamp 1644511149
transform 1 0 23920 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1413_
timestamp 1644511149
transform 1 0 24104 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1414_
timestamp 1644511149
transform 1 0 24380 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1415_
timestamp 1644511149
transform 1 0 24288 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1416_
timestamp 1644511149
transform 1 0 24748 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1417_
timestamp 1644511149
transform 1 0 26588 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1418_
timestamp 1644511149
transform 1 0 27140 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1419_
timestamp 1644511149
transform 1 0 27232 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1420_
timestamp 1644511149
transform 1 0 29072 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1421_
timestamp 1644511149
transform 1 0 25668 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1422__9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6072 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1423__10
timestamp 1644511149
transform 1 0 1564 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1424__11
timestamp 1644511149
transform 1 0 15548 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1425__12
timestamp 1644511149
transform 1 0 2576 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1426__13
timestamp 1644511149
transform 1 0 28152 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1427__14
timestamp 1644511149
transform 1 0 5336 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1428__15
timestamp 1644511149
transform 1 0 30728 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1429__16
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1430__17
timestamp 1644511149
transform 1 0 11592 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1431__18
timestamp 1644511149
transform 1 0 13340 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1432__19
timestamp 1644511149
transform 1 0 32936 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1433__20
timestamp 1644511149
transform 1 0 17756 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1434__21
timestamp 1644511149
transform 1 0 12236 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1435__22
timestamp 1644511149
transform 1 0 4416 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1436__23
timestamp 1644511149
transform 1 0 12696 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1437__24
timestamp 1644511149
transform 1 0 9660 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1438__25
timestamp 1644511149
transform 1 0 31464 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1439__26
timestamp 1644511149
transform 1 0 11408 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1440__27
timestamp 1644511149
transform 1 0 5060 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1441__28
timestamp 1644511149
transform 1 0 29900 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1442__29
timestamp 1644511149
transform 1 0 2484 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1443__30
timestamp 1644511149
transform 1 0 10764 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1444__31
timestamp 1644511149
transform 1 0 11592 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1445__32
timestamp 1644511149
transform 1 0 10304 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1446__33
timestamp 1644511149
transform 1 0 31372 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1447__34
timestamp 1644511149
transform 1 0 6716 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1448__35
timestamp 1644511149
transform 1 0 33764 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1449__36
timestamp 1644511149
transform 1 0 3772 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1450__37
timestamp 1644511149
transform 1 0 32292 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1451__38
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1452__39
timestamp 1644511149
transform 1 0 32292 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1453__40
timestamp 1644511149
transform 1 0 12052 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1454__41
timestamp 1644511149
transform 1 0 11408 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1455__42
timestamp 1644511149
transform 1 0 12052 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1456__43
timestamp 1644511149
transform 1 0 4876 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1457__44
timestamp 1644511149
transform 1 0 1840 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1458__45
timestamp 1644511149
transform 1 0 30084 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1459__46
timestamp 1644511149
transform 1 0 11408 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1460__47
timestamp 1644511149
transform 1 0 10764 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1461__48
timestamp 1644511149
transform 1 0 1656 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1462__49
timestamp 1644511149
transform 1 0 14352 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1463__50
timestamp 1644511149
transform 1 0 1656 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1464__51
timestamp 1644511149
transform 1 0 32936 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1465__52
timestamp 1644511149
transform 1 0 2576 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1466__53
timestamp 1644511149
transform 1 0 4324 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1467__54
timestamp 1644511149
transform 1 0 30084 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1468__55
timestamp 1644511149
transform 1 0 10120 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1469__56
timestamp 1644511149
transform 1 0 33764 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1470__57
timestamp 1644511149
transform 1 0 1472 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1471__58
timestamp 1644511149
transform 1 0 10764 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1472__59
timestamp 1644511149
transform 1 0 1472 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1473__60
timestamp 1644511149
transform 1 0 24380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1474__61
timestamp 1644511149
transform 1 0 30820 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1475__62
timestamp 1644511149
transform 1 0 21068 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1476__63
timestamp 1644511149
transform 1 0 10672 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1477__64
timestamp 1644511149
transform 1 0 5520 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1478__65
timestamp 1644511149
transform 1 0 10120 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1479__66
timestamp 1644511149
transform 1 0 12972 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1480__67
timestamp 1644511149
transform 1 0 31004 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1481__68
timestamp 1644511149
transform 1 0 4968 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1482__69
timestamp 1644511149
transform 1 0 2484 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1483__70
timestamp 1644511149
transform 1 0 2208 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1484__71
timestamp 1644511149
transform 1 0 33764 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1485__72
timestamp 1644511149
transform 1 0 12696 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1486__73
timestamp 1644511149
transform 1 0 12052 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1487__74
timestamp 1644511149
transform 1 0 8924 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1488__75
timestamp 1644511149
transform 1 0 10028 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1489__76
timestamp 1644511149
transform 1 0 20148 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1490__77
timestamp 1644511149
transform 1 0 28428 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1491__78
timestamp 1644511149
transform 1 0 9476 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1492__79
timestamp 1644511149
transform 1 0 19504 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1493__80
timestamp 1644511149
transform 1 0 30360 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1494__81
timestamp 1644511149
transform 1 0 1840 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1495__82
timestamp 1644511149
transform 1 0 30728 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1496__83
timestamp 1644511149
transform 1 0 6532 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1497__84
timestamp 1644511149
transform 1 0 6992 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1498__85
timestamp 1644511149
transform 1 0 7820 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1499__86
timestamp 1644511149
transform 1 0 3220 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1500__87
timestamp 1644511149
transform 1 0 30176 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1501__88
timestamp 1644511149
transform 1 0 32384 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1502__89
timestamp 1644511149
transform 1 0 31372 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1503__90
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1504__91
timestamp 1644511149
transform 1 0 7176 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1505__92
timestamp 1644511149
transform 1 0 33764 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1506__93
timestamp 1644511149
transform 1 0 11868 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1507__94
timestamp 1644511149
transform 1 0 8188 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1508__95
timestamp 1644511149
transform 1 0 7912 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1509__96
timestamp 1644511149
transform 1 0 29440 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1510__97
timestamp 1644511149
transform 1 0 6348 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1511__98
timestamp 1644511149
transform 1 0 3864 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1512__99
timestamp 1644511149
transform 1 0 10120 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1513__100
timestamp 1644511149
transform 1 0 9384 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1514__101
timestamp 1644511149
transform 1 0 27508 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1515__102
timestamp 1644511149
transform 1 0 12052 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1516__103
timestamp 1644511149
transform 1 0 11868 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1517__104
timestamp 1644511149
transform 1 0 31372 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1518__105
timestamp 1644511149
transform 1 0 13340 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1519__106
timestamp 1644511149
transform 1 0 4416 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1520__107
timestamp 1644511149
transform 1 0 31648 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1521__108
timestamp 1644511149
transform 1 0 1748 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1522__109
timestamp 1644511149
transform 1 0 33120 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1523__110
timestamp 1644511149
transform 1 0 5612 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1524__111
timestamp 1644511149
transform 1 0 2392 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1525__112
timestamp 1644511149
transform 1 0 2392 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1526__113
timestamp 1644511149
transform 1 0 2576 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1527_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1528_
timestamp 1644511149
transform 1 0 1380 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1529_
timestamp 1644511149
transform 1 0 15456 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1530_
timestamp 1644511149
transform 1 0 1564 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1531_
timestamp 1644511149
transform 1 0 30452 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1532_
timestamp 1644511149
transform 1 0 2300 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1533_
timestamp 1644511149
transform 1 0 32292 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1534_
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1535_
timestamp 1644511149
transform 1 0 32292 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1536_
timestamp 1644511149
transform 1 0 32292 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1537_
timestamp 1644511149
transform 1 0 32292 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1538_
timestamp 1644511149
transform 1 0 16836 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1539_
timestamp 1644511149
transform 1 0 32292 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1540_
timestamp 1644511149
transform 1 0 1472 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1541_
timestamp 1644511149
transform 1 0 17480 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1542_
timestamp 1644511149
transform 1 0 9108 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1543_
timestamp 1644511149
transform 1 0 32292 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1544_
timestamp 1644511149
transform 1 0 32292 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1545_
timestamp 1644511149
transform 1 0 1380 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1546_
timestamp 1644511149
transform 1 0 32292 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1547_
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1548_
timestamp 1644511149
transform 1 0 32292 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1549_
timestamp 1644511149
transform 1 0 20056 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1550_
timestamp 1644511149
transform 1 0 9568 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1551_
timestamp 1644511149
transform 1 0 32292 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1552_
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1553_
timestamp 1644511149
transform 1 0 32292 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1554_
timestamp 1644511149
transform 1 0 2116 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1555_
timestamp 1644511149
transform 1 0 32292 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1556_
timestamp 1644511149
transform 1 0 3864 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1557_
timestamp 1644511149
transform 1 0 32292 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1558_
timestamp 1644511149
transform 1 0 32292 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1559_
timestamp 1644511149
transform 1 0 32292 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1560_
timestamp 1644511149
transform 1 0 22172 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1561_
timestamp 1644511149
transform 1 0 4416 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1562_
timestamp 1644511149
transform 1 0 1380 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1563_
timestamp 1644511149
transform 1 0 32292 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1564_
timestamp 1644511149
transform 1 0 14168 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1565_
timestamp 1644511149
transform 1 0 32292 0 -1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1566_
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1567_
timestamp 1644511149
transform 1 0 14260 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1568_
timestamp 1644511149
transform 1 0 1564 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1569_
timestamp 1644511149
transform 1 0 32292 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1570_
timestamp 1644511149
transform 1 0 1748 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1571_
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1572_
timestamp 1644511149
transform 1 0 29808 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1573_
timestamp 1644511149
transform 1 0 32292 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1574_
timestamp 1644511149
transform 1 0 27508 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1575_
timestamp 1644511149
transform 1 0 32292 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1576_
timestamp 1644511149
transform 1 0 32108 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1577_
timestamp 1644511149
transform 1 0 32292 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1578_
timestamp 1644511149
transform 1 0 1472 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1579_
timestamp 1644511149
transform 1 0 27692 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1580_
timestamp 1644511149
transform 1 0 1472 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1581_
timestamp 1644511149
transform 1 0 23828 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1582_
timestamp 1644511149
transform 1 0 32292 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1583_
timestamp 1644511149
transform 1 0 20792 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1584_
timestamp 1644511149
transform 1 0 25116 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1585_
timestamp 1644511149
transform 1 0 5152 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1586_
timestamp 1644511149
transform 1 0 26956 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1587_
timestamp 1644511149
transform 1 0 11960 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1588_
timestamp 1644511149
transform 1 0 32292 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1589_
timestamp 1644511149
transform 1 0 2576 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1590_
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1591_
timestamp 1644511149
transform 1 0 1380 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1592_
timestamp 1644511149
transform 1 0 32292 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1593_
timestamp 1644511149
transform 1 0 32292 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1594_
timestamp 1644511149
transform 1 0 32292 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1595_
timestamp 1644511149
transform 1 0 8556 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1596_
timestamp 1644511149
transform 1 0 29716 0 -1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1597_
timestamp 1644511149
transform 1 0 19412 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1598_
timestamp 1644511149
transform 1 0 29624 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1599_
timestamp 1644511149
transform 1 0 29532 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1600_
timestamp 1644511149
transform 1 0 19412 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1601_
timestamp 1644511149
transform 1 0 32108 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1602_
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1603_
timestamp 1644511149
transform 1 0 32292 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1604_
timestamp 1644511149
transform 1 0 6532 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1605_
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1606_
timestamp 1644511149
transform 1 0 7728 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1607_
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1608_
timestamp 1644511149
transform 1 0 32292 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1609_
timestamp 1644511149
transform 1 0 32292 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1610_
timestamp 1644511149
transform 1 0 32292 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1611_
timestamp 1644511149
transform 1 0 2024 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1612_
timestamp 1644511149
transform 1 0 7176 0 -1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1613_
timestamp 1644511149
transform 1 0 32292 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1614_
timestamp 1644511149
transform 1 0 9108 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1615_
timestamp 1644511149
transform 1 0 24472 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1616_
timestamp 1644511149
transform 1 0 8924 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1617_
timestamp 1644511149
transform 1 0 32292 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1618_
timestamp 1644511149
transform 1 0 3772 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1619_
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1620_
timestamp 1644511149
transform 1 0 15456 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1621_
timestamp 1644511149
transform 1 0 16652 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1622_
timestamp 1644511149
transform 1 0 32292 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1623_
timestamp 1644511149
transform 1 0 32292 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1624_
timestamp 1644511149
transform 1 0 19412 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1625_
timestamp 1644511149
transform 1 0 29716 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1626_
timestamp 1644511149
transform 1 0 32292 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1627_
timestamp 1644511149
transform 1 0 2576 0 -1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1628_
timestamp 1644511149
transform 1 0 31648 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1629_
timestamp 1644511149
transform 1 0 1748 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1630_
timestamp 1644511149
transform 1 0 29716 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1631_
timestamp 1644511149
transform 1 0 4232 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1632_
timestamp 1644511149
transform 1 0 1472 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1633_
timestamp 1644511149
transform 1 0 1472 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1634_
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24748 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_wb_clk_i
timestamp 1644511149
transform 1 0 14996 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 15824 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_0_0_wb_clk_i
timestamp 1644511149
transform 1 0 15088 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 31372 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_2_0_wb_clk_i
timestamp 1644511149
transform 1 0 15364 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_3_0_wb_clk_i
timestamp 1644511149
transform 1 0 15088 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_0_0_wb_clk_i
timestamp 1644511149
transform 1 0 15364 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_2_0_wb_clk_i
timestamp 1644511149
transform 1 0 30820 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_3_0_wb_clk_i
timestamp 1644511149
transform 1 0 32108 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_4_0_wb_clk_i
timestamp 1644511149
transform 1 0 14536 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_5_0_wb_clk_i
timestamp 1644511149
transform 1 0 18400 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_6_0_wb_clk_i
timestamp 1644511149
transform 1 0 14628 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_7_0_wb_clk_i
timestamp 1644511149
transform 1 0 24380 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input1
timestamp 1644511149
transform 1 0 1380 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1644511149
transform 1 0 10764 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input3
timestamp 1644511149
transform 1 0 1380 0 1 39168
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input4
timestamp 1644511149
transform 1 0 33304 0 -1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1644511149
transform 1 0 18124 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1644511149
transform -1 0 12236 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1644511149
transform 1 0 4968 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1644511149
transform 1 0 33856 0 1 9792
box -38 -48 406 592
<< labels >>
rlabel metal3 s 0 35988 800 36228 6 active
port 0 nsew signal input
rlabel metal2 s 11582 0 11694 800 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 18666 41200 18778 42000 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 0 38708 800 38948 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 35200 35988 36000 36228 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 18022 0 18134 800 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 11582 41200 11694 42000 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 35200 37348 36000 37588 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 35200 6068 36000 6308 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 5142 41200 5254 42000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 6430 41200 6542 42000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 33478 0 33590 800 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 0 12188 800 12428 6 io_in[1]
port 12 nsew signal input
rlabel metal3 s 0 22388 800 22628 6 io_in[20]
port 13 nsew signal input
rlabel metal3 s 0 14908 800 15148 6 io_in[21]
port 14 nsew signal input
rlabel metal3 s 35200 15588 36000 15828 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 4498 41200 4610 42000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 1922 41200 2034 42000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 28970 0 29082 800 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 28326 0 28438 800 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 35200 11508 36000 11748 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 25750 0 25862 800 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 35410 41200 35522 42000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 12870 0 12982 800 6 io_in[2]
port 23 nsew signal input
rlabel metal3 s 35200 18308 36000 18548 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 0 34628 800 34868 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 23818 0 23930 800 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 0 20348 800 20588 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 26394 41200 26506 42000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 30902 41200 31014 42000 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 35200 27148 36000 27388 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 31546 41200 31658 42000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 19310 41200 19422 42000 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 35200 26468 36000 26708 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 35200 40068 36000 40308 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 0 23748 800 23988 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 0 16268 800 16508 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 35200 29188 36000 29428 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 3210 41200 3322 42000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 20598 0 20710 800 6 io_oeb[0]
port 39 nsew signal tristate
rlabel metal3 s 0 13548 800 13788 6 io_oeb[10]
port 40 nsew signal tristate
rlabel metal3 s 35200 25108 36000 25348 6 io_oeb[11]
port 41 nsew signal tristate
rlabel metal3 s 35200 14228 36000 14468 6 io_oeb[12]
port 42 nsew signal tristate
rlabel metal3 s 35200 13548 36000 13788 6 io_oeb[13]
port 43 nsew signal tristate
rlabel metal3 s 0 3348 800 3588 6 io_oeb[14]
port 44 nsew signal tristate
rlabel metal2 s 7718 41200 7830 42000 6 io_oeb[15]
port 45 nsew signal tristate
rlabel metal3 s 35200 4708 36000 4948 6 io_oeb[16]
port 46 nsew signal tristate
rlabel metal2 s 10294 0 10406 800 6 io_oeb[17]
port 47 nsew signal tristate
rlabel metal2 s 25106 41200 25218 42000 6 io_oeb[18]
port 48 nsew signal tristate
rlabel metal2 s 8362 41200 8474 42000 6 io_oeb[19]
port 49 nsew signal tristate
rlabel metal2 s 30258 0 30370 800 6 io_oeb[1]
port 50 nsew signal tristate
rlabel metal3 s 35200 19668 36000 19908 6 io_oeb[20]
port 51 nsew signal tristate
rlabel metal3 s 0 40748 800 40988 6 io_oeb[21]
port 52 nsew signal tristate
rlabel metal2 s 3854 0 3966 800 6 io_oeb[22]
port 53 nsew signal tristate
rlabel metal2 s 16090 41200 16202 42000 6 io_oeb[23]
port 54 nsew signal tristate
rlabel metal2 s 17378 41200 17490 42000 6 io_oeb[24]
port 55 nsew signal tristate
rlabel metal3 s 35200 628 36000 868 6 io_oeb[25]
port 56 nsew signal tristate
rlabel metal3 s 35200 33268 36000 33508 6 io_oeb[26]
port 57 nsew signal tristate
rlabel metal2 s 19954 41200 20066 42000 6 io_oeb[27]
port 58 nsew signal tristate
rlabel metal2 s 32834 0 32946 800 6 io_oeb[28]
port 59 nsew signal tristate
rlabel metal3 s 35200 27828 36000 28068 6 io_oeb[29]
port 60 nsew signal tristate
rlabel metal2 s 28970 41200 29082 42000 6 io_oeb[2]
port 61 nsew signal tristate
rlabel metal3 s 0 41428 800 41668 6 io_oeb[30]
port 62 nsew signal tristate
rlabel metal2 s 32190 0 32302 800 6 io_oeb[31]
port 63 nsew signal tristate
rlabel metal3 s 0 18988 800 19228 6 io_oeb[32]
port 64 nsew signal tristate
rlabel metal3 s 35200 1988 36000 2228 6 io_oeb[33]
port 65 nsew signal tristate
rlabel metal2 s 5786 41200 5898 42000 6 io_oeb[34]
port 66 nsew signal tristate
rlabel metal3 s 0 16948 800 17188 6 io_oeb[35]
port 67 nsew signal tristate
rlabel metal3 s 0 8788 800 9028 6 io_oeb[36]
port 68 nsew signal tristate
rlabel metal3 s 0 14228 800 14468 6 io_oeb[37]
port 69 nsew signal tristate
rlabel metal2 s 19954 0 20066 800 6 io_oeb[3]
port 70 nsew signal tristate
rlabel metal3 s 35200 3348 36000 3588 6 io_oeb[4]
port 71 nsew signal tristate
rlabel metal3 s 0 25108 800 25348 6 io_oeb[5]
port 72 nsew signal tristate
rlabel metal3 s 35200 16948 36000 17188 6 io_oeb[6]
port 73 nsew signal tristate
rlabel metal2 s 7074 41200 7186 42000 6 io_oeb[7]
port 74 nsew signal tristate
rlabel metal2 s 3210 0 3322 800 6 io_oeb[8]
port 75 nsew signal tristate
rlabel metal2 s 8362 0 8474 800 6 io_oeb[9]
port 76 nsew signal tristate
rlabel metal3 s 35200 39388 36000 39628 6 io_out[0]
port 77 nsew signal tristate
rlabel metal3 s 35200 24428 36000 24668 6 io_out[10]
port 78 nsew signal tristate
rlabel metal3 s 0 1988 800 2228 6 io_out[11]
port 79 nsew signal tristate
rlabel metal3 s 0 5388 800 5628 6 io_out[12]
port 80 nsew signal tristate
rlabel metal2 s 30902 0 31014 800 6 io_out[13]
port 81 nsew signal tristate
rlabel metal3 s 35200 33948 36000 34188 6 io_out[14]
port 82 nsew signal tristate
rlabel metal3 s 0 31908 800 32148 6 io_out[15]
port 83 nsew signal tristate
rlabel metal3 s 35200 23748 36000 23988 6 io_out[16]
port 84 nsew signal tristate
rlabel metal2 s 32834 41200 32946 42000 6 io_out[17]
port 85 nsew signal tristate
rlabel metal3 s 35200 -52 36000 188 6 io_out[18]
port 86 nsew signal tristate
rlabel metal3 s 0 18308 800 18548 6 io_out[19]
port 87 nsew signal tristate
rlabel metal2 s 22530 41200 22642 42000 6 io_out[1]
port 88 nsew signal tristate
rlabel metal2 s 28326 41200 28438 42000 6 io_out[20]
port 89 nsew signal tristate
rlabel metal3 s 0 31228 800 31468 6 io_out[21]
port 90 nsew signal tristate
rlabel metal2 s 24462 0 24574 800 6 io_out[22]
port 91 nsew signal tristate
rlabel metal3 s 35200 20348 36000 20588 6 io_out[23]
port 92 nsew signal tristate
rlabel metal2 s 21242 0 21354 800 6 io_out[24]
port 93 nsew signal tristate
rlabel metal2 s 25750 41200 25862 42000 6 io_out[25]
port 94 nsew signal tristate
rlabel metal3 s 0 4028 800 4268 6 io_out[26]
port 95 nsew signal tristate
rlabel metal2 s 27038 41200 27150 42000 6 io_out[27]
port 96 nsew signal tristate
rlabel metal2 s 13514 0 13626 800 6 io_out[28]
port 97 nsew signal tristate
rlabel metal3 s 35200 4028 36000 4268 6 io_out[29]
port 98 nsew signal tristate
rlabel metal2 s 5142 0 5254 800 6 io_out[2]
port 99 nsew signal tristate
rlabel metal3 s 0 4708 800 4948 6 io_out[30]
port 100 nsew signal tristate
rlabel metal3 s 0 10828 800 11068 6 io_out[31]
port 101 nsew signal tristate
rlabel metal3 s 0 36668 800 36908 6 io_out[32]
port 102 nsew signal tristate
rlabel metal3 s 35200 8788 36000 9028 6 io_out[33]
port 103 nsew signal tristate
rlabel metal3 s 35200 34628 36000 34868 6 io_out[34]
port 104 nsew signal tristate
rlabel metal3 s 35200 32588 36000 32828 6 io_out[35]
port 105 nsew signal tristate
rlabel metal2 s 9006 41200 9118 42000 6 io_out[36]
port 106 nsew signal tristate
rlabel metal3 s 35200 38028 36000 38268 6 io_out[37]
port 107 nsew signal tristate
rlabel metal3 s 0 33948 800 34188 6 io_out[3]
port 108 nsew signal tristate
rlabel metal3 s 35200 25788 36000 26028 6 io_out[4]
port 109 nsew signal tristate
rlabel metal2 s 14802 41200 14914 42000 6 io_out[5]
port 110 nsew signal tristate
rlabel metal2 s 34122 41200 34234 42000 6 io_out[6]
port 111 nsew signal tristate
rlabel metal3 s 0 15588 800 15828 6 io_out[7]
port 112 nsew signal tristate
rlabel metal2 s 14802 0 14914 800 6 io_out[8]
port 113 nsew signal tristate
rlabel metal3 s 0 11508 800 11748 6 io_out[9]
port 114 nsew signal tristate
rlabel metal3 s 35200 9468 36000 9708 6 la1_data_in[0]
port 115 nsew signal input
rlabel metal2 s 16734 0 16846 800 6 la1_data_in[10]
port 116 nsew signal input
rlabel metal3 s 35200 7428 36000 7668 6 la1_data_in[11]
port 117 nsew signal input
rlabel metal3 s 0 29188 800 29428 6 la1_data_in[12]
port 118 nsew signal input
rlabel metal2 s 26394 0 26506 800 6 la1_data_in[13]
port 119 nsew signal input
rlabel metal3 s 0 10148 800 10388 6 la1_data_in[14]
port 120 nsew signal input
rlabel metal2 s 9650 41200 9762 42000 6 la1_data_in[15]
port 121 nsew signal input
rlabel metal2 s 21242 41200 21354 42000 6 la1_data_in[16]
port 122 nsew signal input
rlabel metal2 s 15446 41200 15558 42000 6 la1_data_in[17]
port 123 nsew signal input
rlabel metal2 s 34122 0 34234 800 6 la1_data_in[18]
port 124 nsew signal input
rlabel metal2 s 10938 41200 11050 42000 6 la1_data_in[19]
port 125 nsew signal input
rlabel metal2 s 15446 0 15558 800 6 la1_data_in[1]
port 126 nsew signal input
rlabel metal3 s 0 28508 800 28748 6 la1_data_in[20]
port 127 nsew signal input
rlabel metal2 s 34766 41200 34878 42000 6 la1_data_in[21]
port 128 nsew signal input
rlabel metal3 s 35200 10148 36000 10388 6 la1_data_in[22]
port 129 nsew signal input
rlabel metal3 s 0 628 800 868 6 la1_data_in[23]
port 130 nsew signal input
rlabel metal2 s 10938 0 11050 800 6 la1_data_in[24]
port 131 nsew signal input
rlabel metal3 s 0 29868 800 30108 6 la1_data_in[25]
port 132 nsew signal input
rlabel metal3 s 35200 5388 36000 5628 6 la1_data_in[26]
port 133 nsew signal input
rlabel metal2 s 22530 0 22642 800 6 la1_data_in[27]
port 134 nsew signal input
rlabel metal3 s 0 25788 800 26028 6 la1_data_in[28]
port 135 nsew signal input
rlabel metal3 s 0 39388 800 39628 6 la1_data_in[29]
port 136 nsew signal input
rlabel metal2 s 9006 0 9118 800 6 la1_data_in[2]
port 137 nsew signal input
rlabel metal2 s 1278 0 1390 800 6 la1_data_in[30]
port 138 nsew signal input
rlabel metal2 s 29614 0 29726 800 6 la1_data_in[31]
port 139 nsew signal input
rlabel metal3 s 0 24428 800 24668 6 la1_data_in[3]
port 140 nsew signal input
rlabel metal2 s 30258 41200 30370 42000 6 la1_data_in[4]
port 141 nsew signal input
rlabel metal3 s 35200 22388 36000 22628 6 la1_data_in[5]
port 142 nsew signal input
rlabel metal2 s 12226 41200 12338 42000 6 la1_data_in[6]
port 143 nsew signal input
rlabel metal3 s 0 17628 800 17868 6 la1_data_in[7]
port 144 nsew signal input
rlabel metal2 s 12870 41200 12982 42000 6 la1_data_in[8]
port 145 nsew signal input
rlabel metal3 s 0 27148 800 27388 6 la1_data_in[9]
port 146 nsew signal input
rlabel metal2 s 6430 0 6542 800 6 la1_data_out[0]
port 147 nsew signal tristate
rlabel metal3 s 35200 12188 36000 12428 6 la1_data_out[10]
port 148 nsew signal tristate
rlabel metal2 s 17378 0 17490 800 6 la1_data_out[11]
port 149 nsew signal tristate
rlabel metal3 s 35200 38708 36000 38948 6 la1_data_out[12]
port 150 nsew signal tristate
rlabel metal2 s 634 41200 746 42000 6 la1_data_out[13]
port 151 nsew signal tristate
rlabel metal2 s 18022 41200 18134 42000 6 la1_data_out[14]
port 152 nsew signal tristate
rlabel metal3 s 0 1308 800 1548 6 la1_data_out[15]
port 153 nsew signal tristate
rlabel metal3 s 35200 16268 36000 16508 6 la1_data_out[16]
port 154 nsew signal tristate
rlabel metal3 s 35200 31228 36000 31468 6 la1_data_out[17]
port 155 nsew signal tristate
rlabel metal2 s 1278 41200 1390 42000 6 la1_data_out[18]
port 156 nsew signal tristate
rlabel metal3 s 35200 23068 36000 23308 6 la1_data_out[19]
port 157 nsew signal tristate
rlabel metal3 s 0 35308 800 35548 6 la1_data_out[1]
port 158 nsew signal tristate
rlabel metal3 s 0 8108 800 8348 6 la1_data_out[20]
port 159 nsew signal tristate
rlabel metal3 s 35200 36668 36000 36908 6 la1_data_out[21]
port 160 nsew signal tristate
rlabel metal2 s 20598 41200 20710 42000 6 la1_data_out[22]
port 161 nsew signal tristate
rlabel metal2 s 9650 0 9762 800 6 la1_data_out[23]
port 162 nsew signal tristate
rlabel metal3 s 35200 17628 36000 17868 6 la1_data_out[24]
port 163 nsew signal tristate
rlabel metal3 s 0 2668 800 2908 6 la1_data_out[25]
port 164 nsew signal tristate
rlabel metal3 s 35200 6748 36000 6988 6 la1_data_out[26]
port 165 nsew signal tristate
rlabel metal3 s 0 37348 800 37588 6 la1_data_out[27]
port 166 nsew signal tristate
rlabel metal2 s 34766 0 34878 800 6 la1_data_out[28]
port 167 nsew signal tristate
rlabel metal2 s 4498 0 4610 800 6 la1_data_out[29]
port 168 nsew signal tristate
rlabel metal2 s 16090 0 16202 800 6 la1_data_out[2]
port 169 nsew signal tristate
rlabel metal3 s 35200 12868 36000 13108 6 la1_data_out[30]
port 170 nsew signal tristate
rlabel metal3 s 35200 40748 36000 40988 6 la1_data_out[31]
port 171 nsew signal tristate
rlabel metal3 s 0 7428 800 7668 6 la1_data_out[3]
port 172 nsew signal tristate
rlabel metal2 s 35410 0 35522 800 6 la1_data_out[4]
port 173 nsew signal tristate
rlabel metal2 s 2566 0 2678 800 6 la1_data_out[5]
port 174 nsew signal tristate
rlabel metal3 s 35200 18988 36000 19228 6 la1_data_out[6]
port 175 nsew signal tristate
rlabel metal2 s 634 0 746 800 6 la1_data_out[7]
port 176 nsew signal tristate
rlabel metal3 s 35200 31908 36000 32148 6 la1_data_out[8]
port 177 nsew signal tristate
rlabel metal2 s 33478 41200 33590 42000 6 la1_data_out[9]
port 178 nsew signal tristate
rlabel metal3 s 35200 2668 36000 2908 6 la1_oenb[0]
port 179 nsew signal input
rlabel metal2 s 32190 41200 32302 42000 6 la1_oenb[10]
port 180 nsew signal input
rlabel metal3 s 0 21708 800 21948 6 la1_oenb[11]
port 181 nsew signal input
rlabel metal3 s 0 23068 800 23308 6 la1_oenb[12]
port 182 nsew signal input
rlabel metal2 s 23174 0 23286 800 6 la1_oenb[13]
port 183 nsew signal input
rlabel metal2 s -10 0 102 800 6 la1_oenb[14]
port 184 nsew signal input
rlabel metal2 s 27682 0 27794 800 6 la1_oenb[15]
port 185 nsew signal input
rlabel metal3 s 0 27828 800 28068 6 la1_oenb[16]
port 186 nsew signal input
rlabel metal2 s -10 41200 102 42000 6 la1_oenb[17]
port 187 nsew signal input
rlabel metal2 s 14158 41200 14270 42000 6 la1_oenb[18]
port 188 nsew signal input
rlabel metal3 s 0 21028 800 21268 6 la1_oenb[19]
port 189 nsew signal input
rlabel metal2 s 7074 0 7186 800 6 la1_oenb[1]
port 190 nsew signal input
rlabel metal2 s 1922 0 2034 800 6 la1_oenb[20]
port 191 nsew signal input
rlabel metal2 s 21886 41200 21998 42000 6 la1_oenb[21]
port 192 nsew signal input
rlabel metal2 s 13514 41200 13626 42000 6 la1_oenb[22]
port 193 nsew signal input
rlabel metal2 s 19310 0 19422 800 6 la1_oenb[23]
port 194 nsew signal input
rlabel metal2 s 27682 41200 27794 42000 6 la1_oenb[24]
port 195 nsew signal input
rlabel metal3 s 35200 10828 36000 11068 6 la1_oenb[25]
port 196 nsew signal input
rlabel metal3 s 0 30548 800 30788 6 la1_oenb[26]
port 197 nsew signal input
rlabel metal3 s 35200 30548 36000 30788 6 la1_oenb[27]
port 198 nsew signal input
rlabel metal2 s 7718 0 7830 800 6 la1_oenb[28]
port 199 nsew signal input
rlabel metal2 s 14158 0 14270 800 6 la1_oenb[29]
port 200 nsew signal input
rlabel metal3 s 0 6748 800 6988 6 la1_oenb[2]
port 201 nsew signal input
rlabel metal3 s 35200 29868 36000 30108 6 la1_oenb[30]
port 202 nsew signal input
rlabel metal2 s 21886 0 21998 800 6 la1_oenb[31]
port 203 nsew signal input
rlabel metal2 s 24462 41200 24574 42000 6 la1_oenb[3]
port 204 nsew signal input
rlabel metal2 s 23818 41200 23930 42000 6 la1_oenb[4]
port 205 nsew signal input
rlabel metal3 s 0 38028 800 38268 6 la1_oenb[5]
port 206 nsew signal input
rlabel metal2 s 2566 41200 2678 42000 6 la1_oenb[6]
port 207 nsew signal input
rlabel metal2 s 27038 0 27150 800 6 la1_oenb[7]
port 208 nsew signal input
rlabel metal3 s 0 9468 800 9708 6 la1_oenb[8]
port 209 nsew signal input
rlabel metal3 s 0 32588 800 32828 6 la1_oenb[9]
port 210 nsew signal input
rlabel metal4 s 6576 2128 6896 39760 6 vccd1
port 211 nsew power input
rlabel metal4 s 17840 2128 18160 39760 6 vccd1
port 211 nsew power input
rlabel metal4 s 29104 2128 29424 39760 6 vccd1
port 211 nsew power input
rlabel metal4 s 12208 2128 12528 39760 6 vssd1
port 212 nsew ground input
rlabel metal4 s 23472 2128 23792 39760 6 vssd1
port 212 nsew ground input
rlabel metal3 s 35200 21028 36000 21268 6 wb_clk_i
port 213 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 36000 42000
<< end >>
