always @(*) begin
    if(active) begin
        // active properties here
    end
    if(!active) begin
        // inactive properties here
    end
end
